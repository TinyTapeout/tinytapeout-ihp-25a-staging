module tt_um_murmann_group (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire \my_decimation_filter.Y[0] ;
 wire \my_decimation_filter.Y[10] ;
 wire \my_decimation_filter.Y[11] ;
 wire \my_decimation_filter.Y[12] ;
 wire \my_decimation_filter.Y[13] ;
 wire \my_decimation_filter.Y[14] ;
 wire \my_decimation_filter.Y[15] ;
 wire \my_decimation_filter.Y[1] ;
 wire \my_decimation_filter.Y[2] ;
 wire \my_decimation_filter.Y[3] ;
 wire \my_decimation_filter.Y[4] ;
 wire \my_decimation_filter.Y[5] ;
 wire \my_decimation_filter.Y[6] ;
 wire \my_decimation_filter.Y[7] ;
 wire \my_decimation_filter.Y[8] ;
 wire \my_decimation_filter.Y[9] ;
 wire \my_decimation_filter.comb_1[0] ;
 wire \my_decimation_filter.comb_1[10] ;
 wire \my_decimation_filter.comb_1[11] ;
 wire \my_decimation_filter.comb_1[12] ;
 wire \my_decimation_filter.comb_1[13] ;
 wire \my_decimation_filter.comb_1[14] ;
 wire \my_decimation_filter.comb_1[15] ;
 wire \my_decimation_filter.comb_1[1] ;
 wire \my_decimation_filter.comb_1[2] ;
 wire \my_decimation_filter.comb_1[3] ;
 wire \my_decimation_filter.comb_1[4] ;
 wire \my_decimation_filter.comb_1[5] ;
 wire \my_decimation_filter.comb_1[6] ;
 wire \my_decimation_filter.comb_1[7] ;
 wire \my_decimation_filter.comb_1[8] ;
 wire \my_decimation_filter.comb_1[9] ;
 wire \my_decimation_filter.comb_2[0] ;
 wire \my_decimation_filter.comb_2[10] ;
 wire \my_decimation_filter.comb_2[11] ;
 wire \my_decimation_filter.comb_2[12] ;
 wire \my_decimation_filter.comb_2[13] ;
 wire \my_decimation_filter.comb_2[14] ;
 wire \my_decimation_filter.comb_2[15] ;
 wire \my_decimation_filter.comb_2[1] ;
 wire \my_decimation_filter.comb_2[2] ;
 wire \my_decimation_filter.comb_2[3] ;
 wire \my_decimation_filter.comb_2[4] ;
 wire \my_decimation_filter.comb_2[5] ;
 wire \my_decimation_filter.comb_2[6] ;
 wire \my_decimation_filter.comb_2[7] ;
 wire \my_decimation_filter.comb_2[8] ;
 wire \my_decimation_filter.comb_2[9] ;
 wire \my_decimation_filter.decimation_count[0] ;
 wire \my_decimation_filter.decimation_count[1] ;
 wire \my_decimation_filter.decimation_count[2] ;
 wire \my_decimation_filter.decimation_count[3] ;
 wire \my_decimation_filter.decimation_count[4] ;
 wire \my_decimation_filter.decimation_count[5] ;
 wire \my_decimation_filter.decimation_count[6] ;
 wire \my_decimation_filter.input_accumulator[0] ;
 wire \my_decimation_filter.input_accumulator[10] ;
 wire \my_decimation_filter.input_accumulator[11] ;
 wire \my_decimation_filter.input_accumulator[12] ;
 wire \my_decimation_filter.input_accumulator[13] ;
 wire \my_decimation_filter.input_accumulator[14] ;
 wire \my_decimation_filter.input_accumulator[15] ;
 wire \my_decimation_filter.input_accumulator[1] ;
 wire \my_decimation_filter.input_accumulator[2] ;
 wire \my_decimation_filter.input_accumulator[3] ;
 wire \my_decimation_filter.input_accumulator[4] ;
 wire \my_decimation_filter.input_accumulator[5] ;
 wire \my_decimation_filter.input_accumulator[6] ;
 wire \my_decimation_filter.input_accumulator[7] ;
 wire \my_decimation_filter.input_accumulator[8] ;
 wire \my_decimation_filter.input_accumulator[9] ;
 wire \my_decimation_filter.reset_d ;
 wire \my_decimation_filter.type_dec_d ;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire clknet_0_clk;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;

 sg13g2_inv_1 _0577_ (.Y(_0094_),
    .A(net184));
 sg13g2_inv_1 _0578_ (.Y(_0095_),
    .A(net157));
 sg13g2_inv_1 _0579_ (.Y(_0096_),
    .A(net219));
 sg13g2_inv_1 _0580_ (.Y(_0097_),
    .A(net244));
 sg13g2_inv_1 _0581_ (.Y(_0098_),
    .A(net257));
 sg13g2_inv_1 _0582_ (.Y(_0099_),
    .A(net199));
 sg13g2_inv_1 _0583_ (.Y(_0100_),
    .A(net249));
 sg13g2_inv_1 _0584_ (.Y(_0101_),
    .A(net210));
 sg13g2_inv_1 _0585_ (.Y(_0102_),
    .A(net246));
 sg13g2_inv_1 _0586_ (.Y(_0103_),
    .A(net213));
 sg13g2_inv_1 _0587_ (.Y(_0104_),
    .A(net171));
 sg13g2_inv_1 _0588_ (.Y(_0105_),
    .A(net228));
 sg13g2_inv_1 _0589_ (.Y(_0106_),
    .A(net241));
 sg13g2_inv_1 _0590_ (.Y(_0107_),
    .A(net252));
 sg13g2_inv_1 _0591_ (.Y(_0108_),
    .A(net174));
 sg13g2_inv_1 _0592_ (.Y(_0109_),
    .A(net254));
 sg13g2_inv_1 _0593_ (.Y(_0110_),
    .A(net215));
 sg13g2_inv_1 _0594_ (.Y(_0111_),
    .A(net226));
 sg13g2_inv_1 _0595_ (.Y(_0112_),
    .A(net159));
 sg13g2_inv_1 _0596_ (.Y(_0113_),
    .A(\my_decimation_filter.comb_2[13] ));
 sg13g2_inv_1 _0597_ (.Y(_0114_),
    .A(\my_decimation_filter.comb_2[11] ));
 sg13g2_inv_1 _0598_ (.Y(_0115_),
    .A(\my_decimation_filter.comb_2[5] ));
 sg13g2_inv_1 _0599_ (.Y(_0116_),
    .A(net176));
 sg13g2_inv_1 _0600_ (.Y(_0117_),
    .A(\my_decimation_filter.input_accumulator[5] ));
 sg13g2_inv_1 _0601_ (.Y(_0118_),
    .A(\my_decimation_filter.input_accumulator[13] ));
 sg13g2_nor2_1 _0602_ (.A(net1),
    .B(net143),
    .Y(_0006_));
 sg13g2_and3_1 _0603_ (.X(_0119_),
    .A(net144),
    .B(net147),
    .C(net152));
 sg13g2_and3_1 _0604_ (.X(_0120_),
    .A(\my_decimation_filter.decimation_count[2] ),
    .B(\my_decimation_filter.decimation_count[1] ),
    .C(\my_decimation_filter.decimation_count[0] ));
 sg13g2_and2_1 _0605_ (.A(net240),
    .B(_0119_),
    .X(_0121_));
 sg13g2_and2_1 _0606_ (.A(net248),
    .B(_0121_),
    .X(_0122_));
 sg13g2_nor2_1 _0607_ (.A(\my_decimation_filter.decimation_count[5] ),
    .B(\my_decimation_filter.decimation_count[4] ),
    .Y(_0123_));
 sg13g2_and3_1 _0608_ (.X(_0124_),
    .A(_0000_),
    .B(_0122_),
    .C(_0123_));
 sg13g2_nand3_1 _0609_ (.B(_0122_),
    .C(_0123_),
    .A(_0000_),
    .Y(_0125_));
 sg13g2_xor2_1 _0610_ (.B(\my_decimation_filter.type_dec_d ),
    .A(net3),
    .X(_0126_));
 sg13g2_nor2_1 _0611_ (.A(net1),
    .B(\my_decimation_filter.reset_d ),
    .Y(_0127_));
 sg13g2_nor2_1 _0612_ (.A(_0126_),
    .B(_0127_),
    .Y(_0128_));
 sg13g2_and2_1 _0613_ (.A(net119),
    .B(net136),
    .X(_0129_));
 sg13g2_nand2_1 _0614_ (.Y(_0130_),
    .A(net119),
    .B(net136));
 sg13g2_nor3_1 _0615_ (.A(net143),
    .B(_0126_),
    .C(_0127_),
    .Y(_0131_));
 sg13g2_nand2b_1 _0616_ (.Y(_0132_),
    .B(net138),
    .A_N(net142));
 sg13g2_nor2_1 _0617_ (.A(net126),
    .B(_0132_),
    .Y(_0133_));
 sg13g2_nand2_1 _0618_ (.Y(_0134_),
    .A(net120),
    .B(net132));
 sg13g2_nand2_1 _0619_ (.Y(_0135_),
    .A(net256),
    .B(net2));
 sg13g2_o21ai_1 _0620_ (.B1(net112),
    .Y(_0136_),
    .A1(net256),
    .A2(net2));
 sg13g2_nor2b_1 _0621_ (.A(_0136_),
    .B_N(_0135_),
    .Y(_0007_));
 sg13g2_nor2_1 _0622_ (.A(net103),
    .B(_0135_),
    .Y(_0137_));
 sg13g2_and2_1 _0623_ (.A(net103),
    .B(_0135_),
    .X(_0138_));
 sg13g2_nor3_1 _0624_ (.A(net110),
    .B(_0137_),
    .C(net104),
    .Y(_0008_));
 sg13g2_and2_1 _0625_ (.A(net233),
    .B(_0137_),
    .X(_0139_));
 sg13g2_nor2_1 _0626_ (.A(net233),
    .B(_0137_),
    .Y(_0140_));
 sg13g2_nor3_1 _0627_ (.A(net110),
    .B(_0139_),
    .C(net234),
    .Y(_0009_));
 sg13g2_and2_1 _0628_ (.A(net222),
    .B(_0139_),
    .X(_0141_));
 sg13g2_nor2_1 _0629_ (.A(net222),
    .B(_0139_),
    .Y(_0142_));
 sg13g2_nor3_1 _0630_ (.A(net109),
    .B(_0141_),
    .C(net223),
    .Y(_0010_));
 sg13g2_nor2b_1 _0631_ (.A(net150),
    .B_N(_0141_),
    .Y(_0143_));
 sg13g2_nor2b_1 _0632_ (.A(_0141_),
    .B_N(net150),
    .Y(_0144_));
 sg13g2_nor3_1 _0633_ (.A(net109),
    .B(_0143_),
    .C(net151),
    .Y(_0011_));
 sg13g2_xnor2_1 _0634_ (.Y(_0145_),
    .A(net173),
    .B(_0143_));
 sg13g2_nor2_1 _0635_ (.A(net109),
    .B(_0145_),
    .Y(_0012_));
 sg13g2_and2_1 _0636_ (.A(\my_decimation_filter.input_accumulator[4] ),
    .B(net173),
    .X(_0146_));
 sg13g2_a21oi_1 _0637_ (.A1(_0141_),
    .A2(_0146_),
    .Y(_0147_),
    .B1(net204));
 sg13g2_and3_1 _0638_ (.X(_0148_),
    .A(net204),
    .B(_0141_),
    .C(_0146_));
 sg13g2_nor3_1 _0639_ (.A(net109),
    .B(net205),
    .C(_0148_),
    .Y(_0013_));
 sg13g2_and2_1 _0640_ (.A(net258),
    .B(_0148_),
    .X(_0149_));
 sg13g2_o21ai_1 _0641_ (.B1(net112),
    .Y(_0150_),
    .A1(net258),
    .A2(_0148_));
 sg13g2_nor2_1 _0642_ (.A(_0149_),
    .B(_0150_),
    .Y(_0014_));
 sg13g2_nor2b_1 _0643_ (.A(_0149_),
    .B_N(net153),
    .Y(_0151_));
 sg13g2_nor2b_1 _0644_ (.A(net153),
    .B_N(_0149_),
    .Y(_0152_));
 sg13g2_nor3_1 _0645_ (.A(net110),
    .B(net154),
    .C(_0152_),
    .Y(_0015_));
 sg13g2_xnor2_1 _0646_ (.Y(_0153_),
    .A(net170),
    .B(_0152_));
 sg13g2_nor2_1 _0647_ (.A(net110),
    .B(_0153_),
    .Y(_0016_));
 sg13g2_and2_1 _0648_ (.A(\my_decimation_filter.input_accumulator[8] ),
    .B(net170),
    .X(_0154_));
 sg13g2_a21oi_1 _0649_ (.A1(_0149_),
    .A2(_0154_),
    .Y(_0155_),
    .B1(net178));
 sg13g2_and3_1 _0650_ (.X(_0156_),
    .A(net178),
    .B(_0149_),
    .C(_0154_));
 sg13g2_nor3_1 _0651_ (.A(_0134_),
    .B(net179),
    .C(_0156_),
    .Y(_0017_));
 sg13g2_nand2_1 _0652_ (.Y(_0157_),
    .A(net259),
    .B(_0156_));
 sg13g2_o21ai_1 _0653_ (.B1(net113),
    .Y(_0158_),
    .A1(net259),
    .A2(_0156_));
 sg13g2_nor2b_1 _0654_ (.A(_0158_),
    .B_N(_0157_),
    .Y(_0018_));
 sg13g2_nor2_1 _0655_ (.A(net106),
    .B(_0157_),
    .Y(_0159_));
 sg13g2_a21oi_1 _0656_ (.A1(net106),
    .A2(_0157_),
    .Y(_0160_),
    .B1(net111));
 sg13g2_nor2b_1 _0657_ (.A(_0159_),
    .B_N(net107),
    .Y(_0019_));
 sg13g2_o21ai_1 _0658_ (.B1(net113),
    .Y(_0161_),
    .A1(net238),
    .A2(_0159_));
 sg13g2_a21oi_1 _0659_ (.A1(net238),
    .A2(_0159_),
    .Y(_0020_),
    .B1(_0161_));
 sg13g2_nand4_1 _0660_ (.B(\my_decimation_filter.input_accumulator[12] ),
    .C(\my_decimation_filter.input_accumulator[13] ),
    .A(\my_decimation_filter.input_accumulator[11] ),
    .Y(_0162_),
    .D(_0156_));
 sg13g2_nor2_1 _0661_ (.A(net101),
    .B(_0162_),
    .Y(_0163_));
 sg13g2_o21ai_1 _0662_ (.B1(net112),
    .Y(_0164_),
    .A1(net101),
    .A2(_0162_));
 sg13g2_a21oi_1 _0663_ (.A1(net101),
    .A2(_0162_),
    .Y(_0021_),
    .B1(_0164_));
 sg13g2_xnor2_1 _0664_ (.Y(_0165_),
    .A(net208),
    .B(_0163_));
 sg13g2_nor2_1 _0665_ (.A(net111),
    .B(net209),
    .Y(_0022_));
 sg13g2_o21ai_1 _0666_ (.B1(net133),
    .Y(_0166_),
    .A1(net144),
    .A2(net152));
 sg13g2_a21oi_1 _0667_ (.A1(net144),
    .A2(net152),
    .Y(_0023_),
    .B1(_0166_));
 sg13g2_a21oi_1 _0668_ (.A1(net144),
    .A2(\my_decimation_filter.decimation_count[0] ),
    .Y(_0167_),
    .B1(net147));
 sg13g2_nor3_1 _0669_ (.A(_0119_),
    .B(_0132_),
    .C(net148),
    .Y(_0024_));
 sg13g2_o21ai_1 _0670_ (.B1(net133),
    .Y(_0168_),
    .A1(net240),
    .A2(_0119_));
 sg13g2_nor2_1 _0671_ (.A(_0121_),
    .B(_0168_),
    .Y(_0025_));
 sg13g2_o21ai_1 _0672_ (.B1(net133),
    .Y(_0169_),
    .A1(net248),
    .A2(_0121_));
 sg13g2_nor2_1 _0673_ (.A(_0122_),
    .B(_0169_),
    .Y(_0026_));
 sg13g2_and2_1 _0674_ (.A(net191),
    .B(_0122_),
    .X(_0170_));
 sg13g2_nor2_1 _0675_ (.A(net191),
    .B(_0122_),
    .Y(_0171_));
 sg13g2_nor3_1 _0676_ (.A(net111),
    .B(_0170_),
    .C(net192),
    .Y(_0027_));
 sg13g2_nand4_1 _0677_ (.B(\my_decimation_filter.decimation_count[4] ),
    .C(\my_decimation_filter.decimation_count[3] ),
    .A(net145),
    .Y(_0172_),
    .D(_0120_));
 sg13g2_o21ai_1 _0678_ (.B1(net133),
    .Y(_0173_),
    .A1(net145),
    .A2(_0170_));
 sg13g2_a21oi_1 _0679_ (.A1(net145),
    .A2(_0170_),
    .Y(_0028_),
    .B1(_0173_));
 sg13g2_xnor2_1 _0680_ (.Y(_0174_),
    .A(_0000_),
    .B(_0172_));
 sg13g2_o21ai_1 _0681_ (.B1(net133),
    .Y(_0175_),
    .A1(net164),
    .A2(net144));
 sg13g2_a21oi_1 _0682_ (.A1(net144),
    .A2(_0174_),
    .Y(_0029_),
    .B1(_0175_));
 sg13g2_o21ai_1 _0683_ (.B1(net132),
    .Y(_0176_),
    .A1(\my_decimation_filter.comb_2[0] ),
    .A2(net125));
 sg13g2_a21oi_1 _0684_ (.A1(_0112_),
    .A2(net125),
    .Y(_0030_),
    .B1(_0176_));
 sg13g2_o21ai_1 _0685_ (.B1(net131),
    .Y(_0177_),
    .A1(net230),
    .A2(net124));
 sg13g2_a21oi_1 _0686_ (.A1(_0111_),
    .A2(net124),
    .Y(_0031_),
    .B1(_0177_));
 sg13g2_o21ai_1 _0687_ (.B1(net130),
    .Y(_0178_),
    .A1(net243),
    .A2(net124));
 sg13g2_a21oi_1 _0688_ (.A1(_0110_),
    .A2(net124),
    .Y(_0032_),
    .B1(_0178_));
 sg13g2_o21ai_1 _0689_ (.B1(net130),
    .Y(_0179_),
    .A1(\my_decimation_filter.comb_1[3] ),
    .A2(net119));
 sg13g2_a21oi_1 _0690_ (.A1(_0116_),
    .A2(net119),
    .Y(_0033_),
    .B1(_0179_));
 sg13g2_o21ai_1 _0691_ (.B1(net129),
    .Y(_0180_),
    .A1(net182),
    .A2(net123));
 sg13g2_a21oi_1 _0692_ (.A1(_0108_),
    .A2(net123),
    .Y(_0034_),
    .B1(_0180_));
 sg13g2_o21ai_1 _0693_ (.B1(net129),
    .Y(_0181_),
    .A1(\my_decimation_filter.comb_2[5] ),
    .A2(net123));
 sg13g2_a21oi_1 _0694_ (.A1(_0106_),
    .A2(net123),
    .Y(_0035_),
    .B1(_0181_));
 sg13g2_o21ai_1 _0695_ (.B1(net129),
    .Y(_0182_),
    .A1(\my_decimation_filter.comb_2[6] ),
    .A2(net123));
 sg13g2_a21oi_1 _0696_ (.A1(_0105_),
    .A2(net123),
    .Y(_0036_),
    .B1(_0182_));
 sg13g2_o21ai_1 _0697_ (.B1(net129),
    .Y(_0183_),
    .A1(\my_decimation_filter.comb_2[7] ),
    .A2(net123));
 sg13g2_a21oi_1 _0698_ (.A1(_0104_),
    .A2(net123),
    .Y(_0037_),
    .B1(_0183_));
 sg13g2_o21ai_1 _0699_ (.B1(net134),
    .Y(_0184_),
    .A1(net237),
    .A2(net128));
 sg13g2_a21oi_1 _0700_ (.A1(_0103_),
    .A2(net128),
    .Y(_0038_),
    .B1(_0184_));
 sg13g2_o21ai_1 _0701_ (.B1(net134),
    .Y(_0185_),
    .A1(net253),
    .A2(net127));
 sg13g2_a21oi_1 _0702_ (.A1(_0102_),
    .A2(net127),
    .Y(_0039_),
    .B1(_0185_));
 sg13g2_o21ai_1 _0703_ (.B1(net133),
    .Y(_0186_),
    .A1(\my_decimation_filter.comb_2[10] ),
    .A2(net127));
 sg13g2_a21oi_1 _0704_ (.A1(_0101_),
    .A2(net127),
    .Y(_0040_),
    .B1(_0186_));
 sg13g2_o21ai_1 _0705_ (.B1(net133),
    .Y(_0187_),
    .A1(net251),
    .A2(net127));
 sg13g2_a21oi_1 _0706_ (.A1(_0100_),
    .A2(net126),
    .Y(_0041_),
    .B1(_0187_));
 sg13g2_o21ai_1 _0707_ (.B1(net135),
    .Y(_0188_),
    .A1(net203),
    .A2(net126));
 sg13g2_a21oi_1 _0708_ (.A1(_0099_),
    .A2(net126),
    .Y(_0042_),
    .B1(_0188_));
 sg13g2_o21ai_1 _0709_ (.B1(net133),
    .Y(_0189_),
    .A1(\my_decimation_filter.comb_2[13] ),
    .A2(net126));
 sg13g2_a21oi_1 _0710_ (.A1(_0097_),
    .A2(net126),
    .Y(_0043_),
    .B1(_0189_));
 sg13g2_o21ai_1 _0711_ (.B1(net132),
    .Y(_0190_),
    .A1(net232),
    .A2(net128));
 sg13g2_a21oi_1 _0712_ (.A1(_0096_),
    .A2(net128),
    .Y(_0044_),
    .B1(_0190_));
 sg13g2_o21ai_1 _0713_ (.B1(net132),
    .Y(_0191_),
    .A1(net163),
    .A2(net128));
 sg13g2_a21oi_1 _0714_ (.A1(_0095_),
    .A2(net128),
    .Y(_0045_),
    .B1(_0191_));
 sg13g2_o21ai_1 _0715_ (.B1(net132),
    .Y(_0192_),
    .A1(net188),
    .A2(net122));
 sg13g2_a21oi_1 _0716_ (.A1(_0112_),
    .A2(net122),
    .Y(_0046_),
    .B1(net189));
 sg13g2_o21ai_1 _0717_ (.B1(net131),
    .Y(_0193_),
    .A1(\my_decimation_filter.Y[1] ),
    .A2(net119));
 sg13g2_a21oi_1 _0718_ (.A1(_0111_),
    .A2(net119),
    .Y(_0047_),
    .B1(_0193_));
 sg13g2_o21ai_1 _0719_ (.B1(net130),
    .Y(_0194_),
    .A1(\my_decimation_filter.Y[2] ),
    .A2(net118));
 sg13g2_a21oi_1 _0720_ (.A1(_0110_),
    .A2(net118),
    .Y(_0048_),
    .B1(_0194_));
 sg13g2_o21ai_1 _0721_ (.B1(net130),
    .Y(_0195_),
    .A1(\my_decimation_filter.comb_1[3] ),
    .A2(net124));
 sg13g2_a21oi_1 _0722_ (.A1(_0109_),
    .A2(net125),
    .Y(_0049_),
    .B1(_0195_));
 sg13g2_o21ai_1 _0723_ (.B1(net129),
    .Y(_0196_),
    .A1(\my_decimation_filter.Y[4] ),
    .A2(net118));
 sg13g2_a21oi_1 _0724_ (.A1(_0108_),
    .A2(net118),
    .Y(_0050_),
    .B1(_0196_));
 sg13g2_o21ai_1 _0725_ (.B1(net129),
    .Y(_0197_),
    .A1(net241),
    .A2(net124));
 sg13g2_a21oi_1 _0726_ (.A1(_0107_),
    .A2(net124),
    .Y(_0051_),
    .B1(_0197_));
 sg13g2_o21ai_1 _0727_ (.B1(net129),
    .Y(_0198_),
    .A1(net231),
    .A2(net118));
 sg13g2_a21oi_1 _0728_ (.A1(_0105_),
    .A2(net118),
    .Y(_0052_),
    .B1(_0198_));
 sg13g2_o21ai_1 _0729_ (.B1(net129),
    .Y(_0199_),
    .A1(net183),
    .A2(net118));
 sg13g2_a21oi_1 _0730_ (.A1(_0104_),
    .A2(net118),
    .Y(_0053_),
    .B1(_0199_));
 sg13g2_o21ai_1 _0731_ (.B1(net134),
    .Y(_0200_),
    .A1(\my_decimation_filter.Y[8] ),
    .A2(net120));
 sg13g2_a21oi_1 _0732_ (.A1(_0103_),
    .A2(net120),
    .Y(_0054_),
    .B1(_0200_));
 sg13g2_o21ai_1 _0733_ (.B1(net134),
    .Y(_0201_),
    .A1(\my_decimation_filter.Y[9] ),
    .A2(net120));
 sg13g2_a21oi_1 _0734_ (.A1(_0102_),
    .A2(net121),
    .Y(_0055_),
    .B1(_0201_));
 sg13g2_o21ai_1 _0735_ (.B1(net134),
    .Y(_0202_),
    .A1(net221),
    .A2(net121));
 sg13g2_a21oi_1 _0736_ (.A1(_0101_),
    .A2(net121),
    .Y(_0056_),
    .B1(_0202_));
 sg13g2_o21ai_1 _0737_ (.B1(net134),
    .Y(_0203_),
    .A1(\my_decimation_filter.Y[11] ),
    .A2(net121));
 sg13g2_a21oi_1 _0738_ (.A1(_0100_),
    .A2(net121),
    .Y(_0057_),
    .B1(_0203_));
 sg13g2_o21ai_1 _0739_ (.B1(net135),
    .Y(_0204_),
    .A1(\my_decimation_filter.Y[12] ),
    .A2(net121));
 sg13g2_a21oi_1 _0740_ (.A1(_0099_),
    .A2(net121),
    .Y(_0058_),
    .B1(_0204_));
 sg13g2_o21ai_1 _0741_ (.B1(net134),
    .Y(_0205_),
    .A1(net244),
    .A2(net126));
 sg13g2_a21oi_1 _0742_ (.A1(_0098_),
    .A2(net126),
    .Y(_0059_),
    .B1(_0205_));
 sg13g2_o21ai_1 _0743_ (.B1(net132),
    .Y(_0206_),
    .A1(\my_decimation_filter.Y[14] ),
    .A2(net120));
 sg13g2_a21oi_1 _0744_ (.A1(_0096_),
    .A2(net120),
    .Y(_0060_),
    .B1(_0206_));
 sg13g2_o21ai_1 _0745_ (.B1(net132),
    .Y(_0207_),
    .A1(\my_decimation_filter.Y[15] ),
    .A2(net120));
 sg13g2_a21oi_1 _0746_ (.A1(_0095_),
    .A2(net120),
    .Y(_0061_),
    .B1(_0207_));
 sg13g2_or2_1 _0747_ (.X(_0208_),
    .B(net256),
    .A(net188));
 sg13g2_nand2_1 _0748_ (.Y(_0209_),
    .A(net188),
    .B(net256));
 sg13g2_and3_1 _0749_ (.X(_0062_),
    .A(net112),
    .B(_0208_),
    .C(_0209_));
 sg13g2_nand2_1 _0750_ (.Y(_0210_),
    .A(net269),
    .B(net261));
 sg13g2_nor2_1 _0751_ (.A(\my_decimation_filter.Y[1] ),
    .B(net261),
    .Y(_0211_));
 sg13g2_xnor2_1 _0752_ (.Y(_0212_),
    .A(\my_decimation_filter.Y[1] ),
    .B(net261));
 sg13g2_xnor2_1 _0753_ (.Y(_0213_),
    .A(_0209_),
    .B(net262));
 sg13g2_nor2_1 _0754_ (.A(net109),
    .B(_0213_),
    .Y(_0063_));
 sg13g2_and2_1 _0755_ (.A(\my_decimation_filter.Y[2] ),
    .B(net272),
    .X(_0214_));
 sg13g2_xor2_1 _0756_ (.B(net233),
    .A(\my_decimation_filter.Y[2] ),
    .X(_0215_));
 sg13g2_o21ai_1 _0757_ (.B1(_0210_),
    .Y(_0216_),
    .A1(_0209_),
    .A2(_0211_));
 sg13g2_xnor2_1 _0758_ (.Y(_0217_),
    .A(_0215_),
    .B(_0216_));
 sg13g2_nor2_1 _0759_ (.A(net109),
    .B(net270),
    .Y(_0064_));
 sg13g2_a21oi_1 _0760_ (.A1(_0215_),
    .A2(_0216_),
    .Y(_0218_),
    .B1(_0214_));
 sg13g2_nand2_1 _0761_ (.Y(_0219_),
    .A(\my_decimation_filter.Y[3] ),
    .B(net279));
 sg13g2_xnor2_1 _0762_ (.Y(_0220_),
    .A(\my_decimation_filter.Y[3] ),
    .B(net222));
 sg13g2_xnor2_1 _0763_ (.Y(_0221_),
    .A(_0218_),
    .B(_0220_));
 sg13g2_nor2_1 _0764_ (.A(net110),
    .B(net273),
    .Y(_0065_));
 sg13g2_xor2_1 _0765_ (.B(net278),
    .A(\my_decimation_filter.Y[4] ),
    .X(_0222_));
 sg13g2_o21ai_1 _0766_ (.B1(_0219_),
    .Y(_0223_),
    .A1(_0218_),
    .A2(_0220_));
 sg13g2_nor2_1 _0767_ (.A(_0222_),
    .B(_0223_),
    .Y(_0224_));
 sg13g2_and2_1 _0768_ (.A(_0222_),
    .B(_0223_),
    .X(_0225_));
 sg13g2_nor3_1 _0769_ (.A(net109),
    .B(_0224_),
    .C(_0225_),
    .Y(_0066_));
 sg13g2_xor2_1 _0770_ (.B(\my_decimation_filter.input_accumulator[5] ),
    .A(\my_decimation_filter.Y[5] ),
    .X(_0226_));
 sg13g2_a21o_1 _0771_ (.A2(net278),
    .A1(\my_decimation_filter.Y[4] ),
    .B1(_0226_),
    .X(_0227_));
 sg13g2_and2_1 _0772_ (.A(_0225_),
    .B(_0226_),
    .X(_0228_));
 sg13g2_nand3_1 _0773_ (.B(_0223_),
    .C(_0226_),
    .A(_0222_),
    .Y(_0229_));
 sg13g2_nand3_1 _0774_ (.B(net278),
    .C(_0226_),
    .A(\my_decimation_filter.Y[4] ),
    .Y(_0230_));
 sg13g2_o21ai_1 _0775_ (.B1(_0230_),
    .Y(_0231_),
    .A1(_0225_),
    .A2(_0227_));
 sg13g2_nor3_1 _0776_ (.A(net109),
    .B(_0228_),
    .C(_0231_),
    .Y(_0067_));
 sg13g2_nand2_1 _0777_ (.Y(_0232_),
    .A(\my_decimation_filter.Y[6] ),
    .B(net204));
 sg13g2_nor2_1 _0778_ (.A(\my_decimation_filter.Y[6] ),
    .B(net266),
    .Y(_0233_));
 sg13g2_xnor2_1 _0779_ (.Y(_0234_),
    .A(net231),
    .B(net204));
 sg13g2_o21ai_1 _0780_ (.B1(_0230_),
    .Y(_0235_),
    .A1(_0107_),
    .A2(_0117_));
 sg13g2_nor2_1 _0781_ (.A(_0228_),
    .B(_0235_),
    .Y(_0236_));
 sg13g2_o21ai_1 _0782_ (.B1(net112),
    .Y(_0237_),
    .A1(_0234_),
    .A2(_0236_));
 sg13g2_a21oi_1 _0783_ (.A1(_0234_),
    .A2(_0236_),
    .Y(_0068_),
    .B1(_0237_));
 sg13g2_nor2_1 _0784_ (.A(net183),
    .B(net258),
    .Y(_0238_));
 sg13g2_nand2_1 _0785_ (.Y(_0239_),
    .A(\my_decimation_filter.Y[7] ),
    .B(net258));
 sg13g2_nor2b_1 _0786_ (.A(_0238_),
    .B_N(_0239_),
    .Y(_0240_));
 sg13g2_o21ai_1 _0787_ (.B1(_0232_),
    .Y(_0241_),
    .A1(_0233_),
    .A2(_0236_));
 sg13g2_o21ai_1 _0788_ (.B1(net112),
    .Y(_0242_),
    .A1(_0240_),
    .A2(_0241_));
 sg13g2_a21oi_1 _0789_ (.A1(_0240_),
    .A2(net267),
    .Y(_0069_),
    .B1(_0242_));
 sg13g2_o21ai_1 _0790_ (.B1(_0239_),
    .Y(_0243_),
    .A1(_0232_),
    .A2(_0238_));
 sg13g2_nor2_1 _0791_ (.A(_0235_),
    .B(_0243_),
    .Y(_0244_));
 sg13g2_a221oi_1 _0792_ (.B2(_0229_),
    .C1(_0238_),
    .B1(_0244_),
    .A1(_0233_),
    .Y(_0245_),
    .A2(_0239_));
 sg13g2_and2_1 _0793_ (.A(\my_decimation_filter.Y[8] ),
    .B(\my_decimation_filter.input_accumulator[8] ),
    .X(_0246_));
 sg13g2_xor2_1 _0794_ (.B(net271),
    .A(\my_decimation_filter.Y[8] ),
    .X(_0247_));
 sg13g2_o21ai_1 _0795_ (.B1(net112),
    .Y(_0248_),
    .A1(_0245_),
    .A2(_0247_));
 sg13g2_a21oi_1 _0796_ (.A1(_0245_),
    .A2(_0247_),
    .Y(_0070_),
    .B1(_0248_));
 sg13g2_a21o_1 _0797_ (.A2(_0247_),
    .A1(_0245_),
    .B1(_0246_),
    .X(_0249_));
 sg13g2_and2_1 _0798_ (.A(net260),
    .B(net170),
    .X(_0250_));
 sg13g2_xor2_1 _0799_ (.B(net280),
    .A(\my_decimation_filter.Y[9] ),
    .X(_0251_));
 sg13g2_a21oi_1 _0800_ (.A1(_0249_),
    .A2(_0251_),
    .Y(_0252_),
    .B1(net111));
 sg13g2_o21ai_1 _0801_ (.B1(_0252_),
    .Y(_0253_),
    .A1(_0249_),
    .A2(_0251_));
 sg13g2_inv_1 _0802_ (.Y(_0071_),
    .A(_0253_));
 sg13g2_nand2_1 _0803_ (.Y(_0254_),
    .A(net221),
    .B(net178));
 sg13g2_xnor2_1 _0804_ (.Y(_0255_),
    .A(net221),
    .B(net178));
 sg13g2_a21oi_1 _0805_ (.A1(_0249_),
    .A2(_0251_),
    .Y(_0256_),
    .B1(_0250_));
 sg13g2_or2_1 _0806_ (.X(_0257_),
    .B(_0256_),
    .A(_0255_));
 sg13g2_nand2_1 _0807_ (.Y(_0258_),
    .A(net113),
    .B(_0257_));
 sg13g2_a21oi_1 _0808_ (.A1(_0255_),
    .A2(_0256_),
    .Y(_0072_),
    .B1(_0258_));
 sg13g2_nand2_1 _0809_ (.Y(_0259_),
    .A(\my_decimation_filter.Y[11] ),
    .B(\my_decimation_filter.input_accumulator[11] ));
 sg13g2_nor2_1 _0810_ (.A(\my_decimation_filter.Y[11] ),
    .B(\my_decimation_filter.input_accumulator[11] ),
    .Y(_0260_));
 sg13g2_xnor2_1 _0811_ (.Y(_0261_),
    .A(\my_decimation_filter.Y[11] ),
    .B(net259));
 sg13g2_a21oi_1 _0812_ (.A1(_0254_),
    .A2(_0257_),
    .Y(_0262_),
    .B1(_0261_));
 sg13g2_and3_1 _0813_ (.X(_0263_),
    .A(_0254_),
    .B(_0257_),
    .C(_0261_));
 sg13g2_nor3_1 _0814_ (.A(net111),
    .B(_0262_),
    .C(_0263_),
    .Y(_0073_));
 sg13g2_nor2_1 _0815_ (.A(_0255_),
    .B(_0261_),
    .Y(_0264_));
 sg13g2_and3_1 _0816_ (.X(_0265_),
    .A(_0247_),
    .B(_0251_),
    .C(_0264_));
 sg13g2_a21o_1 _0817_ (.A2(_0251_),
    .A1(_0246_),
    .B1(_0250_),
    .X(_0266_));
 sg13g2_o21ai_1 _0818_ (.B1(_0259_),
    .Y(_0267_),
    .A1(_0254_),
    .A2(_0260_));
 sg13g2_a221oi_1 _0819_ (.B2(_0264_),
    .C1(_0267_),
    .B1(_0266_),
    .A1(_0245_),
    .Y(_0268_),
    .A2(_0265_));
 sg13g2_nand2_1 _0820_ (.Y(_0269_),
    .A(\my_decimation_filter.Y[12] ),
    .B(net275));
 sg13g2_xnor2_1 _0821_ (.Y(_0270_),
    .A(\my_decimation_filter.Y[12] ),
    .B(net275));
 sg13g2_xnor2_1 _0822_ (.Y(_0271_),
    .A(_0268_),
    .B(_0270_));
 sg13g2_nor2_1 _0823_ (.A(net111),
    .B(_0271_),
    .Y(_0074_));
 sg13g2_xnor2_1 _0824_ (.Y(_0272_),
    .A(\my_decimation_filter.Y[13] ),
    .B(\my_decimation_filter.input_accumulator[13] ));
 sg13g2_o21ai_1 _0825_ (.B1(net276),
    .Y(_0273_),
    .A1(_0268_),
    .A2(_0270_));
 sg13g2_xor2_1 _0826_ (.B(_0273_),
    .A(_0272_),
    .X(_0274_));
 sg13g2_nor2_1 _0827_ (.A(net111),
    .B(net277),
    .Y(_0075_));
 sg13g2_nor2_1 _0828_ (.A(_0270_),
    .B(_0272_),
    .Y(_0275_));
 sg13g2_inv_1 _0829_ (.Y(_0276_),
    .A(_0275_));
 sg13g2_a21oi_1 _0830_ (.A1(_0098_),
    .A2(_0118_),
    .Y(_0277_),
    .B1(_0269_));
 sg13g2_a21oi_1 _0831_ (.A1(net257),
    .A2(\my_decimation_filter.input_accumulator[13] ),
    .Y(_0278_),
    .B1(_0277_));
 sg13g2_o21ai_1 _0832_ (.B1(_0278_),
    .Y(_0279_),
    .A1(_0268_),
    .A2(_0276_));
 sg13g2_and2_1 _0833_ (.A(\my_decimation_filter.Y[14] ),
    .B(\my_decimation_filter.input_accumulator[14] ),
    .X(_0280_));
 sg13g2_xor2_1 _0834_ (.B(net263),
    .A(\my_decimation_filter.Y[14] ),
    .X(_0281_));
 sg13g2_o21ai_1 _0835_ (.B1(net113),
    .Y(_0282_),
    .A1(_0279_),
    .A2(_0281_));
 sg13g2_a21oi_1 _0836_ (.A1(_0279_),
    .A2(net264),
    .Y(_0076_),
    .B1(_0282_));
 sg13g2_a21o_1 _0837_ (.A2(_0281_),
    .A1(_0279_),
    .B1(_0280_),
    .X(_0283_));
 sg13g2_xor2_1 _0838_ (.B(net208),
    .A(net274),
    .X(_0284_));
 sg13g2_nand2_1 _0839_ (.Y(_0285_),
    .A(_0283_),
    .B(_0284_));
 sg13g2_or2_1 _0840_ (.X(_0286_),
    .B(_0284_),
    .A(_0283_));
 sg13g2_and3_1 _0841_ (.X(_0077_),
    .A(net112),
    .B(_0285_),
    .C(_0286_));
 sg13g2_nor2_1 _0842_ (.A(net217),
    .B(net114),
    .Y(_0287_));
 sg13g2_nor2b_1 _0843_ (.A(\my_decimation_filter.comb_1[0] ),
    .B_N(\my_decimation_filter.comb_2[0] ),
    .Y(_0288_));
 sg13g2_xor2_1 _0844_ (.B(\my_decimation_filter.comb_2[0] ),
    .A(net159),
    .X(_0289_));
 sg13g2_nor4_2 _0845_ (.A(net144),
    .B(net1),
    .C(\my_decimation_filter.reset_d ),
    .Y(_0290_),
    .D(\my_decimation_filter.type_dec_d ));
 sg13g2_a221oi_1 _0846_ (.B2(net188),
    .C1(net117),
    .B1(net139),
    .A1(net137),
    .Y(_0291_),
    .A2(_0289_));
 sg13g2_nor3_1 _0847_ (.A(net142),
    .B(_0287_),
    .C(_0291_),
    .Y(_0078_));
 sg13g2_nand2b_1 _0848_ (.Y(_0292_),
    .B(\my_decimation_filter.comb_1[1] ),
    .A_N(\my_decimation_filter.comb_2[1] ));
 sg13g2_xor2_1 _0849_ (.B(\my_decimation_filter.comb_2[1] ),
    .A(\my_decimation_filter.comb_1[1] ),
    .X(_0293_));
 sg13g2_nor2_1 _0850_ (.A(_0288_),
    .B(_0293_),
    .Y(_0294_));
 sg13g2_nand2_1 _0851_ (.Y(_0295_),
    .A(_0288_),
    .B(_0293_));
 sg13g2_nor2b_1 _0852_ (.A(_0294_),
    .B_N(net137),
    .Y(_0296_));
 sg13g2_a221oi_1 _0853_ (.B2(_0296_),
    .C1(net117),
    .B1(_0295_),
    .A1(\my_decimation_filter.Y[1] ),
    .Y(_0297_),
    .A2(net139));
 sg13g2_nor2_1 _0854_ (.A(net193),
    .B(net114),
    .Y(_0298_));
 sg13g2_nor3_1 _0855_ (.A(net141),
    .B(_0297_),
    .C(_0298_),
    .Y(_0079_));
 sg13g2_nor2_1 _0856_ (.A(_0110_),
    .B(\my_decimation_filter.comb_2[2] ),
    .Y(_0299_));
 sg13g2_xnor2_1 _0857_ (.Y(_0300_),
    .A(\my_decimation_filter.comb_1[2] ),
    .B(\my_decimation_filter.comb_2[2] ));
 sg13g2_o21ai_1 _0858_ (.B1(_0292_),
    .Y(_0301_),
    .A1(_0288_),
    .A2(_0293_));
 sg13g2_xor2_1 _0859_ (.B(_0301_),
    .A(_0300_),
    .X(_0302_));
 sg13g2_a221oi_1 _0860_ (.B2(net136),
    .C1(net117),
    .B1(_0302_),
    .A1(\my_decimation_filter.Y[2] ),
    .Y(_0303_),
    .A2(net139));
 sg13g2_nor2_1 _0861_ (.A(net195),
    .B(net114),
    .Y(_0304_));
 sg13g2_nor3_1 _0862_ (.A(net141),
    .B(_0303_),
    .C(_0304_),
    .Y(_0080_));
 sg13g2_a21oi_1 _0863_ (.A1(_0300_),
    .A2(_0301_),
    .Y(_0305_),
    .B1(_0299_));
 sg13g2_nor2_1 _0864_ (.A(\my_decimation_filter.comb_1[3] ),
    .B(_0116_),
    .Y(_0306_));
 sg13g2_xnor2_1 _0865_ (.Y(_0307_),
    .A(\my_decimation_filter.comb_1[3] ),
    .B(\my_decimation_filter.comb_2[3] ));
 sg13g2_xnor2_1 _0866_ (.Y(_0308_),
    .A(_0305_),
    .B(_0307_));
 sg13g2_a221oi_1 _0867_ (.B2(net136),
    .C1(net117),
    .B1(_0308_),
    .A1(\my_decimation_filter.Y[3] ),
    .Y(_0309_),
    .A2(net139));
 sg13g2_nor2_1 _0868_ (.A(net201),
    .B(net114),
    .Y(_0310_));
 sg13g2_nor3_1 _0869_ (.A(net141),
    .B(_0309_),
    .C(_0310_),
    .Y(_0081_));
 sg13g2_nor2b_1 _0870_ (.A(\my_decimation_filter.comb_2[4] ),
    .B_N(\my_decimation_filter.comb_1[4] ),
    .Y(_0311_));
 sg13g2_xor2_1 _0871_ (.B(\my_decimation_filter.comb_2[4] ),
    .A(\my_decimation_filter.comb_1[4] ),
    .X(_0312_));
 sg13g2_a221oi_1 _0872_ (.B2(_0301_),
    .C1(_0299_),
    .B1(_0300_),
    .A1(\my_decimation_filter.comb_1[3] ),
    .Y(_0313_),
    .A2(_0116_));
 sg13g2_o21ai_1 _0873_ (.B1(_0312_),
    .Y(_0314_),
    .A1(_0306_),
    .A2(_0313_));
 sg13g2_nor3_1 _0874_ (.A(_0306_),
    .B(_0312_),
    .C(_0313_),
    .Y(_0315_));
 sg13g2_nor2b_1 _0875_ (.A(_0315_),
    .B_N(net136),
    .Y(_0316_));
 sg13g2_a221oi_1 _0876_ (.B2(_0316_),
    .C1(net117),
    .B1(_0314_),
    .A1(\my_decimation_filter.Y[4] ),
    .Y(_0317_),
    .A2(net139));
 sg13g2_nor2_1 _0877_ (.A(net180),
    .B(net114),
    .Y(_0318_));
 sg13g2_nor3_1 _0878_ (.A(net141),
    .B(_0317_),
    .C(_0318_),
    .Y(_0082_));
 sg13g2_xnor2_1 _0879_ (.Y(_0319_),
    .A(\my_decimation_filter.comb_1[5] ),
    .B(\my_decimation_filter.comb_2[5] ));
 sg13g2_inv_1 _0880_ (.Y(_0320_),
    .A(_0319_));
 sg13g2_nor2_1 _0881_ (.A(_0311_),
    .B(_0315_),
    .Y(_0321_));
 sg13g2_xnor2_1 _0882_ (.Y(_0322_),
    .A(_0319_),
    .B(_0321_));
 sg13g2_a221oi_1 _0883_ (.B2(net136),
    .C1(net117),
    .B1(_0322_),
    .A1(\my_decimation_filter.Y[5] ),
    .Y(_0323_),
    .A2(net139));
 sg13g2_nor2_1 _0884_ (.A(net206),
    .B(net114),
    .Y(_0324_));
 sg13g2_nor3_1 _0885_ (.A(net141),
    .B(_0323_),
    .C(_0324_),
    .Y(_0083_));
 sg13g2_nand2b_1 _0886_ (.Y(_0325_),
    .B(\my_decimation_filter.comb_1[6] ),
    .A_N(\my_decimation_filter.comb_2[6] ));
 sg13g2_nor2b_1 _0887_ (.A(\my_decimation_filter.comb_1[6] ),
    .B_N(\my_decimation_filter.comb_2[6] ),
    .Y(_0326_));
 sg13g2_xnor2_1 _0888_ (.Y(_0327_),
    .A(\my_decimation_filter.comb_1[6] ),
    .B(\my_decimation_filter.comb_2[6] ));
 sg13g2_nor4_2 _0889_ (.A(_0306_),
    .B(_0312_),
    .C(_0313_),
    .Y(_0328_),
    .D(_0320_));
 sg13g2_a21oi_1 _0890_ (.A1(\my_decimation_filter.comb_1[5] ),
    .A2(_0115_),
    .Y(_0329_),
    .B1(_0311_));
 sg13g2_a21oi_1 _0891_ (.A1(_0106_),
    .A2(\my_decimation_filter.comb_2[5] ),
    .Y(_0330_),
    .B1(_0329_));
 sg13g2_nor2_1 _0892_ (.A(_0328_),
    .B(_0330_),
    .Y(_0331_));
 sg13g2_xnor2_1 _0893_ (.Y(_0332_),
    .A(_0327_),
    .B(_0331_));
 sg13g2_a221oi_1 _0894_ (.B2(net136),
    .C1(net117),
    .B1(_0332_),
    .A1(\my_decimation_filter.Y[6] ),
    .Y(_0333_),
    .A2(net139));
 sg13g2_nor2_1 _0895_ (.A(net197),
    .B(net114),
    .Y(_0334_));
 sg13g2_nor3_1 _0896_ (.A(net141),
    .B(_0333_),
    .C(_0334_),
    .Y(_0084_));
 sg13g2_nor2b_1 _0897_ (.A(\my_decimation_filter.comb_1[7] ),
    .B_N(\my_decimation_filter.comb_2[7] ),
    .Y(_0335_));
 sg13g2_nand2b_1 _0898_ (.Y(_0336_),
    .B(\my_decimation_filter.comb_1[7] ),
    .A_N(\my_decimation_filter.comb_2[7] ));
 sg13g2_nand2b_1 _0899_ (.Y(_0337_),
    .B(_0336_),
    .A_N(_0335_));
 sg13g2_o21ai_1 _0900_ (.B1(_0325_),
    .Y(_0338_),
    .A1(_0326_),
    .A2(_0331_));
 sg13g2_xnor2_1 _0901_ (.Y(_0339_),
    .A(_0337_),
    .B(_0338_));
 sg13g2_a221oi_1 _0902_ (.B2(net136),
    .C1(net117),
    .B1(_0339_),
    .A1(net183),
    .Y(_0340_),
    .A2(net139));
 sg13g2_nor2_1 _0903_ (.A(net212),
    .B(net114),
    .Y(_0341_));
 sg13g2_nor3_1 _0904_ (.A(net141),
    .B(_0340_),
    .C(_0341_),
    .Y(_0085_));
 sg13g2_nor2_1 _0905_ (.A(_0103_),
    .B(\my_decimation_filter.comb_2[8] ),
    .Y(_0342_));
 sg13g2_xnor2_1 _0906_ (.Y(_0343_),
    .A(\my_decimation_filter.comb_1[8] ),
    .B(\my_decimation_filter.comb_2[8] ));
 sg13g2_o21ai_1 _0907_ (.B1(_0336_),
    .Y(_0344_),
    .A1(_0325_),
    .A2(_0335_));
 sg13g2_or2_1 _0908_ (.X(_0345_),
    .B(_0344_),
    .A(_0330_));
 sg13g2_a21oi_1 _0909_ (.A1(_0326_),
    .A2(_0336_),
    .Y(_0346_),
    .B1(_0335_));
 sg13g2_o21ai_1 _0910_ (.B1(_0346_),
    .Y(_0347_),
    .A1(_0328_),
    .A2(_0345_));
 sg13g2_inv_1 _0911_ (.Y(_0348_),
    .A(_0347_));
 sg13g2_xnor2_1 _0912_ (.Y(_0349_),
    .A(_0343_),
    .B(_0347_));
 sg13g2_a221oi_1 _0913_ (.B2(net138),
    .C1(net116),
    .B1(_0349_),
    .A1(\my_decimation_filter.Y[8] ),
    .Y(_0350_),
    .A2(net140));
 sg13g2_nor2_1 _0914_ (.A(net155),
    .B(net115),
    .Y(_0351_));
 sg13g2_nor3_1 _0915_ (.A(net142),
    .B(_0350_),
    .C(_0351_),
    .Y(_0086_));
 sg13g2_nand2_1 _0916_ (.Y(_0352_),
    .A(_0102_),
    .B(\my_decimation_filter.comb_2[9] ));
 sg13g2_nor2_1 _0917_ (.A(_0102_),
    .B(\my_decimation_filter.comb_2[9] ),
    .Y(_0353_));
 sg13g2_xnor2_1 _0918_ (.Y(_0354_),
    .A(\my_decimation_filter.comb_1[9] ),
    .B(\my_decimation_filter.comb_2[9] ));
 sg13g2_a21oi_1 _0919_ (.A1(_0343_),
    .A2(_0348_),
    .Y(_0355_),
    .B1(_0342_));
 sg13g2_xnor2_1 _0920_ (.Y(_0356_),
    .A(_0354_),
    .B(_0355_));
 sg13g2_a221oi_1 _0921_ (.B2(net138),
    .C1(net116),
    .B1(_0356_),
    .A1(\my_decimation_filter.Y[9] ),
    .Y(_0357_),
    .A2(net140));
 sg13g2_nor2_1 _0922_ (.A(net166),
    .B(net115),
    .Y(_0358_));
 sg13g2_nor3_1 _0923_ (.A(net142),
    .B(_0357_),
    .C(_0358_),
    .Y(_0087_));
 sg13g2_nor2_1 _0924_ (.A(_0101_),
    .B(\my_decimation_filter.comb_2[10] ),
    .Y(_0359_));
 sg13g2_xor2_1 _0925_ (.B(\my_decimation_filter.comb_2[10] ),
    .A(\my_decimation_filter.comb_1[10] ),
    .X(_0360_));
 sg13g2_a21oi_1 _0926_ (.A1(_0342_),
    .A2(_0352_),
    .Y(_0361_),
    .B1(_0353_));
 sg13g2_inv_1 _0927_ (.Y(_0362_),
    .A(_0361_));
 sg13g2_nand2_1 _0928_ (.Y(_0363_),
    .A(_0343_),
    .B(_0354_));
 sg13g2_or2_1 _0929_ (.X(_0364_),
    .B(_0363_),
    .A(_0347_));
 sg13g2_a21oi_1 _0930_ (.A1(_0361_),
    .A2(_0364_),
    .Y(_0365_),
    .B1(_0360_));
 sg13g2_nand3_1 _0931_ (.B(_0361_),
    .C(_0364_),
    .A(_0360_),
    .Y(_0366_));
 sg13g2_nand3b_1 _0932_ (.B(_0366_),
    .C(net138),
    .Y(_0367_),
    .A_N(_0365_));
 sg13g2_a21oi_1 _0933_ (.A1(\my_decimation_filter.Y[10] ),
    .A2(net140),
    .Y(_0368_),
    .B1(_0129_));
 sg13g2_a221oi_1 _0934_ (.B2(_0368_),
    .C1(net142),
    .B1(_0367_),
    .A1(_0094_),
    .Y(_0088_),
    .A2(net116));
 sg13g2_xnor2_1 _0935_ (.Y(_0369_),
    .A(\my_decimation_filter.comb_1[11] ),
    .B(\my_decimation_filter.comb_2[11] ));
 sg13g2_nor2_1 _0936_ (.A(_0359_),
    .B(_0365_),
    .Y(_0370_));
 sg13g2_xnor2_1 _0937_ (.Y(_0371_),
    .A(_0369_),
    .B(_0370_));
 sg13g2_a221oi_1 _0938_ (.B2(net138),
    .C1(net116),
    .B1(_0371_),
    .A1(\my_decimation_filter.Y[11] ),
    .Y(_0372_),
    .A2(net140));
 sg13g2_nor2_1 _0939_ (.A(net168),
    .B(net115),
    .Y(_0373_));
 sg13g2_nor3_1 _0940_ (.A(net143),
    .B(_0372_),
    .C(_0373_),
    .Y(_0089_));
 sg13g2_nor2b_1 _0941_ (.A(_0360_),
    .B_N(_0369_),
    .Y(_0374_));
 sg13g2_nand2b_1 _0942_ (.Y(_0375_),
    .B(_0374_),
    .A_N(_0363_));
 sg13g2_o21ai_1 _0943_ (.B1(_0359_),
    .Y(_0376_),
    .A1(\my_decimation_filter.comb_1[11] ),
    .A2(_0114_));
 sg13g2_o21ai_1 _0944_ (.B1(_0376_),
    .Y(_0377_),
    .A1(_0100_),
    .A2(\my_decimation_filter.comb_2[11] ));
 sg13g2_a21oi_1 _0945_ (.A1(_0362_),
    .A2(_0374_),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_o21ai_1 _0946_ (.B1(_0378_),
    .Y(_0379_),
    .A1(_0347_),
    .A2(_0375_));
 sg13g2_nor2_1 _0947_ (.A(_0099_),
    .B(\my_decimation_filter.comb_2[12] ),
    .Y(_0380_));
 sg13g2_xnor2_1 _0948_ (.Y(_0381_),
    .A(\my_decimation_filter.comb_1[12] ),
    .B(\my_decimation_filter.comb_2[12] ));
 sg13g2_xor2_1 _0949_ (.B(_0381_),
    .A(_0379_),
    .X(_0382_));
 sg13g2_a221oi_1 _0950_ (.B2(net138),
    .C1(net116),
    .B1(_0382_),
    .A1(\my_decimation_filter.Y[12] ),
    .Y(_0383_),
    .A2(net140));
 sg13g2_nor2_1 _0951_ (.A(net235),
    .B(net115),
    .Y(_0384_));
 sg13g2_nor3_1 _0952_ (.A(net143),
    .B(_0383_),
    .C(_0384_),
    .Y(_0090_));
 sg13g2_xnor2_1 _0953_ (.Y(_0385_),
    .A(\my_decimation_filter.comb_1[13] ),
    .B(\my_decimation_filter.comb_2[13] ));
 sg13g2_a21oi_1 _0954_ (.A1(_0379_),
    .A2(_0381_),
    .Y(_0386_),
    .B1(_0380_));
 sg13g2_xnor2_1 _0955_ (.Y(_0387_),
    .A(_0385_),
    .B(_0386_));
 sg13g2_a221oi_1 _0956_ (.B2(net138),
    .C1(net116),
    .B1(_0387_),
    .A1(\my_decimation_filter.Y[13] ),
    .Y(_0388_),
    .A2(net140));
 sg13g2_nor2_1 _0957_ (.A(net224),
    .B(net115),
    .Y(_0389_));
 sg13g2_nor3_1 _0958_ (.A(net142),
    .B(_0388_),
    .C(_0389_),
    .Y(_0091_));
 sg13g2_nand2b_1 _0959_ (.Y(_0390_),
    .B(\my_decimation_filter.comb_1[14] ),
    .A_N(\my_decimation_filter.comb_2[14] ));
 sg13g2_nor2b_1 _0960_ (.A(\my_decimation_filter.comb_1[14] ),
    .B_N(\my_decimation_filter.comb_2[14] ),
    .Y(_0391_));
 sg13g2_xnor2_1 _0961_ (.Y(_0392_),
    .A(\my_decimation_filter.comb_1[14] ),
    .B(\my_decimation_filter.comb_2[14] ));
 sg13g2_and2_1 _0962_ (.A(_0381_),
    .B(_0385_),
    .X(_0393_));
 sg13g2_o21ai_1 _0963_ (.B1(_0380_),
    .Y(_0394_),
    .A1(\my_decimation_filter.comb_1[13] ),
    .A2(_0113_));
 sg13g2_o21ai_1 _0964_ (.B1(_0394_),
    .Y(_0395_),
    .A1(_0097_),
    .A2(\my_decimation_filter.comb_2[13] ));
 sg13g2_a21oi_2 _0965_ (.B1(_0395_),
    .Y(_0396_),
    .A2(_0393_),
    .A1(_0379_));
 sg13g2_xnor2_1 _0966_ (.Y(_0397_),
    .A(_0392_),
    .B(_0396_));
 sg13g2_a221oi_1 _0967_ (.B2(net137),
    .C1(net116),
    .B1(_0397_),
    .A1(\my_decimation_filter.Y[14] ),
    .Y(_0398_),
    .A2(net140));
 sg13g2_nor2_1 _0968_ (.A(net161),
    .B(net115),
    .Y(_0399_));
 sg13g2_nor3_1 _0969_ (.A(net142),
    .B(_0398_),
    .C(_0399_),
    .Y(_0092_));
 sg13g2_o21ai_1 _0970_ (.B1(_0390_),
    .Y(_0400_),
    .A1(_0391_),
    .A2(_0396_));
 sg13g2_xor2_1 _0971_ (.B(\my_decimation_filter.comb_2[15] ),
    .A(\my_decimation_filter.comb_1[15] ),
    .X(_0401_));
 sg13g2_xnor2_1 _0972_ (.Y(_0402_),
    .A(_0400_),
    .B(_0401_));
 sg13g2_a221oi_1 _0973_ (.B2(net137),
    .C1(net116),
    .B1(_0402_),
    .A1(\my_decimation_filter.Y[15] ),
    .Y(_0403_),
    .A2(net140));
 sg13g2_nor2_1 _0974_ (.A(net186),
    .B(net115),
    .Y(_0404_));
 sg13g2_nor3_1 _0975_ (.A(net141),
    .B(_0403_),
    .C(_0404_),
    .Y(_0093_));
 sg13g2_dfrbp_1 _0976_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net64),
    .D(_0006_),
    .Q_N(_0487_),
    .Q(\my_decimation_filter.reset_d ));
 sg13g2_dfrbp_1 _0977_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net5),
    .D(net144),
    .Q_N(_0486_),
    .Q(\my_decimation_filter.type_dec_d ));
 sg13g2_dfrbp_1 _0978_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net39),
    .D(_0007_),
    .Q_N(_0485_),
    .Q(\my_decimation_filter.input_accumulator[0] ));
 sg13g2_dfrbp_1 _0979_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net38),
    .D(net105),
    .Q_N(_0001_),
    .Q(\my_decimation_filter.input_accumulator[1] ));
 sg13g2_dfrbp_1 _0980_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net37),
    .D(_0009_),
    .Q_N(_0484_),
    .Q(\my_decimation_filter.input_accumulator[2] ));
 sg13g2_dfrbp_1 _0981_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net36),
    .D(_0010_),
    .Q_N(_0483_),
    .Q(\my_decimation_filter.input_accumulator[3] ));
 sg13g2_dfrbp_1 _0982_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net35),
    .D(_0011_),
    .Q_N(_0002_),
    .Q(\my_decimation_filter.input_accumulator[4] ));
 sg13g2_dfrbp_1 _0983_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net34),
    .D(_0012_),
    .Q_N(_0482_),
    .Q(\my_decimation_filter.input_accumulator[5] ));
 sg13g2_dfrbp_1 _0984_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net33),
    .D(_0013_),
    .Q_N(_0481_),
    .Q(\my_decimation_filter.input_accumulator[6] ));
 sg13g2_dfrbp_1 _0985_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net32),
    .D(_0014_),
    .Q_N(_0480_),
    .Q(\my_decimation_filter.input_accumulator[7] ));
 sg13g2_dfrbp_1 _0986_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net31),
    .D(_0015_),
    .Q_N(_0003_),
    .Q(\my_decimation_filter.input_accumulator[8] ));
 sg13g2_dfrbp_1 _0987_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net30),
    .D(_0016_),
    .Q_N(_0479_),
    .Q(\my_decimation_filter.input_accumulator[9] ));
 sg13g2_dfrbp_1 _0988_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net29),
    .D(_0017_),
    .Q_N(_0478_),
    .Q(\my_decimation_filter.input_accumulator[10] ));
 sg13g2_dfrbp_1 _0989_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net28),
    .D(_0018_),
    .Q_N(_0477_),
    .Q(\my_decimation_filter.input_accumulator[11] ));
 sg13g2_dfrbp_1 _0990_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net27),
    .D(net108),
    .Q_N(_0004_),
    .Q(\my_decimation_filter.input_accumulator[12] ));
 sg13g2_dfrbp_1 _0991_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net26),
    .D(net239),
    .Q_N(_0476_),
    .Q(\my_decimation_filter.input_accumulator[13] ));
 sg13g2_dfrbp_1 _0992_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net25),
    .D(net102),
    .Q_N(_0005_),
    .Q(\my_decimation_filter.input_accumulator[14] ));
 sg13g2_dfrbp_1 _0993_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net24),
    .D(_0022_),
    .Q_N(_0475_),
    .Q(\my_decimation_filter.input_accumulator[15] ));
 sg13g2_dfrbp_1 _0994_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net23),
    .D(_0023_),
    .Q_N(_0474_),
    .Q(\my_decimation_filter.decimation_count[0] ));
 sg13g2_dfrbp_1 _0995_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net21),
    .D(net149),
    .Q_N(_0473_),
    .Q(\my_decimation_filter.decimation_count[1] ));
 sg13g2_dfrbp_1 _0996_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net19),
    .D(_0025_),
    .Q_N(_0472_),
    .Q(\my_decimation_filter.decimation_count[2] ));
 sg13g2_dfrbp_1 _0997_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net17),
    .D(_0026_),
    .Q_N(_0471_),
    .Q(\my_decimation_filter.decimation_count[3] ));
 sg13g2_dfrbp_1 _0998_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net15),
    .D(_0027_),
    .Q_N(_0470_),
    .Q(\my_decimation_filter.decimation_count[4] ));
 sg13g2_dfrbp_1 _0999_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net13),
    .D(net146),
    .Q_N(_0469_),
    .Q(\my_decimation_filter.decimation_count[5] ));
 sg13g2_dfrbp_1 _1000_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net11),
    .D(net165),
    .Q_N(_0000_),
    .Q(\my_decimation_filter.decimation_count[6] ));
 sg13g2_dfrbp_1 _1001_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net9),
    .D(net160),
    .Q_N(_0468_),
    .Q(\my_decimation_filter.comb_2[0] ));
 sg13g2_dfrbp_1 _1002_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net7),
    .D(_0031_),
    .Q_N(_0467_),
    .Q(\my_decimation_filter.comb_2[1] ));
 sg13g2_dfrbp_1 _1003_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net4),
    .D(_0032_),
    .Q_N(_0466_),
    .Q(\my_decimation_filter.comb_2[2] ));
 sg13g2_dfrbp_1 _1004_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net91),
    .D(net177),
    .Q_N(_0465_),
    .Q(\my_decimation_filter.comb_2[3] ));
 sg13g2_dfrbp_1 _1005_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net89),
    .D(_0034_),
    .Q_N(_0464_),
    .Q(\my_decimation_filter.comb_2[4] ));
 sg13g2_dfrbp_1 _1006_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net87),
    .D(net242),
    .Q_N(_0463_),
    .Q(\my_decimation_filter.comb_2[5] ));
 sg13g2_dfrbp_1 _1007_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net85),
    .D(net229),
    .Q_N(_0462_),
    .Q(\my_decimation_filter.comb_2[6] ));
 sg13g2_dfrbp_1 _1008_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net83),
    .D(net172),
    .Q_N(_0461_),
    .Q(\my_decimation_filter.comb_2[7] ));
 sg13g2_dfrbp_1 _1009_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net81),
    .D(_0038_),
    .Q_N(_0460_),
    .Q(\my_decimation_filter.comb_2[8] ));
 sg13g2_dfrbp_1 _1010_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net79),
    .D(_0039_),
    .Q_N(_0459_),
    .Q(\my_decimation_filter.comb_2[9] ));
 sg13g2_dfrbp_1 _1011_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net77),
    .D(net211),
    .Q_N(_0458_),
    .Q(\my_decimation_filter.comb_2[10] ));
 sg13g2_dfrbp_1 _1012_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net75),
    .D(_0041_),
    .Q_N(_0457_),
    .Q(\my_decimation_filter.comb_2[11] ));
 sg13g2_dfrbp_1 _1013_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net73),
    .D(_0042_),
    .Q_N(_0456_),
    .Q(\my_decimation_filter.comb_2[12] ));
 sg13g2_dfrbp_1 _1014_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net71),
    .D(net245),
    .Q_N(_0455_),
    .Q(\my_decimation_filter.comb_2[13] ));
 sg13g2_dfrbp_1 _1015_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net69),
    .D(_0044_),
    .Q_N(_0454_),
    .Q(\my_decimation_filter.comb_2[14] ));
 sg13g2_dfrbp_1 _1016_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net67),
    .D(_0045_),
    .Q_N(_0453_),
    .Q(\my_decimation_filter.comb_2[15] ));
 sg13g2_dfrbp_1 _1017_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net65),
    .D(net190),
    .Q_N(_0452_),
    .Q(\my_decimation_filter.comb_1[0] ));
 sg13g2_dfrbp_1 _1018_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net63),
    .D(net227),
    .Q_N(_0451_),
    .Q(\my_decimation_filter.comb_1[1] ));
 sg13g2_dfrbp_1 _1019_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net61),
    .D(net216),
    .Q_N(_0450_),
    .Q(\my_decimation_filter.comb_1[2] ));
 sg13g2_dfrbp_1 _1020_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net59),
    .D(net255),
    .Q_N(_0449_),
    .Q(\my_decimation_filter.comb_1[3] ));
 sg13g2_dfrbp_1 _1021_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net57),
    .D(net175),
    .Q_N(_0448_),
    .Q(\my_decimation_filter.comb_1[4] ));
 sg13g2_dfrbp_1 _1022_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net55),
    .D(_0051_),
    .Q_N(_0447_),
    .Q(\my_decimation_filter.comb_1[5] ));
 sg13g2_dfrbp_1 _1023_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net53),
    .D(_0052_),
    .Q_N(_0446_),
    .Q(\my_decimation_filter.comb_1[6] ));
 sg13g2_dfrbp_1 _1024_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net51),
    .D(_0053_),
    .Q_N(_0445_),
    .Q(\my_decimation_filter.comb_1[7] ));
 sg13g2_dfrbp_1 _1025_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net49),
    .D(net214),
    .Q_N(_0444_),
    .Q(\my_decimation_filter.comb_1[8] ));
 sg13g2_dfrbp_1 _1026_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net47),
    .D(net247),
    .Q_N(_0443_),
    .Q(\my_decimation_filter.comb_1[9] ));
 sg13g2_dfrbp_1 _1027_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net45),
    .D(_0056_),
    .Q_N(_0442_),
    .Q(\my_decimation_filter.comb_1[10] ));
 sg13g2_dfrbp_1 _1028_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net43),
    .D(net250),
    .Q_N(_0441_),
    .Q(\my_decimation_filter.comb_1[11] ));
 sg13g2_dfrbp_1 _1029_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net41),
    .D(net200),
    .Q_N(_0440_),
    .Q(\my_decimation_filter.comb_1[12] ));
 sg13g2_dfrbp_1 _1030_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net22),
    .D(_0059_),
    .Q_N(_0439_),
    .Q(\my_decimation_filter.comb_1[13] ));
 sg13g2_dfrbp_1 _1031_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net18),
    .D(net220),
    .Q_N(_0438_),
    .Q(\my_decimation_filter.comb_1[14] ));
 sg13g2_dfrbp_1 _1032_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net14),
    .D(net158),
    .Q_N(_0437_),
    .Q(\my_decimation_filter.comb_1[15] ));
 sg13g2_dfrbp_1 _1033_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net10),
    .D(_0062_),
    .Q_N(_0436_),
    .Q(\my_decimation_filter.Y[0] ));
 sg13g2_dfrbp_1 _1034_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net8),
    .D(_0063_),
    .Q_N(_0435_),
    .Q(\my_decimation_filter.Y[1] ));
 sg13g2_dfrbp_1 _1035_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net6),
    .D(_0064_),
    .Q_N(_0434_),
    .Q(\my_decimation_filter.Y[2] ));
 sg13g2_dfrbp_1 _1036_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net92),
    .D(_0065_),
    .Q_N(_0433_),
    .Q(\my_decimation_filter.Y[3] ));
 sg13g2_dfrbp_1 _1037_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net90),
    .D(_0066_),
    .Q_N(_0432_),
    .Q(\my_decimation_filter.Y[4] ));
 sg13g2_dfrbp_1 _1038_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net88),
    .D(_0067_),
    .Q_N(_0431_),
    .Q(\my_decimation_filter.Y[5] ));
 sg13g2_dfrbp_1 _1039_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net86),
    .D(_0068_),
    .Q_N(_0430_),
    .Q(\my_decimation_filter.Y[6] ));
 sg13g2_dfrbp_1 _1040_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net84),
    .D(net268),
    .Q_N(_0429_),
    .Q(\my_decimation_filter.Y[7] ));
 sg13g2_dfrbp_1 _1041_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net82),
    .D(_0070_),
    .Q_N(_0428_),
    .Q(\my_decimation_filter.Y[8] ));
 sg13g2_dfrbp_1 _1042_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net80),
    .D(_0071_),
    .Q_N(_0427_),
    .Q(\my_decimation_filter.Y[9] ));
 sg13g2_dfrbp_1 _1043_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net78),
    .D(_0072_),
    .Q_N(_0426_),
    .Q(\my_decimation_filter.Y[10] ));
 sg13g2_dfrbp_1 _1044_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net76),
    .D(_0073_),
    .Q_N(_0425_),
    .Q(\my_decimation_filter.Y[11] ));
 sg13g2_dfrbp_1 _1045_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net74),
    .D(_0074_),
    .Q_N(_0424_),
    .Q(\my_decimation_filter.Y[12] ));
 sg13g2_dfrbp_1 _1046_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net72),
    .D(_0075_),
    .Q_N(_0423_),
    .Q(\my_decimation_filter.Y[13] ));
 sg13g2_dfrbp_1 _1047_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net70),
    .D(net265),
    .Q_N(_0422_),
    .Q(\my_decimation_filter.Y[14] ));
 sg13g2_dfrbp_1 _1048_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net68),
    .D(_0077_),
    .Q_N(_0421_),
    .Q(\my_decimation_filter.Y[15] ));
 sg13g2_dfrbp_1 _1049_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net66),
    .D(net218),
    .Q_N(_0420_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _1050_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net62),
    .D(net194),
    .Q_N(_0419_),
    .Q(uio_out[1]));
 sg13g2_dfrbp_1 _1051_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net58),
    .D(net196),
    .Q_N(_0418_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _1052_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net54),
    .D(net202),
    .Q_N(_0417_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _1053_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net50),
    .D(net181),
    .Q_N(_0416_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _1054_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net46),
    .D(net207),
    .Q_N(_0415_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _1055_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net42),
    .D(net198),
    .Q_N(_0414_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _1056_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net20),
    .D(_0085_),
    .Q_N(_0413_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _1057_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net12),
    .D(net156),
    .Q_N(_0412_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1058_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net60),
    .D(net167),
    .Q_N(_0411_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1059_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net52),
    .D(net185),
    .Q_N(_0410_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1060_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net44),
    .D(net169),
    .Q_N(_0409_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1061_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net16),
    .D(net236),
    .Q_N(_0408_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1062_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net56),
    .D(net225),
    .Q_N(_0407_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1063_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net40),
    .D(net162),
    .Q_N(_0406_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1064_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net48),
    .D(net187),
    .Q_N(_0405_),
    .Q(uo_out[7]));
 sg13g2_tiehi _0977__5 (.L_HI(net5));
 sg13g2_tiehi _1035__6 (.L_HI(net6));
 sg13g2_tiehi _1002__7 (.L_HI(net7));
 sg13g2_tiehi _1034__8 (.L_HI(net8));
 sg13g2_tiehi _1001__9 (.L_HI(net9));
 sg13g2_tiehi _1033__10 (.L_HI(net10));
 sg13g2_tiehi _1000__11 (.L_HI(net11));
 sg13g2_tiehi _1057__12 (.L_HI(net12));
 sg13g2_tiehi _0999__13 (.L_HI(net13));
 sg13g2_tiehi _1032__14 (.L_HI(net14));
 sg13g2_tiehi _0998__15 (.L_HI(net15));
 sg13g2_tiehi _1061__16 (.L_HI(net16));
 sg13g2_tiehi _0997__17 (.L_HI(net17));
 sg13g2_tiehi _1031__18 (.L_HI(net18));
 sg13g2_tiehi _0996__19 (.L_HI(net19));
 sg13g2_tiehi _1056__20 (.L_HI(net20));
 sg13g2_tiehi _0995__21 (.L_HI(net21));
 sg13g2_tiehi _1030__22 (.L_HI(net22));
 sg13g2_tiehi _0994__23 (.L_HI(net23));
 sg13g2_tiehi _0993__24 (.L_HI(net24));
 sg13g2_tiehi _0992__25 (.L_HI(net25));
 sg13g2_tiehi _0991__26 (.L_HI(net26));
 sg13g2_tiehi _0990__27 (.L_HI(net27));
 sg13g2_tiehi _0989__28 (.L_HI(net28));
 sg13g2_tiehi _0988__29 (.L_HI(net29));
 sg13g2_tiehi _0987__30 (.L_HI(net30));
 sg13g2_tiehi _0986__31 (.L_HI(net31));
 sg13g2_tiehi _0985__32 (.L_HI(net32));
 sg13g2_tiehi _0984__33 (.L_HI(net33));
 sg13g2_tiehi _0983__34 (.L_HI(net34));
 sg13g2_tiehi _0982__35 (.L_HI(net35));
 sg13g2_tiehi _0981__36 (.L_HI(net36));
 sg13g2_tiehi _0980__37 (.L_HI(net37));
 sg13g2_tiehi _0979__38 (.L_HI(net38));
 sg13g2_tiehi _0978__39 (.L_HI(net39));
 sg13g2_tiehi _1063__40 (.L_HI(net40));
 sg13g2_tiehi _1029__41 (.L_HI(net41));
 sg13g2_tiehi _1055__42 (.L_HI(net42));
 sg13g2_tiehi _1028__43 (.L_HI(net43));
 sg13g2_tiehi _1060__44 (.L_HI(net44));
 sg13g2_tiehi _1027__45 (.L_HI(net45));
 sg13g2_tiehi _1054__46 (.L_HI(net46));
 sg13g2_tiehi _1026__47 (.L_HI(net47));
 sg13g2_tiehi _1064__48 (.L_HI(net48));
 sg13g2_tiehi _1025__49 (.L_HI(net49));
 sg13g2_tiehi _1053__50 (.L_HI(net50));
 sg13g2_tiehi _1024__51 (.L_HI(net51));
 sg13g2_tiehi _1059__52 (.L_HI(net52));
 sg13g2_tiehi _1023__53 (.L_HI(net53));
 sg13g2_tiehi _1052__54 (.L_HI(net54));
 sg13g2_tiehi _1022__55 (.L_HI(net55));
 sg13g2_tiehi _1062__56 (.L_HI(net56));
 sg13g2_tiehi _1021__57 (.L_HI(net57));
 sg13g2_tiehi _1051__58 (.L_HI(net58));
 sg13g2_tiehi _1020__59 (.L_HI(net59));
 sg13g2_tiehi _1058__60 (.L_HI(net60));
 sg13g2_tiehi _1019__61 (.L_HI(net61));
 sg13g2_tiehi _1050__62 (.L_HI(net62));
 sg13g2_tiehi _1018__63 (.L_HI(net63));
 sg13g2_tiehi _0976__64 (.L_HI(net64));
 sg13g2_tiehi _1017__65 (.L_HI(net65));
 sg13g2_tiehi _1049__66 (.L_HI(net66));
 sg13g2_tiehi _1016__67 (.L_HI(net67));
 sg13g2_tiehi _1048__68 (.L_HI(net68));
 sg13g2_tiehi _1015__69 (.L_HI(net69));
 sg13g2_tiehi _1047__70 (.L_HI(net70));
 sg13g2_tiehi _1014__71 (.L_HI(net71));
 sg13g2_tiehi _1046__72 (.L_HI(net72));
 sg13g2_tiehi _1013__73 (.L_HI(net73));
 sg13g2_tiehi _1045__74 (.L_HI(net74));
 sg13g2_tiehi _1012__75 (.L_HI(net75));
 sg13g2_tiehi _1044__76 (.L_HI(net76));
 sg13g2_tiehi _1011__77 (.L_HI(net77));
 sg13g2_tiehi _1043__78 (.L_HI(net78));
 sg13g2_tiehi _1010__79 (.L_HI(net79));
 sg13g2_tiehi _1042__80 (.L_HI(net80));
 sg13g2_tiehi _1009__81 (.L_HI(net81));
 sg13g2_tiehi _1041__82 (.L_HI(net82));
 sg13g2_tiehi _1008__83 (.L_HI(net83));
 sg13g2_tiehi _1040__84 (.L_HI(net84));
 sg13g2_tiehi _1007__85 (.L_HI(net85));
 sg13g2_tiehi _1039__86 (.L_HI(net86));
 sg13g2_tiehi _1006__87 (.L_HI(net87));
 sg13g2_tiehi _1038__88 (.L_HI(net88));
 sg13g2_tiehi _1005__89 (.L_HI(net89));
 sg13g2_tiehi _1037__90 (.L_HI(net90));
 sg13g2_tiehi _1004__91 (.L_HI(net91));
 sg13g2_tiehi _1036__92 (.L_HI(net92));
 sg13g2_tiehi tt_um_murmann_group_93 (.L_HI(net93));
 sg13g2_tiehi tt_um_murmann_group_94 (.L_HI(net94));
 sg13g2_tiehi tt_um_murmann_group_95 (.L_HI(net95));
 sg13g2_tiehi tt_um_murmann_group_96 (.L_HI(net96));
 sg13g2_tiehi tt_um_murmann_group_97 (.L_HI(net97));
 sg13g2_tiehi tt_um_murmann_group_98 (.L_HI(net98));
 sg13g2_tiehi tt_um_murmann_group_99 (.L_HI(net99));
 sg13g2_tiehi tt_um_murmann_group_100 (.L_HI(net100));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 fanout109 (.A(net110),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(net111),
    .X(net110));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(_0134_));
 sg13g2_buf_2 fanout112 (.A(_0133_),
    .X(net112));
 sg13g2_buf_1 fanout113 (.A(_0133_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0130_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_0130_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_0129_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_0129_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(net119),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(net122),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(net122),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(net122),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_0125_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(net124),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(net125),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_0124_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(net128),
    .X(net126));
 sg13g2_buf_1 fanout127 (.A(net128),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_0124_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(net131),
    .X(net129));
 sg13g2_buf_1 fanout130 (.A(net131),
    .X(net130));
 sg13g2_buf_1 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(net135),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(net135),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_0131_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_1 fanout137 (.A(net138),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_0128_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_0290_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_0290_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(net142),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(ui_in[2]),
    .X(net142));
 sg13g2_buf_1 fanout143 (.A(ui_in[2]),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(net3),
    .X(net144));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_tiehi _1003__4 (.L_HI(net4));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0005_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0021_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0001_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0138_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0008_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0004_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0160_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0019_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold9 (.A(\my_decimation_filter.decimation_count[5] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0028_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold11 (.A(\my_decimation_filter.decimation_count[1] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0167_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0024_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0002_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0144_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold16 (.A(\my_decimation_filter.decimation_count[0] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0003_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0151_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold19 (.A(uo_out[0]),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0086_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold21 (.A(\my_decimation_filter.comb_1[15] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0061_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold23 (.A(\my_decimation_filter.comb_1[0] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0030_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold25 (.A(uo_out[6]),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0092_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold27 (.A(\my_decimation_filter.comb_2[15] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold28 (.A(\my_decimation_filter.decimation_count[6] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0029_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold30 (.A(uo_out[1]),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0087_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold32 (.A(uo_out[3]),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0089_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold34 (.A(\my_decimation_filter.input_accumulator[9] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold35 (.A(\my_decimation_filter.comb_1[7] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0037_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold37 (.A(\my_decimation_filter.input_accumulator[5] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold38 (.A(\my_decimation_filter.comb_1[4] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0050_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold40 (.A(\my_decimation_filter.comb_2[3] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0033_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold42 (.A(\my_decimation_filter.input_accumulator[10] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0155_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold44 (.A(uio_out[4]),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0082_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold46 (.A(\my_decimation_filter.comb_2[4] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold47 (.A(\my_decimation_filter.Y[7] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold48 (.A(uo_out[2]),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0088_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold50 (.A(uo_out[7]),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0093_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold52 (.A(\my_decimation_filter.Y[0] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0192_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0046_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold55 (.A(\my_decimation_filter.decimation_count[4] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0171_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold57 (.A(uio_out[1]),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0079_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold59 (.A(uio_out[2]),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0080_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold61 (.A(uio_out[6]),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0084_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold63 (.A(\my_decimation_filter.comb_1[12] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0058_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold65 (.A(uio_out[3]),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0081_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold67 (.A(\my_decimation_filter.comb_2[12] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold68 (.A(\my_decimation_filter.input_accumulator[6] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0147_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold70 (.A(uio_out[5]),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0083_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold72 (.A(\my_decimation_filter.input_accumulator[15] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0165_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold74 (.A(\my_decimation_filter.comb_1[10] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0040_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold76 (.A(uio_out[7]),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold77 (.A(\my_decimation_filter.comb_1[8] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0054_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold79 (.A(\my_decimation_filter.comb_1[2] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0048_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold81 (.A(uio_out[0]),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0078_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold83 (.A(\my_decimation_filter.comb_1[14] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0060_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold85 (.A(\my_decimation_filter.Y[10] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold86 (.A(\my_decimation_filter.input_accumulator[3] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0142_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold88 (.A(uo_out[5]),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0091_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold90 (.A(\my_decimation_filter.comb_1[1] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0047_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold92 (.A(\my_decimation_filter.comb_1[6] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0036_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold94 (.A(\my_decimation_filter.comb_2[1] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold95 (.A(\my_decimation_filter.Y[6] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold96 (.A(\my_decimation_filter.comb_2[14] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold97 (.A(\my_decimation_filter.input_accumulator[2] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0140_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold99 (.A(uo_out[4]),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0090_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold101 (.A(\my_decimation_filter.comb_2[8] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold102 (.A(\my_decimation_filter.input_accumulator[13] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0020_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold104 (.A(\my_decimation_filter.decimation_count[2] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold105 (.A(\my_decimation_filter.comb_1[5] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0035_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold107 (.A(\my_decimation_filter.comb_2[2] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold108 (.A(\my_decimation_filter.comb_1[13] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0043_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold110 (.A(\my_decimation_filter.comb_1[9] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0055_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold112 (.A(\my_decimation_filter.decimation_count[3] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold113 (.A(\my_decimation_filter.comb_1[11] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0057_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold115 (.A(\my_decimation_filter.comb_2[11] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold116 (.A(\my_decimation_filter.Y[5] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold117 (.A(\my_decimation_filter.comb_2[9] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold118 (.A(\my_decimation_filter.Y[3] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0049_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold120 (.A(\my_decimation_filter.input_accumulator[0] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold121 (.A(\my_decimation_filter.Y[13] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold122 (.A(\my_decimation_filter.input_accumulator[7] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold123 (.A(\my_decimation_filter.input_accumulator[11] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold124 (.A(\my_decimation_filter.Y[9] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold125 (.A(\my_decimation_filter.input_accumulator[1] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0212_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold127 (.A(\my_decimation_filter.input_accumulator[14] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0281_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0076_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold130 (.A(\my_decimation_filter.input_accumulator[6] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0241_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0069_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold133 (.A(\my_decimation_filter.Y[1] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0217_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold135 (.A(\my_decimation_filter.input_accumulator[8] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold136 (.A(\my_decimation_filter.input_accumulator[2] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0221_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold138 (.A(\my_decimation_filter.Y[15] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold139 (.A(\my_decimation_filter.input_accumulator[12] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0269_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0274_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold142 (.A(\my_decimation_filter.input_accumulator[4] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold143 (.A(\my_decimation_filter.input_accumulator[3] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold144 (.A(\my_decimation_filter.input_accumulator[9] ),
    .X(net280));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_4 FILLER_18_203 ();
 sg13g2_fill_1 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_211 ();
 sg13g2_fill_2 FILLER_18_218 ();
 sg13g2_fill_1 FILLER_18_220 ();
 sg13g2_decap_8 FILLER_18_230 ();
 sg13g2_decap_8 FILLER_18_237 ();
 sg13g2_decap_4 FILLER_18_244 ();
 sg13g2_fill_2 FILLER_18_248 ();
 sg13g2_decap_8 FILLER_18_276 ();
 sg13g2_decap_8 FILLER_18_283 ();
 sg13g2_decap_8 FILLER_18_290 ();
 sg13g2_decap_8 FILLER_18_297 ();
 sg13g2_decap_8 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_decap_8 FILLER_18_318 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_decap_8 FILLER_18_332 ();
 sg13g2_decap_8 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_4 FILLER_19_56 ();
 sg13g2_decap_4 FILLER_19_64 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_4 FILLER_19_119 ();
 sg13g2_fill_1 FILLER_19_123 ();
 sg13g2_decap_8 FILLER_19_128 ();
 sg13g2_decap_8 FILLER_19_135 ();
 sg13g2_decap_8 FILLER_19_142 ();
 sg13g2_decap_8 FILLER_19_149 ();
 sg13g2_decap_8 FILLER_19_156 ();
 sg13g2_decap_8 FILLER_19_163 ();
 sg13g2_decap_4 FILLER_19_170 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_decap_8 FILLER_19_180 ();
 sg13g2_decap_8 FILLER_19_187 ();
 sg13g2_fill_2 FILLER_19_194 ();
 sg13g2_fill_1 FILLER_19_196 ();
 sg13g2_fill_1 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_267 ();
 sg13g2_fill_2 FILLER_19_274 ();
 sg13g2_fill_1 FILLER_19_302 ();
 sg13g2_fill_2 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_fill_2 FILLER_20_58 ();
 sg13g2_fill_1 FILLER_20_60 ();
 sg13g2_fill_1 FILLER_20_69 ();
 sg13g2_fill_2 FILLER_20_80 ();
 sg13g2_fill_1 FILLER_20_82 ();
 sg13g2_fill_1 FILLER_20_100 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_4 FILLER_20_112 ();
 sg13g2_fill_1 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_143 ();
 sg13g2_decap_8 FILLER_20_150 ();
 sg13g2_decap_4 FILLER_20_157 ();
 sg13g2_fill_2 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_233 ();
 sg13g2_fill_1 FILLER_20_246 ();
 sg13g2_fill_2 FILLER_20_252 ();
 sg13g2_fill_1 FILLER_20_254 ();
 sg13g2_fill_1 FILLER_20_260 ();
 sg13g2_decap_8 FILLER_20_265 ();
 sg13g2_decap_8 FILLER_20_276 ();
 sg13g2_fill_1 FILLER_20_283 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_4 FILLER_21_28 ();
 sg13g2_fill_1 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_66 ();
 sg13g2_fill_1 FILLER_21_68 ();
 sg13g2_fill_2 FILLER_21_88 ();
 sg13g2_fill_1 FILLER_21_90 ();
 sg13g2_fill_1 FILLER_21_117 ();
 sg13g2_fill_2 FILLER_21_185 ();
 sg13g2_decap_4 FILLER_21_204 ();
 sg13g2_fill_2 FILLER_21_222 ();
 sg13g2_fill_1 FILLER_21_245 ();
 sg13g2_fill_1 FILLER_21_258 ();
 sg13g2_fill_2 FILLER_21_271 ();
 sg13g2_fill_1 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_331 ();
 sg13g2_decap_8 FILLER_21_338 ();
 sg13g2_decap_8 FILLER_21_345 ();
 sg13g2_decap_8 FILLER_21_352 ();
 sg13g2_decap_8 FILLER_21_359 ();
 sg13g2_decap_8 FILLER_21_366 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_fill_1 FILLER_22_28 ();
 sg13g2_fill_2 FILLER_22_109 ();
 sg13g2_fill_1 FILLER_22_111 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_fill_1 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_210 ();
 sg13g2_decap_4 FILLER_22_225 ();
 sg13g2_fill_1 FILLER_22_237 ();
 sg13g2_decap_8 FILLER_22_251 ();
 sg13g2_fill_2 FILLER_22_258 ();
 sg13g2_fill_1 FILLER_22_260 ();
 sg13g2_fill_1 FILLER_22_274 ();
 sg13g2_fill_2 FILLER_22_302 ();
 sg13g2_fill_1 FILLER_22_313 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_2 FILLER_23_73 ();
 sg13g2_fill_2 FILLER_23_89 ();
 sg13g2_fill_1 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_122 ();
 sg13g2_fill_1 FILLER_23_124 ();
 sg13g2_fill_2 FILLER_23_152 ();
 sg13g2_fill_2 FILLER_23_173 ();
 sg13g2_fill_1 FILLER_23_193 ();
 sg13g2_fill_2 FILLER_23_203 ();
 sg13g2_fill_2 FILLER_23_214 ();
 sg13g2_fill_1 FILLER_23_216 ();
 sg13g2_decap_8 FILLER_23_230 ();
 sg13g2_fill_2 FILLER_23_242 ();
 sg13g2_fill_2 FILLER_23_248 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_fill_1 FILLER_23_260 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_decap_8 FILLER_23_355 ();
 sg13g2_decap_8 FILLER_23_362 ();
 sg13g2_decap_8 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_376 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_46 ();
 sg13g2_fill_1 FILLER_24_48 ();
 sg13g2_fill_2 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_150 ();
 sg13g2_fill_1 FILLER_24_152 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_decap_4 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_decap_8 FILLER_24_361 ();
 sg13g2_decap_8 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_14 ();
 sg13g2_fill_1 FILLER_25_138 ();
 sg13g2_decap_8 FILLER_25_165 ();
 sg13g2_fill_2 FILLER_25_181 ();
 sg13g2_fill_1 FILLER_25_183 ();
 sg13g2_fill_2 FILLER_25_201 ();
 sg13g2_decap_4 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_217 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_1 FILLER_25_282 ();
 sg13g2_fill_2 FILLER_25_343 ();
 sg13g2_fill_1 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_25 ();
 sg13g2_decap_4 FILLER_26_30 ();
 sg13g2_fill_1 FILLER_26_34 ();
 sg13g2_fill_1 FILLER_26_39 ();
 sg13g2_decap_4 FILLER_26_57 ();
 sg13g2_fill_1 FILLER_26_78 ();
 sg13g2_fill_1 FILLER_26_97 ();
 sg13g2_fill_2 FILLER_26_141 ();
 sg13g2_decap_4 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_203 ();
 sg13g2_fill_2 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_254 ();
 sg13g2_fill_1 FILLER_26_311 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_fill_1 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_352 ();
 sg13g2_decap_8 FILLER_26_359 ();
 sg13g2_decap_8 FILLER_26_366 ();
 sg13g2_decap_8 FILLER_26_373 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_23 ();
 sg13g2_fill_1 FILLER_27_50 ();
 sg13g2_fill_1 FILLER_27_55 ();
 sg13g2_fill_2 FILLER_27_116 ();
 sg13g2_fill_2 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_146 ();
 sg13g2_fill_2 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_269 ();
 sg13g2_fill_1 FILLER_27_271 ();
 sg13g2_fill_1 FILLER_27_277 ();
 sg13g2_fill_1 FILLER_27_291 ();
 sg13g2_fill_2 FILLER_27_318 ();
 sg13g2_fill_1 FILLER_27_349 ();
 sg13g2_decap_8 FILLER_27_354 ();
 sg13g2_decap_8 FILLER_27_361 ();
 sg13g2_decap_8 FILLER_27_368 ();
 sg13g2_decap_8 FILLER_27_375 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_68 ();
 sg13g2_fill_1 FILLER_28_80 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_129 ();
 sg13g2_fill_2 FILLER_28_195 ();
 sg13g2_decap_4 FILLER_28_227 ();
 sg13g2_fill_1 FILLER_28_283 ();
 sg13g2_decap_4 FILLER_28_293 ();
 sg13g2_fill_2 FILLER_28_297 ();
 sg13g2_fill_2 FILLER_28_309 ();
 sg13g2_fill_1 FILLER_28_321 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_4 FILLER_29_14 ();
 sg13g2_fill_1 FILLER_29_18 ();
 sg13g2_fill_2 FILLER_29_50 ();
 sg13g2_fill_1 FILLER_29_61 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_fill_2 FILLER_29_178 ();
 sg13g2_fill_1 FILLER_29_203 ();
 sg13g2_fill_1 FILLER_29_258 ();
 sg13g2_fill_2 FILLER_29_273 ();
 sg13g2_fill_1 FILLER_29_279 ();
 sg13g2_decap_4 FILLER_29_299 ();
 sg13g2_decap_4 FILLER_29_359 ();
 sg13g2_fill_2 FILLER_29_368 ();
 sg13g2_fill_1 FILLER_29_393 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_23 ();
 sg13g2_fill_2 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_34 ();
 sg13g2_fill_1 FILLER_30_36 ();
 sg13g2_fill_2 FILLER_30_75 ();
 sg13g2_fill_2 FILLER_30_82 ();
 sg13g2_fill_1 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_100 ();
 sg13g2_fill_2 FILLER_30_122 ();
 sg13g2_fill_2 FILLER_30_137 ();
 sg13g2_fill_1 FILLER_30_139 ();
 sg13g2_fill_2 FILLER_30_145 ();
 sg13g2_fill_2 FILLER_30_213 ();
 sg13g2_fill_1 FILLER_30_215 ();
 sg13g2_fill_2 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_330 ();
 sg13g2_fill_1 FILLER_30_367 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_11 ();
 sg13g2_fill_1 FILLER_31_85 ();
 sg13g2_fill_2 FILLER_31_95 ();
 sg13g2_fill_1 FILLER_31_97 ();
 sg13g2_fill_2 FILLER_31_119 ();
 sg13g2_fill_1 FILLER_31_151 ();
 sg13g2_decap_4 FILLER_31_201 ();
 sg13g2_fill_2 FILLER_31_219 ();
 sg13g2_decap_4 FILLER_31_259 ();
 sg13g2_fill_1 FILLER_31_279 ();
 sg13g2_fill_2 FILLER_31_302 ();
 sg13g2_fill_1 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_357 ();
 sg13g2_fill_1 FILLER_31_359 ();
 sg13g2_fill_1 FILLER_31_367 ();
 sg13g2_fill_1 FILLER_31_372 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_16 ();
 sg13g2_fill_2 FILLER_32_43 ();
 sg13g2_fill_2 FILLER_32_73 ();
 sg13g2_fill_1 FILLER_32_88 ();
 sg13g2_fill_2 FILLER_32_116 ();
 sg13g2_fill_1 FILLER_32_118 ();
 sg13g2_fill_1 FILLER_32_132 ();
 sg13g2_fill_2 FILLER_32_158 ();
 sg13g2_fill_2 FILLER_32_173 ();
 sg13g2_fill_2 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_199 ();
 sg13g2_fill_1 FILLER_32_206 ();
 sg13g2_decap_4 FILLER_32_235 ();
 sg13g2_fill_2 FILLER_32_254 ();
 sg13g2_decap_8 FILLER_32_261 ();
 sg13g2_fill_2 FILLER_32_268 ();
 sg13g2_decap_4 FILLER_32_288 ();
 sg13g2_fill_2 FILLER_32_292 ();
 sg13g2_decap_8 FILLER_32_320 ();
 sg13g2_decap_4 FILLER_32_327 ();
 sg13g2_fill_2 FILLER_32_335 ();
 sg13g2_fill_1 FILLER_32_374 ();
 sg13g2_fill_2 FILLER_32_380 ();
 sg13g2_fill_1 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_4 FILLER_33_21 ();
 sg13g2_fill_2 FILLER_33_25 ();
 sg13g2_fill_1 FILLER_33_31 ();
 sg13g2_fill_1 FILLER_33_69 ();
 sg13g2_fill_1 FILLER_33_80 ();
 sg13g2_fill_1 FILLER_33_96 ();
 sg13g2_fill_1 FILLER_33_116 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_fill_2 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_180 ();
 sg13g2_fill_2 FILLER_33_213 ();
 sg13g2_decap_4 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_246 ();
 sg13g2_fill_2 FILLER_33_251 ();
 sg13g2_fill_2 FILLER_33_280 ();
 sg13g2_fill_1 FILLER_33_282 ();
 sg13g2_fill_1 FILLER_33_374 ();
 sg13g2_fill_1 FILLER_33_392 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_54 ();
 sg13g2_fill_2 FILLER_34_82 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_fill_2 FILLER_34_196 ();
 sg13g2_decap_4 FILLER_34_211 ();
 sg13g2_fill_2 FILLER_34_215 ();
 sg13g2_fill_1 FILLER_34_297 ();
 sg13g2_fill_2 FILLER_34_307 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_4 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_18 ();
 sg13g2_fill_1 FILLER_35_102 ();
 sg13g2_fill_2 FILLER_35_108 ();
 sg13g2_fill_2 FILLER_35_118 ();
 sg13g2_fill_1 FILLER_35_144 ();
 sg13g2_fill_2 FILLER_35_186 ();
 sg13g2_fill_1 FILLER_35_188 ();
 sg13g2_decap_4 FILLER_35_229 ();
 sg13g2_decap_4 FILLER_35_241 ();
 sg13g2_fill_2 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_347 ();
 sg13g2_fill_2 FILLER_35_379 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_21 ();
 sg13g2_fill_2 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_58 ();
 sg13g2_fill_1 FILLER_36_77 ();
 sg13g2_fill_2 FILLER_36_92 ();
 sg13g2_fill_1 FILLER_36_108 ();
 sg13g2_fill_2 FILLER_36_134 ();
 sg13g2_fill_1 FILLER_36_168 ();
 sg13g2_fill_1 FILLER_36_174 ();
 sg13g2_fill_2 FILLER_36_189 ();
 sg13g2_fill_1 FILLER_36_191 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_255 ();
 sg13g2_fill_2 FILLER_36_270 ();
 sg13g2_fill_2 FILLER_36_294 ();
 sg13g2_fill_1 FILLER_36_301 ();
 sg13g2_fill_1 FILLER_36_307 ();
 sg13g2_fill_2 FILLER_36_331 ();
 sg13g2_fill_1 FILLER_36_333 ();
 sg13g2_fill_2 FILLER_36_351 ();
 sg13g2_fill_2 FILLER_36_361 ();
 sg13g2_fill_1 FILLER_36_377 ();
 sg13g2_fill_1 FILLER_36_391 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_21 ();
 sg13g2_fill_2 FILLER_37_60 ();
 sg13g2_fill_2 FILLER_37_135 ();
 sg13g2_fill_2 FILLER_37_276 ();
 sg13g2_fill_1 FILLER_37_343 ();
 sg13g2_fill_2 FILLER_37_361 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_fill_1 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_77 ();
 sg13g2_fill_2 FILLER_38_181 ();
 sg13g2_fill_2 FILLER_38_218 ();
 sg13g2_fill_1 FILLER_38_220 ();
 sg13g2_fill_1 FILLER_38_255 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_fill_2 FILLER_38_321 ();
 sg13g2_fill_1 FILLER_38_323 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net93;
 assign uio_oe[1] = net94;
 assign uio_oe[2] = net95;
 assign uio_oe[3] = net96;
 assign uio_oe[4] = net97;
 assign uio_oe[5] = net98;
 assign uio_oe[6] = net99;
 assign uio_oe[7] = net100;
endmodule

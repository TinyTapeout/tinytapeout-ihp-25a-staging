module tt_um_vga_glyph_mode (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire clknet_0_clk;
 wire \a[0] ;
 wire \a[1] ;
 wire b;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \div3.in[0] ;
 wire \div3.in[1] ;
 wire \div3.in[2] ;
 wire \div3.in[3] ;
 wire \div3.in[4] ;
 wire \div3.in[5] ;
 wire \div3.in[6] ;
 wire \div3.out[0] ;
 wire \div3.out[1] ;
 wire \div3.out[2] ;
 wire \div3.out[3] ;
 wire \div3.out[4] ;
 wire \div3.out[5] ;
 wire \g_x[0] ;
 wire \g_x[1] ;
 wire \g_x[2] ;
 wire hsync;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;

 sg13g2_inv_2 _1127_ (.Y(_0167_),
    .A(net91));
 sg13g2_inv_1 _1128_ (.Y(_0175_),
    .A(\hvsync_gen.hpos[9] ));
 sg13g2_inv_1 _1129_ (.Y(_0182_),
    .A(net82));
 sg13g2_inv_1 _1130_ (.Y(_0189_),
    .A(\g_x[0] ));
 sg13g2_inv_1 _1131_ (.Y(_0197_),
    .A(\g_x[1] ));
 sg13g2_inv_1 _1132_ (.Y(_0202_),
    .A(net60));
 sg13g2_inv_1 _1133_ (.Y(_0203_),
    .A(net429));
 sg13g2_inv_1 _1134_ (.Y(_0204_),
    .A(net2));
 sg13g2_inv_1 _1135_ (.Y(_0205_),
    .A(\div3.in[2] ));
 sg13g2_inv_1 _1136_ (.Y(_0206_),
    .A(\hvsync_gen.vpos[9] ));
 sg13g2_inv_1 _1137_ (.Y(_0207_),
    .A(\counter[3] ));
 sg13g2_inv_2 _1138_ (.Y(_0208_),
    .A(net428));
 sg13g2_inv_1 _1139_ (.Y(_0209_),
    .A(net64));
 sg13g2_inv_1 _1140_ (.Y(_0210_),
    .A(_0031_));
 sg13g2_nor2_1 _1141_ (.A(\div3.out[0] ),
    .B(\div3.in[0] ),
    .Y(_0211_));
 sg13g2_xor2_1 _1142_ (.B(\div3.in[0] ),
    .A(\div3.out[0] ),
    .X(_0212_));
 sg13g2_xnor2_1 _1143_ (.Y(_0213_),
    .A(\div3.out[0] ),
    .B(\div3.in[0] ));
 sg13g2_xor2_1 _1144_ (.B(\div3.out[1] ),
    .A(\div3.in[1] ),
    .X(_0214_));
 sg13g2_and2_2 _1145_ (.A(_0212_),
    .B(_0214_),
    .X(_0215_));
 sg13g2_nand2_2 _1146_ (.Y(_0216_),
    .A(_0212_),
    .B(_0214_));
 sg13g2_xor2_1 _1147_ (.B(\div3.out[3] ),
    .A(\hvsync_gen.hpos[7] ),
    .X(_0217_));
 sg13g2_nor2_1 _1148_ (.A(\hvsync_gen.hpos[8] ),
    .B(\hvsync_gen.hpos[7] ),
    .Y(_0218_));
 sg13g2_xor2_1 _1149_ (.B(\hvsync_gen.hpos[7] ),
    .A(\hvsync_gen.hpos[8] ),
    .X(_0219_));
 sg13g2_xnor2_1 _1150_ (.Y(_0220_),
    .A(_0029_),
    .B(_0219_));
 sg13g2_xnor2_1 _1151_ (.Y(_0221_),
    .A(net423),
    .B(net428));
 sg13g2_xor2_1 _1152_ (.B(net427),
    .A(net424),
    .X(_0222_));
 sg13g2_nand2_1 _1153_ (.Y(_0223_),
    .A(net426),
    .B(\hvsync_gen.hpos[6] ));
 sg13g2_or2_1 _1154_ (.X(_0224_),
    .B(\hvsync_gen.hpos[6] ),
    .A(net426));
 sg13g2_xor2_1 _1155_ (.B(\hvsync_gen.hpos[6] ),
    .A(net426),
    .X(_0225_));
 sg13g2_xnor2_1 _1156_ (.Y(_0226_),
    .A(_0221_),
    .B(_0225_));
 sg13g2_xor2_1 _1157_ (.B(_0226_),
    .A(_0220_),
    .X(_0227_));
 sg13g2_xnor2_1 _1158_ (.Y(_0228_),
    .A(_0220_),
    .B(_0226_));
 sg13g2_mux2_1 _1159_ (.A0(_0026_),
    .A1(_0025_),
    .S(_0228_),
    .X(_0229_));
 sg13g2_xor2_1 _1160_ (.B(_0229_),
    .A(_0029_),
    .X(_0230_));
 sg13g2_nor2b_1 _1161_ (.A(_0230_),
    .B_N(_0033_),
    .Y(_0231_));
 sg13g2_nor2_1 _1162_ (.A(\hvsync_gen.hpos[9] ),
    .B(_0229_),
    .Y(_0232_));
 sg13g2_nor2_1 _1163_ (.A(_0231_),
    .B(_0232_),
    .Y(_0233_));
 sg13g2_mux2_1 _1164_ (.A0(_0024_),
    .A1(_0025_),
    .S(_0227_),
    .X(_0234_));
 sg13g2_xor2_1 _1165_ (.B(_0234_),
    .A(_0019_),
    .X(_0235_));
 sg13g2_nor2b_1 _1166_ (.A(_0235_),
    .B_N(_0034_),
    .Y(_0236_));
 sg13g2_xnor2_1 _1167_ (.Y(_0237_),
    .A(_0034_),
    .B(_0235_));
 sg13g2_nor2b_1 _1168_ (.A(_0233_),
    .B_N(_0237_),
    .Y(_0238_));
 sg13g2_mux2_1 _1169_ (.A0(_0026_),
    .A1(_0027_),
    .S(_0227_),
    .X(_0239_));
 sg13g2_nand2b_1 _1170_ (.Y(_0240_),
    .B(_0239_),
    .A_N(_0020_));
 sg13g2_xnor2_1 _1171_ (.Y(_0241_),
    .A(_0033_),
    .B(_0230_));
 sg13g2_nand2_1 _1172_ (.Y(_0242_),
    .A(_0240_),
    .B(_0241_));
 sg13g2_xnor2_1 _1173_ (.Y(_0243_),
    .A(_0020_),
    .B(_0239_));
 sg13g2_nand3b_1 _1174_ (.B(\counter[3] ),
    .C(_0228_),
    .Y(_0244_),
    .A_N(net423));
 sg13g2_o21ai_1 _1175_ (.B1(net423),
    .Y(_0245_),
    .A1(_0207_),
    .A2(_0227_));
 sg13g2_nand3_1 _1176_ (.B(_0244_),
    .C(_0245_),
    .A(_0031_),
    .Y(_0246_));
 sg13g2_nand3_1 _1177_ (.B(_0018_),
    .C(_0228_),
    .A(\counter[3] ),
    .Y(_0247_));
 sg13g2_a21oi_1 _1178_ (.A1(_0246_),
    .A2(_0247_),
    .Y(_0248_),
    .B1(_0243_));
 sg13g2_nand3_1 _1179_ (.B(_0246_),
    .C(_0247_),
    .A(_0243_),
    .Y(_0249_));
 sg13g2_nor2b_1 _1180_ (.A(_0248_),
    .B_N(_0249_),
    .Y(_0250_));
 sg13g2_a21oi_1 _1181_ (.A1(_0032_),
    .A2(_0249_),
    .Y(_0251_),
    .B1(_0248_));
 sg13g2_xnor2_1 _1182_ (.Y(_0252_),
    .A(_0240_),
    .B(_0241_));
 sg13g2_o21ai_1 _1183_ (.B1(_0242_),
    .Y(_0253_),
    .A1(_0251_),
    .A2(_0252_));
 sg13g2_xnor2_1 _1184_ (.Y(_0254_),
    .A(_0233_),
    .B(_0237_));
 sg13g2_a21oi_1 _1185_ (.A1(_0253_),
    .A2(_0254_),
    .Y(_0255_),
    .B1(_0238_));
 sg13g2_nor2_1 _1186_ (.A(net426),
    .B(_0234_),
    .Y(_0256_));
 sg13g2_nor2_1 _1187_ (.A(_0236_),
    .B(_0256_),
    .Y(_0257_));
 sg13g2_mux2_1 _1188_ (.A0(_0024_),
    .A1(_0023_),
    .S(_0228_),
    .X(_0258_));
 sg13g2_xor2_1 _1189_ (.B(_0258_),
    .A(_0016_),
    .X(_0259_));
 sg13g2_nor2b_1 _1190_ (.A(_0259_),
    .B_N(_0007_),
    .Y(_0260_));
 sg13g2_xnor2_1 _1191_ (.Y(_0261_),
    .A(_0007_),
    .B(_0259_));
 sg13g2_o21ai_1 _1192_ (.B1(_0261_),
    .Y(_0262_),
    .A1(_0236_),
    .A2(_0256_));
 sg13g2_xnor2_1 _1193_ (.Y(_0263_),
    .A(_0257_),
    .B(_0261_));
 sg13g2_inv_1 _1194_ (.Y(_0264_),
    .A(_0263_));
 sg13g2_xnor2_1 _1195_ (.Y(_0265_),
    .A(_0255_),
    .B(_0263_));
 sg13g2_and2_1 _1196_ (.A(_0208_),
    .B(_0265_),
    .X(_0266_));
 sg13g2_nor2_1 _1197_ (.A(\hvsync_gen.hpos[7] ),
    .B(_0258_),
    .Y(_0267_));
 sg13g2_nor2_1 _1198_ (.A(_0260_),
    .B(_0267_),
    .Y(_0268_));
 sg13g2_mux2_1 _1199_ (.A0(_0022_),
    .A1(_0023_),
    .S(_0227_),
    .X(_0269_));
 sg13g2_xor2_1 _1200_ (.B(_0269_),
    .A(_0019_),
    .X(_0270_));
 sg13g2_nand2b_1 _1201_ (.Y(_0271_),
    .B(_0030_),
    .A_N(_0270_));
 sg13g2_xnor2_1 _1202_ (.Y(_0272_),
    .A(_0030_),
    .B(_0270_));
 sg13g2_nor2b_1 _1203_ (.A(_0268_),
    .B_N(_0272_),
    .Y(_0273_));
 sg13g2_xnor2_1 _1204_ (.Y(_0274_),
    .A(_0268_),
    .B(_0272_));
 sg13g2_o21ai_1 _1205_ (.B1(_0262_),
    .Y(_0275_),
    .A1(_0255_),
    .A2(_0264_));
 sg13g2_xor2_1 _1206_ (.B(_0275_),
    .A(_0274_),
    .X(_0276_));
 sg13g2_a21oi_1 _1207_ (.A1(net427),
    .A2(_0276_),
    .Y(_0277_),
    .B1(_0266_));
 sg13g2_a21oi_2 _1208_ (.B1(_0273_),
    .Y(_0278_),
    .A2(_0275_),
    .A1(_0274_));
 sg13g2_o21ai_1 _1209_ (.B1(_0271_),
    .Y(_0279_),
    .A1(net426),
    .A2(_0269_));
 sg13g2_mux2_1 _1210_ (.A0(\counter[8] ),
    .A1(\counter[9] ),
    .S(_0228_),
    .X(_0280_));
 sg13g2_xnor2_1 _1211_ (.Y(_0281_),
    .A(\hvsync_gen.hpos[6] ),
    .B(_0280_));
 sg13g2_xnor2_1 _1212_ (.Y(_0282_),
    .A(_0279_),
    .B(_0281_));
 sg13g2_xnor2_1 _1213_ (.Y(_0283_),
    .A(_0278_),
    .B(_0282_));
 sg13g2_xor2_1 _1214_ (.B(_0282_),
    .A(_0278_),
    .X(_0284_));
 sg13g2_nor2_1 _1215_ (.A(net427),
    .B(_0284_),
    .Y(_0285_));
 sg13g2_nor3_1 _1216_ (.A(_0167_),
    .B(net427),
    .C(_0284_),
    .Y(_0286_));
 sg13g2_nor2_1 _1217_ (.A(net425),
    .B(_0277_),
    .Y(_0287_));
 sg13g2_o21ai_1 _1218_ (.B1(_0217_),
    .Y(_0288_),
    .A1(_0286_),
    .A2(_0287_));
 sg13g2_xor2_1 _1219_ (.B(\div3.out[1] ),
    .A(net427),
    .X(_0289_));
 sg13g2_inv_1 _1220_ (.Y(_0290_),
    .A(_0289_));
 sg13g2_nor3_1 _1221_ (.A(_0217_),
    .B(_0286_),
    .C(_0287_),
    .Y(_0291_));
 sg13g2_or3_1 _1222_ (.A(_0217_),
    .B(_0286_),
    .C(_0287_),
    .X(_0292_));
 sg13g2_nand3_1 _1223_ (.B(_0289_),
    .C(_0292_),
    .A(_0288_),
    .Y(_0293_));
 sg13g2_o21ai_1 _1224_ (.B1(_0288_),
    .Y(_0294_),
    .A1(_0290_),
    .A2(_0291_));
 sg13g2_and2_1 _1225_ (.A(_0208_),
    .B(_0276_),
    .X(_0295_));
 sg13g2_a21oi_1 _1226_ (.A1(net427),
    .A2(_0283_),
    .Y(_0296_),
    .B1(_0295_));
 sg13g2_nor2b_1 _1227_ (.A(net425),
    .B_N(\div3.out[2] ),
    .Y(_0297_));
 sg13g2_nand2b_1 _1228_ (.Y(_0298_),
    .B(_0297_),
    .A_N(_0296_));
 sg13g2_xnor2_1 _1229_ (.Y(_0299_),
    .A(net425),
    .B(\div3.out[2] ));
 sg13g2_o21ai_1 _1230_ (.B1(_0299_),
    .Y(_0300_),
    .A1(net425),
    .A2(_0296_));
 sg13g2_xor2_1 _1231_ (.B(\hvsync_gen.hpos[9] ),
    .A(\div3.out[0] ),
    .X(_0301_));
 sg13g2_nand3_1 _1232_ (.B(_0300_),
    .C(_0301_),
    .A(_0298_),
    .Y(_0302_));
 sg13g2_a21o_1 _1233_ (.A2(_0300_),
    .A1(_0298_),
    .B1(_0301_),
    .X(_0303_));
 sg13g2_nand3_1 _1234_ (.B(_0302_),
    .C(_0303_),
    .A(_0294_),
    .Y(_0304_));
 sg13g2_xor2_1 _1235_ (.B(\div3.out[4] ),
    .A(\hvsync_gen.hpos[6] ),
    .X(_0305_));
 sg13g2_xnor2_1 _1236_ (.Y(_0306_),
    .A(_0253_),
    .B(_0254_));
 sg13g2_inv_1 _1237_ (.Y(_0307_),
    .A(_0306_));
 sg13g2_mux4_1 _1238_ (.S0(\a[1] ),
    .A0(_0265_),
    .A1(_0283_),
    .A2(_0307_),
    .A3(_0276_),
    .S1(_0208_),
    .X(_0308_));
 sg13g2_nand2_1 _1239_ (.Y(_0309_),
    .A(_0305_),
    .B(_0308_));
 sg13g2_xnor2_1 _1240_ (.Y(_0310_),
    .A(_0305_),
    .B(_0308_));
 sg13g2_o21ai_1 _1241_ (.B1(_0309_),
    .Y(_0311_),
    .A1(_0299_),
    .A2(_0310_));
 sg13g2_a21o_1 _1242_ (.A2(_0292_),
    .A1(_0288_),
    .B1(_0289_),
    .X(_0312_));
 sg13g2_nand3_1 _1243_ (.B(_0311_),
    .C(_0312_),
    .A(_0293_),
    .Y(_0313_));
 sg13g2_a21oi_1 _1244_ (.A1(_0302_),
    .A2(_0303_),
    .Y(_0314_),
    .B1(_0294_));
 sg13g2_a21o_1 _1245_ (.A2(_0303_),
    .A1(_0302_),
    .B1(_0294_),
    .X(_0315_));
 sg13g2_o21ai_1 _1246_ (.B1(_0304_),
    .Y(_0316_),
    .A1(_0313_),
    .A2(_0314_));
 sg13g2_and2_1 _1247_ (.A(_0298_),
    .B(_0302_),
    .X(_0317_));
 sg13g2_a21oi_1 _1248_ (.A1(_0019_),
    .A2(_0285_),
    .Y(_0318_),
    .B1(_0289_));
 sg13g2_nand3_1 _1249_ (.B(\div3.out[1] ),
    .C(_0285_),
    .A(_0019_),
    .Y(_0319_));
 sg13g2_nand2b_1 _1250_ (.Y(_0320_),
    .B(_0319_),
    .A_N(_0318_));
 sg13g2_xor2_1 _1251_ (.B(\div3.out[5] ),
    .A(\hvsync_gen.hpos[8] ),
    .X(_0321_));
 sg13g2_nand2b_1 _1252_ (.Y(_0322_),
    .B(_0321_),
    .A_N(_0320_));
 sg13g2_xnor2_1 _1253_ (.Y(_0323_),
    .A(_0320_),
    .B(_0321_));
 sg13g2_nor2b_1 _1254_ (.A(_0317_),
    .B_N(_0323_),
    .Y(_0324_));
 sg13g2_xnor2_1 _1255_ (.Y(_0325_),
    .A(_0317_),
    .B(_0323_));
 sg13g2_xnor2_1 _1256_ (.Y(_0326_),
    .A(_0316_),
    .B(_0325_));
 sg13g2_a21oi_1 _1257_ (.A1(_0304_),
    .A2(_0315_),
    .Y(_0327_),
    .B1(_0313_));
 sg13g2_nand3_1 _1258_ (.B(_0313_),
    .C(_0315_),
    .A(_0304_),
    .Y(_0328_));
 sg13g2_nor2b_2 _1259_ (.A(_0327_),
    .B_N(_0328_),
    .Y(_0329_));
 sg13g2_and2_1 _1260_ (.A(_0326_),
    .B(_0329_),
    .X(_0330_));
 sg13g2_xor2_1 _1261_ (.B(_0329_),
    .A(_0326_),
    .X(_0331_));
 sg13g2_a21o_1 _1262_ (.A2(_0312_),
    .A1(_0293_),
    .B1(_0311_),
    .X(_0332_));
 sg13g2_nand2_1 _1263_ (.Y(_0333_),
    .A(_0313_),
    .B(_0332_));
 sg13g2_xor2_1 _1264_ (.B(_0310_),
    .A(_0299_),
    .X(_0334_));
 sg13g2_a21oi_1 _1265_ (.A1(_0313_),
    .A2(_0332_),
    .Y(_0335_),
    .B1(_0334_));
 sg13g2_a21o_1 _1266_ (.A2(_0332_),
    .A1(_0313_),
    .B1(_0334_),
    .X(_0336_));
 sg13g2_nand3b_1 _1267_ (.B(_0328_),
    .C(_0333_),
    .Y(_0337_),
    .A_N(_0327_));
 sg13g2_nand2_1 _1268_ (.Y(_0338_),
    .A(_0336_),
    .B(_0337_));
 sg13g2_xor2_1 _1269_ (.B(_0338_),
    .A(_0331_),
    .X(_0339_));
 sg13g2_and2_1 _1270_ (.A(_0215_),
    .B(_0339_),
    .X(_0340_));
 sg13g2_nand4_1 _1271_ (.B(_0313_),
    .C(_0315_),
    .A(_0304_),
    .Y(_0341_),
    .D(_0332_));
 sg13g2_and3_1 _1272_ (.X(_0342_),
    .A(_0336_),
    .B(_0337_),
    .C(_0341_));
 sg13g2_nand3_1 _1273_ (.B(_0337_),
    .C(_0341_),
    .A(_0336_),
    .Y(_0343_));
 sg13g2_and2_1 _1274_ (.A(_0329_),
    .B(_0335_),
    .X(_0344_));
 sg13g2_nand2_1 _1275_ (.Y(_0345_),
    .A(_0329_),
    .B(_0335_));
 sg13g2_a21oi_2 _1276_ (.B1(_0216_),
    .Y(_0346_),
    .A2(_0345_),
    .A1(_0343_));
 sg13g2_o21ai_1 _1277_ (.B1(_0215_),
    .Y(_0347_),
    .A1(_0342_),
    .A2(_0344_));
 sg13g2_xnor2_1 _1278_ (.Y(_0348_),
    .A(_0333_),
    .B(_0334_));
 sg13g2_xnor2_1 _1279_ (.Y(_0349_),
    .A(_0211_),
    .B(_0214_));
 sg13g2_nor2b_1 _1280_ (.A(_0349_),
    .B_N(_0348_),
    .Y(_0350_));
 sg13g2_nor2_2 _1281_ (.A(_0213_),
    .B(_0334_),
    .Y(_0351_));
 sg13g2_xnor2_1 _1282_ (.Y(_0352_),
    .A(_0348_),
    .B(_0349_));
 sg13g2_a21oi_2 _1283_ (.B1(_0350_),
    .Y(_0353_),
    .A2(_0352_),
    .A1(_0351_));
 sg13g2_nor3_2 _1284_ (.A(_0215_),
    .B(_0342_),
    .C(_0344_),
    .Y(_0354_));
 sg13g2_nand3_1 _1285_ (.B(_0343_),
    .C(_0345_),
    .A(_0216_),
    .Y(_0355_));
 sg13g2_nor3_2 _1286_ (.A(_0346_),
    .B(_0353_),
    .C(_0354_),
    .Y(_0356_));
 sg13g2_or3_1 _1287_ (.A(_0346_),
    .B(_0353_),
    .C(_0354_),
    .X(_0357_));
 sg13g2_o21ai_1 _1288_ (.B1(_0347_),
    .Y(_0358_),
    .A1(_0353_),
    .A2(_0354_));
 sg13g2_xnor2_1 _1289_ (.Y(_0359_),
    .A(_0216_),
    .B(_0339_));
 sg13g2_a21oi_1 _1290_ (.A1(_0358_),
    .A2(_0359_),
    .Y(_0360_),
    .B1(_0340_));
 sg13g2_a21oi_1 _1291_ (.A1(_0331_),
    .A2(_0338_),
    .Y(_0361_),
    .B1(_0330_));
 sg13g2_a21oi_2 _1292_ (.B1(_0324_),
    .Y(_0362_),
    .A2(_0325_),
    .A1(_0316_));
 sg13g2_xnor2_1 _1293_ (.Y(_0363_),
    .A(\div3.out[0] ),
    .B(net424));
 sg13g2_and3_1 _1294_ (.X(_0364_),
    .A(_0319_),
    .B(_0322_),
    .C(_0363_));
 sg13g2_a21oi_2 _1295_ (.B1(_0363_),
    .Y(_0365_),
    .A2(_0322_),
    .A1(_0319_));
 sg13g2_a21oi_1 _1296_ (.A1(_0362_),
    .A2(_0364_),
    .Y(_0366_),
    .B1(_0365_));
 sg13g2_a21o_1 _1297_ (.A2(_0364_),
    .A1(_0362_),
    .B1(_0365_),
    .X(_0367_));
 sg13g2_or3_1 _1298_ (.A(_0362_),
    .B(_0364_),
    .C(_0365_),
    .X(_0368_));
 sg13g2_and3_1 _1299_ (.X(_0369_),
    .A(_0326_),
    .B(_0366_),
    .C(_0368_));
 sg13g2_nand3_1 _1300_ (.B(_0366_),
    .C(_0368_),
    .A(_0326_),
    .Y(_0370_));
 sg13g2_a21oi_1 _1301_ (.A1(_0366_),
    .A2(_0368_),
    .Y(_0371_),
    .B1(_0326_));
 sg13g2_or3_1 _1302_ (.A(_0361_),
    .B(_0369_),
    .C(_0371_),
    .X(_0372_));
 sg13g2_o21ai_1 _1303_ (.B1(_0361_),
    .Y(_0373_),
    .A1(_0369_),
    .A2(_0371_));
 sg13g2_and3_1 _1304_ (.X(_0374_),
    .A(_0215_),
    .B(_0372_),
    .C(_0373_));
 sg13g2_nand3_1 _1305_ (.B(_0372_),
    .C(_0373_),
    .A(_0215_),
    .Y(_0375_));
 sg13g2_a21oi_1 _1306_ (.A1(_0372_),
    .A2(_0373_),
    .Y(_0376_),
    .B1(_0215_));
 sg13g2_or3_1 _1307_ (.A(_0360_),
    .B(_0374_),
    .C(_0376_),
    .X(_0377_));
 sg13g2_o21ai_1 _1308_ (.B1(_0360_),
    .Y(_0378_),
    .A1(_0374_),
    .A2(_0376_));
 sg13g2_and2_1 _1309_ (.A(_0377_),
    .B(_0378_),
    .X(_0379_));
 sg13g2_nand2_2 _1310_ (.Y(_0380_),
    .A(_0377_),
    .B(_0378_));
 sg13g2_xor2_1 _1311_ (.B(_0352_),
    .A(_0351_),
    .X(_0381_));
 sg13g2_xnor2_1 _1312_ (.Y(_0382_),
    .A(_0351_),
    .B(_0352_));
 sg13g2_and2_2 _1313_ (.A(net422),
    .B(net419),
    .X(_0383_));
 sg13g2_nand2_1 _1314_ (.Y(_0384_),
    .A(net422),
    .B(net419));
 sg13g2_nor2_2 _1315_ (.A(net384),
    .B(_0383_),
    .Y(_0385_));
 sg13g2_xnor2_1 _1316_ (.Y(_0386_),
    .A(_0212_),
    .B(_0334_));
 sg13g2_xnor2_1 _1317_ (.Y(_0387_),
    .A(_0213_),
    .B(_0334_));
 sg13g2_nand2b_1 _1318_ (.Y(_0388_),
    .B(net403),
    .A_N(net421));
 sg13g2_nor2_2 _1319_ (.A(net421),
    .B(net420),
    .Y(_0389_));
 sg13g2_or2_2 _1320_ (.X(_0390_),
    .B(net419),
    .A(net422));
 sg13g2_nor2_2 _1321_ (.A(net407),
    .B(_0390_),
    .Y(_0391_));
 sg13g2_nand2_2 _1322_ (.Y(_0392_),
    .A(net405),
    .B(_0389_));
 sg13g2_nand2_2 _1323_ (.Y(_0393_),
    .A(_0385_),
    .B(_0392_));
 sg13g2_a221oi_1 _1324_ (.B2(_0347_),
    .C1(_0350_),
    .B1(_0355_),
    .A1(_0351_),
    .Y(_0394_),
    .A2(_0352_));
 sg13g2_o21ai_1 _1325_ (.B1(_0353_),
    .Y(_0395_),
    .A1(_0346_),
    .A2(_0354_));
 sg13g2_nor2_1 _1326_ (.A(_0356_),
    .B(_0394_),
    .Y(_0396_));
 sg13g2_nand2_1 _1327_ (.Y(_0397_),
    .A(net383),
    .B(net381));
 sg13g2_nor2_2 _1328_ (.A(\hvsync_gen.vpos[1] ),
    .B(net406),
    .Y(_0398_));
 sg13g2_nand2b_2 _1329_ (.Y(_0399_),
    .B(net407),
    .A_N(net419));
 sg13g2_nor2_2 _1330_ (.A(_0352_),
    .B(_0399_),
    .Y(_0400_));
 sg13g2_nand2_2 _1331_ (.Y(_0401_),
    .A(net388),
    .B(_0398_));
 sg13g2_nor2b_2 _1332_ (.A(net421),
    .B_N(net418),
    .Y(_0402_));
 sg13g2_nand2b_2 _1333_ (.Y(_0403_),
    .B(net418),
    .A_N(net421));
 sg13g2_nor2b_2 _1334_ (.A(net418),
    .B_N(net421),
    .Y(_0404_));
 sg13g2_nand2b_2 _1335_ (.Y(_0405_),
    .B(net421),
    .A_N(net418));
 sg13g2_nand2_1 _1336_ (.Y(_0406_),
    .A(net384),
    .B(_0405_));
 sg13g2_nor2_2 _1337_ (.A(_0402_),
    .B(_0404_),
    .Y(_0407_));
 sg13g2_nand2_2 _1338_ (.Y(_0408_),
    .A(_0403_),
    .B(_0405_));
 sg13g2_nor2_1 _1339_ (.A(net409),
    .B(_0408_),
    .Y(_0409_));
 sg13g2_nand2_2 _1340_ (.Y(_0410_),
    .A(net405),
    .B(_0407_));
 sg13g2_o21ai_1 _1341_ (.B1(net390),
    .Y(_0411_),
    .A1(_0398_),
    .A2(_0409_));
 sg13g2_and2_1 _1342_ (.A(net362),
    .B(_0411_),
    .X(_0412_));
 sg13g2_xor2_1 _1343_ (.B(_0359_),
    .A(_0358_),
    .X(_0413_));
 sg13g2_xnor2_1 _1344_ (.Y(_0414_),
    .A(_0358_),
    .B(_0359_));
 sg13g2_and2_1 _1345_ (.A(net420),
    .B(net408),
    .X(_0415_));
 sg13g2_nand2_2 _1346_ (.Y(_0416_),
    .A(net418),
    .B(net407));
 sg13g2_nand2_2 _1347_ (.Y(_0417_),
    .A(_0383_),
    .B(net408));
 sg13g2_nor2_2 _1348_ (.A(net420),
    .B(net409),
    .Y(_0418_));
 sg13g2_nand2b_2 _1349_ (.Y(_0419_),
    .B(net403),
    .A_N(net418));
 sg13g2_nand2_2 _1350_ (.Y(_0420_),
    .A(net404),
    .B(_0404_));
 sg13g2_and2_2 _1351_ (.A(net418),
    .B(net403),
    .X(_0421_));
 sg13g2_nand2_2 _1352_ (.Y(_0422_),
    .A(net418),
    .B(net403));
 sg13g2_nor2_2 _1353_ (.A(_0398_),
    .B(_0421_),
    .Y(_0423_));
 sg13g2_nand2_2 _1354_ (.Y(_0424_),
    .A(_0399_),
    .B(net402));
 sg13g2_nand2_1 _1355_ (.Y(_0425_),
    .A(net422),
    .B(_0423_));
 sg13g2_nand2_1 _1356_ (.Y(_0426_),
    .A(net387),
    .B(_0425_));
 sg13g2_nand2_2 _1357_ (.Y(_0427_),
    .A(net398),
    .B(net406));
 sg13g2_nand2_2 _1358_ (.Y(_0428_),
    .A(net395),
    .B(_0417_));
 sg13g2_and2_1 _1359_ (.A(net395),
    .B(_0417_),
    .X(_0429_));
 sg13g2_nand2_2 _1360_ (.Y(_0430_),
    .A(_0392_),
    .B(net379));
 sg13g2_and2_1 _1361_ (.A(net371),
    .B(_0430_),
    .X(_0431_));
 sg13g2_a221oi_1 _1362_ (.B2(_0431_),
    .C1(net345),
    .B1(_0426_),
    .A1(_0393_),
    .Y(_0432_),
    .A2(_0412_));
 sg13g2_nor2_1 _1363_ (.A(net373),
    .B(net357),
    .Y(_0433_));
 sg13g2_nand2_2 _1364_ (.Y(_0434_),
    .A(net365),
    .B(net349));
 sg13g2_nor2_1 _1365_ (.A(net420),
    .B(net401),
    .Y(_0435_));
 sg13g2_inv_1 _1366_ (.Y(_0436_),
    .A(_0435_));
 sg13g2_o21ai_1 _1367_ (.B1(net386),
    .Y(_0437_),
    .A1(_0389_),
    .A2(_0398_));
 sg13g2_nand2_1 _1368_ (.Y(_0438_),
    .A(_0430_),
    .B(_0437_));
 sg13g2_nor2_2 _1369_ (.A(net409),
    .B(_0389_),
    .Y(_0439_));
 sg13g2_nand2_2 _1370_ (.Y(_0440_),
    .A(net404),
    .B(_0390_));
 sg13g2_nor2_1 _1371_ (.A(net397),
    .B(_0439_),
    .Y(_0441_));
 sg13g2_and2_1 _1372_ (.A(net419),
    .B(net396),
    .X(_0442_));
 sg13g2_nor2_1 _1373_ (.A(net367),
    .B(_0442_),
    .Y(_0443_));
 sg13g2_nor4_1 _1374_ (.A(net367),
    .B(net355),
    .C(_0441_),
    .D(_0442_),
    .Y(_0444_));
 sg13g2_a21o_1 _1375_ (.A2(_0438_),
    .A1(net342),
    .B1(_0444_),
    .X(_0445_));
 sg13g2_o21ai_1 _1376_ (.B1(net331),
    .Y(_0446_),
    .A1(_0432_),
    .A2(_0445_));
 sg13g2_o21ai_1 _1377_ (.B1(_0375_),
    .Y(_0447_),
    .A1(_0360_),
    .A2(_0376_));
 sg13g2_nand2_1 _1378_ (.Y(_0448_),
    .A(_0362_),
    .B(_0365_));
 sg13g2_and2_1 _1379_ (.A(_0368_),
    .B(_0448_),
    .X(_0449_));
 sg13g2_o21ai_1 _1380_ (.B1(_0370_),
    .Y(_0450_),
    .A1(_0361_),
    .A2(_0371_));
 sg13g2_xor2_1 _1381_ (.B(_0450_),
    .A(_0449_),
    .X(_0451_));
 sg13g2_and2_1 _1382_ (.A(_0215_),
    .B(_0451_),
    .X(_0452_));
 sg13g2_xnor2_1 _1383_ (.Y(_0453_),
    .A(_0216_),
    .B(_0451_));
 sg13g2_xor2_1 _1384_ (.B(_0453_),
    .A(_0447_),
    .X(_0454_));
 sg13g2_xnor2_1 _1385_ (.Y(_0455_),
    .A(_0447_),
    .B(_0453_));
 sg13g2_nor2_1 _1386_ (.A(net365),
    .B(net359),
    .Y(_0456_));
 sg13g2_nand2_2 _1387_ (.Y(_0457_),
    .A(net393),
    .B(_0421_));
 sg13g2_nor2_2 _1388_ (.A(net415),
    .B(net407),
    .Y(_0458_));
 sg13g2_nand2_2 _1389_ (.Y(_0459_),
    .A(_0383_),
    .B(net403));
 sg13g2_nand2_1 _1390_ (.Y(_0460_),
    .A(net393),
    .B(_0458_));
 sg13g2_o21ai_1 _1391_ (.B1(_0460_),
    .Y(_0461_),
    .A1(_0406_),
    .A2(_0421_));
 sg13g2_nand3_1 _1392_ (.B(net347),
    .C(_0461_),
    .A(net369),
    .Y(_0462_));
 sg13g2_nand2_1 _1393_ (.Y(_0463_),
    .A(net386),
    .B(_0403_));
 sg13g2_nand3_1 _1394_ (.B(_0403_),
    .C(_0424_),
    .A(net387),
    .Y(_0464_));
 sg13g2_a21oi_1 _1395_ (.A1(_0428_),
    .A2(_0464_),
    .Y(_0465_),
    .B1(_0434_));
 sg13g2_nor2_2 _1396_ (.A(net396),
    .B(net408),
    .Y(_0466_));
 sg13g2_nand2_2 _1397_ (.Y(_0467_),
    .A(net389),
    .B(net406));
 sg13g2_nor2_2 _1398_ (.A(net395),
    .B(_0389_),
    .Y(_0468_));
 sg13g2_nor2_2 _1399_ (.A(net405),
    .B(_0390_),
    .Y(_0469_));
 sg13g2_nand2_2 _1400_ (.Y(_0470_),
    .A(net407),
    .B(_0389_));
 sg13g2_nor2_2 _1401_ (.A(net401),
    .B(_0469_),
    .Y(_0471_));
 sg13g2_nand2_2 _1402_ (.Y(_0472_),
    .A(net407),
    .B(_0390_));
 sg13g2_nor2_1 _1403_ (.A(_0439_),
    .B(_0469_),
    .Y(_0473_));
 sg13g2_and2_1 _1404_ (.A(net391),
    .B(_0473_),
    .X(_0474_));
 sg13g2_and2_2 _1405_ (.A(_0352_),
    .B(net409),
    .X(_0475_));
 sg13g2_nand2_2 _1406_ (.Y(_0476_),
    .A(_0352_),
    .B(net409));
 sg13g2_nor2_2 _1407_ (.A(net389),
    .B(_0399_),
    .Y(_0477_));
 sg13g2_nand2_2 _1408_ (.Y(_0478_),
    .A(net397),
    .B(_0398_));
 sg13g2_nor3_1 _1409_ (.A(net377),
    .B(_0474_),
    .C(_0477_),
    .Y(_0479_));
 sg13g2_nor2_2 _1410_ (.A(net397),
    .B(_0418_),
    .Y(_0480_));
 sg13g2_nand4_1 _1411_ (.B(_0388_),
    .C(_0419_),
    .A(net384),
    .Y(_0481_),
    .D(_0472_));
 sg13g2_nor2_2 _1412_ (.A(net405),
    .B(_0405_),
    .Y(_0482_));
 sg13g2_nand2_1 _1413_ (.Y(_0483_),
    .A(net407),
    .B(_0404_));
 sg13g2_nand3_1 _1414_ (.B(_0403_),
    .C(_0483_),
    .A(net394),
    .Y(_0484_));
 sg13g2_nand4_1 _1415_ (.B(net380),
    .C(_0481_),
    .A(net382),
    .Y(_0485_),
    .D(_0484_));
 sg13g2_nand2_1 _1416_ (.Y(_0486_),
    .A(net356),
    .B(_0485_));
 sg13g2_o21ai_1 _1417_ (.B1(_0462_),
    .Y(_0487_),
    .A1(_0479_),
    .A2(_0486_));
 sg13g2_o21ai_1 _1418_ (.B1(net334),
    .Y(_0488_),
    .A1(_0465_),
    .A2(_0487_));
 sg13g2_and3_1 _1419_ (.X(_0489_),
    .A(_0446_),
    .B(net329),
    .C(_0488_));
 sg13g2_a21oi_2 _1420_ (.B1(_0452_),
    .Y(_0490_),
    .A2(_0453_),
    .A1(_0447_));
 sg13g2_nand2_1 _1421_ (.Y(_0491_),
    .A(_0367_),
    .B(_0449_));
 sg13g2_nor2_1 _1422_ (.A(_0372_),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_o21ai_1 _1423_ (.B1(_0449_),
    .Y(_0493_),
    .A1(_0367_),
    .A2(_0450_));
 sg13g2_or2_1 _1424_ (.X(_0494_),
    .B(_0493_),
    .A(_0492_));
 sg13g2_xnor2_1 _1425_ (.Y(_0495_),
    .A(_0216_),
    .B(_0494_));
 sg13g2_nor2_1 _1426_ (.A(_0490_),
    .B(_0495_),
    .Y(_0496_));
 sg13g2_xor2_1 _1427_ (.B(_0495_),
    .A(_0490_),
    .X(_0497_));
 sg13g2_xnor2_1 _1428_ (.Y(_0498_),
    .A(_0490_),
    .B(_0495_));
 sg13g2_nor2_2 _1429_ (.A(net364),
    .B(net352),
    .Y(_0499_));
 sg13g2_nand2_2 _1430_ (.Y(_0500_),
    .A(net369),
    .B(net356));
 sg13g2_nor2_1 _1431_ (.A(net407),
    .B(_0403_),
    .Y(_0501_));
 sg13g2_nand2_2 _1432_ (.Y(_0502_),
    .A(net403),
    .B(_0402_));
 sg13g2_nand2_2 _1433_ (.Y(_0503_),
    .A(_0399_),
    .B(_0502_));
 sg13g2_nor2_2 _1434_ (.A(net390),
    .B(_0398_),
    .Y(_0504_));
 sg13g2_nor2_1 _1435_ (.A(net400),
    .B(_0383_),
    .Y(_0505_));
 sg13g2_nand2_2 _1436_ (.Y(_0506_),
    .A(net384),
    .B(net415));
 sg13g2_nor2_1 _1437_ (.A(_0415_),
    .B(_0506_),
    .Y(_0507_));
 sg13g2_a21oi_1 _1438_ (.A1(_0502_),
    .A2(net378),
    .Y(_0508_),
    .B1(_0507_));
 sg13g2_nor2_2 _1439_ (.A(net399),
    .B(_0459_),
    .Y(_0509_));
 sg13g2_nand2_1 _1440_ (.Y(_0510_),
    .A(net386),
    .B(_0458_));
 sg13g2_nor2_1 _1441_ (.A(net420),
    .B(net391),
    .Y(_0511_));
 sg13g2_nand2b_1 _1442_ (.Y(_0512_),
    .B(net400),
    .A_N(net420));
 sg13g2_nand2_1 _1443_ (.Y(_0513_),
    .A(net396),
    .B(_0389_));
 sg13g2_nor2_2 _1444_ (.A(net389),
    .B(_0416_),
    .Y(_0514_));
 sg13g2_nor2_1 _1445_ (.A(net385),
    .B(_0421_),
    .Y(_0515_));
 sg13g2_nand2_1 _1446_ (.Y(_0516_),
    .A(net398),
    .B(_0422_));
 sg13g2_nand3_1 _1447_ (.B(_0407_),
    .C(net402),
    .A(net393),
    .Y(_0517_));
 sg13g2_o21ai_1 _1448_ (.B1(net356),
    .Y(_0518_),
    .A1(net369),
    .A2(_0509_));
 sg13g2_o21ai_1 _1449_ (.B1(_0518_),
    .Y(_0519_),
    .A1(net361),
    .A2(_0517_));
 sg13g2_o21ai_1 _1450_ (.B1(_0519_),
    .Y(_0520_),
    .A1(_0500_),
    .A2(_0508_));
 sg13g2_nand2_2 _1451_ (.Y(_0521_),
    .A(net402),
    .B(net379));
 sg13g2_a22oi_1 _1452_ (.Y(_0522_),
    .B1(net379),
    .B2(net402),
    .A2(_0424_),
    .A1(net385));
 sg13g2_nor2_1 _1453_ (.A(net399),
    .B(_0482_),
    .Y(_0523_));
 sg13g2_nand2_2 _1454_ (.Y(_0524_),
    .A(net388),
    .B(_0459_));
 sg13g2_nand3_1 _1455_ (.B(_0459_),
    .C(_0483_),
    .A(net385),
    .Y(_0525_));
 sg13g2_nand2_1 _1456_ (.Y(_0526_),
    .A(_0476_),
    .B(_0525_));
 sg13g2_a21oi_1 _1457_ (.A1(net370),
    .A2(_0526_),
    .Y(_0527_),
    .B1(net346));
 sg13g2_o21ai_1 _1458_ (.B1(_0527_),
    .Y(_0528_),
    .A1(net370),
    .A2(_0522_));
 sg13g2_nand2_1 _1459_ (.Y(_0529_),
    .A(net404),
    .B(_0408_));
 sg13g2_and2_1 _1460_ (.A(net395),
    .B(_0529_),
    .X(_0530_));
 sg13g2_nor2_2 _1461_ (.A(net403),
    .B(_0403_),
    .Y(_0531_));
 sg13g2_nor2_1 _1462_ (.A(_0525_),
    .B(_0531_),
    .Y(_0532_));
 sg13g2_nor3_1 _1463_ (.A(net368),
    .B(_0530_),
    .C(_0532_),
    .Y(_0533_));
 sg13g2_nor4_2 _1464_ (.A(net386),
    .B(_0458_),
    .C(_0482_),
    .Y(_0534_),
    .D(_0531_));
 sg13g2_nor2_1 _1465_ (.A(_0383_),
    .B(net406),
    .Y(_0535_));
 sg13g2_nand2_2 _1466_ (.Y(_0536_),
    .A(net416),
    .B(net408));
 sg13g2_nor2_2 _1467_ (.A(net400),
    .B(_0535_),
    .Y(_0537_));
 sg13g2_nand2_1 _1468_ (.Y(_0538_),
    .A(net384),
    .B(_0536_));
 sg13g2_nor3_2 _1469_ (.A(_0356_),
    .B(_0394_),
    .C(_0537_),
    .Y(_0539_));
 sg13g2_nand2b_1 _1470_ (.Y(_0540_),
    .B(_0539_),
    .A_N(_0534_));
 sg13g2_nand2b_1 _1471_ (.Y(_0541_),
    .B(_0540_),
    .A_N(_0533_));
 sg13g2_a21oi_1 _1472_ (.A1(net345),
    .A2(_0541_),
    .Y(_0542_),
    .B1(net331));
 sg13g2_a221oi_1 _1473_ (.B2(_0542_),
    .C1(net329),
    .B1(_0528_),
    .A1(net331),
    .Y(_0543_),
    .A2(_0520_));
 sg13g2_nor3_1 _1474_ (.A(_0489_),
    .B(_0497_),
    .C(_0543_),
    .Y(_0544_));
 sg13g2_xnor2_1 _1475_ (.Y(_0545_),
    .A(_0216_),
    .B(_0492_));
 sg13g2_inv_1 _1476_ (.Y(_0546_),
    .A(_0545_));
 sg13g2_and2_1 _1477_ (.A(_0494_),
    .B(_0545_),
    .X(_0547_));
 sg13g2_inv_1 _1478_ (.Y(_0548_),
    .A(_0547_));
 sg13g2_mux2_2 _1479_ (.A0(_0548_),
    .A1(_0545_),
    .S(_0496_),
    .X(_0549_));
 sg13g2_mux2_1 _1480_ (.A0(_0547_),
    .A1(_0546_),
    .S(_0496_),
    .X(_0550_));
 sg13g2_and3_1 _1481_ (.X(_0551_),
    .A(net342),
    .B(_0457_),
    .C(_0463_));
 sg13g2_and3_1 _1482_ (.X(_0552_),
    .A(net382),
    .B(net380),
    .C(_0517_));
 sg13g2_nand2_1 _1483_ (.Y(_0553_),
    .A(net388),
    .B(_0422_));
 sg13g2_nand2_2 _1484_ (.Y(_0554_),
    .A(net402),
    .B(_0537_));
 sg13g2_nand2_1 _1485_ (.Y(_0555_),
    .A(net393),
    .B(_0420_));
 sg13g2_nand3_1 _1486_ (.B(_0416_),
    .C(_0420_),
    .A(net393),
    .Y(_0556_));
 sg13g2_nor2_2 _1487_ (.A(net394),
    .B(_0391_),
    .Y(_0557_));
 sg13g2_o21ai_1 _1488_ (.B1(_0556_),
    .Y(_0558_),
    .A1(_0391_),
    .A2(_0506_));
 sg13g2_a221oi_1 _1489_ (.B2(net361),
    .C1(net347),
    .B1(_0558_),
    .A1(_0552_),
    .Y(_0559_),
    .A2(_0554_));
 sg13g2_nand2_1 _1490_ (.Y(_0560_),
    .A(net394),
    .B(_0472_));
 sg13g2_and3_1 _1491_ (.X(_0561_),
    .A(_0437_),
    .B(net341),
    .C(_0560_));
 sg13g2_nor4_1 _1492_ (.A(net331),
    .B(_0551_),
    .C(_0559_),
    .D(_0561_),
    .Y(_0562_));
 sg13g2_nand2_1 _1493_ (.Y(_0563_),
    .A(net400),
    .B(_0440_));
 sg13g2_nor2_1 _1494_ (.A(net405),
    .B(_0404_),
    .Y(_0564_));
 sg13g2_nor3_1 _1495_ (.A(net388),
    .B(_0439_),
    .C(_0564_),
    .Y(_0565_));
 sg13g2_a21oi_2 _1496_ (.B1(_0565_),
    .Y(_0566_),
    .A2(net380),
    .A1(net382));
 sg13g2_nor2_2 _1497_ (.A(_0352_),
    .B(net406),
    .Y(_0567_));
 sg13g2_nand2_1 _1498_ (.Y(_0568_),
    .A(_0390_),
    .B(_0567_));
 sg13g2_nor2_2 _1499_ (.A(net384),
    .B(_0419_),
    .Y(_0569_));
 sg13g2_nor2_2 _1500_ (.A(net386),
    .B(_0420_),
    .Y(_0570_));
 sg13g2_nand2_1 _1501_ (.Y(_0571_),
    .A(net421),
    .B(_0569_));
 sg13g2_nor3_1 _1502_ (.A(net361),
    .B(_0509_),
    .C(_0531_),
    .Y(_0572_));
 sg13g2_a221oi_1 _1503_ (.B2(_0572_),
    .C1(net347),
    .B1(_0571_),
    .A1(_0566_),
    .Y(_0573_),
    .A2(_0568_));
 sg13g2_nand2_1 _1504_ (.Y(_0574_),
    .A(net398),
    .B(_0423_));
 sg13g2_and4_2 _1505_ (.A(net382),
    .B(net380),
    .C(_0463_),
    .D(_0467_),
    .X(_0575_));
 sg13g2_and3_1 _1506_ (.X(_0576_),
    .A(net349),
    .B(_0574_),
    .C(_0575_));
 sg13g2_nand2_1 _1507_ (.Y(_0577_),
    .A(_0385_),
    .B(_0416_));
 sg13g2_nand2_1 _1508_ (.Y(_0578_),
    .A(_0417_),
    .B(_0468_));
 sg13g2_and3_1 _1509_ (.X(_0579_),
    .A(net342),
    .B(_0577_),
    .C(_0578_));
 sg13g2_nor4_1 _1510_ (.A(net334),
    .B(_0573_),
    .C(_0576_),
    .D(_0579_),
    .Y(_0580_));
 sg13g2_nor3_1 _1511_ (.A(net328),
    .B(_0562_),
    .C(_0580_),
    .Y(_0581_));
 sg13g2_nand2_1 _1512_ (.Y(_0582_),
    .A(net415),
    .B(_0466_));
 sg13g2_nor2_2 _1513_ (.A(net390),
    .B(_0536_),
    .Y(_0583_));
 sg13g2_nor2_1 _1514_ (.A(net365),
    .B(_0583_),
    .Y(_0584_));
 sg13g2_nor3_1 _1515_ (.A(net362),
    .B(net355),
    .C(_0583_),
    .Y(_0585_));
 sg13g2_nand2_1 _1516_ (.Y(_0586_),
    .A(net343),
    .B(_0574_));
 sg13g2_a22oi_1 _1517_ (.Y(_0587_),
    .B1(_0557_),
    .B2(_0417_),
    .A2(_0423_),
    .A1(net395));
 sg13g2_a22oi_1 _1518_ (.Y(_0588_),
    .B1(_0587_),
    .B2(net342),
    .A2(_0585_),
    .A1(_0582_));
 sg13g2_nor2_1 _1519_ (.A(_0400_),
    .B(net351),
    .Y(_0589_));
 sg13g2_nor2_1 _1520_ (.A(net373),
    .B(_0504_),
    .Y(_0590_));
 sg13g2_nand2b_1 _1521_ (.Y(_0591_),
    .B(net364),
    .A_N(net378));
 sg13g2_a22oi_1 _1522_ (.Y(_0592_),
    .B1(_0405_),
    .B2(net378),
    .A2(net381),
    .A1(net383));
 sg13g2_nand2_2 _1523_ (.Y(_0593_),
    .A(_0459_),
    .B(net378));
 sg13g2_and3_1 _1524_ (.X(_0594_),
    .A(net376),
    .B(_0436_),
    .C(_0593_));
 sg13g2_a22oi_1 _1525_ (.Y(_0595_),
    .B1(_0594_),
    .B2(net358),
    .A2(_0592_),
    .A1(_0589_));
 sg13g2_nand3_1 _1526_ (.B(_0588_),
    .C(_0595_),
    .A(net331),
    .Y(_0596_));
 sg13g2_nand2_1 _1527_ (.Y(_0597_),
    .A(net415),
    .B(_0388_));
 sg13g2_a22oi_1 _1528_ (.Y(_0598_),
    .B1(_0597_),
    .B2(net395),
    .A2(_0557_),
    .A1(_0472_));
 sg13g2_a21oi_2 _1529_ (.B1(net400),
    .Y(_0599_),
    .A2(net381),
    .A1(net383));
 sg13g2_a21o_1 _1530_ (.A2(_0598_),
    .A1(net370),
    .B1(_0599_),
    .X(_0600_));
 sg13g2_nor2_1 _1531_ (.A(net384),
    .B(_0470_),
    .Y(_0601_));
 sg13g2_nand2_1 _1532_ (.Y(_0602_),
    .A(net399),
    .B(_0469_));
 sg13g2_a21oi_2 _1533_ (.B1(_0601_),
    .Y(_0603_),
    .A2(net380),
    .A1(net382));
 sg13g2_nand3_1 _1534_ (.B(net404),
    .C(_0405_),
    .A(net387),
    .Y(_0604_));
 sg13g2_a21oi_1 _1535_ (.A1(_0385_),
    .A2(_0416_),
    .Y(_0605_),
    .B1(_0468_));
 sg13g2_a22oi_1 _1536_ (.Y(_0606_),
    .B1(_0605_),
    .B2(net370),
    .A2(_0604_),
    .A1(_0603_));
 sg13g2_mux2_1 _1537_ (.A0(_0600_),
    .A1(_0606_),
    .S(net346),
    .X(_0607_));
 sg13g2_a21oi_1 _1538_ (.A1(net335),
    .A2(_0607_),
    .Y(_0608_),
    .B1(net329));
 sg13g2_a21o_1 _1539_ (.A2(_0608_),
    .A1(_0596_),
    .B1(net326),
    .X(_0609_));
 sg13g2_o21ai_1 _1540_ (.B1(_0549_),
    .Y(_0610_),
    .A1(_0581_),
    .A2(_0609_));
 sg13g2_a22oi_1 _1541_ (.Y(_0611_),
    .B1(_0440_),
    .B2(_0537_),
    .A2(_0395_),
    .A1(_0357_));
 sg13g2_nand2_2 _1542_ (.Y(_0612_),
    .A(net394),
    .B(_0470_));
 sg13g2_and2_2 _1543_ (.A(net374),
    .B(_0612_),
    .X(_0613_));
 sg13g2_nor3_1 _1544_ (.A(_0439_),
    .B(_0611_),
    .C(_0613_),
    .Y(_0614_));
 sg13g2_nand2_1 _1545_ (.Y(_0615_),
    .A(net399),
    .B(_0536_));
 sg13g2_nor2_2 _1546_ (.A(net405),
    .B(_0407_),
    .Y(_0616_));
 sg13g2_nor2_1 _1547_ (.A(net391),
    .B(_0616_),
    .Y(_0617_));
 sg13g2_nor3_2 _1548_ (.A(net387),
    .B(_0418_),
    .C(_0616_),
    .Y(_0618_));
 sg13g2_nand2_2 _1549_ (.Y(_0619_),
    .A(net390),
    .B(_0469_));
 sg13g2_a21oi_1 _1550_ (.A1(net415),
    .A2(_0466_),
    .Y(_0620_),
    .B1(_0618_));
 sg13g2_nand3_1 _1551_ (.B(_0619_),
    .C(_0620_),
    .A(net342),
    .Y(_0621_));
 sg13g2_nand3_1 _1552_ (.B(_0478_),
    .C(_0513_),
    .A(net341),
    .Y(_0622_));
 sg13g2_nand2_1 _1553_ (.Y(_0623_),
    .A(_0621_),
    .B(_0622_));
 sg13g2_a21o_1 _1554_ (.A2(_0614_),
    .A1(net355),
    .B1(_0623_),
    .X(_0624_));
 sg13g2_a21oi_1 _1555_ (.A1(net325),
    .A2(_0624_),
    .Y(_0625_),
    .B1(\g_x[0] ));
 sg13g2_o21ai_1 _1556_ (.B1(_0625_),
    .Y(_0626_),
    .A1(_0544_),
    .A2(_0610_));
 sg13g2_a21oi_1 _1557_ (.A1(net394),
    .A2(_0597_),
    .Y(_0627_),
    .B1(net368));
 sg13g2_a21oi_1 _1558_ (.A1(net361),
    .A2(_0466_),
    .Y(_0628_),
    .B1(net345));
 sg13g2_o21ai_1 _1559_ (.B1(_0628_),
    .Y(_0629_),
    .A1(_0594_),
    .A2(_0627_));
 sg13g2_nor2_1 _1560_ (.A(_0469_),
    .B(_0524_),
    .Y(_0630_));
 sg13g2_nor4_2 _1561_ (.A(net364),
    .B(net358),
    .C(_0477_),
    .Y(_0631_),
    .D(_0630_));
 sg13g2_a21oi_1 _1562_ (.A1(net342),
    .A2(_0530_),
    .Y(_0632_),
    .B1(_0631_));
 sg13g2_a21o_1 _1563_ (.A2(_0632_),
    .A1(_0629_),
    .B1(net335),
    .X(_0633_));
 sg13g2_a21oi_1 _1564_ (.A1(_0430_),
    .A2(_0539_),
    .Y(_0634_),
    .B1(net346));
 sg13g2_nand3b_1 _1565_ (.B(net368),
    .C(_0521_),
    .Y(_0635_),
    .A_N(_0557_));
 sg13g2_nand2_1 _1566_ (.Y(_0636_),
    .A(net387),
    .B(_0597_));
 sg13g2_a21oi_1 _1567_ (.A1(_0603_),
    .A2(_0636_),
    .Y(_0637_),
    .B1(net356));
 sg13g2_a21oi_1 _1568_ (.A1(_0635_),
    .A2(_0637_),
    .Y(_0638_),
    .B1(_0634_));
 sg13g2_a21oi_1 _1569_ (.A1(net335),
    .A2(_0638_),
    .Y(_0639_),
    .B1(net329));
 sg13g2_o21ai_1 _1570_ (.B1(net388),
    .Y(_0640_),
    .A1(_0458_),
    .A2(_0531_));
 sg13g2_o21ai_1 _1571_ (.B1(_0640_),
    .Y(_0641_),
    .A1(_0407_),
    .A2(_0516_));
 sg13g2_nor3_1 _1572_ (.A(net363),
    .B(net349),
    .C(_0641_),
    .Y(_0642_));
 sg13g2_o21ai_1 _1573_ (.B1(_0575_),
    .Y(_0643_),
    .A1(_0383_),
    .A2(_0427_));
 sg13g2_a21oi_1 _1574_ (.A1(net382),
    .A2(net380),
    .Y(_0644_),
    .B1(_0480_));
 sg13g2_a21oi_1 _1575_ (.A1(_0521_),
    .A2(_0644_),
    .Y(_0645_),
    .B1(net358));
 sg13g2_a21oi_1 _1576_ (.A1(_0554_),
    .A2(_0602_),
    .Y(_0646_),
    .B1(net374));
 sg13g2_a221oi_1 _1577_ (.B2(net358),
    .C1(_0642_),
    .B1(_0646_),
    .A1(_0643_),
    .Y(_0647_),
    .A2(_0645_));
 sg13g2_nand2_1 _1578_ (.Y(_0648_),
    .A(_0552_),
    .B(_0568_));
 sg13g2_a21oi_1 _1579_ (.A1(net395),
    .A2(_0425_),
    .Y(_0649_),
    .B1(_0503_));
 sg13g2_or2_1 _1580_ (.X(_0650_),
    .B(_0649_),
    .A(net368));
 sg13g2_a21o_1 _1581_ (.A2(_0650_),
    .A1(_0648_),
    .B1(net345),
    .X(_0651_));
 sg13g2_nand2_1 _1582_ (.Y(_0652_),
    .A(_0506_),
    .B(_0560_));
 sg13g2_nor2_1 _1583_ (.A(net393),
    .B(_0407_),
    .Y(_0653_));
 sg13g2_nand2_1 _1584_ (.Y(_0654_),
    .A(net391),
    .B(_0408_));
 sg13g2_nor4_1 _1585_ (.A(net368),
    .B(_0569_),
    .C(_0601_),
    .D(_0653_),
    .Y(_0655_));
 sg13g2_a22oi_1 _1586_ (.Y(_0656_),
    .B1(_0655_),
    .B2(net345),
    .A2(_0652_),
    .A1(net341));
 sg13g2_nand3_1 _1587_ (.B(_0651_),
    .C(_0656_),
    .A(net335),
    .Y(_0657_));
 sg13g2_a21oi_1 _1588_ (.A1(net331),
    .A2(_0647_),
    .Y(_0658_),
    .B1(net328));
 sg13g2_a22oi_1 _1589_ (.Y(_0659_),
    .B1(_0657_),
    .B2(_0658_),
    .A2(_0639_),
    .A1(_0633_));
 sg13g2_or4_1 _1590_ (.A(net370),
    .B(net346),
    .C(_0440_),
    .D(_0442_),
    .X(_0660_));
 sg13g2_nor2_1 _1591_ (.A(_0402_),
    .B(_0525_),
    .Y(_0661_));
 sg13g2_nor2_1 _1592_ (.A(net379),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_o21ai_1 _1593_ (.B1(_0480_),
    .Y(_0663_),
    .A1(_0014_),
    .A2(net404));
 sg13g2_nand2_1 _1594_ (.Y(_0664_),
    .A(_0470_),
    .B(_0515_));
 sg13g2_nand3_1 _1595_ (.B(_0663_),
    .C(_0664_),
    .A(net341),
    .Y(_0665_));
 sg13g2_a22oi_1 _1596_ (.Y(_0666_),
    .B1(net402),
    .B2(_0483_),
    .A2(_0403_),
    .A1(net394));
 sg13g2_a22oi_1 _1597_ (.Y(_0667_),
    .B1(_0666_),
    .B2(_0499_),
    .A2(_0662_),
    .A1(net344));
 sg13g2_nand4_1 _1598_ (.B(_0660_),
    .C(_0665_),
    .A(net335),
    .Y(_0668_),
    .D(_0667_));
 sg13g2_nand2_2 _1599_ (.Y(_0669_),
    .A(net386),
    .B(_0391_));
 sg13g2_nand2_1 _1600_ (.Y(_0670_),
    .A(net420),
    .B(net389));
 sg13g2_nor2_2 _1601_ (.A(net400),
    .B(_0398_),
    .Y(_0671_));
 sg13g2_nand2_1 _1602_ (.Y(_0672_),
    .A(net387),
    .B(_0399_));
 sg13g2_nand2_2 _1603_ (.Y(_0673_),
    .A(_0405_),
    .B(_0671_));
 sg13g2_nand3_1 _1604_ (.B(_0478_),
    .C(_0673_),
    .A(net370),
    .Y(_0674_));
 sg13g2_o21ai_1 _1605_ (.B1(net395),
    .Y(_0675_),
    .A1(net408),
    .A2(_0402_));
 sg13g2_a21oi_1 _1606_ (.A1(_0412_),
    .A2(_0675_),
    .Y(_0676_),
    .B1(net345));
 sg13g2_a221oi_1 _1607_ (.B2(_0669_),
    .C1(net355),
    .B1(_0603_),
    .A1(_0428_),
    .Y(_0677_),
    .A2(_0539_));
 sg13g2_a21o_1 _1608_ (.A2(_0676_),
    .A1(_0674_),
    .B1(_0677_),
    .X(_0678_));
 sg13g2_a21oi_1 _1609_ (.A1(net331),
    .A2(_0678_),
    .Y(_0679_),
    .B1(net328));
 sg13g2_nor2_2 _1610_ (.A(net391),
    .B(_0440_),
    .Y(_0680_));
 sg13g2_nor2_2 _1611_ (.A(net377),
    .B(_0680_),
    .Y(_0681_));
 sg13g2_o21ai_1 _1612_ (.B1(_0484_),
    .Y(_0682_),
    .A1(_0525_),
    .A2(_0531_));
 sg13g2_a221oi_1 _1613_ (.B2(net371),
    .C1(net348),
    .B1(_0682_),
    .A1(_0619_),
    .Y(_0683_),
    .A2(_0681_));
 sg13g2_a21oi_1 _1614_ (.A1(net341),
    .A2(_0475_),
    .Y(_0684_),
    .B1(_0683_));
 sg13g2_a221oi_1 _1615_ (.B2(_0442_),
    .C1(net370),
    .B1(_0536_),
    .A1(net415),
    .Y(_0685_),
    .A2(_0466_));
 sg13g2_nor2b_1 _1616_ (.A(_0685_),
    .B_N(_0527_),
    .Y(_0686_));
 sg13g2_nand2_1 _1617_ (.Y(_0687_),
    .A(_0425_),
    .B(_0468_));
 sg13g2_a221oi_1 _1618_ (.B2(net362),
    .C1(net355),
    .B1(_0687_),
    .A1(_0443_),
    .Y(_0688_),
    .A2(_0472_));
 sg13g2_o21ai_1 _1619_ (.B1(net335),
    .Y(_0689_),
    .A1(_0686_),
    .A2(_0688_));
 sg13g2_o21ai_1 _1620_ (.B1(_0689_),
    .Y(_0690_),
    .A1(net335),
    .A2(_0684_));
 sg13g2_a221oi_1 _1621_ (.B2(net328),
    .C1(_0497_),
    .B1(_0690_),
    .A1(_0668_),
    .Y(_0691_),
    .A2(_0679_));
 sg13g2_o21ai_1 _1622_ (.B1(_0549_),
    .Y(_0692_),
    .A1(net326),
    .A2(_0659_));
 sg13g2_o21ai_1 _1623_ (.B1(net342),
    .Y(_0693_),
    .A1(_0507_),
    .A2(_0618_));
 sg13g2_inv_1 _1624_ (.Y(_0694_),
    .A(_0693_));
 sg13g2_nor2_1 _1625_ (.A(_0385_),
    .B(_0475_),
    .Y(_0695_));
 sg13g2_a221oi_1 _1626_ (.B2(_0557_),
    .C1(_0475_),
    .B1(_0417_),
    .A1(net396),
    .Y(_0696_),
    .A2(net415));
 sg13g2_a22oi_1 _1627_ (.Y(_0697_),
    .B1(_0696_),
    .B2(net362),
    .A2(_0513_),
    .A1(net345));
 sg13g2_a21oi_1 _1628_ (.A1(_0434_),
    .A2(_0697_),
    .Y(_0698_),
    .B1(_0694_));
 sg13g2_a21oi_1 _1629_ (.A1(net325),
    .A2(_0698_),
    .Y(_0699_),
    .B1(_0189_));
 sg13g2_o21ai_1 _1630_ (.B1(_0699_),
    .Y(_0700_),
    .A1(_0691_),
    .A2(_0692_));
 sg13g2_a21o_1 _1631_ (.A2(_0700_),
    .A1(_0626_),
    .B1(\g_x[1] ),
    .X(_0701_));
 sg13g2_nand2_1 _1632_ (.Y(_0702_),
    .A(net362),
    .B(_0570_));
 sg13g2_a21oi_1 _1633_ (.A1(net363),
    .A2(_0570_),
    .Y(_0703_),
    .B1(net349));
 sg13g2_nor2_1 _1634_ (.A(net376),
    .B(_0583_),
    .Y(_0704_));
 sg13g2_or2_1 _1635_ (.X(_0705_),
    .B(_0583_),
    .A(net375));
 sg13g2_nor2_1 _1636_ (.A(net361),
    .B(_0534_),
    .Y(_0706_));
 sg13g2_a22oi_1 _1637_ (.Y(_0707_),
    .B1(_0706_),
    .B2(_0401_),
    .A2(_0583_),
    .A1(net362));
 sg13g2_nor4_2 _1638_ (.A(_0356_),
    .B(_0394_),
    .C(_0466_),
    .Y(_0708_),
    .D(_0505_));
 sg13g2_and2_2 _1639_ (.A(net363),
    .B(_0553_),
    .X(_0709_));
 sg13g2_nor3_1 _1640_ (.A(net390),
    .B(_0439_),
    .C(_0535_),
    .Y(_0710_));
 sg13g2_nor3_2 _1641_ (.A(_0356_),
    .B(_0394_),
    .C(_0710_),
    .Y(_0711_));
 sg13g2_o21ai_1 _1642_ (.B1(_0537_),
    .Y(_0712_),
    .A1(net409),
    .A2(_0402_));
 sg13g2_a221oi_1 _1643_ (.B2(net404),
    .C1(net369),
    .B1(_0653_),
    .A1(net393),
    .Y(_0713_),
    .A2(_0421_));
 sg13g2_a21o_1 _1644_ (.A2(_0712_),
    .A1(_0711_),
    .B1(_0713_),
    .X(_0714_));
 sg13g2_a22oi_1 _1645_ (.Y(_0715_),
    .B1(_0709_),
    .B2(_0430_),
    .A2(_0708_),
    .A1(_0695_));
 sg13g2_mux4_1 _1646_ (.S0(net347),
    .A0(_0702_),
    .A1(_0707_),
    .A2(_0714_),
    .A3(_0715_),
    .S1(_0380_),
    .X(_0716_));
 sg13g2_nand2_1 _1647_ (.Y(_0717_),
    .A(_0471_),
    .B(_0529_));
 sg13g2_and3_1 _1648_ (.X(_0718_),
    .A(net374),
    .B(_0481_),
    .C(_0615_));
 sg13g2_nor2_1 _1649_ (.A(_0402_),
    .B(_0574_),
    .Y(_0719_));
 sg13g2_nand3_1 _1650_ (.B(net380),
    .C(_0569_),
    .A(net382),
    .Y(_0720_));
 sg13g2_o21ai_1 _1651_ (.B1(_0720_),
    .Y(_0721_),
    .A1(net374),
    .A2(_0719_));
 sg13g2_o21ai_1 _1652_ (.B1(net358),
    .Y(_0722_),
    .A1(_0718_),
    .A2(_0721_));
 sg13g2_a22oi_1 _1653_ (.Y(_0723_),
    .B1(_0717_),
    .B2(_0456_),
    .A2(_0476_),
    .A1(net344));
 sg13g2_nand3_1 _1654_ (.B(_0722_),
    .C(_0723_),
    .A(net333),
    .Y(_0724_));
 sg13g2_nor3_1 _1655_ (.A(net376),
    .B(net350),
    .C(_0509_),
    .Y(_0725_));
 sg13g2_nand2_1 _1656_ (.Y(_0726_),
    .A(_0464_),
    .B(_0555_));
 sg13g2_o21ai_1 _1657_ (.B1(_0708_),
    .Y(_0727_),
    .A1(net390),
    .A2(_0418_));
 sg13g2_a21oi_1 _1658_ (.A1(_0599_),
    .A2(_0616_),
    .Y(_0728_),
    .B1(net356));
 sg13g2_a221oi_1 _1659_ (.B2(_0728_),
    .C1(_0725_),
    .B1(_0727_),
    .A1(_0499_),
    .Y(_0729_),
    .A2(_0726_));
 sg13g2_a21oi_1 _1660_ (.A1(net334),
    .A2(_0729_),
    .Y(_0730_),
    .B1(net329));
 sg13g2_a221oi_1 _1661_ (.B2(_0730_),
    .C1(_0497_),
    .B1(_0724_),
    .A1(net329),
    .Y(_0731_),
    .A2(_0716_));
 sg13g2_nand2_1 _1662_ (.Y(_0732_),
    .A(net401),
    .B(_0503_));
 sg13g2_nand3_1 _1663_ (.B(net357),
    .C(_0732_),
    .A(net375),
    .Y(_0733_));
 sg13g2_nand2_1 _1664_ (.Y(_0734_),
    .A(_0393_),
    .B(_0467_));
 sg13g2_a221oi_1 _1665_ (.B2(_0385_),
    .C1(_0466_),
    .B1(_0392_),
    .A1(net388),
    .Y(_0735_),
    .A2(_0390_));
 sg13g2_nand3b_1 _1666_ (.B(net373),
    .C(net352),
    .Y(_0736_),
    .A_N(_0735_));
 sg13g2_nand3b_1 _1667_ (.B(_0733_),
    .C(_0736_),
    .Y(_0737_),
    .A_N(_0681_));
 sg13g2_and2_1 _1668_ (.A(net353),
    .B(_0611_),
    .X(_0738_));
 sg13g2_nor2_1 _1669_ (.A(net353),
    .B(_0711_),
    .Y(_0739_));
 sg13g2_nor2_2 _1670_ (.A(_0458_),
    .B(_0672_),
    .Y(_0740_));
 sg13g2_or2_1 _1671_ (.X(_0741_),
    .B(_0740_),
    .A(net375));
 sg13g2_and3_1 _1672_ (.X(_0742_),
    .A(net375),
    .B(net353),
    .C(_0563_));
 sg13g2_a221oi_1 _1673_ (.B2(_0741_),
    .C1(_0742_),
    .B1(_0739_),
    .A1(_0512_),
    .Y(_0743_),
    .A2(_0738_));
 sg13g2_mux2_1 _1674_ (.A0(_0737_),
    .A1(_0743_),
    .S(net337),
    .X(_0744_));
 sg13g2_o21ai_1 _1675_ (.B1(_0640_),
    .Y(_0745_),
    .A1(_0482_),
    .A2(_0516_));
 sg13g2_nand2_1 _1676_ (.Y(_0746_),
    .A(net391),
    .B(_0416_));
 sg13g2_nor2_1 _1677_ (.A(net397),
    .B(_0415_),
    .Y(_0747_));
 sg13g2_nor2_1 _1678_ (.A(net399),
    .B(_0440_),
    .Y(_0748_));
 sg13g2_nor2_1 _1679_ (.A(_0400_),
    .B(_0748_),
    .Y(_0749_));
 sg13g2_or4_1 _1680_ (.A(net364),
    .B(_0400_),
    .C(net378),
    .D(_0748_),
    .X(_0750_));
 sg13g2_a221oi_1 _1681_ (.B2(net351),
    .C1(_0566_),
    .B1(_0750_),
    .A1(_0499_),
    .Y(_0751_),
    .A2(_0745_));
 sg13g2_o21ai_1 _1682_ (.B1(_0406_),
    .Y(_0752_),
    .A1(_0501_),
    .A2(_0612_));
 sg13g2_nand2b_1 _1683_ (.Y(_0753_),
    .B(_0499_),
    .A_N(_0474_));
 sg13g2_nor2_1 _1684_ (.A(_0509_),
    .B(_0719_),
    .Y(_0754_));
 sg13g2_nand3_1 _1685_ (.B(net402),
    .C(_0589_),
    .A(net364),
    .Y(_0755_));
 sg13g2_a22oi_1 _1686_ (.Y(_0756_),
    .B1(_0754_),
    .B2(net340),
    .A2(_0752_),
    .A1(net343));
 sg13g2_nand4_1 _1687_ (.B(_0753_),
    .C(_0755_),
    .A(net336),
    .Y(_0757_),
    .D(_0756_));
 sg13g2_a21oi_1 _1688_ (.A1(net332),
    .A2(_0751_),
    .Y(_0758_),
    .B1(net327));
 sg13g2_a221oi_1 _1689_ (.B2(_0758_),
    .C1(_0498_),
    .B1(_0757_),
    .A1(net327),
    .Y(_0759_),
    .A2(_0744_));
 sg13g2_o21ai_1 _1690_ (.B1(_0549_),
    .Y(_0760_),
    .A1(_0731_),
    .A2(_0759_));
 sg13g2_a21oi_1 _1691_ (.A1(_0619_),
    .A2(_0695_),
    .Y(_0761_),
    .B1(net371));
 sg13g2_o21ai_1 _1692_ (.B1(net355),
    .Y(_0762_),
    .A1(_0613_),
    .A2(_0761_));
 sg13g2_nor3_1 _1693_ (.A(net397),
    .B(_0536_),
    .C(_0761_),
    .Y(_0763_));
 sg13g2_o21ai_1 _1694_ (.B1(net342),
    .Y(_0764_),
    .A1(_0618_),
    .A2(_0747_));
 sg13g2_o21ai_1 _1695_ (.B1(_0764_),
    .Y(_0765_),
    .A1(_0762_),
    .A2(_0763_));
 sg13g2_a21oi_1 _1696_ (.A1(net341),
    .A2(_0478_),
    .Y(_0766_),
    .B1(_0765_));
 sg13g2_nand2_1 _1697_ (.Y(_0767_),
    .A(net325),
    .B(_0766_));
 sg13g2_and4_1 _1698_ (.A(\g_x[0] ),
    .B(\g_x[1] ),
    .C(_0760_),
    .D(_0767_),
    .X(_0768_));
 sg13g2_or3_1 _1699_ (.A(net364),
    .B(_0514_),
    .C(_0735_),
    .X(_0769_));
 sg13g2_nand3_1 _1700_ (.B(_0591_),
    .C(_0769_),
    .A(net332),
    .Y(_0770_));
 sg13g2_nand3_1 _1701_ (.B(net379),
    .C(_0440_),
    .A(net373),
    .Y(_0771_));
 sg13g2_or3_1 _1702_ (.A(net373),
    .B(_0514_),
    .C(_0748_),
    .X(_0772_));
 sg13g2_nand3_1 _1703_ (.B(_0771_),
    .C(_0772_),
    .A(net336),
    .Y(_0773_));
 sg13g2_nand3_1 _1704_ (.B(_0770_),
    .C(_0773_),
    .A(net351),
    .Y(_0774_));
 sg13g2_nor2_1 _1705_ (.A(net375),
    .B(_0671_),
    .Y(_0775_));
 sg13g2_o21ai_1 _1706_ (.B1(net398),
    .Y(_0776_),
    .A1(_0389_),
    .A2(_0398_));
 sg13g2_a22oi_1 _1707_ (.Y(_0777_),
    .B1(_0775_),
    .B2(_0776_),
    .A2(_0593_),
    .A1(_0575_));
 sg13g2_a22oi_1 _1708_ (.Y(_0778_),
    .B1(_0746_),
    .B2(_0431_),
    .A2(_0740_),
    .A1(net365));
 sg13g2_mux2_1 _1709_ (.A0(_0777_),
    .A1(_0778_),
    .S(net336),
    .X(_0779_));
 sg13g2_a21oi_1 _1710_ (.A1(net357),
    .A2(_0779_),
    .Y(_0780_),
    .B1(net330));
 sg13g2_a221oi_1 _1711_ (.B2(net379),
    .C1(net361),
    .B1(_0419_),
    .A1(net384),
    .Y(_0781_),
    .A2(net415));
 sg13g2_a21oi_1 _1712_ (.A1(_0420_),
    .A2(_0752_),
    .Y(_0782_),
    .B1(net368));
 sg13g2_o21ai_1 _1713_ (.B1(net335),
    .Y(_0783_),
    .A1(_0781_),
    .A2(_0782_));
 sg13g2_a221oi_1 _1714_ (.B2(_0502_),
    .C1(net368),
    .B1(net379),
    .A1(net385),
    .Y(_0784_),
    .A2(_0420_));
 sg13g2_a221oi_1 _1715_ (.B2(_0557_),
    .C1(net361),
    .B1(_0416_),
    .A1(_0385_),
    .Y(_0785_),
    .A2(net403));
 sg13g2_o21ai_1 _1716_ (.B1(net331),
    .Y(_0786_),
    .A1(_0784_),
    .A2(_0785_));
 sg13g2_nand3_1 _1717_ (.B(_0783_),
    .C(_0786_),
    .A(net345),
    .Y(_0787_));
 sg13g2_o21ai_1 _1718_ (.B1(_0611_),
    .Y(_0788_),
    .A1(_0428_),
    .A2(_0439_));
 sg13g2_nand2_1 _1719_ (.Y(_0789_),
    .A(_0390_),
    .B(net379));
 sg13g2_nand2_1 _1720_ (.Y(_0790_),
    .A(net374),
    .B(_0789_));
 sg13g2_o21ai_1 _1721_ (.B1(_0788_),
    .Y(_0791_),
    .A1(_0480_),
    .A2(_0790_));
 sg13g2_o21ai_1 _1722_ (.B1(_0603_),
    .Y(_0792_),
    .A1(net394),
    .A2(_0424_));
 sg13g2_o21ai_1 _1723_ (.B1(net369),
    .Y(_0793_),
    .A1(_0404_),
    .A2(_0516_));
 sg13g2_a21o_1 _1724_ (.A2(_0793_),
    .A1(_0792_),
    .B1(net334),
    .X(_0794_));
 sg13g2_a21oi_1 _1725_ (.A1(net334),
    .A2(_0791_),
    .Y(_0795_),
    .B1(net347));
 sg13g2_a21oi_1 _1726_ (.A1(_0794_),
    .A2(_0795_),
    .Y(_0796_),
    .B1(net328));
 sg13g2_a221oi_1 _1727_ (.B2(_0796_),
    .C1(net326),
    .B1(_0787_),
    .A1(_0774_),
    .Y(_0797_),
    .A2(_0780_));
 sg13g2_nand3_1 _1728_ (.B(net340),
    .C(_0475_),
    .A(_0408_),
    .Y(_0798_));
 sg13g2_nand2_1 _1729_ (.Y(_0799_),
    .A(net363),
    .B(_0467_));
 sg13g2_nand2b_1 _1730_ (.Y(_0800_),
    .B(net364),
    .A_N(_0471_));
 sg13g2_nor2_1 _1731_ (.A(_0471_),
    .B(_0705_),
    .Y(_0801_));
 sg13g2_nor2_1 _1732_ (.A(_0511_),
    .B(_0740_),
    .Y(_0802_));
 sg13g2_a221oi_1 _1733_ (.B2(_0499_),
    .C1(net338),
    .B1(_0802_),
    .A1(net359),
    .Y(_0803_),
    .A2(_0801_));
 sg13g2_and3_2 _1734_ (.X(_0804_),
    .A(net383),
    .B(net381),
    .C(_0619_));
 sg13g2_a221oi_1 _1735_ (.B2(_0555_),
    .C1(net349),
    .B1(_0804_),
    .A1(_0521_),
    .Y(_0805_),
    .A2(_0709_));
 sg13g2_nand2_1 _1736_ (.Y(_0806_),
    .A(_0436_),
    .B(_0473_));
 sg13g2_a22oi_1 _1737_ (.Y(_0807_),
    .B1(_0806_),
    .B2(net340),
    .A2(_0654_),
    .A1(net344));
 sg13g2_nand2b_1 _1738_ (.Y(_0808_),
    .B(_0807_),
    .A_N(_0805_));
 sg13g2_a221oi_1 _1739_ (.B2(net338),
    .C1(net330),
    .B1(_0808_),
    .A1(_0798_),
    .Y(_0809_),
    .A2(_0803_));
 sg13g2_nand2_1 _1740_ (.Y(_0810_),
    .A(_0593_),
    .B(_0804_));
 sg13g2_a21oi_1 _1741_ (.A1(net398),
    .A2(_0502_),
    .Y(_0811_),
    .B1(_0523_));
 sg13g2_a21oi_1 _1742_ (.A1(net374),
    .A2(_0811_),
    .Y(_0812_),
    .B1(_0509_));
 sg13g2_a22oi_1 _1743_ (.Y(_0813_),
    .B1(_0812_),
    .B2(_0703_),
    .A2(_0810_),
    .A1(net349));
 sg13g2_a221oi_1 _1744_ (.B2(_0671_),
    .C1(_0434_),
    .B1(_0459_),
    .A1(net400),
    .Y(_0814_),
    .A2(net406));
 sg13g2_nor3_1 _1745_ (.A(net333),
    .B(_0813_),
    .C(_0814_),
    .Y(_0815_));
 sg13g2_nand3_1 _1746_ (.B(_0411_),
    .C(_0563_),
    .A(net365),
    .Y(_0816_));
 sg13g2_nand3_1 _1747_ (.B(_0478_),
    .C(_0636_),
    .A(net371),
    .Y(_0817_));
 sg13g2_nand3_1 _1748_ (.B(_0816_),
    .C(_0817_),
    .A(net359),
    .Y(_0818_));
 sg13g2_nor2_1 _1749_ (.A(net398),
    .B(_0564_),
    .Y(_0819_));
 sg13g2_or2_1 _1750_ (.X(_0820_),
    .B(_0564_),
    .A(net398));
 sg13g2_nand2b_1 _1751_ (.Y(_0821_),
    .B(_0820_),
    .A_N(_0385_));
 sg13g2_a22oi_1 _1752_ (.Y(_0822_),
    .B1(_0821_),
    .B2(net340),
    .A2(_0646_),
    .A1(net349));
 sg13g2_a21oi_1 _1753_ (.A1(_0818_),
    .A2(_0822_),
    .Y(_0823_),
    .B1(net338));
 sg13g2_nor3_1 _1754_ (.A(net327),
    .B(_0815_),
    .C(_0823_),
    .Y(_0824_));
 sg13g2_nor3_1 _1755_ (.A(_0497_),
    .B(_0809_),
    .C(_0824_),
    .Y(_0825_));
 sg13g2_or3_1 _1756_ (.A(net325),
    .B(_0797_),
    .C(_0825_),
    .X(_0826_));
 sg13g2_nor2_1 _1757_ (.A(_0585_),
    .B(_0694_),
    .Y(_0827_));
 sg13g2_and3_1 _1758_ (.X(_0828_),
    .A(net325),
    .B(_0762_),
    .C(_0827_));
 sg13g2_nor3_1 _1759_ (.A(\g_x[0] ),
    .B(_0197_),
    .C(_0828_),
    .Y(_0829_));
 sg13g2_a21oi_1 _1760_ (.A1(_0826_),
    .A2(_0829_),
    .Y(_0830_),
    .B1(_0768_));
 sg13g2_a21oi_2 _1761_ (.B1(_0202_),
    .Y(_0831_),
    .A2(_0830_),
    .A1(_0701_));
 sg13g2_nand3_1 _1762_ (.B(_0467_),
    .C(_0602_),
    .A(net375),
    .Y(_0832_));
 sg13g2_nand2_1 _1763_ (.Y(_0833_),
    .A(net365),
    .B(_0671_));
 sg13g2_nand3_1 _1764_ (.B(_0832_),
    .C(_0833_),
    .A(net357),
    .Y(_0834_));
 sg13g2_o21ai_1 _1765_ (.B1(net375),
    .Y(_0835_),
    .A1(_0474_),
    .A2(_0477_));
 sg13g2_nand3_1 _1766_ (.B(_0512_),
    .C(_0673_),
    .A(net365),
    .Y(_0836_));
 sg13g2_nand3_1 _1767_ (.B(_0835_),
    .C(_0836_),
    .A(net353),
    .Y(_0837_));
 sg13g2_nand3_1 _1768_ (.B(_0834_),
    .C(_0837_),
    .A(net337),
    .Y(_0838_));
 sg13g2_nand3_1 _1769_ (.B(_0401_),
    .C(_0602_),
    .A(net377),
    .Y(_0839_));
 sg13g2_nand4_1 _1770_ (.B(net361),
    .C(_0472_),
    .A(_0388_),
    .Y(_0840_),
    .D(_0515_));
 sg13g2_nand3_1 _1771_ (.B(_0839_),
    .C(_0840_),
    .A(net360),
    .Y(_0841_));
 sg13g2_nand4_1 _1772_ (.B(_0586_),
    .C(_0736_),
    .A(net332),
    .Y(_0842_),
    .D(_0841_));
 sg13g2_a21oi_1 _1773_ (.A1(_0838_),
    .A2(_0842_),
    .Y(_0843_),
    .B1(net330));
 sg13g2_a221oi_1 _1774_ (.B2(_0804_),
    .C1(net349),
    .B1(_0789_),
    .A1(_0524_),
    .Y(_0844_),
    .A2(_0592_));
 sg13g2_o21ai_1 _1775_ (.B1(net340),
    .Y(_0845_),
    .A1(_0583_),
    .A2(_0740_));
 sg13g2_nand2_1 _1776_ (.Y(_0846_),
    .A(_0506_),
    .B(_0612_));
 sg13g2_a21oi_1 _1777_ (.A1(net343),
    .A2(_0846_),
    .Y(_0847_),
    .B1(_0844_));
 sg13g2_a21oi_1 _1778_ (.A1(_0845_),
    .A2(_0847_),
    .Y(_0848_),
    .B1(net332));
 sg13g2_nor2_1 _1779_ (.A(net399),
    .B(_0616_),
    .Y(_0849_));
 sg13g2_nand3_1 _1780_ (.B(_0401_),
    .C(_0457_),
    .A(net373),
    .Y(_0850_));
 sg13g2_o21ai_1 _1781_ (.B1(_0850_),
    .Y(_0851_),
    .A1(_0591_),
    .A2(_0849_));
 sg13g2_a21oi_1 _1782_ (.A1(_0566_),
    .A2(_0670_),
    .Y(_0852_),
    .B1(net351));
 sg13g2_a221oi_1 _1783_ (.B2(_0771_),
    .C1(net336),
    .B1(_0852_),
    .A1(net352),
    .Y(_0853_),
    .A2(_0851_));
 sg13g2_nor3_1 _1784_ (.A(net328),
    .B(_0848_),
    .C(_0853_),
    .Y(_0854_));
 sg13g2_nor3_1 _1785_ (.A(net326),
    .B(_0843_),
    .C(_0854_),
    .Y(_0855_));
 sg13g2_nand4_1 _1786_ (.B(net356),
    .C(_0510_),
    .A(net362),
    .Y(_0856_),
    .D(_0571_));
 sg13g2_o21ai_1 _1787_ (.B1(_0856_),
    .Y(_0857_),
    .A1(_0500_),
    .A2(_0811_));
 sg13g2_a21oi_1 _1788_ (.A1(_0612_),
    .A2(_0804_),
    .Y(_0858_),
    .B1(net358));
 sg13g2_nor3_1 _1789_ (.A(net373),
    .B(_0569_),
    .C(_0748_),
    .Y(_0859_));
 sg13g2_nor2b_1 _1790_ (.A(_0859_),
    .B_N(_0858_),
    .Y(_0860_));
 sg13g2_or3_1 _1791_ (.A(net333),
    .B(_0857_),
    .C(_0860_),
    .X(_0861_));
 sg13g2_nand3_1 _1792_ (.B(_0459_),
    .C(_0536_),
    .A(net400),
    .Y(_0862_));
 sg13g2_nand3_1 _1793_ (.B(_0820_),
    .C(_0862_),
    .A(net376),
    .Y(_0863_));
 sg13g2_a22oi_1 _1794_ (.Y(_0864_),
    .B1(_0863_),
    .B2(_0705_),
    .A2(_0819_),
    .A1(net402));
 sg13g2_and2_1 _1795_ (.A(net363),
    .B(_0437_),
    .X(_0865_));
 sg13g2_a221oi_1 _1796_ (.B2(_0865_),
    .C1(net350),
    .B1(_0862_),
    .A1(_0584_),
    .Y(_0866_),
    .A2(_0669_));
 sg13g2_o21ai_1 _1797_ (.B1(net333),
    .Y(_0867_),
    .A1(net357),
    .A2(_0864_));
 sg13g2_o21ai_1 _1798_ (.B1(_0861_),
    .Y(_0868_),
    .A1(_0866_),
    .A2(_0867_));
 sg13g2_nor2_1 _1799_ (.A(net365),
    .B(_0567_),
    .Y(_0869_));
 sg13g2_nand2_1 _1800_ (.Y(_0870_),
    .A(_0471_),
    .B(_0502_));
 sg13g2_a221oi_1 _1801_ (.B2(_0704_),
    .C1(net350),
    .B1(_0870_),
    .A1(_0484_),
    .Y(_0871_),
    .A2(_0869_));
 sg13g2_a21oi_1 _1802_ (.A1(net375),
    .A2(_0570_),
    .Y(_0872_),
    .B1(net359));
 sg13g2_o21ai_1 _1803_ (.B1(net333),
    .Y(_0873_),
    .A1(_0871_),
    .A2(_0872_));
 sg13g2_a221oi_1 _1804_ (.B2(net389),
    .C1(_0719_),
    .B1(_0423_),
    .A1(net383),
    .Y(_0874_),
    .A2(net381));
 sg13g2_a21o_1 _1805_ (.A2(_0804_),
    .A1(_0457_),
    .B1(_0874_),
    .X(_0875_));
 sg13g2_a22oi_1 _1806_ (.Y(_0876_),
    .B1(_0875_),
    .B2(net357),
    .A2(_0858_),
    .A1(_0800_));
 sg13g2_a21oi_1 _1807_ (.A1(net337),
    .A2(_0876_),
    .Y(_0877_),
    .B1(net330));
 sg13g2_a221oi_1 _1808_ (.B2(_0877_),
    .C1(_0497_),
    .B1(_0873_),
    .A1(net330),
    .Y(_0878_),
    .A2(_0868_));
 sg13g2_or3_1 _1809_ (.A(_0550_),
    .B(_0855_),
    .C(_0878_),
    .X(_0879_));
 sg13g2_nor2_2 _1810_ (.A(net371),
    .B(_0696_),
    .Y(_0880_));
 sg13g2_o21ai_1 _1811_ (.B1(net359),
    .Y(_0881_),
    .A1(_0869_),
    .A2(_0880_));
 sg13g2_nor2b_1 _1812_ (.A(_0880_),
    .B_N(_0680_),
    .Y(_0882_));
 sg13g2_a21oi_1 _1813_ (.A1(_0476_),
    .A2(_0802_),
    .Y(_0883_),
    .B1(_0434_));
 sg13g2_nand2b_1 _1814_ (.Y(_0884_),
    .B(net340),
    .A_N(_0514_));
 sg13g2_o21ai_1 _1815_ (.B1(_0884_),
    .Y(_0885_),
    .A1(_0881_),
    .A2(_0882_));
 sg13g2_nor2_1 _1816_ (.A(_0883_),
    .B(_0885_),
    .Y(_0886_));
 sg13g2_a21oi_1 _1817_ (.A1(net325),
    .A2(_0886_),
    .Y(_0887_),
    .B1(\g_x[0] ));
 sg13g2_nand3b_1 _1818_ (.B(net393),
    .C(_0419_),
    .Y(_0888_),
    .A_N(_0531_));
 sg13g2_nand3_1 _1819_ (.B(_0709_),
    .C(_0888_),
    .A(net347),
    .Y(_0889_));
 sg13g2_nand2_1 _1820_ (.Y(_0890_),
    .A(_0457_),
    .B(_0525_));
 sg13g2_o21ai_1 _1821_ (.B1(_0484_),
    .Y(_0891_),
    .A1(_0406_),
    .A2(_0423_));
 sg13g2_a22oi_1 _1822_ (.Y(_0892_),
    .B1(_0891_),
    .B2(_0499_),
    .A2(_0890_),
    .A1(net341));
 sg13g2_nand3_1 _1823_ (.B(_0889_),
    .C(_0892_),
    .A(_0856_),
    .Y(_0893_));
 sg13g2_o21ai_1 _1824_ (.B1(_0430_),
    .Y(_0894_),
    .A1(_0421_),
    .A2(_0820_));
 sg13g2_nand3_1 _1825_ (.B(_0538_),
    .C(_0560_),
    .A(net368),
    .Y(_0895_));
 sg13g2_o21ai_1 _1826_ (.B1(_0895_),
    .Y(_0896_),
    .A1(net369),
    .A2(_0894_));
 sg13g2_nand2_1 _1827_ (.Y(_0897_),
    .A(_0410_),
    .B(_0537_));
 sg13g2_a21oi_1 _1828_ (.A1(_0411_),
    .A2(_0577_),
    .Y(_0898_),
    .B1(net371));
 sg13g2_a21oi_1 _1829_ (.A1(_0711_),
    .A2(_0897_),
    .Y(_0899_),
    .B1(_0898_));
 sg13g2_mux2_1 _1830_ (.A0(_0896_),
    .A1(_0899_),
    .S(net355),
    .X(_0900_));
 sg13g2_o21ai_1 _1831_ (.B1(net329),
    .Y(_0901_),
    .A1(net339),
    .A2(_0900_));
 sg13g2_a21oi_1 _1832_ (.A1(net334),
    .A2(_0893_),
    .Y(_0902_),
    .B1(_0901_));
 sg13g2_o21ai_1 _1833_ (.B1(_0709_),
    .Y(_0903_),
    .A1(_0418_),
    .A2(_0428_));
 sg13g2_a22oi_1 _1834_ (.Y(_0904_),
    .B1(_0505_),
    .B2(_0392_),
    .A2(net378),
    .A1(_0502_));
 sg13g2_a21oi_1 _1835_ (.A1(net376),
    .A2(_0904_),
    .Y(_0905_),
    .B1(net350));
 sg13g2_a221oi_1 _1836_ (.B2(_0905_),
    .C1(net334),
    .B1(_0903_),
    .A1(net350),
    .Y(_0906_),
    .A2(_0720_));
 sg13g2_nor3_1 _1837_ (.A(net370),
    .B(_0530_),
    .C(_0661_),
    .Y(_0907_));
 sg13g2_a21oi_1 _1838_ (.A1(_0672_),
    .A2(_0706_),
    .Y(_0908_),
    .B1(_0907_));
 sg13g2_a221oi_1 _1839_ (.B2(net390),
    .C1(_0511_),
    .B1(_0409_),
    .A1(net383),
    .Y(_0909_),
    .A2(net381));
 sg13g2_a221oi_1 _1840_ (.B2(_0523_),
    .C1(net363),
    .B1(_0502_),
    .A1(_0392_),
    .Y(_0910_),
    .A2(_0429_));
 sg13g2_o21ai_1 _1841_ (.B1(net359),
    .Y(_0911_),
    .A1(_0909_),
    .A2(_0910_));
 sg13g2_o21ai_1 _1842_ (.B1(_0911_),
    .Y(_0912_),
    .A1(net356),
    .A2(_0908_));
 sg13g2_a21oi_1 _1843_ (.A1(net334),
    .A2(_0912_),
    .Y(_0913_),
    .B1(_0906_));
 sg13g2_o21ai_1 _1844_ (.B1(net326),
    .Y(_0914_),
    .A1(net329),
    .A2(_0913_));
 sg13g2_o21ai_1 _1845_ (.B1(_0506_),
    .Y(_0915_),
    .A1(_0404_),
    .A2(_0427_));
 sg13g2_nand2_1 _1846_ (.Y(_0916_),
    .A(net363),
    .B(_0915_));
 sg13g2_a21oi_1 _1847_ (.A1(_0510_),
    .A2(_0552_),
    .Y(_0917_),
    .B1(net347));
 sg13g2_nand2_1 _1848_ (.Y(_0918_),
    .A(_0916_),
    .B(_0917_));
 sg13g2_o21ai_1 _1849_ (.B1(_0578_),
    .Y(_0919_),
    .A1(net416),
    .A2(_0476_));
 sg13g2_nor3_1 _1850_ (.A(net376),
    .B(_0435_),
    .C(_0680_),
    .Y(_0920_));
 sg13g2_a22oi_1 _1851_ (.Y(_0921_),
    .B1(_0920_),
    .B2(net353),
    .A2(_0919_),
    .A1(net340));
 sg13g2_nand3_1 _1852_ (.B(_0918_),
    .C(_0921_),
    .A(net336),
    .Y(_0922_));
 sg13g2_o21ai_1 _1853_ (.B1(_0556_),
    .Y(_0923_),
    .A1(_0524_),
    .A2(_0531_));
 sg13g2_nand2_1 _1854_ (.Y(_0924_),
    .A(net374),
    .B(_0923_));
 sg13g2_a221oi_1 _1855_ (.B2(net398),
    .C1(net405),
    .B1(_0407_),
    .A1(net382),
    .Y(_0925_),
    .A2(net380));
 sg13g2_a21o_1 _1856_ (.A2(_0575_),
    .A1(_0460_),
    .B1(_0925_),
    .X(_0926_));
 sg13g2_a22oi_1 _1857_ (.Y(_0927_),
    .B1(_0926_),
    .B2(net351),
    .A2(_0924_),
    .A1(_0852_));
 sg13g2_a21oi_1 _1858_ (.A1(net332),
    .A2(_0927_),
    .Y(_0928_),
    .B1(net328));
 sg13g2_nor2_1 _1859_ (.A(_0468_),
    .B(_0617_),
    .Y(_0929_));
 sg13g2_o21ai_1 _1860_ (.B1(_0426_),
    .Y(_0930_),
    .A1(net387),
    .A2(_0415_));
 sg13g2_nor4_1 _1861_ (.A(net366),
    .B(_0400_),
    .C(net360),
    .D(_0929_),
    .Y(_0931_));
 sg13g2_a221oi_1 _1862_ (.B2(net343),
    .C1(_0931_),
    .B1(_0930_),
    .A1(net359),
    .Y(_0932_),
    .A2(_0832_));
 sg13g2_a221oi_1 _1863_ (.B2(_0504_),
    .C1(_0567_),
    .B1(_0405_),
    .A1(_0357_),
    .Y(_0933_),
    .A2(_0395_));
 sg13g2_and4_1 _1864_ (.A(_0357_),
    .B(_0395_),
    .C(_0746_),
    .D(_0862_),
    .X(_0934_));
 sg13g2_nor3_1 _1865_ (.A(net353),
    .B(_0933_),
    .C(_0934_),
    .Y(_0935_));
 sg13g2_nand2_1 _1866_ (.Y(_0936_),
    .A(_0410_),
    .B(net378));
 sg13g2_a221oi_1 _1867_ (.B2(_0936_),
    .C1(_0935_),
    .B1(_0738_),
    .A1(net340),
    .Y(_0937_),
    .A2(_0734_));
 sg13g2_mux2_1 _1868_ (.A0(_0932_),
    .A1(_0937_),
    .S(net332),
    .X(_0938_));
 sg13g2_a221oi_1 _1869_ (.B2(net327),
    .C1(net326),
    .B1(_0938_),
    .A1(_0922_),
    .Y(_0939_),
    .A2(_0928_));
 sg13g2_nor2_1 _1870_ (.A(_0550_),
    .B(_0939_),
    .Y(_0940_));
 sg13g2_o21ai_1 _1871_ (.B1(_0940_),
    .Y(_0941_),
    .A1(_0902_),
    .A2(_0914_));
 sg13g2_a221oi_1 _1872_ (.B2(net390),
    .C1(_0509_),
    .B1(_0535_),
    .A1(net383),
    .Y(_0942_),
    .A2(net381));
 sg13g2_o21ai_1 _1873_ (.B1(net347),
    .Y(_0943_),
    .A1(_0443_),
    .A2(_0942_));
 sg13g2_o21ai_1 _1874_ (.B1(net355),
    .Y(_0944_),
    .A1(_0613_),
    .A2(_0880_));
 sg13g2_and2_1 _1875_ (.A(_0943_),
    .B(_0944_),
    .X(_0945_));
 sg13g2_a21oi_1 _1876_ (.A1(net325),
    .A2(_0945_),
    .Y(_0946_),
    .B1(_0189_));
 sg13g2_a221oi_1 _1877_ (.B2(_0946_),
    .C1(_0197_),
    .B1(_0941_),
    .A1(_0879_),
    .Y(_0947_),
    .A2(_0887_));
 sg13g2_a221oi_1 _1878_ (.B2(_0644_),
    .C1(net358),
    .B1(_0615_),
    .A1(_0401_),
    .Y(_0948_),
    .A2(_0613_));
 sg13g2_nor3_1 _1879_ (.A(net333),
    .B(_0857_),
    .C(_0948_),
    .Y(_0949_));
 sg13g2_a221oi_1 _1880_ (.B2(_0865_),
    .C1(net350),
    .B1(_0593_),
    .A1(_0554_),
    .Y(_0950_),
    .A2(_0584_));
 sg13g2_a221oi_1 _1881_ (.B2(_0593_),
    .C1(net359),
    .B1(_0708_),
    .A1(_0436_),
    .Y(_0951_),
    .A2(_0704_));
 sg13g2_nor3_1 _1882_ (.A(net337),
    .B(_0950_),
    .C(_0951_),
    .Y(_0952_));
 sg13g2_or3_1 _1883_ (.A(net327),
    .B(_0949_),
    .C(_0952_),
    .X(_0953_));
 sg13g2_a21o_1 _1884_ (.A2(_0403_),
    .A1(net397),
    .B1(_0441_),
    .X(_0954_));
 sg13g2_a221oi_1 _1885_ (.B2(net376),
    .C1(net350),
    .B1(_0954_),
    .A1(_0619_),
    .Y(_0955_),
    .A2(_0681_));
 sg13g2_nor2_1 _1886_ (.A(net337),
    .B(_0955_),
    .Y(_0956_));
 sg13g2_o21ai_1 _1887_ (.B1(net352),
    .Y(_0957_),
    .A1(net373),
    .A2(_0630_));
 sg13g2_nor2_1 _1888_ (.A(_0613_),
    .B(_0957_),
    .Y(_0958_));
 sg13g2_and3_1 _1889_ (.X(_0959_),
    .A(net357),
    .B(_0524_),
    .C(_0590_));
 sg13g2_a21oi_1 _1890_ (.A1(_0393_),
    .A2(_0672_),
    .Y(_0960_),
    .B1(_0500_));
 sg13g2_nor4_1 _1891_ (.A(net332),
    .B(_0958_),
    .C(_0959_),
    .D(_0960_),
    .Y(_0961_));
 sg13g2_o21ai_1 _1892_ (.B1(net327),
    .Y(_0962_),
    .A1(_0956_),
    .A2(_0961_));
 sg13g2_nand3_1 _1893_ (.B(_0953_),
    .C(_0962_),
    .A(net326),
    .Y(_0963_));
 sg13g2_nor2_1 _1894_ (.A(_0407_),
    .B(_0553_),
    .Y(_0964_));
 sg13g2_o21ai_1 _1895_ (.B1(net343),
    .Y(_0965_),
    .A1(_0514_),
    .A2(_0964_));
 sg13g2_nand2b_1 _1896_ (.Y(_0966_),
    .B(_0739_),
    .A_N(_0775_));
 sg13g2_nand3_1 _1897_ (.B(_0613_),
    .C(_0749_),
    .A(net351),
    .Y(_0967_));
 sg13g2_nand4_1 _1898_ (.B(_0965_),
    .C(_0966_),
    .A(net336),
    .Y(_0968_),
    .D(_0967_));
 sg13g2_o21ai_1 _1899_ (.B1(net388),
    .Y(_0969_),
    .A1(net405),
    .A2(_0402_));
 sg13g2_a21o_1 _1900_ (.A2(_0969_),
    .A1(_0593_),
    .B1(net363),
    .X(_0970_));
 sg13g2_a22oi_1 _1901_ (.Y(_0971_),
    .B1(_0703_),
    .B2(_0970_),
    .A2(net343),
    .A1(_0427_));
 sg13g2_a21o_1 _1902_ (.A2(_0971_),
    .A1(_0736_),
    .B1(net336),
    .X(_0972_));
 sg13g2_nand3_1 _1903_ (.B(_0968_),
    .C(_0972_),
    .A(net327),
    .Y(_0973_));
 sg13g2_o21ai_1 _1904_ (.B1(_0725_),
    .Y(_0974_),
    .A1(net388),
    .A2(_0502_));
 sg13g2_nand2b_1 _1905_ (.Y(_0975_),
    .B(_0499_),
    .A_N(_0630_));
 sg13g2_a22oi_1 _1906_ (.Y(_0976_),
    .B1(_0846_),
    .B2(net343),
    .A2(_0718_),
    .A1(net351));
 sg13g2_nor4_1 _1907_ (.A(_0400_),
    .B(net357),
    .C(net378),
    .D(_0603_),
    .Y(_0977_));
 sg13g2_nand3_1 _1908_ (.B(_0521_),
    .C(_0640_),
    .A(net374),
    .Y(_0978_));
 sg13g2_a221oi_1 _1909_ (.B2(_0978_),
    .C1(net351),
    .B1(_0799_),
    .A1(_0566_),
    .Y(_0979_),
    .A2(_0670_));
 sg13g2_o21ai_1 _1910_ (.B1(net332),
    .Y(_0980_),
    .A1(_0977_),
    .A2(_0979_));
 sg13g2_nand4_1 _1911_ (.B(_0974_),
    .C(_0975_),
    .A(net336),
    .Y(_0981_),
    .D(_0976_));
 sg13g2_a21o_1 _1912_ (.A2(_0981_),
    .A1(_0980_),
    .B1(net327),
    .X(_0982_));
 sg13g2_a21oi_1 _1913_ (.A1(_0973_),
    .A2(_0982_),
    .Y(_0983_),
    .B1(net326));
 sg13g2_nand3b_1 _1914_ (.B(_0549_),
    .C(_0963_),
    .Y(_0984_),
    .A_N(_0983_));
 sg13g2_or2_1 _1915_ (.X(_0985_),
    .B(\g_x[1] ),
    .A(_0021_));
 sg13g2_nand2_1 _1916_ (.Y(_0986_),
    .A(net343),
    .B(_0862_));
 sg13g2_nand3_1 _1917_ (.B(_0884_),
    .C(_0986_),
    .A(_0881_),
    .Y(_0987_));
 sg13g2_a21oi_1 _1918_ (.A1(net325),
    .A2(_0987_),
    .Y(_0988_),
    .B1(_0985_));
 sg13g2_a21o_1 _1919_ (.A2(_0988_),
    .A1(_0984_),
    .B1(\g_x[2] ),
    .X(_0989_));
 sg13g2_nand4_1 _1920_ (.B(\div3.in[4] ),
    .C(\div3.in[5] ),
    .A(\div3.in[3] ),
    .Y(_0990_),
    .D(net64));
 sg13g2_o21ai_1 _1921_ (.B1(_0990_),
    .Y(_0991_),
    .A1(_0029_),
    .A2(_0218_));
 sg13g2_nor2_1 _1922_ (.A(\hvsync_gen.vpos[9] ),
    .B(_0991_),
    .Y(_0992_));
 sg13g2_o21ai_1 _1923_ (.B1(_0992_),
    .Y(_0993_),
    .A1(_0947_),
    .A2(_0989_));
 sg13g2_nor2_2 _1924_ (.A(net424),
    .B(net427),
    .Y(_0994_));
 sg13g2_nand2b_1 _1925_ (.Y(_0995_),
    .B(_0994_),
    .A_N(_0224_));
 sg13g2_xnor2_1 _1926_ (.Y(_0996_),
    .A(_0225_),
    .B(_0994_));
 sg13g2_mux2_1 _1927_ (.A0(_0017_),
    .A1(_0016_),
    .S(_0222_),
    .X(_0997_));
 sg13g2_a21oi_1 _1928_ (.A1(net424),
    .A2(_0208_),
    .Y(_0998_),
    .B1(_0996_));
 sg13g2_o21ai_1 _1929_ (.B1(_0995_),
    .Y(_0999_),
    .A1(_0223_),
    .A2(_0994_));
 sg13g2_a21oi_1 _1930_ (.A1(_0996_),
    .A2(_0997_),
    .Y(_1000_),
    .B1(_0999_));
 sg13g2_nand2b_1 _1931_ (.Y(_1001_),
    .B(_1000_),
    .A_N(_0998_));
 sg13g2_o21ai_1 _1932_ (.B1(_1001_),
    .Y(_1002_),
    .A1(_0015_),
    .A2(_0995_));
 sg13g2_inv_1 _1933_ (.Y(_1003_),
    .A(_1002_));
 sg13g2_or2_1 _1934_ (.X(_1004_),
    .B(_0995_),
    .A(_0016_));
 sg13g2_nand2_1 _1935_ (.Y(_1005_),
    .A(_0018_),
    .B(_0221_));
 sg13g2_nand2_1 _1936_ (.Y(_1006_),
    .A(_0017_),
    .B(_0222_));
 sg13g2_nand3_1 _1937_ (.B(_1005_),
    .C(_1006_),
    .A(_0996_),
    .Y(_1007_));
 sg13g2_o21ai_1 _1938_ (.B1(_1004_),
    .Y(_1008_),
    .A1(_0999_),
    .A2(_1007_));
 sg13g2_a21oi_1 _1939_ (.A1(_0017_),
    .A2(_0994_),
    .Y(_1009_),
    .B1(_0224_));
 sg13g2_xor2_1 _1940_ (.B(_0225_),
    .A(_0015_),
    .X(_1010_));
 sg13g2_or2_1 _1941_ (.X(_1011_),
    .B(_0995_),
    .A(_0018_));
 sg13g2_o21ai_1 _1942_ (.B1(_1010_),
    .Y(_1012_),
    .A1(_0306_),
    .A2(_1011_));
 sg13g2_a221oi_1 _1943_ (.B2(_0266_),
    .C1(_1012_),
    .B1(_1009_),
    .A1(_0276_),
    .Y(_1013_),
    .A2(_1008_));
 sg13g2_o21ai_1 _1944_ (.B1(_1013_),
    .Y(_1014_),
    .A1(_0284_),
    .A2(_1003_));
 sg13g2_inv_1 _1945_ (.Y(_1015_),
    .A(_1014_));
 sg13g2_xor2_1 _1946_ (.B(_0252_),
    .A(_0251_),
    .X(_1016_));
 sg13g2_inv_1 _1947_ (.Y(_1017_),
    .A(_1016_));
 sg13g2_nand2_1 _1948_ (.Y(_1018_),
    .A(_0208_),
    .B(_1016_));
 sg13g2_o21ai_1 _1949_ (.B1(_1018_),
    .Y(_1019_),
    .A1(_0208_),
    .A2(_0306_));
 sg13g2_inv_1 _1950_ (.Y(_1020_),
    .A(_1019_));
 sg13g2_nor2_1 _1951_ (.A(net425),
    .B(_1019_),
    .Y(_1021_));
 sg13g2_a21oi_2 _1952_ (.B1(_1021_),
    .Y(_1022_),
    .A2(_0277_),
    .A1(net425));
 sg13g2_xnor2_1 _1953_ (.Y(_1023_),
    .A(_0032_),
    .B(_0250_));
 sg13g2_inv_1 _1954_ (.Y(_1024_),
    .A(_1023_));
 sg13g2_a21oi_1 _1955_ (.A1(_0244_),
    .A2(_0245_),
    .Y(_1025_),
    .B1(_0210_));
 sg13g2_nand3_1 _1956_ (.B(_0244_),
    .C(_0245_),
    .A(_0210_),
    .Y(_1026_));
 sg13g2_nor2b_1 _1957_ (.A(_1025_),
    .B_N(_1026_),
    .Y(_1027_));
 sg13g2_nand2b_1 _1958_ (.Y(_1028_),
    .B(_0208_),
    .A_N(_1027_));
 sg13g2_a21oi_1 _1959_ (.A1(net427),
    .A2(_1024_),
    .Y(_1029_),
    .B1(net425));
 sg13g2_a22oi_1 _1960_ (.Y(_1030_),
    .B1(_1028_),
    .B2(_1029_),
    .A2(_1020_),
    .A1(net425));
 sg13g2_and2_1 _1961_ (.A(_1022_),
    .B(_1030_),
    .X(_1031_));
 sg13g2_nor2_1 _1962_ (.A(net1),
    .B(_1031_),
    .Y(_1032_));
 sg13g2_mux4_1 _1963_ (.S0(_0208_),
    .A0(_0265_),
    .A1(_0307_),
    .A2(_1016_),
    .A3(_1024_),
    .S1(_0167_),
    .X(_1033_));
 sg13g2_nor2_1 _1964_ (.A(_1022_),
    .B(_1033_),
    .Y(_1034_));
 sg13g2_or2_1 _1965_ (.X(_1035_),
    .B(_1033_),
    .A(_1022_));
 sg13g2_nor2_1 _1966_ (.A(_1022_),
    .B(_1030_),
    .Y(_1036_));
 sg13g2_nor2_1 _1967_ (.A(_1030_),
    .B(_1033_),
    .Y(_1037_));
 sg13g2_nor2_1 _1968_ (.A(_1030_),
    .B(_1035_),
    .Y(_1038_));
 sg13g2_nand4_1 _1969_ (.B(_1023_),
    .C(_1027_),
    .A(_1017_),
    .Y(_1039_),
    .D(_1038_));
 sg13g2_nand2b_1 _1970_ (.Y(_1040_),
    .B(_1033_),
    .A_N(_1022_));
 sg13g2_o21ai_1 _1971_ (.B1(net2),
    .Y(_1041_),
    .A1(_1032_),
    .A2(_1036_));
 sg13g2_o21ai_1 _1972_ (.B1(_1041_),
    .Y(_1042_),
    .A1(net2),
    .A2(_1040_));
 sg13g2_nor2b_1 _1973_ (.A(_1042_),
    .B_N(_1039_),
    .Y(_1043_));
 sg13g2_nor4_2 _1974_ (.A(_0831_),
    .B(_0993_),
    .C(_1014_),
    .Y(uo_out[6]),
    .D(_1043_));
 sg13g2_nand2_1 _1975_ (.Y(_1044_),
    .A(net2),
    .B(_1039_));
 sg13g2_and2_1 _1976_ (.A(_1022_),
    .B(_1033_),
    .X(_1045_));
 sg13g2_nor2_1 _1977_ (.A(net429),
    .B(_1045_),
    .Y(_1046_));
 sg13g2_nand2_1 _1978_ (.Y(_1047_),
    .A(_1030_),
    .B(_1033_));
 sg13g2_nor2_1 _1979_ (.A(_1034_),
    .B(_1036_),
    .Y(_1048_));
 sg13g2_nand2b_1 _1980_ (.Y(_1049_),
    .B(_1048_),
    .A_N(_1046_));
 sg13g2_a22oi_1 _1981_ (.Y(_1050_),
    .B1(_1049_),
    .B2(net2),
    .A2(_1044_),
    .A1(_1034_));
 sg13g2_nor4_2 _1982_ (.A(_0831_),
    .B(_0993_),
    .C(_1014_),
    .Y(uo_out[2]),
    .D(_1050_));
 sg13g2_nor2_1 _1983_ (.A(_1037_),
    .B(_1048_),
    .Y(_1051_));
 sg13g2_a21oi_1 _1984_ (.A1(net429),
    .A2(_1051_),
    .Y(_1052_),
    .B1(_1032_));
 sg13g2_o21ai_1 _1985_ (.B1(_1039_),
    .Y(_1053_),
    .A1(net2),
    .A2(_1052_));
 sg13g2_a21oi_1 _1986_ (.A1(net429),
    .A2(_1030_),
    .Y(_1054_),
    .B1(_0204_));
 sg13g2_o21ai_1 _1987_ (.B1(_1022_),
    .Y(_1055_),
    .A1(_0203_),
    .A2(_1033_));
 sg13g2_and3_1 _1988_ (.X(_1056_),
    .A(_1035_),
    .B(_1054_),
    .C(_1055_));
 sg13g2_o21ai_1 _1989_ (.B1(_1015_),
    .Y(_1057_),
    .A1(_1053_),
    .A2(_1056_));
 sg13g2_nor3_2 _1990_ (.A(_0831_),
    .B(_0993_),
    .C(_1057_),
    .Y(uo_out[5]));
 sg13g2_or2_1 _1991_ (.X(_1058_),
    .B(_1046_),
    .A(_1038_));
 sg13g2_nor2_1 _1992_ (.A(_0203_),
    .B(_1045_),
    .Y(_1059_));
 sg13g2_nand2_1 _1993_ (.Y(_1060_),
    .A(_1048_),
    .B(_1059_));
 sg13g2_o21ai_1 _1994_ (.B1(_1060_),
    .Y(_1061_),
    .A1(net429),
    .A2(_1035_));
 sg13g2_a22oi_1 _1995_ (.Y(_1062_),
    .B1(_1061_),
    .B2(net2),
    .A2(_1058_),
    .A1(_1044_));
 sg13g2_nor4_2 _1996_ (.A(_0831_),
    .B(_0993_),
    .C(_1014_),
    .Y(uo_out[1]),
    .D(_1062_));
 sg13g2_o21ai_1 _1997_ (.B1(_1031_),
    .Y(_1063_),
    .A1(_0204_),
    .A2(_1033_));
 sg13g2_o21ai_1 _1998_ (.B1(_1063_),
    .Y(_1064_),
    .A1(_0204_),
    .A2(_1022_));
 sg13g2_nand3b_1 _1999_ (.B(_1064_),
    .C(net429),
    .Y(_1065_),
    .A_N(_1037_));
 sg13g2_o21ai_1 _2000_ (.B1(_1065_),
    .Y(_1066_),
    .A1(net429),
    .A2(_1051_));
 sg13g2_a21o_1 _2001_ (.A2(_1066_),
    .A1(_1039_),
    .B1(_1014_),
    .X(_1067_));
 sg13g2_nor3_2 _2002_ (.A(_0831_),
    .B(_0993_),
    .C(_1067_),
    .Y(uo_out[4]));
 sg13g2_nand4_1 _2003_ (.B(net2),
    .C(_1040_),
    .A(net429),
    .Y(_1068_),
    .D(_1047_));
 sg13g2_a22oi_1 _2004_ (.Y(_1069_),
    .B1(_1059_),
    .B2(_0204_),
    .A2(_1038_),
    .A1(_0203_));
 sg13g2_nand3_1 _2005_ (.B(_1068_),
    .C(_1069_),
    .A(_1039_),
    .Y(_1070_));
 sg13g2_nand2_1 _2006_ (.Y(_1071_),
    .A(_1015_),
    .B(_1070_));
 sg13g2_nor3_2 _2007_ (.A(_0831_),
    .B(_0993_),
    .C(_1071_),
    .Y(uo_out[0]));
 sg13g2_nor3_2 _2008_ (.A(_0189_),
    .B(_0197_),
    .C(_0202_),
    .Y(_1072_));
 sg13g2_and2_1 _2009_ (.A(net428),
    .B(_1072_),
    .X(_1073_));
 sg13g2_nand2_1 _2010_ (.Y(_1074_),
    .A(net428),
    .B(_1072_));
 sg13g2_nor2_2 _2011_ (.A(_0167_),
    .B(_1074_),
    .Y(_1075_));
 sg13g2_nor3_1 _2012_ (.A(net423),
    .B(\hvsync_gen.hpos[6] ),
    .C(\hvsync_gen.hpos[7] ),
    .Y(_1076_));
 sg13g2_nand4_1 _2013_ (.B(\hvsync_gen.hpos[8] ),
    .C(_1075_),
    .A(\hvsync_gen.hpos[9] ),
    .Y(_1077_),
    .D(_1076_));
 sg13g2_and2_1 _2014_ (.A(net431),
    .B(_1077_),
    .X(_1078_));
 sg13g2_nand2_2 _2015_ (.Y(_0066_),
    .A(net431),
    .B(_1077_));
 sg13g2_nor4_1 _2016_ (.A(\div3.in[4] ),
    .B(_0206_),
    .C(\div3.in[5] ),
    .D(\div3.in[6] ),
    .Y(_0067_));
 sg13g2_nor3_1 _2017_ (.A(\div3.in[2] ),
    .B(\div3.in[3] ),
    .C(_0390_),
    .Y(_0068_));
 sg13g2_nand4_1 _2018_ (.B(\div3.in[0] ),
    .C(_0067_),
    .A(\div3.in[1] ),
    .Y(_0069_),
    .D(_0068_));
 sg13g2_nand2_1 _2019_ (.Y(_0070_),
    .A(net430),
    .B(_0069_));
 sg13g2_nor2_2 _2020_ (.A(_1077_),
    .B(_0070_),
    .Y(_0071_));
 sg13g2_or2_2 _2021_ (.X(_0072_),
    .B(_0070_),
    .A(_1077_));
 sg13g2_nand3_1 _2022_ (.B(\div3.in[0] ),
    .C(_0383_),
    .A(\div3.in[1] ),
    .Y(_0073_));
 sg13g2_nor2_1 _2023_ (.A(_0205_),
    .B(_0073_),
    .Y(_0074_));
 sg13g2_nand4_1 _2024_ (.B(\div3.in[4] ),
    .C(\div3.in[5] ),
    .A(\div3.in[3] ),
    .Y(_0075_),
    .D(_0074_));
 sg13g2_xor2_1 _2025_ (.B(_0075_),
    .A(_0008_),
    .X(_0076_));
 sg13g2_nand2_1 _2026_ (.Y(_0077_),
    .A(_0071_),
    .B(_0076_));
 sg13g2_o21ai_1 _2027_ (.B1(_0077_),
    .Y(_0078_),
    .A1(_0008_),
    .A2(_0066_));
 sg13g2_nand2_1 _2028_ (.Y(_0079_),
    .A(\div3.in[3] ),
    .B(_0074_));
 sg13g2_nor2_1 _2029_ (.A(_0009_),
    .B(_0079_),
    .Y(_0080_));
 sg13g2_a21o_1 _2030_ (.A2(_0080_),
    .A1(_0066_),
    .B1(\div3.in[5] ),
    .X(_0081_));
 sg13g2_nand2_1 _2031_ (.Y(_0082_),
    .A(_0066_),
    .B(_0070_));
 sg13g2_nand3_1 _2032_ (.B(_0066_),
    .C(_0080_),
    .A(\div3.in[5] ),
    .Y(_0083_));
 sg13g2_nand3_1 _2033_ (.B(_0082_),
    .C(_0083_),
    .A(_0081_),
    .Y(_0084_));
 sg13g2_inv_1 _2034_ (.Y(_0062_),
    .A(_0084_));
 sg13g2_nand2_1 _2035_ (.Y(_0085_),
    .A(net84),
    .B(net413));
 sg13g2_xnor2_1 _2036_ (.Y(_0086_),
    .A(_0009_),
    .B(_0079_));
 sg13g2_o21ai_1 _2037_ (.B1(_0085_),
    .Y(_0061_),
    .A1(_0072_),
    .A2(_0086_));
 sg13g2_inv_1 _2038_ (.Y(_0087_),
    .A(net411));
 sg13g2_nand2_1 _2039_ (.Y(_0088_),
    .A(\div3.in[2] ),
    .B(net413));
 sg13g2_nor2_1 _2040_ (.A(_0011_),
    .B(_0073_),
    .Y(_0089_));
 sg13g2_xnor2_1 _2041_ (.Y(_0090_),
    .A(_0011_),
    .B(_0073_));
 sg13g2_o21ai_1 _2042_ (.B1(_0088_),
    .Y(_0059_),
    .A1(_0072_),
    .A2(_0090_));
 sg13g2_inv_1 _2043_ (.Y(_0091_),
    .A(_0059_));
 sg13g2_nand2_1 _2044_ (.Y(_0092_),
    .A(net73),
    .B(net413));
 sg13g2_nor2_1 _2045_ (.A(_0013_),
    .B(net416),
    .Y(_0093_));
 sg13g2_xor2_1 _2046_ (.B(_0093_),
    .A(net89),
    .X(_0094_));
 sg13g2_o21ai_1 _2047_ (.B1(_0092_),
    .Y(_0058_),
    .A1(_0072_),
    .A2(net90));
 sg13g2_nand2_1 _2048_ (.Y(_0095_),
    .A(\div3.in[0] ),
    .B(net413));
 sg13g2_xnor2_1 _2049_ (.Y(_0096_),
    .A(net78),
    .B(net416));
 sg13g2_o21ai_1 _2050_ (.B1(_0095_),
    .Y(_0057_),
    .A1(_0072_),
    .A2(_0096_));
 sg13g2_nand2_1 _2051_ (.Y(_0097_),
    .A(_0058_),
    .B(_0057_));
 sg13g2_nand2_1 _2052_ (.Y(_0098_),
    .A(_0091_),
    .B(_0097_));
 sg13g2_nand2_1 _2053_ (.Y(_0099_),
    .A(\div3.in[3] ),
    .B(net413));
 sg13g2_xor2_1 _2054_ (.B(_0089_),
    .A(_0010_),
    .X(_0100_));
 sg13g2_o21ai_1 _2055_ (.B1(_0099_),
    .Y(_0060_),
    .A1(_0072_),
    .A2(_0100_));
 sg13g2_inv_1 _2056_ (.Y(_0101_),
    .A(net410));
 sg13g2_a21oi_1 _2057_ (.A1(_0059_),
    .A2(_0058_),
    .Y(_0102_),
    .B1(net410));
 sg13g2_inv_1 _2058_ (.Y(_0103_),
    .A(_0102_));
 sg13g2_nor2_1 _2059_ (.A(_0058_),
    .B(_0057_),
    .Y(_0104_));
 sg13g2_a21oi_1 _2060_ (.A1(_0059_),
    .A2(_0097_),
    .Y(_0105_),
    .B1(_0104_));
 sg13g2_a22oi_1 _2061_ (.Y(_0106_),
    .B1(_0105_),
    .B2(_0060_),
    .A2(_0102_),
    .A1(_0098_));
 sg13g2_nor2_1 _2062_ (.A(net411),
    .B(_0106_),
    .Y(_0107_));
 sg13g2_a21oi_1 _2063_ (.A1(_0059_),
    .A2(_0058_),
    .Y(_0108_),
    .B1(_0101_));
 sg13g2_or2_1 _2064_ (.X(_0109_),
    .B(_0058_),
    .A(_0059_));
 sg13g2_inv_1 _2065_ (.Y(_0110_),
    .A(_0109_));
 sg13g2_o21ai_1 _2066_ (.B1(_0109_),
    .Y(_0111_),
    .A1(_0091_),
    .A2(_0104_));
 sg13g2_a22oi_1 _2067_ (.Y(_0112_),
    .B1(_0111_),
    .B2(_0101_),
    .A2(_0108_),
    .A1(_0098_));
 sg13g2_nor2_1 _2068_ (.A(_0087_),
    .B(_0112_),
    .Y(_0113_));
 sg13g2_nor2_1 _2069_ (.A(_0107_),
    .B(_0113_),
    .Y(_0114_));
 sg13g2_nor2_1 _2070_ (.A(_0062_),
    .B(_0114_),
    .Y(_0115_));
 sg13g2_and2_1 _2071_ (.A(_0101_),
    .B(_0105_),
    .X(_0116_));
 sg13g2_a21oi_1 _2072_ (.A1(_0060_),
    .A2(_0111_),
    .Y(_0117_),
    .B1(_0116_));
 sg13g2_nor3_1 _2073_ (.A(_0084_),
    .B(net411),
    .C(_0117_),
    .Y(_0118_));
 sg13g2_nor2_1 _2074_ (.A(_0084_),
    .B(_0087_),
    .Y(_0119_));
 sg13g2_nor2b_1 _2075_ (.A(_0106_),
    .B_N(_0119_),
    .Y(_0120_));
 sg13g2_nor3_1 _2076_ (.A(_0115_),
    .B(_0118_),
    .C(_0120_),
    .Y(_0121_));
 sg13g2_a21oi_1 _2077_ (.A1(net411),
    .A2(_0111_),
    .Y(_0122_),
    .B1(_0107_));
 sg13g2_nand2_1 _2078_ (.Y(_0123_),
    .A(_0078_),
    .B(_0062_));
 sg13g2_inv_1 _2079_ (.Y(_0065_),
    .A(_0123_));
 sg13g2_nor2_1 _2080_ (.A(_0122_),
    .B(_0123_),
    .Y(_0124_));
 sg13g2_and2_1 _2081_ (.A(_0078_),
    .B(_0084_),
    .X(_0125_));
 sg13g2_nand2_1 _2082_ (.Y(_0126_),
    .A(_0078_),
    .B(_0084_));
 sg13g2_nand2_1 _2083_ (.Y(_0127_),
    .A(_0087_),
    .B(_0125_));
 sg13g2_nor2_1 _2084_ (.A(_0112_),
    .B(_0127_),
    .Y(_0128_));
 sg13g2_nand2_1 _2085_ (.Y(_0129_),
    .A(net411),
    .B(_0125_));
 sg13g2_nor2_1 _2086_ (.A(_0117_),
    .B(_0129_),
    .Y(_0130_));
 sg13g2_nor3_1 _2087_ (.A(_0124_),
    .B(_0128_),
    .C(_0130_),
    .Y(_0131_));
 sg13g2_o21ai_1 _2088_ (.B1(_0131_),
    .Y(_0000_),
    .A1(_0078_),
    .A2(_0121_));
 sg13g2_a21oi_2 _2089_ (.B1(net412),
    .Y(_0132_),
    .A2(net410),
    .A1(_0059_));
 sg13g2_a22oi_1 _2090_ (.Y(_0133_),
    .B1(_0132_),
    .B2(_0103_),
    .A2(_0109_),
    .A1(net412));
 sg13g2_nor2b_1 _2091_ (.A(_0132_),
    .B_N(_0108_),
    .Y(_0134_));
 sg13g2_nor3_1 _2092_ (.A(_0062_),
    .B(_0133_),
    .C(_0134_),
    .Y(_0135_));
 sg13g2_o21ai_1 _2093_ (.B1(net412),
    .Y(_0136_),
    .A1(_0091_),
    .A2(_0101_));
 sg13g2_nor3_1 _2094_ (.A(_0084_),
    .B(_0102_),
    .C(_0136_),
    .Y(_0137_));
 sg13g2_nor2_1 _2095_ (.A(_0059_),
    .B(net410),
    .Y(_0138_));
 sg13g2_a21oi_1 _2096_ (.A1(net410),
    .A2(_0109_),
    .Y(_0139_),
    .B1(_0138_));
 sg13g2_nor3_1 _2097_ (.A(_0084_),
    .B(net411),
    .C(_0139_),
    .Y(_0140_));
 sg13g2_nor3_1 _2098_ (.A(_0135_),
    .B(_0137_),
    .C(_0140_),
    .Y(_0141_));
 sg13g2_nor3_1 _2099_ (.A(_0108_),
    .B(_0110_),
    .C(_0127_),
    .Y(_0142_));
 sg13g2_nor2_1 _2100_ (.A(_0123_),
    .B(_0133_),
    .Y(_0143_));
 sg13g2_nor2_1 _2101_ (.A(_0129_),
    .B(_0139_),
    .Y(_0144_));
 sg13g2_nor3_1 _2102_ (.A(_0142_),
    .B(_0143_),
    .C(_0144_),
    .Y(_0145_));
 sg13g2_o21ai_1 _2103_ (.B1(_0145_),
    .Y(_0001_),
    .A1(_0078_),
    .A2(_0141_));
 sg13g2_or2_1 _2104_ (.X(_0146_),
    .B(_0084_),
    .A(_0078_));
 sg13g2_nand2b_1 _2105_ (.Y(_0147_),
    .B(_0136_),
    .A_N(_0146_));
 sg13g2_a21oi_1 _2106_ (.A1(_0129_),
    .A2(_0147_),
    .Y(_0148_),
    .B1(_0138_));
 sg13g2_a21oi_1 _2107_ (.A1(net411),
    .A2(net410),
    .Y(_0149_),
    .B1(_0062_));
 sg13g2_or2_1 _2108_ (.X(_0150_),
    .B(_0149_),
    .A(_0078_));
 sg13g2_nand2b_1 _2109_ (.Y(_0151_),
    .B(_0150_),
    .A_N(_0132_));
 sg13g2_nand2_1 _2110_ (.Y(_0152_),
    .A(_0126_),
    .B(_0151_));
 sg13g2_o21ai_1 _2111_ (.B1(_0125_),
    .Y(_0153_),
    .A1(net411),
    .A2(net410));
 sg13g2_a21o_1 _2112_ (.A2(_0153_),
    .A1(_0152_),
    .B1(_0148_),
    .X(_0002_));
 sg13g2_o21ai_1 _2113_ (.B1(_0153_),
    .Y(_0003_),
    .A1(_0119_),
    .A2(_0150_));
 sg13g2_o21ai_1 _2114_ (.B1(_0126_),
    .Y(_0004_),
    .A1(_0087_),
    .A2(_0146_));
 sg13g2_nor3_1 _2115_ (.A(\div3.in[0] ),
    .B(\div3.in[2] ),
    .C(net62),
    .Y(_0154_));
 sg13g2_nand3_1 _2116_ (.B(net73),
    .C(_0154_),
    .A(net419),
    .Y(_0155_));
 sg13g2_nor2_1 _2117_ (.A(_0990_),
    .B(net74),
    .Y(_0006_));
 sg13g2_nand3_1 _2118_ (.B(net423),
    .C(\hvsync_gen.hpos[6] ),
    .A(net426),
    .Y(_0156_));
 sg13g2_a21oi_1 _2119_ (.A1(_0182_),
    .A2(_0156_),
    .Y(_0157_),
    .B1(net68));
 sg13g2_nor3_1 _2120_ (.A(\hvsync_gen.hpos[8] ),
    .B(net423),
    .C(_0224_),
    .Y(_0158_));
 sg13g2_nor4_1 _2121_ (.A(_0175_),
    .B(_0218_),
    .C(net69),
    .D(_0158_),
    .Y(_0005_));
 sg13g2_and2_1 _2122_ (.A(net430),
    .B(_0028_),
    .X(_0035_));
 sg13g2_o21ai_1 _2123_ (.B1(net430),
    .Y(_0159_),
    .A1(\counter[1] ),
    .A2(\counter[0] ));
 sg13g2_a21oi_1 _2124_ (.A1(\counter[1] ),
    .A2(\counter[0] ),
    .Y(_0036_),
    .B1(_0159_));
 sg13g2_a21oi_1 _2125_ (.A1(\counter[1] ),
    .A2(\counter[0] ),
    .Y(_0160_),
    .B1(\counter[2] ));
 sg13g2_nand3_1 _2126_ (.B(\counter[0] ),
    .C(\counter[2] ),
    .A(\counter[1] ),
    .Y(_0161_));
 sg13g2_nand2_1 _2127_ (.Y(_0162_),
    .A(net430),
    .B(_0161_));
 sg13g2_nor2_1 _2128_ (.A(_0160_),
    .B(_0162_),
    .Y(_0037_));
 sg13g2_nor2_1 _2129_ (.A(_0207_),
    .B(_0161_),
    .Y(_0163_));
 sg13g2_o21ai_1 _2130_ (.B1(net430),
    .Y(_0164_),
    .A1(_0207_),
    .A2(_0161_));
 sg13g2_a21oi_1 _2131_ (.A1(_0207_),
    .A2(_0161_),
    .Y(_0038_),
    .B1(_0164_));
 sg13g2_o21ai_1 _2132_ (.B1(net430),
    .Y(_0165_),
    .A1(\counter[4] ),
    .A2(_0163_));
 sg13g2_a21oi_1 _2133_ (.A1(\counter[4] ),
    .A2(_0163_),
    .Y(_0039_),
    .B1(_0165_));
 sg13g2_nor3_1 _2134_ (.A(_0207_),
    .B(_0026_),
    .C(_0161_),
    .Y(_0166_));
 sg13g2_o21ai_1 _2135_ (.B1(net430),
    .Y(_0168_),
    .A1(\counter[5] ),
    .A2(_0166_));
 sg13g2_a21oi_1 _2136_ (.A1(\counter[5] ),
    .A2(_0166_),
    .Y(_0040_),
    .B1(_0168_));
 sg13g2_nand3_1 _2137_ (.B(\counter[5] ),
    .C(_0163_),
    .A(\counter[4] ),
    .Y(_0169_));
 sg13g2_inv_1 _2138_ (.Y(_0170_),
    .A(_0169_));
 sg13g2_and2_1 _2139_ (.A(\counter[6] ),
    .B(_0170_),
    .X(_0171_));
 sg13g2_o21ai_1 _2140_ (.B1(net430),
    .Y(_0172_),
    .A1(\counter[6] ),
    .A2(_0170_));
 sg13g2_nor2_1 _2141_ (.A(_0171_),
    .B(_0172_),
    .Y(_0041_));
 sg13g2_nor2_1 _2142_ (.A(_0024_),
    .B(_0169_),
    .Y(_0173_));
 sg13g2_o21ai_1 _2143_ (.B1(net431),
    .Y(_0174_),
    .A1(\counter[7] ),
    .A2(_0173_));
 sg13g2_a21oi_1 _2144_ (.A1(\counter[7] ),
    .A2(_0173_),
    .Y(_0042_),
    .B1(_0174_));
 sg13g2_and2_1 _2145_ (.A(\counter[7] ),
    .B(_0171_),
    .X(_0176_));
 sg13g2_o21ai_1 _2146_ (.B1(net431),
    .Y(_0177_),
    .A1(\counter[8] ),
    .A2(_0176_));
 sg13g2_a21oi_1 _2147_ (.A1(\counter[8] ),
    .A2(_0176_),
    .Y(_0043_),
    .B1(_0177_));
 sg13g2_nor2b_1 _2148_ (.A(_0022_),
    .B_N(_0176_),
    .Y(_0178_));
 sg13g2_o21ai_1 _2149_ (.B1(net431),
    .Y(_0179_),
    .A1(\counter[9] ),
    .A2(_0178_));
 sg13g2_a21oi_1 _2150_ (.A1(\counter[9] ),
    .A2(_0178_),
    .Y(_0044_),
    .B1(_0179_));
 sg13g2_and2_1 _2151_ (.A(net57),
    .B(net414),
    .X(_0045_));
 sg13g2_o21ai_1 _2152_ (.B1(net414),
    .Y(_0180_),
    .A1(\g_x[0] ),
    .A2(net66));
 sg13g2_a21oi_1 _2153_ (.A1(\g_x[0] ),
    .A2(net66),
    .Y(_0046_),
    .B1(_0180_));
 sg13g2_a21oi_1 _2154_ (.A1(\g_x[0] ),
    .A2(\g_x[1] ),
    .Y(_0181_),
    .B1(net60));
 sg13g2_nor3_1 _2155_ (.A(_1072_),
    .B(_0066_),
    .C(net61),
    .Y(_0047_));
 sg13g2_o21ai_1 _2156_ (.B1(net431),
    .Y(_0183_),
    .A1(net428),
    .A2(_1072_));
 sg13g2_nor2_1 _2157_ (.A(_1073_),
    .B(_0183_),
    .Y(_0048_));
 sg13g2_o21ai_1 _2158_ (.B1(net431),
    .Y(_0184_),
    .A1(net426),
    .A2(_1073_));
 sg13g2_nor2_1 _2159_ (.A(_1075_),
    .B(_0184_),
    .Y(_0049_));
 sg13g2_nor2_1 _2160_ (.A(_0019_),
    .B(_1074_),
    .Y(_0185_));
 sg13g2_xnor2_1 _2161_ (.Y(_0186_),
    .A(net423),
    .B(_0185_));
 sg13g2_nor2_1 _2162_ (.A(_0066_),
    .B(net88),
    .Y(_0050_));
 sg13g2_nand2_1 _2163_ (.Y(_0187_),
    .A(net424),
    .B(_1075_));
 sg13g2_a21oi_1 _2164_ (.A1(net423),
    .A2(_1075_),
    .Y(_0188_),
    .B1(net80));
 sg13g2_nor2_1 _2165_ (.A(_1074_),
    .B(_0156_),
    .Y(_0190_));
 sg13g2_nor3_1 _2166_ (.A(_0066_),
    .B(net81),
    .C(_0190_),
    .Y(_0051_));
 sg13g2_nor2_1 _2167_ (.A(net71),
    .B(_0187_),
    .Y(_0191_));
 sg13g2_o21ai_1 _2168_ (.B1(net414),
    .Y(_0192_),
    .A1(\hvsync_gen.hpos[7] ),
    .A2(_0191_));
 sg13g2_a21oi_1 _2169_ (.A1(\hvsync_gen.hpos[7] ),
    .A2(_0191_),
    .Y(_0052_),
    .B1(_0192_));
 sg13g2_nand2_1 _2170_ (.Y(_0193_),
    .A(\hvsync_gen.hpos[7] ),
    .B(_0190_));
 sg13g2_o21ai_1 _2171_ (.B1(net414),
    .Y(_0194_),
    .A1(_0182_),
    .A2(_0193_));
 sg13g2_a21oi_1 _2172_ (.A1(_0182_),
    .A2(_0193_),
    .Y(_0053_),
    .B1(_0194_));
 sg13g2_nor2_1 _2173_ (.A(_0015_),
    .B(_0193_),
    .Y(_0195_));
 sg13g2_o21ai_1 _2174_ (.B1(net414),
    .Y(_0196_),
    .A1(net76),
    .A2(_0195_));
 sg13g2_a21oi_1 _2175_ (.A1(net76),
    .A2(_0195_),
    .Y(_0054_),
    .B1(_0196_));
 sg13g2_a22oi_1 _2176_ (.Y(_0198_),
    .B1(_0071_),
    .B2(net58),
    .A2(net413),
    .A1(net421));
 sg13g2_inv_1 _2177_ (.Y(_0055_),
    .A(net59));
 sg13g2_a22oi_1 _2178_ (.Y(_0199_),
    .B1(_0071_),
    .B2(_0408_),
    .A2(net413),
    .A1(net419));
 sg13g2_inv_1 _2179_ (.Y(_0056_),
    .A(_0199_));
 sg13g2_o21ai_1 _2180_ (.B1(_0077_),
    .Y(_0063_),
    .A1(_0209_),
    .A2(_0066_));
 sg13g2_nor3_1 _2181_ (.A(_0008_),
    .B(net413),
    .C(_0075_),
    .Y(_0200_));
 sg13g2_o21ai_1 _2182_ (.B1(_0082_),
    .Y(_0201_),
    .A1(net62),
    .A2(_0200_));
 sg13g2_a21oi_1 _2183_ (.A1(net62),
    .A2(_0200_),
    .Y(_0064_),
    .B1(_0201_));
 sg13g2_dfrbp_1 _2184_ (.CLK(net417),
    .RESET_B(net39),
    .D(_0035_),
    .Q_N(_0028_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _2185_ (.CLK(net417),
    .RESET_B(net46),
    .D(_0036_),
    .Q_N(_1087_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _2186_ (.CLK(net417),
    .RESET_B(net45),
    .D(_0037_),
    .Q_N(_1086_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _2187_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net44),
    .D(_0038_),
    .Q_N(_0027_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _2188_ (.CLK(net417),
    .RESET_B(net43),
    .D(_0039_),
    .Q_N(_0026_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _2189_ (.CLK(net417),
    .RESET_B(net42),
    .D(_0040_),
    .Q_N(_0025_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _2190_ (.CLK(net417),
    .RESET_B(net41),
    .D(_0041_),
    .Q_N(_0024_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _2191_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net40),
    .D(_0042_),
    .Q_N(_0023_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _2192_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net38),
    .D(_0043_),
    .Q_N(_0022_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _2193_ (.CLK(net417),
    .RESET_B(net37),
    .D(_0044_),
    .Q_N(_1085_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 _2194_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net36),
    .D(_0045_),
    .Q_N(_0021_),
    .Q(\g_x[0] ));
 sg13g2_dfrbp_1 _2195_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net35),
    .D(net67),
    .Q_N(_1084_),
    .Q(\g_x[1] ));
 sg13g2_dfrbp_1 _2196_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net34),
    .D(_0047_),
    .Q_N(_1083_),
    .Q(\g_x[2] ));
 sg13g2_dfrbp_1 _2197_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net33),
    .D(_0048_),
    .Q_N(_0020_),
    .Q(\a[0] ));
 sg13g2_dfrbp_1 _2198_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net32),
    .D(_0049_),
    .Q_N(_0019_),
    .Q(\a[1] ));
 sg13g2_dfrbp_1 _2199_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net31),
    .D(_0050_),
    .Q_N(_0018_),
    .Q(b));
 sg13g2_dfrbp_1 _2200_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net30),
    .D(_0051_),
    .Q_N(_0017_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _2201_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net29),
    .D(net72),
    .Q_N(_0016_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _2202_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net28),
    .D(net83),
    .Q_N(_0015_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _2203_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net50),
    .D(net77),
    .Q_N(_0029_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _2204_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net27),
    .D(net70),
    .Q_N(_1082_),
    .Q(hsync));
 sg13g2_dfrbp_1 _2205_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net26),
    .D(_0055_),
    .Q_N(_0014_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _2206_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net24),
    .D(_0056_),
    .Q_N(_1081_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _2207_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net22),
    .D(net79),
    .Q_N(_0013_),
    .Q(\div3.in[0] ));
 sg13g2_dfrbp_1 _2208_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net20),
    .D(_0058_),
    .Q_N(_0012_),
    .Q(\div3.in[1] ));
 sg13g2_dfrbp_1 _2209_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net51),
    .D(_0059_),
    .Q_N(_0011_),
    .Q(\div3.in[2] ));
 sg13g2_dfrbp_1 _2210_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net48),
    .D(net410),
    .Q_N(_0010_),
    .Q(\div3.in[3] ));
 sg13g2_dfrbp_1 _2211_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net25),
    .D(net412),
    .Q_N(_0009_),
    .Q(\div3.in[4] ));
 sg13g2_dfrbp_1 _2212_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net21),
    .D(_0062_),
    .Q_N(_1080_),
    .Q(\div3.in[5] ));
 sg13g2_dfrbp_1 _2213_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net49),
    .D(net65),
    .Q_N(_0008_),
    .Q(\div3.in[6] ));
 sg13g2_dfrbp_1 _2214_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net52),
    .D(net63),
    .Q_N(_1088_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _2215_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net23),
    .D(net75),
    .Q_N(_1079_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 _2216_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net53),
    .D(_0065_),
    .Q_N(_0030_),
    .Q(\div3.out[5] ));
 sg13g2_dfrbp_1 _2217_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net54),
    .D(_0000_),
    .Q_N(_0031_),
    .Q(\div3.out[0] ));
 sg13g2_dfrbp_1 _2218_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net55),
    .D(_0001_),
    .Q_N(_0032_),
    .Q(\div3.out[1] ));
 sg13g2_dfrbp_1 _2219_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net56),
    .D(_0002_),
    .Q_N(_0033_),
    .Q(\div3.out[2] ));
 sg13g2_dfrbp_1 _2220_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net19),
    .D(_0003_),
    .Q_N(_0034_),
    .Q(\div3.out[3] ));
 sg13g2_dfrbp_1 _2221_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net47),
    .D(_0004_),
    .Q_N(_0007_),
    .Q(\div3.out[4] ));
 sg13g2_tiehi _2208__20 (.L_HI(net20));
 sg13g2_tiehi _2212__21 (.L_HI(net21));
 sg13g2_tiehi _2207__22 (.L_HI(net22));
 sg13g2_tiehi _2215__23 (.L_HI(net23));
 sg13g2_tiehi _2206__24 (.L_HI(net24));
 sg13g2_tiehi _2211__25 (.L_HI(net25));
 sg13g2_tiehi _2205__26 (.L_HI(net26));
 sg13g2_tiehi _2204__27 (.L_HI(net27));
 sg13g2_tiehi _2202__28 (.L_HI(net28));
 sg13g2_tiehi _2201__29 (.L_HI(net29));
 sg13g2_tiehi _2200__30 (.L_HI(net30));
 sg13g2_tiehi _2199__31 (.L_HI(net31));
 sg13g2_tiehi _2198__32 (.L_HI(net32));
 sg13g2_tiehi _2197__33 (.L_HI(net33));
 sg13g2_tiehi _2196__34 (.L_HI(net34));
 sg13g2_tiehi _2195__35 (.L_HI(net35));
 sg13g2_tiehi _2194__36 (.L_HI(net36));
 sg13g2_tiehi _2193__37 (.L_HI(net37));
 sg13g2_tiehi _2192__38 (.L_HI(net38));
 sg13g2_tiehi _2184__39 (.L_HI(net39));
 sg13g2_tiehi _2191__40 (.L_HI(net40));
 sg13g2_tiehi _2190__41 (.L_HI(net41));
 sg13g2_tiehi _2189__42 (.L_HI(net42));
 sg13g2_tiehi _2188__43 (.L_HI(net43));
 sg13g2_tiehi _2187__44 (.L_HI(net44));
 sg13g2_tiehi _2186__45 (.L_HI(net45));
 sg13g2_tiehi _2185__46 (.L_HI(net46));
 sg13g2_tiehi _2221__47 (.L_HI(net47));
 sg13g2_tiehi _2210__48 (.L_HI(net48));
 sg13g2_tiehi _2213__49 (.L_HI(net49));
 sg13g2_tiehi _2203__50 (.L_HI(net50));
 sg13g2_tiehi _2209__51 (.L_HI(net51));
 sg13g2_tiehi _2214__52 (.L_HI(net52));
 sg13g2_tiehi _2216__53 (.L_HI(net53));
 sg13g2_tiehi _2217__54 (.L_HI(net54));
 sg13g2_tiehi _2218__55 (.L_HI(net55));
 sg13g2_tiehi _2219__56 (.L_HI(net56));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_vga_glyph_mode_4 (.L_LO(net4));
 sg13g2_tielo tt_um_vga_glyph_mode_5 (.L_LO(net5));
 sg13g2_tielo tt_um_vga_glyph_mode_6 (.L_LO(net6));
 sg13g2_tielo tt_um_vga_glyph_mode_7 (.L_LO(net7));
 sg13g2_tielo tt_um_vga_glyph_mode_8 (.L_LO(net8));
 sg13g2_tielo tt_um_vga_glyph_mode_9 (.L_LO(net9));
 sg13g2_tielo tt_um_vga_glyph_mode_10 (.L_LO(net10));
 sg13g2_tielo tt_um_vga_glyph_mode_11 (.L_LO(net11));
 sg13g2_tielo tt_um_vga_glyph_mode_12 (.L_LO(net12));
 sg13g2_tielo tt_um_vga_glyph_mode_13 (.L_LO(net13));
 sg13g2_tielo tt_um_vga_glyph_mode_14 (.L_LO(net14));
 sg13g2_tielo tt_um_vga_glyph_mode_15 (.L_LO(net15));
 sg13g2_tielo tt_um_vga_glyph_mode_16 (.L_LO(net16));
 sg13g2_tielo tt_um_vga_glyph_mode_17 (.L_LO(net17));
 sg13g2_tielo tt_um_vga_glyph_mode_18 (.L_LO(net18));
 sg13g2_tiehi _2220__19 (.L_HI(net19));
 sg13g2_buf_1 _2276_ (.A(net417),
    .X(uo_out[3]));
 sg13g2_buf_1 _2277_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout325 (.A(_0550_),
    .X(net325));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(_0498_));
 sg13g2_buf_2 fanout327 (.A(net328),
    .X(net327));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(_0455_));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(_0454_));
 sg13g2_buf_2 fanout330 (.A(_0454_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_0380_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(net333),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_0380_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(net339),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(net339),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(net338),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(net338),
    .X(net337));
 sg13g2_buf_1 fanout338 (.A(net339),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_0379_),
    .X(net339));
 sg13g2_buf_4 fanout340 (.X(net340),
    .A(net341));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(_0456_));
 sg13g2_buf_2 fanout342 (.A(net344),
    .X(net342));
 sg13g2_buf_4 fanout343 (.X(net343),
    .A(net344));
 sg13g2_buf_2 fanout344 (.A(_0433_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(net348),
    .X(net345));
 sg13g2_buf_1 fanout346 (.A(net348),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(net348),
    .X(net347));
 sg13g2_buf_1 fanout348 (.A(net354),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(net354),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(net354),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(net353),
    .X(net351));
 sg13g2_buf_1 fanout352 (.A(net353),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(net354),
    .X(net353));
 sg13g2_buf_1 fanout354 (.A(_0414_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(net356),
    .X(net355));
 sg13g2_buf_4 fanout356 (.X(net356),
    .A(_0413_));
 sg13g2_buf_2 fanout357 (.A(net358),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(net360),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(net360),
    .X(net359));
 sg13g2_buf_1 fanout360 (.A(_0413_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(net362),
    .X(net361));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(net367));
 sg13g2_buf_2 fanout363 (.A(net366),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(net366),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(net366),
    .X(net365));
 sg13g2_buf_1 fanout366 (.A(net367),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_0397_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(net372),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(net372),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(net372),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(net372),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_0396_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(net377),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(net377),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(net376),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(net377),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_0396_),
    .X(net377));
 sg13g2_buf_4 fanout378 (.X(net378),
    .A(_0504_));
 sg13g2_buf_4 fanout379 (.X(net379),
    .A(_0429_));
 sg13g2_buf_2 fanout380 (.A(net381),
    .X(net380));
 sg13g2_buf_4 fanout381 (.X(net381),
    .A(_0395_));
 sg13g2_buf_2 fanout382 (.A(net383),
    .X(net382));
 sg13g2_buf_4 fanout383 (.X(net383),
    .A(_0357_));
 sg13g2_buf_2 fanout384 (.A(net386),
    .X(net384));
 sg13g2_buf_1 fanout385 (.A(net386),
    .X(net385));
 sg13g2_buf_4 fanout386 (.X(net386),
    .A(net387));
 sg13g2_buf_4 fanout387 (.X(net387),
    .A(net392));
 sg13g2_buf_2 fanout388 (.A(net392),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(net392),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(net391),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(net392),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_0382_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(net394),
    .X(net393));
 sg13g2_buf_4 fanout394 (.X(net394),
    .A(_0381_));
 sg13g2_buf_2 fanout395 (.A(net397),
    .X(net395));
 sg13g2_buf_1 fanout396 (.A(net397),
    .X(net396));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(_0381_));
 sg13g2_buf_2 fanout398 (.A(net399),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(net401),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(net401),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_0381_),
    .X(net401));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(_0422_));
 sg13g2_buf_4 fanout403 (.X(net403),
    .A(net404));
 sg13g2_buf_4 fanout404 (.X(net404),
    .A(_0387_));
 sg13g2_buf_4 fanout405 (.X(net405),
    .A(net406));
 sg13g2_buf_4 fanout406 (.X(net406),
    .A(_0387_));
 sg13g2_buf_4 fanout407 (.X(net407),
    .A(net409));
 sg13g2_buf_2 fanout408 (.A(net409),
    .X(net408));
 sg13g2_buf_4 fanout409 (.X(net409),
    .A(_0386_));
 sg13g2_buf_2 fanout410 (.A(_0060_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(net412),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(net85),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_1078_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_1078_),
    .X(net414));
 sg13g2_buf_4 fanout415 (.X(net415),
    .A(_0384_));
 sg13g2_buf_2 fanout416 (.A(_0384_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(\hvsync_gen.vsync ),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(net419),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(net420),
    .X(net419));
 sg13g2_buf_4 fanout420 (.X(net420),
    .A(\hvsync_gen.vpos[1] ));
 sg13g2_buf_4 fanout421 (.X(net421),
    .A(\hvsync_gen.vpos[0] ));
 sg13g2_buf_1 fanout422 (.A(\hvsync_gen.vpos[0] ),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(net87),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(b),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(net426),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(\a[1] ),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(net428),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(net86),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(net1),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(net431),
    .X(net430));
 sg13g2_buf_4 fanout431 (.X(net431),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_tielo tt_um_vga_glyph_mode_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0021_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0014_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0198_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold4 (.A(\g_x[2] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0181_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold6 (.A(\hvsync_gen.vpos[9] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0064_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold8 (.A(\div3.in[6] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0063_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold10 (.A(\g_x[1] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0046_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0029_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0157_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0005_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0017_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0052_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold17 (.A(\div3.in[1] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0155_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0006_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold20 (.A(\hvsync_gen.hpos[9] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0054_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0013_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0057_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold24 (.A(\hvsync_gen.hpos[6] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0188_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold26 (.A(\hvsync_gen.hpos[8] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0053_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold28 (.A(\div3.in[4] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0061_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold30 (.A(\a[0] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold31 (.A(b),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0186_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0012_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0094_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold35 (.A(\a[1] ),
    .X(net91));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_4 FILLER_2_266 ();
 sg13g2_decap_4 FILLER_2_274 ();
 sg13g2_fill_1 FILLER_2_278 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_4 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_144 ();
 sg13g2_decap_8 FILLER_3_151 ();
 sg13g2_decap_4 FILLER_3_158 ();
 sg13g2_fill_1 FILLER_3_162 ();
 sg13g2_decap_8 FILLER_3_169 ();
 sg13g2_decap_8 FILLER_3_176 ();
 sg13g2_decap_8 FILLER_3_183 ();
 sg13g2_decap_8 FILLER_3_190 ();
 sg13g2_decap_8 FILLER_3_197 ();
 sg13g2_decap_8 FILLER_3_204 ();
 sg13g2_fill_1 FILLER_3_211 ();
 sg13g2_decap_8 FILLER_3_220 ();
 sg13g2_decap_8 FILLER_3_243 ();
 sg13g2_decap_8 FILLER_3_250 ();
 sg13g2_fill_1 FILLER_3_257 ();
 sg13g2_fill_2 FILLER_3_302 ();
 sg13g2_fill_1 FILLER_3_304 ();
 sg13g2_fill_2 FILLER_3_310 ();
 sg13g2_fill_1 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_324 ();
 sg13g2_fill_2 FILLER_3_331 ();
 sg13g2_decap_8 FILLER_3_341 ();
 sg13g2_decap_8 FILLER_3_348 ();
 sg13g2_decap_8 FILLER_3_355 ();
 sg13g2_decap_8 FILLER_3_362 ();
 sg13g2_decap_8 FILLER_3_369 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_fill_2 FILLER_4_126 ();
 sg13g2_fill_1 FILLER_4_128 ();
 sg13g2_decap_4 FILLER_4_152 ();
 sg13g2_fill_1 FILLER_4_156 ();
 sg13g2_fill_2 FILLER_4_179 ();
 sg13g2_fill_2 FILLER_4_196 ();
 sg13g2_fill_1 FILLER_4_228 ();
 sg13g2_fill_2 FILLER_4_234 ();
 sg13g2_fill_1 FILLER_4_236 ();
 sg13g2_fill_1 FILLER_4_254 ();
 sg13g2_fill_2 FILLER_4_278 ();
 sg13g2_fill_1 FILLER_4_280 ();
 sg13g2_fill_1 FILLER_4_303 ();
 sg13g2_fill_2 FILLER_4_334 ();
 sg13g2_fill_1 FILLER_4_341 ();
 sg13g2_decap_8 FILLER_4_352 ();
 sg13g2_fill_2 FILLER_4_363 ();
 sg13g2_decap_8 FILLER_4_370 ();
 sg13g2_decap_8 FILLER_4_377 ();
 sg13g2_decap_8 FILLER_4_384 ();
 sg13g2_decap_8 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_4 FILLER_5_140 ();
 sg13g2_fill_2 FILLER_5_152 ();
 sg13g2_fill_1 FILLER_5_166 ();
 sg13g2_fill_1 FILLER_5_173 ();
 sg13g2_decap_4 FILLER_5_179 ();
 sg13g2_fill_2 FILLER_5_183 ();
 sg13g2_decap_8 FILLER_5_205 ();
 sg13g2_fill_1 FILLER_5_212 ();
 sg13g2_decap_8 FILLER_5_218 ();
 sg13g2_fill_1 FILLER_5_225 ();
 sg13g2_fill_1 FILLER_5_236 ();
 sg13g2_decap_8 FILLER_5_253 ();
 sg13g2_fill_2 FILLER_5_260 ();
 sg13g2_fill_1 FILLER_5_262 ();
 sg13g2_decap_4 FILLER_5_282 ();
 sg13g2_fill_2 FILLER_5_286 ();
 sg13g2_fill_1 FILLER_5_293 ();
 sg13g2_decap_8 FILLER_5_299 ();
 sg13g2_fill_2 FILLER_5_312 ();
 sg13g2_fill_1 FILLER_5_314 ();
 sg13g2_fill_2 FILLER_5_336 ();
 sg13g2_fill_2 FILLER_5_352 ();
 sg13g2_fill_1 FILLER_5_354 ();
 sg13g2_fill_1 FILLER_5_364 ();
 sg13g2_fill_2 FILLER_5_381 ();
 sg13g2_fill_1 FILLER_5_383 ();
 sg13g2_fill_2 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_4 FILLER_5_403 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_fill_2 FILLER_6_126 ();
 sg13g2_decap_4 FILLER_6_133 ();
 sg13g2_fill_1 FILLER_6_142 ();
 sg13g2_decap_4 FILLER_6_159 ();
 sg13g2_fill_2 FILLER_6_163 ();
 sg13g2_fill_2 FILLER_6_178 ();
 sg13g2_fill_1 FILLER_6_180 ();
 sg13g2_fill_1 FILLER_6_202 ();
 sg13g2_decap_4 FILLER_6_227 ();
 sg13g2_decap_4 FILLER_6_252 ();
 sg13g2_fill_2 FILLER_6_256 ();
 sg13g2_fill_2 FILLER_6_282 ();
 sg13g2_fill_1 FILLER_6_284 ();
 sg13g2_fill_2 FILLER_6_290 ();
 sg13g2_fill_1 FILLER_6_292 ();
 sg13g2_fill_2 FILLER_6_303 ();
 sg13g2_decap_4 FILLER_6_310 ();
 sg13g2_fill_2 FILLER_6_314 ();
 sg13g2_decap_4 FILLER_6_322 ();
 sg13g2_fill_1 FILLER_6_326 ();
 sg13g2_decap_4 FILLER_6_333 ();
 sg13g2_fill_2 FILLER_6_337 ();
 sg13g2_fill_2 FILLER_6_343 ();
 sg13g2_fill_1 FILLER_6_345 ();
 sg13g2_decap_4 FILLER_6_361 ();
 sg13g2_fill_1 FILLER_6_373 ();
 sg13g2_fill_2 FILLER_6_378 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_fill_1 FILLER_7_133 ();
 sg13g2_fill_2 FILLER_7_146 ();
 sg13g2_fill_1 FILLER_7_148 ();
 sg13g2_decap_4 FILLER_7_162 ();
 sg13g2_decap_8 FILLER_7_187 ();
 sg13g2_decap_8 FILLER_7_194 ();
 sg13g2_fill_1 FILLER_7_216 ();
 sg13g2_fill_2 FILLER_7_232 ();
 sg13g2_fill_1 FILLER_7_234 ();
 sg13g2_decap_4 FILLER_7_251 ();
 sg13g2_fill_2 FILLER_7_260 ();
 sg13g2_fill_1 FILLER_7_262 ();
 sg13g2_decap_4 FILLER_7_278 ();
 sg13g2_fill_1 FILLER_7_282 ();
 sg13g2_fill_2 FILLER_7_306 ();
 sg13g2_decap_4 FILLER_7_323 ();
 sg13g2_fill_2 FILLER_7_336 ();
 sg13g2_fill_1 FILLER_7_338 ();
 sg13g2_decap_4 FILLER_7_362 ();
 sg13g2_fill_2 FILLER_7_366 ();
 sg13g2_fill_1 FILLER_7_374 ();
 sg13g2_decap_4 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_4 FILLER_8_119 ();
 sg13g2_decap_4 FILLER_8_135 ();
 sg13g2_fill_1 FILLER_8_154 ();
 sg13g2_fill_1 FILLER_8_161 ();
 sg13g2_fill_2 FILLER_8_170 ();
 sg13g2_fill_1 FILLER_8_182 ();
 sg13g2_decap_4 FILLER_8_202 ();
 sg13g2_fill_2 FILLER_8_226 ();
 sg13g2_decap_8 FILLER_8_251 ();
 sg13g2_fill_1 FILLER_8_258 ();
 sg13g2_fill_2 FILLER_8_265 ();
 sg13g2_fill_2 FILLER_8_281 ();
 sg13g2_fill_2 FILLER_8_287 ();
 sg13g2_fill_1 FILLER_8_289 ();
 sg13g2_decap_4 FILLER_8_304 ();
 sg13g2_fill_2 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_fill_1 FILLER_8_336 ();
 sg13g2_fill_2 FILLER_8_357 ();
 sg13g2_fill_1 FILLER_8_359 ();
 sg13g2_fill_1 FILLER_8_385 ();
 sg13g2_decap_4 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_4 FILLER_9_119 ();
 sg13g2_fill_1 FILLER_9_123 ();
 sg13g2_fill_2 FILLER_9_144 ();
 sg13g2_fill_1 FILLER_9_146 ();
 sg13g2_decap_4 FILLER_9_172 ();
 sg13g2_fill_1 FILLER_9_176 ();
 sg13g2_fill_1 FILLER_9_190 ();
 sg13g2_fill_1 FILLER_9_206 ();
 sg13g2_decap_4 FILLER_9_227 ();
 sg13g2_decap_8 FILLER_9_261 ();
 sg13g2_fill_2 FILLER_9_268 ();
 sg13g2_fill_1 FILLER_9_270 ();
 sg13g2_fill_2 FILLER_9_300 ();
 sg13g2_fill_1 FILLER_9_302 ();
 sg13g2_decap_4 FILLER_9_332 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_fill_1 FILLER_9_359 ();
 sg13g2_fill_2 FILLER_9_365 ();
 sg13g2_fill_1 FILLER_9_367 ();
 sg13g2_fill_2 FILLER_9_379 ();
 sg13g2_fill_1 FILLER_9_381 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_fill_2 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_128 ();
 sg13g2_decap_8 FILLER_10_159 ();
 sg13g2_fill_1 FILLER_10_173 ();
 sg13g2_fill_1 FILLER_10_192 ();
 sg13g2_fill_2 FILLER_10_198 ();
 sg13g2_fill_2 FILLER_10_209 ();
 sg13g2_fill_1 FILLER_10_211 ();
 sg13g2_decap_8 FILLER_10_216 ();
 sg13g2_fill_1 FILLER_10_223 ();
 sg13g2_fill_2 FILLER_10_234 ();
 sg13g2_fill_1 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_275 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_decap_8 FILLER_10_303 ();
 sg13g2_decap_4 FILLER_10_322 ();
 sg13g2_fill_2 FILLER_10_341 ();
 sg13g2_decap_4 FILLER_10_363 ();
 sg13g2_fill_1 FILLER_10_367 ();
 sg13g2_fill_1 FILLER_10_383 ();
 sg13g2_fill_1 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_126 ();
 sg13g2_fill_1 FILLER_11_136 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_fill_1 FILLER_11_179 ();
 sg13g2_fill_2 FILLER_11_213 ();
 sg13g2_fill_1 FILLER_11_215 ();
 sg13g2_fill_2 FILLER_11_241 ();
 sg13g2_fill_1 FILLER_11_243 ();
 sg13g2_decap_4 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_270 ();
 sg13g2_decap_4 FILLER_11_277 ();
 sg13g2_fill_1 FILLER_11_281 ();
 sg13g2_fill_2 FILLER_11_297 ();
 sg13g2_decap_4 FILLER_11_304 ();
 sg13g2_fill_2 FILLER_11_323 ();
 sg13g2_fill_1 FILLER_11_325 ();
 sg13g2_fill_1 FILLER_11_331 ();
 sg13g2_fill_2 FILLER_11_338 ();
 sg13g2_fill_1 FILLER_11_340 ();
 sg13g2_fill_1 FILLER_11_346 ();
 sg13g2_fill_2 FILLER_11_351 ();
 sg13g2_decap_4 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_fill_2 FILLER_12_119 ();
 sg13g2_fill_1 FILLER_12_121 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_fill_2 FILLER_12_170 ();
 sg13g2_fill_1 FILLER_12_172 ();
 sg13g2_decap_4 FILLER_12_188 ();
 sg13g2_fill_2 FILLER_12_197 ();
 sg13g2_fill_1 FILLER_12_199 ();
 sg13g2_decap_8 FILLER_12_213 ();
 sg13g2_fill_2 FILLER_12_220 ();
 sg13g2_decap_8 FILLER_12_240 ();
 sg13g2_decap_4 FILLER_12_247 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_fill_2 FILLER_12_329 ();
 sg13g2_fill_2 FILLER_12_335 ();
 sg13g2_decap_8 FILLER_12_342 ();
 sg13g2_fill_1 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_fill_2 FILLER_12_384 ();
 sg13g2_fill_1 FILLER_12_386 ();
 sg13g2_fill_2 FILLER_12_396 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_fill_2 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_4 FILLER_13_154 ();
 sg13g2_fill_1 FILLER_13_158 ();
 sg13g2_decap_4 FILLER_13_167 ();
 sg13g2_fill_2 FILLER_13_171 ();
 sg13g2_decap_4 FILLER_13_189 ();
 sg13g2_fill_2 FILLER_13_229 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_fill_1 FILLER_13_252 ();
 sg13g2_fill_2 FILLER_13_263 ();
 sg13g2_fill_1 FILLER_13_265 ();
 sg13g2_fill_2 FILLER_13_284 ();
 sg13g2_fill_1 FILLER_13_286 ();
 sg13g2_fill_1 FILLER_13_311 ();
 sg13g2_fill_2 FILLER_13_316 ();
 sg13g2_fill_1 FILLER_13_318 ();
 sg13g2_decap_8 FILLER_13_323 ();
 sg13g2_fill_2 FILLER_13_330 ();
 sg13g2_fill_1 FILLER_13_332 ();
 sg13g2_decap_4 FILLER_13_360 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_4 FILLER_14_119 ();
 sg13g2_fill_1 FILLER_14_123 ();
 sg13g2_decap_4 FILLER_14_141 ();
 sg13g2_fill_1 FILLER_14_167 ();
 sg13g2_fill_2 FILLER_14_181 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_decap_4 FILLER_14_198 ();
 sg13g2_fill_1 FILLER_14_202 ();
 sg13g2_decap_8 FILLER_14_211 ();
 sg13g2_decap_8 FILLER_14_218 ();
 sg13g2_decap_4 FILLER_14_225 ();
 sg13g2_decap_4 FILLER_14_250 ();
 sg13g2_decap_8 FILLER_14_275 ();
 sg13g2_decap_8 FILLER_14_282 ();
 sg13g2_fill_2 FILLER_14_289 ();
 sg13g2_fill_1 FILLER_14_291 ();
 sg13g2_decap_4 FILLER_14_317 ();
 sg13g2_fill_2 FILLER_14_321 ();
 sg13g2_fill_2 FILLER_14_331 ();
 sg13g2_fill_2 FILLER_14_338 ();
 sg13g2_fill_2 FILLER_14_344 ();
 sg13g2_fill_2 FILLER_14_361 ();
 sg13g2_fill_1 FILLER_14_372 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_4 FILLER_15_105 ();
 sg13g2_fill_2 FILLER_15_109 ();
 sg13g2_decap_4 FILLER_15_115 ();
 sg13g2_fill_1 FILLER_15_119 ();
 sg13g2_fill_2 FILLER_15_131 ();
 sg13g2_fill_1 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_fill_2 FILLER_15_155 ();
 sg13g2_decap_4 FILLER_15_171 ();
 sg13g2_fill_2 FILLER_15_192 ();
 sg13g2_fill_1 FILLER_15_194 ();
 sg13g2_fill_2 FILLER_15_203 ();
 sg13g2_decap_4 FILLER_15_247 ();
 sg13g2_decap_8 FILLER_15_265 ();
 sg13g2_decap_4 FILLER_15_272 ();
 sg13g2_fill_2 FILLER_15_290 ();
 sg13g2_fill_1 FILLER_15_316 ();
 sg13g2_fill_2 FILLER_15_337 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_fill_2 FILLER_15_371 ();
 sg13g2_fill_1 FILLER_15_373 ();
 sg13g2_fill_1 FILLER_15_379 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_4 FILLER_16_98 ();
 sg13g2_fill_2 FILLER_16_102 ();
 sg13g2_decap_4 FILLER_16_124 ();
 sg13g2_fill_2 FILLER_16_128 ();
 sg13g2_fill_2 FILLER_16_146 ();
 sg13g2_fill_2 FILLER_16_153 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_fill_1 FILLER_16_175 ();
 sg13g2_fill_2 FILLER_16_194 ();
 sg13g2_fill_2 FILLER_16_205 ();
 sg13g2_fill_1 FILLER_16_212 ();
 sg13g2_decap_4 FILLER_16_218 ();
 sg13g2_fill_2 FILLER_16_222 ();
 sg13g2_fill_1 FILLER_16_229 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_fill_2 FILLER_16_242 ();
 sg13g2_fill_1 FILLER_16_244 ();
 sg13g2_decap_8 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_264 ();
 sg13g2_fill_1 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_316 ();
 sg13g2_fill_1 FILLER_16_318 ();
 sg13g2_decap_4 FILLER_16_327 ();
 sg13g2_fill_1 FILLER_16_331 ();
 sg13g2_decap_4 FILLER_16_349 ();
 sg13g2_fill_1 FILLER_16_353 ();
 sg13g2_fill_2 FILLER_16_360 ();
 sg13g2_fill_1 FILLER_16_367 ();
 sg13g2_decap_4 FILLER_16_374 ();
 sg13g2_fill_2 FILLER_16_378 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_fill_1 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_79 ();
 sg13g2_decap_8 FILLER_17_86 ();
 sg13g2_fill_2 FILLER_17_93 ();
 sg13g2_decap_8 FILLER_17_113 ();
 sg13g2_decap_4 FILLER_17_120 ();
 sg13g2_fill_1 FILLER_17_133 ();
 sg13g2_fill_2 FILLER_17_148 ();
 sg13g2_fill_1 FILLER_17_150 ();
 sg13g2_fill_2 FILLER_17_157 ();
 sg13g2_fill_1 FILLER_17_159 ();
 sg13g2_fill_1 FILLER_17_165 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_fill_2 FILLER_17_177 ();
 sg13g2_fill_2 FILLER_17_189 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_223 ();
 sg13g2_fill_1 FILLER_17_245 ();
 sg13g2_fill_2 FILLER_17_256 ();
 sg13g2_fill_2 FILLER_17_264 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_279 ();
 sg13g2_fill_1 FILLER_17_286 ();
 sg13g2_decap_4 FILLER_17_291 ();
 sg13g2_decap_4 FILLER_17_309 ();
 sg13g2_fill_1 FILLER_17_313 ();
 sg13g2_fill_1 FILLER_17_334 ();
 sg13g2_fill_2 FILLER_17_340 ();
 sg13g2_fill_1 FILLER_17_342 ();
 sg13g2_fill_1 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_fill_2 FILLER_18_42 ();
 sg13g2_fill_1 FILLER_18_44 ();
 sg13g2_decap_4 FILLER_18_71 ();
 sg13g2_fill_1 FILLER_18_75 ();
 sg13g2_fill_2 FILLER_18_85 ();
 sg13g2_fill_1 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_109 ();
 sg13g2_decap_4 FILLER_18_139 ();
 sg13g2_decap_8 FILLER_18_162 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_fill_2 FILLER_18_193 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_205 ();
 sg13g2_fill_2 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_fill_2 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_265 ();
 sg13g2_decap_8 FILLER_18_289 ();
 sg13g2_fill_2 FILLER_18_301 ();
 sg13g2_fill_2 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_321 ();
 sg13g2_decap_4 FILLER_18_335 ();
 sg13g2_fill_2 FILLER_18_344 ();
 sg13g2_fill_2 FILLER_18_350 ();
 sg13g2_fill_1 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_358 ();
 sg13g2_fill_1 FILLER_18_372 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_4 FILLER_19_42 ();
 sg13g2_fill_1 FILLER_19_46 ();
 sg13g2_fill_1 FILLER_19_115 ();
 sg13g2_fill_2 FILLER_19_183 ();
 sg13g2_fill_1 FILLER_19_185 ();
 sg13g2_decap_4 FILLER_19_191 ();
 sg13g2_fill_1 FILLER_19_195 ();
 sg13g2_fill_2 FILLER_19_215 ();
 sg13g2_fill_2 FILLER_19_220 ();
 sg13g2_fill_2 FILLER_19_227 ();
 sg13g2_fill_2 FILLER_19_254 ();
 sg13g2_fill_1 FILLER_19_256 ();
 sg13g2_decap_4 FILLER_19_281 ();
 sg13g2_fill_2 FILLER_19_308 ();
 sg13g2_fill_2 FILLER_19_316 ();
 sg13g2_fill_2 FILLER_19_339 ();
 sg13g2_fill_1 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_4 FILLER_20_35 ();
 sg13g2_fill_1 FILLER_20_65 ();
 sg13g2_fill_1 FILLER_20_83 ();
 sg13g2_fill_1 FILLER_20_100 ();
 sg13g2_fill_2 FILLER_20_116 ();
 sg13g2_fill_2 FILLER_20_127 ();
 sg13g2_fill_1 FILLER_20_129 ();
 sg13g2_fill_1 FILLER_20_143 ();
 sg13g2_decap_8 FILLER_20_148 ();
 sg13g2_decap_8 FILLER_20_155 ();
 sg13g2_decap_8 FILLER_20_162 ();
 sg13g2_fill_2 FILLER_20_169 ();
 sg13g2_fill_1 FILLER_20_171 ();
 sg13g2_fill_2 FILLER_20_210 ();
 sg13g2_decap_4 FILLER_20_217 ();
 sg13g2_fill_2 FILLER_20_221 ();
 sg13g2_fill_2 FILLER_20_230 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_fill_2 FILLER_20_252 ();
 sg13g2_fill_1 FILLER_20_254 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_decap_4 FILLER_20_317 ();
 sg13g2_fill_1 FILLER_20_321 ();
 sg13g2_fill_1 FILLER_20_332 ();
 sg13g2_fill_1 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_fill_1 FILLER_20_379 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_fill_1 FILLER_21_82 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_fill_1 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_227 ();
 sg13g2_fill_1 FILLER_21_236 ();
 sg13g2_fill_2 FILLER_21_250 ();
 sg13g2_decap_4 FILLER_21_260 ();
 sg13g2_decap_8 FILLER_21_271 ();
 sg13g2_decap_8 FILLER_21_278 ();
 sg13g2_decap_4 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_330 ();
 sg13g2_fill_2 FILLER_21_344 ();
 sg13g2_decap_4 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_44 ();
 sg13g2_decap_4 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_57 ();
 sg13g2_fill_2 FILLER_22_116 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_fill_2 FILLER_22_182 ();
 sg13g2_fill_1 FILLER_22_193 ();
 sg13g2_fill_2 FILLER_22_220 ();
 sg13g2_fill_1 FILLER_22_222 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_decap_4 FILLER_22_251 ();
 sg13g2_decap_4 FILLER_22_268 ();
 sg13g2_fill_1 FILLER_22_272 ();
 sg13g2_fill_2 FILLER_22_287 ();
 sg13g2_fill_1 FILLER_22_289 ();
 sg13g2_decap_4 FILLER_22_295 ();
 sg13g2_decap_4 FILLER_22_315 ();
 sg13g2_fill_1 FILLER_22_324 ();
 sg13g2_fill_2 FILLER_22_346 ();
 sg13g2_fill_1 FILLER_22_348 ();
 sg13g2_fill_2 FILLER_22_366 ();
 sg13g2_fill_1 FILLER_22_376 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_fill_2 FILLER_23_68 ();
 sg13g2_fill_2 FILLER_23_114 ();
 sg13g2_fill_1 FILLER_23_116 ();
 sg13g2_fill_2 FILLER_23_168 ();
 sg13g2_fill_1 FILLER_23_170 ();
 sg13g2_fill_2 FILLER_23_215 ();
 sg13g2_fill_2 FILLER_23_257 ();
 sg13g2_fill_1 FILLER_23_259 ();
 sg13g2_fill_2 FILLER_23_268 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_fill_2 FILLER_23_285 ();
 sg13g2_fill_1 FILLER_23_287 ();
 sg13g2_fill_2 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_330 ();
 sg13g2_decap_8 FILLER_23_344 ();
 sg13g2_fill_2 FILLER_23_363 ();
 sg13g2_fill_1 FILLER_23_365 ();
 sg13g2_fill_2 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_fill_1 FILLER_24_32 ();
 sg13g2_fill_1 FILLER_24_45 ();
 sg13g2_decap_8 FILLER_24_55 ();
 sg13g2_fill_2 FILLER_24_80 ();
 sg13g2_fill_2 FILLER_24_87 ();
 sg13g2_fill_1 FILLER_24_89 ();
 sg13g2_fill_2 FILLER_24_94 ();
 sg13g2_fill_2 FILLER_24_204 ();
 sg13g2_fill_1 FILLER_24_206 ();
 sg13g2_decap_8 FILLER_24_233 ();
 sg13g2_fill_2 FILLER_24_240 ();
 sg13g2_decap_8 FILLER_24_246 ();
 sg13g2_decap_4 FILLER_24_253 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_decap_4 FILLER_24_296 ();
 sg13g2_fill_2 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_316 ();
 sg13g2_decap_8 FILLER_24_323 ();
 sg13g2_fill_1 FILLER_24_330 ();
 sg13g2_decap_8 FILLER_24_339 ();
 sg13g2_decap_4 FILLER_24_346 ();
 sg13g2_fill_1 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_66 ();
 sg13g2_decap_4 FILLER_25_82 ();
 sg13g2_fill_1 FILLER_25_86 ();
 sg13g2_fill_2 FILLER_25_113 ();
 sg13g2_fill_1 FILLER_25_141 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_fill_2 FILLER_25_261 ();
 sg13g2_fill_1 FILLER_25_263 ();
 sg13g2_decap_4 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_decap_4 FILLER_25_284 ();
 sg13g2_decap_4 FILLER_25_342 ();
 sg13g2_fill_1 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_32 ();
 sg13g2_fill_1 FILLER_26_54 ();
 sg13g2_fill_2 FILLER_26_78 ();
 sg13g2_decap_8 FILLER_26_85 ();
 sg13g2_decap_8 FILLER_26_92 ();
 sg13g2_fill_2 FILLER_26_108 ();
 sg13g2_fill_1 FILLER_26_110 ();
 sg13g2_fill_1 FILLER_26_115 ();
 sg13g2_fill_1 FILLER_26_124 ();
 sg13g2_fill_2 FILLER_26_174 ();
 sg13g2_fill_2 FILLER_26_210 ();
 sg13g2_fill_1 FILLER_26_231 ();
 sg13g2_fill_2 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_288 ();
 sg13g2_decap_8 FILLER_26_311 ();
 sg13g2_decap_8 FILLER_26_318 ();
 sg13g2_fill_2 FILLER_26_345 ();
 sg13g2_fill_1 FILLER_26_347 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_46 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_fill_2 FILLER_27_61 ();
 sg13g2_decap_4 FILLER_27_85 ();
 sg13g2_fill_1 FILLER_27_96 ();
 sg13g2_fill_1 FILLER_27_132 ();
 sg13g2_fill_1 FILLER_27_154 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_fill_1 FILLER_27_197 ();
 sg13g2_fill_2 FILLER_27_206 ();
 sg13g2_fill_1 FILLER_27_208 ();
 sg13g2_fill_1 FILLER_27_227 ();
 sg13g2_decap_4 FILLER_27_270 ();
 sg13g2_fill_2 FILLER_27_274 ();
 sg13g2_fill_2 FILLER_27_298 ();
 sg13g2_fill_1 FILLER_27_300 ();
 sg13g2_decap_8 FILLER_27_311 ();
 sg13g2_decap_4 FILLER_27_347 ();
 sg13g2_fill_2 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_362 ();
 sg13g2_decap_8 FILLER_27_369 ();
 sg13g2_decap_8 FILLER_27_376 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_decap_8 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_fill_2 FILLER_28_28 ();
 sg13g2_fill_1 FILLER_28_30 ();
 sg13g2_fill_2 FILLER_28_54 ();
 sg13g2_fill_2 FILLER_28_71 ();
 sg13g2_fill_1 FILLER_28_95 ();
 sg13g2_decap_4 FILLER_28_122 ();
 sg13g2_fill_2 FILLER_28_126 ();
 sg13g2_fill_2 FILLER_28_132 ();
 sg13g2_fill_2 FILLER_28_160 ();
 sg13g2_fill_2 FILLER_28_190 ();
 sg13g2_fill_2 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_4 FILLER_28_231 ();
 sg13g2_fill_1 FILLER_28_235 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_fill_1 FILLER_28_259 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_275 ();
 sg13g2_decap_4 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_fill_2 FILLER_28_325 ();
 sg13g2_fill_1 FILLER_28_327 ();
 sg13g2_decap_8 FILLER_28_341 ();
 sg13g2_decap_8 FILLER_28_348 ();
 sg13g2_decap_8 FILLER_28_355 ();
 sg13g2_decap_8 FILLER_28_362 ();
 sg13g2_decap_8 FILLER_28_369 ();
 sg13g2_decap_8 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_28_383 ();
 sg13g2_decap_8 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_4 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_51 ();
 sg13g2_decap_4 FILLER_29_58 ();
 sg13g2_fill_2 FILLER_29_62 ();
 sg13g2_fill_2 FILLER_29_79 ();
 sg13g2_decap_4 FILLER_29_90 ();
 sg13g2_fill_1 FILLER_29_94 ();
 sg13g2_fill_2 FILLER_29_104 ();
 sg13g2_fill_1 FILLER_29_106 ();
 sg13g2_decap_4 FILLER_29_111 ();
 sg13g2_fill_2 FILLER_29_115 ();
 sg13g2_fill_2 FILLER_29_143 ();
 sg13g2_fill_2 FILLER_29_154 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_decap_8 FILLER_29_229 ();
 sg13g2_fill_2 FILLER_29_236 ();
 sg13g2_fill_1 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_247 ();
 sg13g2_fill_2 FILLER_29_254 ();
 sg13g2_fill_1 FILLER_29_256 ();
 sg13g2_decap_4 FILLER_29_262 ();
 sg13g2_decap_4 FILLER_29_271 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_fill_1 FILLER_29_282 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_decap_4 FILLER_29_298 ();
 sg13g2_fill_2 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_316 ();
 sg13g2_decap_8 FILLER_29_323 ();
 sg13g2_decap_8 FILLER_29_330 ();
 sg13g2_decap_8 FILLER_29_337 ();
 sg13g2_decap_8 FILLER_29_344 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_81 ();
 sg13g2_fill_2 FILLER_30_144 ();
 sg13g2_fill_2 FILLER_30_172 ();
 sg13g2_fill_2 FILLER_30_219 ();
 sg13g2_fill_1 FILLER_30_221 ();
 sg13g2_fill_2 FILLER_30_230 ();
 sg13g2_fill_2 FILLER_30_248 ();
 sg13g2_decap_4 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_288 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_4 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_100 ();
 sg13g2_decap_8 FILLER_31_111 ();
 sg13g2_fill_2 FILLER_31_118 ();
 sg13g2_decap_8 FILLER_31_124 ();
 sg13g2_fill_2 FILLER_31_153 ();
 sg13g2_decap_4 FILLER_31_173 ();
 sg13g2_decap_8 FILLER_31_185 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_decap_4 FILLER_31_198 ();
 sg13g2_fill_1 FILLER_31_202 ();
 sg13g2_decap_8 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_214 ();
 sg13g2_decap_8 FILLER_31_227 ();
 sg13g2_decap_4 FILLER_31_234 ();
 sg13g2_fill_2 FILLER_31_238 ();
 sg13g2_fill_2 FILLER_31_248 ();
 sg13g2_fill_1 FILLER_31_258 ();
 sg13g2_decap_8 FILLER_31_286 ();
 sg13g2_decap_4 FILLER_31_293 ();
 sg13g2_decap_8 FILLER_31_302 ();
 sg13g2_decap_8 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_316 ();
 sg13g2_decap_8 FILLER_31_323 ();
 sg13g2_decap_8 FILLER_31_330 ();
 sg13g2_decap_8 FILLER_31_337 ();
 sg13g2_decap_8 FILLER_31_344 ();
 sg13g2_decap_8 FILLER_31_351 ();
 sg13g2_decap_8 FILLER_31_358 ();
 sg13g2_decap_8 FILLER_31_365 ();
 sg13g2_decap_8 FILLER_31_372 ();
 sg13g2_decap_8 FILLER_31_379 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_decap_8 FILLER_31_393 ();
 sg13g2_decap_8 FILLER_31_400 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_fill_1 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_89 ();
 sg13g2_fill_1 FILLER_32_96 ();
 sg13g2_fill_2 FILLER_32_123 ();
 sg13g2_decap_8 FILLER_32_129 ();
 sg13g2_fill_2 FILLER_32_136 ();
 sg13g2_fill_1 FILLER_32_138 ();
 sg13g2_fill_2 FILLER_32_165 ();
 sg13g2_fill_1 FILLER_32_167 ();
 sg13g2_fill_1 FILLER_32_173 ();
 sg13g2_decap_4 FILLER_32_190 ();
 sg13g2_fill_1 FILLER_32_194 ();
 sg13g2_decap_4 FILLER_32_264 ();
 sg13g2_fill_2 FILLER_32_268 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_305 ();
 sg13g2_decap_8 FILLER_32_312 ();
 sg13g2_decap_8 FILLER_32_319 ();
 sg13g2_decap_8 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_347 ();
 sg13g2_decap_8 FILLER_32_354 ();
 sg13g2_decap_8 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_375 ();
 sg13g2_decap_8 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_32_389 ();
 sg13g2_decap_8 FILLER_32_396 ();
 sg13g2_decap_4 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_4 FILLER_33_105 ();
 sg13g2_decap_4 FILLER_33_155 ();
 sg13g2_fill_2 FILLER_33_159 ();
 sg13g2_fill_2 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_179 ();
 sg13g2_decap_8 FILLER_33_195 ();
 sg13g2_decap_4 FILLER_33_202 ();
 sg13g2_decap_4 FILLER_33_227 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_254 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_decap_8 FILLER_33_284 ();
 sg13g2_decap_8 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_decap_8 FILLER_33_305 ();
 sg13g2_decap_8 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_319 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_4 FILLER_34_126 ();
 sg13g2_fill_1 FILLER_34_130 ();
 sg13g2_fill_1 FILLER_34_141 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_fill_2 FILLER_34_154 ();
 sg13g2_fill_1 FILLER_34_156 ();
 sg13g2_decap_4 FILLER_34_175 ();
 sg13g2_fill_2 FILLER_34_179 ();
 sg13g2_decap_8 FILLER_34_201 ();
 sg13g2_decap_8 FILLER_34_208 ();
 sg13g2_fill_2 FILLER_34_215 ();
 sg13g2_decap_8 FILLER_34_222 ();
 sg13g2_decap_8 FILLER_34_229 ();
 sg13g2_fill_2 FILLER_34_236 ();
 sg13g2_decap_8 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_257 ();
 sg13g2_decap_8 FILLER_34_289 ();
 sg13g2_decap_8 FILLER_34_296 ();
 sg13g2_decap_8 FILLER_34_303 ();
 sg13g2_decap_8 FILLER_34_310 ();
 sg13g2_decap_8 FILLER_34_317 ();
 sg13g2_decap_8 FILLER_34_324 ();
 sg13g2_decap_8 FILLER_34_331 ();
 sg13g2_decap_8 FILLER_34_338 ();
 sg13g2_decap_8 FILLER_34_345 ();
 sg13g2_decap_8 FILLER_34_352 ();
 sg13g2_decap_8 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_34_366 ();
 sg13g2_decap_8 FILLER_34_373 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_fill_1 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_111 ();
 sg13g2_fill_1 FILLER_35_169 ();
 sg13g2_fill_2 FILLER_35_175 ();
 sg13g2_decap_4 FILLER_35_181 ();
 sg13g2_fill_1 FILLER_35_185 ();
 sg13g2_fill_1 FILLER_35_206 ();
 sg13g2_decap_8 FILLER_35_211 ();
 sg13g2_decap_8 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_225 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_282 ();
 sg13g2_decap_8 FILLER_35_289 ();
 sg13g2_decap_8 FILLER_35_296 ();
 sg13g2_decap_8 FILLER_35_303 ();
 sg13g2_decap_8 FILLER_35_310 ();
 sg13g2_decap_8 FILLER_35_317 ();
 sg13g2_decap_8 FILLER_35_324 ();
 sg13g2_decap_8 FILLER_35_331 ();
 sg13g2_decap_8 FILLER_35_338 ();
 sg13g2_decap_8 FILLER_35_345 ();
 sg13g2_decap_8 FILLER_35_352 ();
 sg13g2_decap_8 FILLER_35_359 ();
 sg13g2_decap_8 FILLER_35_366 ();
 sg13g2_decap_8 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_380 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_100 ();
 sg13g2_fill_2 FILLER_36_130 ();
 sg13g2_decap_8 FILLER_36_146 ();
 sg13g2_fill_1 FILLER_36_153 ();
 sg13g2_decap_4 FILLER_36_158 ();
 sg13g2_decap_4 FILLER_36_192 ();
 sg13g2_decap_8 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_229 ();
 sg13g2_fill_2 FILLER_36_239 ();
 sg13g2_fill_2 FILLER_36_254 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_282 ();
 sg13g2_decap_8 FILLER_36_289 ();
 sg13g2_decap_8 FILLER_36_296 ();
 sg13g2_decap_8 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_310 ();
 sg13g2_decap_8 FILLER_36_317 ();
 sg13g2_decap_8 FILLER_36_324 ();
 sg13g2_decap_8 FILLER_36_331 ();
 sg13g2_decap_8 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_84 ();
 sg13g2_decap_4 FILLER_37_138 ();
 sg13g2_fill_1 FILLER_37_142 ();
 sg13g2_fill_1 FILLER_37_148 ();
 sg13g2_fill_2 FILLER_37_166 ();
 sg13g2_fill_1 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_178 ();
 sg13g2_fill_1 FILLER_37_190 ();
 sg13g2_decap_8 FILLER_37_215 ();
 sg13g2_fill_2 FILLER_37_222 ();
 sg13g2_fill_2 FILLER_37_255 ();
 sg13g2_decap_8 FILLER_37_288 ();
 sg13g2_decap_8 FILLER_37_295 ();
 sg13g2_decap_8 FILLER_37_302 ();
 sg13g2_decap_8 FILLER_37_309 ();
 sg13g2_decap_8 FILLER_37_316 ();
 sg13g2_decap_8 FILLER_37_323 ();
 sg13g2_decap_8 FILLER_37_330 ();
 sg13g2_decap_8 FILLER_37_337 ();
 sg13g2_decap_8 FILLER_37_344 ();
 sg13g2_decap_8 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_92 ();
 sg13g2_fill_2 FILLER_38_115 ();
 sg13g2_fill_1 FILLER_38_117 ();
 sg13g2_fill_2 FILLER_38_126 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_192 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_229 ();
 sg13g2_fill_2 FILLER_38_247 ();
 sg13g2_fill_1 FILLER_38_249 ();
 sg13g2_decap_4 FILLER_38_253 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_fill_2 FILLER_38_365 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
endmodule

module tt_um_instrumented_ring_oscillator (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net15;
 wire net16;
 wire net26;
 wire net27;
 wire net29;
 wire net30;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net49;
 wire net50;
 wire net52;
 wire net53;
 wire net55;
 wire net56;
 wire net58;
 wire net59;
 wire net61;
 wire net62;
 wire net64;
 wire net65;
 wire net67;
 wire net68;
 wire \iro.connect[0] ;
 wire \iro.connect[10] ;
 wire \iro.connect[11] ;
 wire \iro.connect[12] ;
 wire \iro.connect[13] ;
 wire \iro.connect[14] ;
 wire \iro.connect[15] ;
 wire \iro.connect[16] ;
 wire \iro.connect[17] ;
 wire \iro.connect[18] ;
 wire \iro.connect[19] ;
 wire \iro.connect[1] ;
 wire \iro.connect[20] ;
 wire \iro.connect[21] ;
 wire \iro.connect[22] ;
 wire \iro.connect[23] ;
 wire \iro.connect[24] ;
 wire \iro.connect[2] ;
 wire \iro.connect[3] ;
 wire \iro.connect[4] ;
 wire \iro.connect[5] ;
 wire \iro.connect[6] ;
 wire \iro.connect[7] ;
 wire \iro.connect[8] ;
 wire \iro.connect[9] ;
 wire \iro.enable ;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire \iro.ro0/_0_ ;
 wire \iro.ro0/_1_ ;
 wire \iro.ro0/_2_ ;
 wire \iro.ro0/_3_ ;
 wire \iro.ro1/_0_ ;
 wire \iro.ro1/_1_ ;
 wire \iro.ro1/_2_ ;
 wire \iro.ro1/_3_ ;
 wire \iro.ro10/_0_ ;
 wire \iro.ro10/_1_ ;
 wire \iro.ro10/_2_ ;
 wire \iro.ro10/_3_ ;
 wire \iro.ro11/_0_ ;
 wire \iro.ro11/_1_ ;
 wire \iro.ro11/_2_ ;
 wire \iro.ro11/_3_ ;
 wire \iro.ro12/_0_ ;
 wire \iro.ro12/_1_ ;
 wire \iro.ro12/_2_ ;
 wire \iro.ro12/_3_ ;
 wire \iro.ro13/_0_ ;
 wire \iro.ro13/_1_ ;
 wire \iro.ro13/_2_ ;
 wire \iro.ro13/_3_ ;
 wire \iro.ro14/_0_ ;
 wire \iro.ro14/_1_ ;
 wire \iro.ro14/_2_ ;
 wire \iro.ro14/_3_ ;
 wire \iro.ro15/_0_ ;
 wire \iro.ro15/_1_ ;
 wire \iro.ro15/_2_ ;
 wire \iro.ro15/_3_ ;
 wire \iro.ro16/_0_ ;
 wire \iro.ro16/_1_ ;
 wire \iro.ro16/_2_ ;
 wire \iro.ro16/_3_ ;
 wire \iro.ro17/_0_ ;
 wire \iro.ro17/_1_ ;
 wire \iro.ro17/_2_ ;
 wire \iro.ro17/_3_ ;
 wire \iro.ro18/_0_ ;
 wire \iro.ro18/_1_ ;
 wire \iro.ro18/_2_ ;
 wire \iro.ro18/_3_ ;
 wire \iro.ro19/_0_ ;
 wire \iro.ro19/_1_ ;
 wire \iro.ro19/_2_ ;
 wire \iro.ro19/_3_ ;
 wire \iro.ro2/_0_ ;
 wire \iro.ro2/_1_ ;
 wire \iro.ro2/_2_ ;
 wire \iro.ro2/_3_ ;
 wire \iro.ro20/_0_ ;
 wire \iro.ro20/_1_ ;
 wire \iro.ro20/_2_ ;
 wire \iro.ro20/_3_ ;
 wire \iro.ro21/_0_ ;
 wire \iro.ro21/_1_ ;
 wire \iro.ro21/_2_ ;
 wire \iro.ro21/_3_ ;
 wire \iro.ro22/_0_ ;
 wire \iro.ro22/_1_ ;
 wire \iro.ro22/_2_ ;
 wire \iro.ro22/_3_ ;
 wire \iro.ro23/_0_ ;
 wire \iro.ro23/_1_ ;
 wire \iro.ro23/_2_ ;
 wire \iro.ro23/_3_ ;
 wire \iro.ro24/_0_ ;
 wire \iro.ro24/_1_ ;
 wire \iro.ro24/_2_ ;
 wire \iro.ro24/_3_ ;
 wire \iro.ro3/_0_ ;
 wire \iro.ro3/_1_ ;
 wire \iro.ro3/_2_ ;
 wire \iro.ro3/_3_ ;
 wire \iro.ro4/_0_ ;
 wire \iro.ro4/_1_ ;
 wire \iro.ro4/_2_ ;
 wire \iro.ro4/_3_ ;
 wire \iro.ro5/_0_ ;
 wire \iro.ro5/_1_ ;
 wire \iro.ro5/_2_ ;
 wire \iro.ro5/_3_ ;
 wire \iro.ro6/_0_ ;
 wire \iro.ro6/_1_ ;
 wire \iro.ro6/_2_ ;
 wire \iro.ro6/_3_ ;
 wire \iro.ro7/_0_ ;
 wire \iro.ro7/_1_ ;
 wire \iro.ro7/_2_ ;
 wire \iro.ro7/_3_ ;
 wire \iro.ro8/_0_ ;
 wire \iro.ro8/_1_ ;
 wire \iro.ro8/_2_ ;
 wire \iro.ro8/_3_ ;
 wire \iro.ro9/_0_ ;
 wire \iro.ro9/_1_ ;
 wire \iro.ro9/_2_ ;
 wire \iro.ro9/_3_ ;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net14;
 wire net25;
 wire net28;
 wire net31;
 wire net40;
 wire net48;
 wire net51;
 wire net54;
 wire net57;
 wire net60;
 wire net63;
 wire net66;

 sg13g2_inv_1 _055_ (.Y(_010_),
    .A(net6));
 sg13g2_inv_1 _056_ (.Y(_011_),
    .A(net7));
 sg13g2_nor2_1 _057_ (.A(net6),
    .B(net7),
    .Y(_012_));
 sg13g2_inv_1 _058_ (.Y(_005_),
    .A(_012_));
 sg13g2_a21o_1 _059_ (.A2(net5),
    .A1(net6),
    .B1(net7),
    .X(_007_));
 sg13g2_a21o_1 _060_ (.A2(net4),
    .A1(net6),
    .B1(_007_),
    .X(_006_));
 sg13g2_o21ai_1 _061_ (.B1(net7),
    .Y(_013_),
    .A1(net6),
    .A2(net5));
 sg13g2_inv_1 _062_ (.Y(_000_),
    .A(_013_));
 sg13g2_nor3_1 _063_ (.A(net6),
    .B(net5),
    .C(net4),
    .Y(_014_));
 sg13g2_nor2_1 _064_ (.A(_011_),
    .B(_014_),
    .Y(_009_));
 sg13g2_nand2_1 _065_ (.Y(_015_),
    .A(net5),
    .B(net4));
 sg13g2_nand2_1 _066_ (.Y(_004_),
    .A(_012_),
    .B(_015_));
 sg13g2_nand2b_1 _067_ (.Y(_003_),
    .B(_012_),
    .A_N(net5));
 sg13g2_o21ai_1 _068_ (.B1(_011_),
    .Y(_008_),
    .A1(_010_),
    .A2(_015_));
 sg13g2_nand2_1 _069_ (.Y(_002_),
    .A(_011_),
    .B(_014_));
 sg13g2_a21oi_1 _070_ (.A1(_010_),
    .A2(_015_),
    .Y(_001_),
    .B1(_011_));
 sg13g2_and2_1 _071_ (.A(net2),
    .B(net1),
    .X(\iro.enable ));
 sg13g2_tiehi tt_um_instrumented_ring_oscillator_61 (.L_HI(net69));
 sg13g2_tiehi tt_um_instrumented_ring_oscillator_62 (.L_HI(net70));
 sg13g2_tiehi tt_um_instrumented_ring_oscillator_63 (.L_HI(net71));
 sg13g2_tiehi tt_um_instrumented_ring_oscillator_64 (.L_HI(net72));
 sg13g2_tiehi tt_um_instrumented_ring_oscillator_65 (.L_HI(net73));
 sg13g2_tiehi tt_um_instrumented_ring_oscillator_66 (.L_HI(net74));
 sg13g2_tiehi tt_um_instrumented_ring_oscillator_67 (.L_HI(net75));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_tielo \iro.ro0/_5__10  (.L_LO(net10));
 sg13g2_tielo \iro.ro1/_4__11  (.L_LO(net11));
 sg13g2_tielo \iro.ro1/_5__12  (.L_LO(net12));
 sg13g2_tielo \iro.ro10/_6__13  (.L_LO(net13));
 sg13g2_tielo \iro.ro10/_5__15  (.L_LO(net15));
 sg13g2_tielo \iro.ro11/_6__16  (.L_LO(net16));
 sg13g2_tielo \iro.ro11/_5__18  (.L_LO(net26));
 sg13g2_tielo \iro.ro12/_6__19  (.L_LO(net27));
 sg13g2_tielo \iro.ro12/_5__21  (.L_LO(net29));
 sg13g2_tielo \iro.ro13/_6__22  (.L_LO(net30));
 sg13g2_tielo \iro.ro13/_5__24  (.L_LO(net32));
 sg13g2_tielo \iro.ro14/_5__25  (.L_LO(net33));
 sg13g2_tielo \iro.ro15/_5__26  (.L_LO(net34));
 sg13g2_tielo \iro.ro16/_5__27  (.L_LO(net35));
 sg13g2_tielo \iro.ro17/_5__28  (.L_LO(net36));
 sg13g2_tielo \iro.ro18/_5__29  (.L_LO(net37));
 sg13g2_tielo \iro.ro19/_5__30  (.L_LO(net38));
 sg13g2_tielo \iro.ro2/_6__31  (.L_LO(net39));
 sg13g2_tielo \iro.ro2/_5__33  (.L_LO(net41));
 sg13g2_tielo \iro.ro20/_5__34  (.L_LO(net42));
 sg13g2_tielo \iro.ro21/_5__35  (.L_LO(net43));
 sg13g2_tielo \iro.ro22/_5__36  (.L_LO(net44));
 sg13g2_tielo \iro.ro23/_5__37  (.L_LO(net45));
 sg13g2_tielo \iro.ro24/_5__38  (.L_LO(net46));
 sg13g2_tielo \iro.ro3/_6__39  (.L_LO(net47));
 sg13g2_tielo \iro.ro3/_5__41  (.L_LO(net49));
 sg13g2_tielo \iro.ro4/_6__42  (.L_LO(net50));
 sg13g2_tielo \iro.ro4/_5__44  (.L_LO(net52));
 sg13g2_tielo \iro.ro5/_6__45  (.L_LO(net53));
 sg13g2_tielo \iro.ro5/_5__47  (.L_LO(net55));
 sg13g2_tielo \iro.ro6/_6__48  (.L_LO(net56));
 sg13g2_tielo \iro.ro6/_5__50  (.L_LO(net58));
 sg13g2_tielo \iro.ro7/_6__51  (.L_LO(net59));
 sg13g2_tielo \iro.ro7/_5__53  (.L_LO(net61));
 sg13g2_tielo \iro.ro8/_6__54  (.L_LO(net62));
 sg13g2_tielo \iro.ro8/_5__56  (.L_LO(net64));
 sg13g2_tielo \iro.ro9/_6__57  (.L_LO(net65));
 sg13g2_tielo \iro.ro9/_5__59  (.L_LO(net67));
 sg13g2_tiehi tt_um_instrumented_ring_oscillator_60 (.L_HI(net68));
 sg13g2_buf_1 _119_ (.A(\iro.connect[8] ),
    .X(uio_out[0]));
 sg13g2_buf_1 _120_ (.A(\iro.connect[9] ),
    .X(uio_out[1]));
 sg13g2_buf_1 _121_ (.A(\iro.connect[10] ),
    .X(uio_out[2]));
 sg13g2_buf_1 _122_ (.A(\iro.connect[11] ),
    .X(uio_out[3]));
 sg13g2_buf_1 _123_ (.A(\iro.connect[12] ),
    .X(uio_out[4]));
 sg13g2_buf_1 _124_ (.A(\iro.connect[13] ),
    .X(uio_out[5]));
 sg13g2_buf_1 _125_ (.A(\iro.connect[14] ),
    .X(uio_out[6]));
 sg13g2_buf_1 _126_ (.A(\iro.connect[15] ),
    .X(uio_out[7]));
 sg13g2_buf_1 _127_ (.A(\iro.connect[0] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _128_ (.A(\iro.connect[1] ),
    .X(uo_out[1]));
 sg13g2_buf_1 _129_ (.A(\iro.connect[2] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _130_ (.A(\iro.connect[3] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _131_ (.A(\iro.connect[4] ),
    .X(uo_out[4]));
 sg13g2_buf_1 _132_ (.A(\iro.connect[5] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _133_ (.A(\iro.connect[6] ),
    .X(uo_out[6]));
 sg13g2_buf_1 _134_ (.A(\iro.connect[7] ),
    .X(uo_out[7]));
 sg13g2_inv_1 \iro.ro0/_4_  (.Y(\iro.ro0/_1_ ),
    .A(\iro.connect[24] ));
 sg13g2_nor2_1 \iro.ro0/_5_  (.A(net10),
    .B(net23),
    .Y(\iro.ro0/_2_ ));
 sg13g2_o21ai_1 \iro.ro0/_6_  (.B1(net23),
    .Y(\iro.ro0/_3_ ),
    .A1(\iro.connect[24] ),
    .A2(net8));
 sg13g2_a21oi_1 \iro.ro0/_7_  (.A1(\iro.ro0/_1_ ),
    .A2(net9),
    .Y(\iro.ro0/_0_ ),
    .B1(\iro.ro0/_3_ ));
 sg13g2_nor2_1 \iro.ro0/_8_  (.A(\iro.ro0/_2_ ),
    .B(\iro.ro0/_0_ ),
    .Y(\iro.connect[0] ));
 sg13g2_inv_1 \iro.ro1/_4_  (.Y(\iro.ro1/_1_ ),
    .A(net11));
 sg13g2_nor2_1 \iro.ro1/_5_  (.A(net12),
    .B(net23),
    .Y(\iro.ro1/_2_ ));
 sg13g2_o21ai_1 \iro.ro1/_6_  (.B1(net24),
    .Y(\iro.ro1/_3_ ),
    .A1(\iro.connect[0] ),
    .A2(net3));
 sg13g2_a21oi_1 \iro.ro1/_7_  (.A1(\iro.ro1/_1_ ),
    .A2(net3),
    .Y(\iro.ro1/_0_ ),
    .B1(\iro.ro1/_3_ ));
 sg13g2_nor2_1 \iro.ro1/_8_  (.A(\iro.ro1/_2_ ),
    .B(\iro.ro1/_0_ ),
    .Y(\iro.connect[1] ));
 sg13g2_inv_1 \iro.ro10/_4_  (.Y(\iro.ro10/_1_ ),
    .A(\iro.connect[9] ));
 sg13g2_nor2_1 \iro.ro10/_5_  (.A(net15),
    .B(net18),
    .Y(\iro.ro10/_2_ ));
 sg13g2_o21ai_1 \iro.ro10/_6_  (.B1(net18),
    .Y(\iro.ro10/_3_ ),
    .A1(\iro.connect[9] ),
    .A2(net13));
 sg13g2_a21oi_1 \iro.ro10/_7_  (.A1(\iro.ro10/_1_ ),
    .A2(net14),
    .Y(\iro.ro10/_0_ ),
    .B1(\iro.ro10/_3_ ));
 sg13g2_nor2_1 \iro.ro10/_8_  (.A(\iro.ro10/_2_ ),
    .B(\iro.ro10/_0_ ),
    .Y(\iro.connect[10] ));
 sg13g2_inv_1 \iro.ro11/_4_  (.Y(\iro.ro11/_1_ ),
    .A(\iro.connect[10] ));
 sg13g2_nor2_1 \iro.ro11/_5_  (.A(net26),
    .B(net17),
    .Y(\iro.ro11/_2_ ));
 sg13g2_o21ai_1 \iro.ro11/_6_  (.B1(net18),
    .Y(\iro.ro11/_3_ ),
    .A1(\iro.connect[10] ),
    .A2(net16));
 sg13g2_a21oi_1 \iro.ro11/_7_  (.A1(\iro.ro11/_1_ ),
    .A2(net25),
    .Y(\iro.ro11/_0_ ),
    .B1(\iro.ro11/_3_ ));
 sg13g2_nor2_1 \iro.ro11/_8_  (.A(\iro.ro11/_2_ ),
    .B(\iro.ro11/_0_ ),
    .Y(\iro.connect[11] ));
 sg13g2_inv_1 \iro.ro12/_4_  (.Y(\iro.ro12/_1_ ),
    .A(\iro.connect[11] ));
 sg13g2_nor2_1 \iro.ro12/_5_  (.A(net29),
    .B(net17),
    .Y(\iro.ro12/_2_ ));
 sg13g2_o21ai_1 \iro.ro12/_6_  (.B1(net17),
    .Y(\iro.ro12/_3_ ),
    .A1(\iro.connect[11] ),
    .A2(net27));
 sg13g2_a21oi_1 \iro.ro12/_7_  (.A1(\iro.ro12/_1_ ),
    .A2(net28),
    .Y(\iro.ro12/_0_ ),
    .B1(\iro.ro12/_3_ ));
 sg13g2_nor2_1 \iro.ro12/_8_  (.A(\iro.ro12/_2_ ),
    .B(\iro.ro12/_0_ ),
    .Y(\iro.connect[12] ));
 sg13g2_inv_1 \iro.ro13/_4_  (.Y(\iro.ro13/_1_ ),
    .A(\iro.connect[12] ));
 sg13g2_nor2_1 \iro.ro13/_5_  (.A(net32),
    .B(net17),
    .Y(\iro.ro13/_2_ ));
 sg13g2_o21ai_1 \iro.ro13/_6_  (.B1(net17),
    .Y(\iro.ro13/_3_ ),
    .A1(\iro.connect[12] ),
    .A2(net30));
 sg13g2_a21oi_1 \iro.ro13/_7_  (.A1(\iro.ro13/_1_ ),
    .A2(net31),
    .Y(\iro.ro13/_0_ ),
    .B1(\iro.ro13/_3_ ));
 sg13g2_nor2_1 \iro.ro13/_8_  (.A(\iro.ro13/_2_ ),
    .B(\iro.ro13/_0_ ),
    .Y(\iro.connect[13] ));
 sg13g2_inv_1 \iro.ro14/_4_  (.Y(\iro.ro14/_1_ ),
    .A(\iro.connect[13] ));
 sg13g2_nor2_1 \iro.ro14/_5_  (.A(net33),
    .B(net17),
    .Y(\iro.ro14/_2_ ));
 sg13g2_o21ai_1 \iro.ro14/_6_  (.B1(net17),
    .Y(\iro.ro14/_3_ ),
    .A1(\iro.connect[13] ),
    .A2(_001_));
 sg13g2_a21oi_1 \iro.ro14/_7_  (.A1(\iro.ro14/_1_ ),
    .A2(_001_),
    .Y(\iro.ro14/_0_ ),
    .B1(\iro.ro14/_3_ ));
 sg13g2_nor2_1 \iro.ro14/_8_  (.A(\iro.ro14/_2_ ),
    .B(\iro.ro14/_0_ ),
    .Y(\iro.connect[14] ));
 sg13g2_inv_1 \iro.ro15/_4_  (.Y(\iro.ro15/_1_ ),
    .A(\iro.connect[14] ));
 sg13g2_nor2_1 \iro.ro15/_5_  (.A(net34),
    .B(net18),
    .Y(\iro.ro15/_2_ ));
 sg13g2_o21ai_1 \iro.ro15/_6_  (.B1(net17),
    .Y(\iro.ro15/_3_ ),
    .A1(\iro.connect[12] ),
    .A2(_000_));
 sg13g2_a21oi_1 \iro.ro15/_7_  (.A1(\iro.ro15/_1_ ),
    .A2(_000_),
    .Y(\iro.ro15/_0_ ),
    .B1(\iro.ro15/_3_ ));
 sg13g2_nor2_1 \iro.ro15/_8_  (.A(\iro.ro15/_2_ ),
    .B(\iro.ro15/_0_ ),
    .Y(\iro.connect[15] ));
 sg13g2_inv_1 \iro.ro16/_4_  (.Y(\iro.ro16/_1_ ),
    .A(\iro.connect[15] ));
 sg13g2_nor2_1 \iro.ro16/_5_  (.A(net35),
    .B(net18),
    .Y(\iro.ro16/_2_ ));
 sg13g2_o21ai_1 \iro.ro16/_6_  (.B1(net20),
    .Y(\iro.ro16/_3_ ),
    .A1(\iro.connect[11] ),
    .A2(_009_));
 sg13g2_a21oi_1 \iro.ro16/_7_  (.A1(\iro.ro16/_1_ ),
    .A2(_009_),
    .Y(\iro.ro16/_0_ ),
    .B1(\iro.ro16/_3_ ));
 sg13g2_nor2_1 \iro.ro16/_8_  (.A(\iro.ro16/_2_ ),
    .B(\iro.ro16/_0_ ),
    .Y(\iro.connect[16] ));
 sg13g2_inv_1 \iro.ro17/_4_  (.Y(\iro.ro17/_1_ ),
    .A(\iro.connect[16] ));
 sg13g2_nor2_1 \iro.ro17/_5_  (.A(net36),
    .B(net18),
    .Y(\iro.ro17/_2_ ));
 sg13g2_o21ai_1 \iro.ro17/_6_  (.B1(net18),
    .Y(\iro.ro17/_3_ ),
    .A1(\iro.connect[10] ),
    .A2(net7));
 sg13g2_a21oi_1 \iro.ro17/_7_  (.A1(\iro.ro17/_1_ ),
    .A2(net7),
    .Y(\iro.ro17/_0_ ),
    .B1(\iro.ro17/_3_ ));
 sg13g2_nor2_1 \iro.ro17/_8_  (.A(\iro.ro17/_2_ ),
    .B(\iro.ro17/_0_ ),
    .Y(\iro.connect[17] ));
 sg13g2_inv_1 \iro.ro18/_4_  (.Y(\iro.ro18/_1_ ),
    .A(\iro.connect[17] ));
 sg13g2_nor2_1 \iro.ro18/_5_  (.A(net37),
    .B(net19),
    .Y(\iro.ro18/_2_ ));
 sg13g2_o21ai_1 \iro.ro18/_6_  (.B1(net19),
    .Y(\iro.ro18/_3_ ),
    .A1(\iro.connect[9] ),
    .A2(_008_));
 sg13g2_a21oi_1 \iro.ro18/_7_  (.A1(\iro.ro18/_1_ ),
    .A2(_008_),
    .Y(\iro.ro18/_0_ ),
    .B1(\iro.ro18/_3_ ));
 sg13g2_nor2_1 \iro.ro18/_8_  (.A(\iro.ro18/_2_ ),
    .B(\iro.ro18/_0_ ),
    .Y(\iro.connect[18] ));
 sg13g2_inv_1 \iro.ro19/_4_  (.Y(\iro.ro19/_1_ ),
    .A(\iro.connect[18] ));
 sg13g2_nor2_1 \iro.ro19/_5_  (.A(net38),
    .B(net20),
    .Y(\iro.ro19/_2_ ));
 sg13g2_o21ai_1 \iro.ro19/_6_  (.B1(net19),
    .Y(\iro.ro19/_3_ ),
    .A1(\iro.connect[8] ),
    .A2(_007_));
 sg13g2_a21oi_1 \iro.ro19/_7_  (.A1(\iro.ro19/_1_ ),
    .A2(_007_),
    .Y(\iro.ro19/_0_ ),
    .B1(\iro.ro19/_3_ ));
 sg13g2_nor2_1 \iro.ro19/_8_  (.A(\iro.ro19/_2_ ),
    .B(\iro.ro19/_0_ ),
    .Y(\iro.connect[19] ));
 sg13g2_inv_1 \iro.ro2/_4_  (.Y(\iro.ro2/_1_ ),
    .A(\iro.connect[1] ));
 sg13g2_nor2_1 \iro.ro2/_5_  (.A(net41),
    .B(net23),
    .Y(\iro.ro2/_2_ ));
 sg13g2_o21ai_1 \iro.ro2/_6_  (.B1(net23),
    .Y(\iro.ro2/_3_ ),
    .A1(\iro.connect[1] ),
    .A2(net39));
 sg13g2_a21oi_1 \iro.ro2/_7_  (.A1(\iro.ro2/_1_ ),
    .A2(net40),
    .Y(\iro.ro2/_0_ ),
    .B1(\iro.ro2/_3_ ));
 sg13g2_nor2_1 \iro.ro2/_8_  (.A(\iro.ro2/_2_ ),
    .B(\iro.ro2/_0_ ),
    .Y(\iro.connect[2] ));
 sg13g2_inv_1 \iro.ro20/_4_  (.Y(\iro.ro20/_1_ ),
    .A(\iro.connect[19] ));
 sg13g2_nor2_1 \iro.ro20/_5_  (.A(net42),
    .B(net19),
    .Y(\iro.ro20/_2_ ));
 sg13g2_o21ai_1 \iro.ro20/_6_  (.B1(net19),
    .Y(\iro.ro20/_3_ ),
    .A1(\iro.connect[7] ),
    .A2(_006_));
 sg13g2_a21oi_1 \iro.ro20/_7_  (.A1(\iro.ro20/_1_ ),
    .A2(_006_),
    .Y(\iro.ro20/_0_ ),
    .B1(\iro.ro20/_3_ ));
 sg13g2_nor2_1 \iro.ro20/_8_  (.A(\iro.ro20/_2_ ),
    .B(\iro.ro20/_0_ ),
    .Y(\iro.connect[20] ));
 sg13g2_inv_1 \iro.ro21/_4_  (.Y(\iro.ro21/_1_ ),
    .A(\iro.connect[20] ));
 sg13g2_nor2_1 \iro.ro21/_5_  (.A(net43),
    .B(net21),
    .Y(\iro.ro21/_2_ ));
 sg13g2_o21ai_1 \iro.ro21/_6_  (.B1(net21),
    .Y(\iro.ro21/_3_ ),
    .A1(\iro.connect[6] ),
    .A2(_005_));
 sg13g2_a21oi_1 \iro.ro21/_7_  (.A1(\iro.ro21/_1_ ),
    .A2(_005_),
    .Y(\iro.ro21/_0_ ),
    .B1(\iro.ro21/_3_ ));
 sg13g2_nor2_1 \iro.ro21/_8_  (.A(\iro.ro21/_2_ ),
    .B(\iro.ro21/_0_ ),
    .Y(\iro.connect[21] ));
 sg13g2_inv_1 \iro.ro22/_4_  (.Y(\iro.ro22/_1_ ),
    .A(\iro.connect[21] ));
 sg13g2_nor2_1 \iro.ro22/_5_  (.A(net44),
    .B(net22),
    .Y(\iro.ro22/_2_ ));
 sg13g2_o21ai_1 \iro.ro22/_6_  (.B1(net21),
    .Y(\iro.ro22/_3_ ),
    .A1(\iro.connect[5] ),
    .A2(_004_));
 sg13g2_a21oi_1 \iro.ro22/_7_  (.A1(\iro.ro22/_1_ ),
    .A2(_004_),
    .Y(\iro.ro22/_0_ ),
    .B1(\iro.ro22/_3_ ));
 sg13g2_nor2_1 \iro.ro22/_8_  (.A(\iro.ro22/_2_ ),
    .B(\iro.ro22/_0_ ),
    .Y(\iro.connect[22] ));
 sg13g2_inv_1 \iro.ro23/_4_  (.Y(\iro.ro23/_1_ ),
    .A(\iro.connect[22] ));
 sg13g2_nor2_1 \iro.ro23/_5_  (.A(net45),
    .B(net21),
    .Y(\iro.ro23/_2_ ));
 sg13g2_o21ai_1 \iro.ro23/_6_  (.B1(net22),
    .Y(\iro.ro23/_3_ ),
    .A1(\iro.connect[4] ),
    .A2(_003_));
 sg13g2_a21oi_1 \iro.ro23/_7_  (.A1(\iro.ro23/_1_ ),
    .A2(_003_),
    .Y(\iro.ro23/_0_ ),
    .B1(\iro.ro23/_3_ ));
 sg13g2_nor2_1 \iro.ro23/_8_  (.A(\iro.ro23/_2_ ),
    .B(\iro.ro23/_0_ ),
    .Y(\iro.connect[23] ));
 sg13g2_inv_1 \iro.ro24/_4_  (.Y(\iro.ro24/_1_ ),
    .A(\iro.connect[23] ));
 sg13g2_nor2_1 \iro.ro24/_5_  (.A(net46),
    .B(net23),
    .Y(\iro.ro24/_2_ ));
 sg13g2_o21ai_1 \iro.ro24/_6_  (.B1(net21),
    .Y(\iro.ro24/_3_ ),
    .A1(\iro.connect[3] ),
    .A2(_002_));
 sg13g2_a21oi_1 \iro.ro24/_7_  (.A1(\iro.ro24/_1_ ),
    .A2(_002_),
    .Y(\iro.ro24/_0_ ),
    .B1(\iro.ro24/_3_ ));
 sg13g2_nor2_1 \iro.ro24/_8_  (.A(\iro.ro24/_2_ ),
    .B(\iro.ro24/_0_ ),
    .Y(\iro.connect[24] ));
 sg13g2_inv_1 \iro.ro3/_4_  (.Y(\iro.ro3/_1_ ),
    .A(\iro.connect[2] ));
 sg13g2_nor2_1 \iro.ro3/_5_  (.A(net49),
    .B(net23),
    .Y(\iro.ro3/_2_ ));
 sg13g2_o21ai_1 \iro.ro3/_6_  (.B1(net23),
    .Y(\iro.ro3/_3_ ),
    .A1(\iro.connect[2] ),
    .A2(net47));
 sg13g2_a21oi_1 \iro.ro3/_7_  (.A1(\iro.ro3/_1_ ),
    .A2(net48),
    .Y(\iro.ro3/_0_ ),
    .B1(\iro.ro3/_3_ ));
 sg13g2_nor2_2 \iro.ro3/_8_  (.A(\iro.ro3/_2_ ),
    .B(\iro.ro3/_0_ ),
    .Y(\iro.connect[3] ));
 sg13g2_inv_1 \iro.ro4/_4_  (.Y(\iro.ro4/_1_ ),
    .A(\iro.connect[3] ));
 sg13g2_nor2_1 \iro.ro4/_5_  (.A(net52),
    .B(net22),
    .Y(\iro.ro4/_2_ ));
 sg13g2_o21ai_1 \iro.ro4/_6_  (.B1(net22),
    .Y(\iro.ro4/_3_ ),
    .A1(\iro.connect[3] ),
    .A2(net50));
 sg13g2_a21oi_1 \iro.ro4/_7_  (.A1(\iro.ro4/_1_ ),
    .A2(net51),
    .Y(\iro.ro4/_0_ ),
    .B1(\iro.ro4/_3_ ));
 sg13g2_nor2_1 \iro.ro4/_8_  (.A(\iro.ro4/_2_ ),
    .B(\iro.ro4/_0_ ),
    .Y(\iro.connect[4] ));
 sg13g2_inv_1 \iro.ro5/_4_  (.Y(\iro.ro5/_1_ ),
    .A(\iro.connect[4] ));
 sg13g2_nor2_1 \iro.ro5/_5_  (.A(net55),
    .B(net21),
    .Y(\iro.ro5/_2_ ));
 sg13g2_o21ai_1 \iro.ro5/_6_  (.B1(net22),
    .Y(\iro.ro5/_3_ ),
    .A1(\iro.connect[4] ),
    .A2(net53));
 sg13g2_a21oi_1 \iro.ro5/_7_  (.A1(\iro.ro5/_1_ ),
    .A2(net54),
    .Y(\iro.ro5/_0_ ),
    .B1(\iro.ro5/_3_ ));
 sg13g2_nor2_2 \iro.ro5/_8_  (.A(\iro.ro5/_2_ ),
    .B(\iro.ro5/_0_ ),
    .Y(\iro.connect[5] ));
 sg13g2_inv_1 \iro.ro6/_4_  (.Y(\iro.ro6/_1_ ),
    .A(\iro.connect[5] ));
 sg13g2_nor2_1 \iro.ro6/_5_  (.A(net58),
    .B(net21),
    .Y(\iro.ro6/_2_ ));
 sg13g2_o21ai_1 \iro.ro6/_6_  (.B1(net21),
    .Y(\iro.ro6/_3_ ),
    .A1(\iro.connect[5] ),
    .A2(net56));
 sg13g2_a21oi_1 \iro.ro6/_7_  (.A1(\iro.ro6/_1_ ),
    .A2(net57),
    .Y(\iro.ro6/_0_ ),
    .B1(\iro.ro6/_3_ ));
 sg13g2_nor2_2 \iro.ro6/_8_  (.A(\iro.ro6/_2_ ),
    .B(\iro.ro6/_0_ ),
    .Y(\iro.connect[6] ));
 sg13g2_inv_1 \iro.ro7/_4_  (.Y(\iro.ro7/_1_ ),
    .A(\iro.connect[6] ));
 sg13g2_nor2_1 \iro.ro7/_5_  (.A(net61),
    .B(net20),
    .Y(\iro.ro7/_2_ ));
 sg13g2_o21ai_1 \iro.ro7/_6_  (.B1(net20),
    .Y(\iro.ro7/_3_ ),
    .A1(\iro.connect[6] ),
    .A2(net59));
 sg13g2_a21oi_1 \iro.ro7/_7_  (.A1(\iro.ro7/_1_ ),
    .A2(net60),
    .Y(\iro.ro7/_0_ ),
    .B1(\iro.ro7/_3_ ));
 sg13g2_nor2_2 \iro.ro7/_8_  (.A(\iro.ro7/_2_ ),
    .B(\iro.ro7/_0_ ),
    .Y(\iro.connect[7] ));
 sg13g2_inv_1 \iro.ro8/_4_  (.Y(\iro.ro8/_1_ ),
    .A(\iro.connect[7] ));
 sg13g2_nor2_1 \iro.ro8/_5_  (.A(net64),
    .B(net19),
    .Y(\iro.ro8/_2_ ));
 sg13g2_o21ai_1 \iro.ro8/_6_  (.B1(net19),
    .Y(\iro.ro8/_3_ ),
    .A1(\iro.connect[7] ),
    .A2(net62));
 sg13g2_a21oi_1 \iro.ro8/_7_  (.A1(\iro.ro8/_1_ ),
    .A2(net63),
    .Y(\iro.ro8/_0_ ),
    .B1(\iro.ro8/_3_ ));
 sg13g2_nor2_2 \iro.ro8/_8_  (.A(\iro.ro8/_2_ ),
    .B(\iro.ro8/_0_ ),
    .Y(\iro.connect[8] ));
 sg13g2_inv_1 \iro.ro9/_4_  (.Y(\iro.ro9/_1_ ),
    .A(\iro.connect[8] ));
 sg13g2_nor2_1 \iro.ro9/_5_  (.A(net67),
    .B(net20),
    .Y(\iro.ro9/_2_ ));
 sg13g2_o21ai_1 \iro.ro9/_6_  (.B1(net19),
    .Y(\iro.ro9/_3_ ),
    .A1(\iro.connect[8] ),
    .A2(net65));
 sg13g2_a21oi_1 \iro.ro9/_7_  (.A1(\iro.ro9/_1_ ),
    .A2(net66),
    .Y(\iro.ro9/_0_ ),
    .B1(\iro.ro9/_3_ ));
 sg13g2_nor2_2 \iro.ro9/_8_  (.A(\iro.ro9/_2_ ),
    .B(\iro.ro9/_0_ ),
    .Y(\iro.connect[9] ));
 sg13g2_buf_2 fanout17 (.A(net18),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(net20),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(net20),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(\iro.enable ),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(net24),
    .X(net21));
 sg13g2_buf_1 fanout22 (.A(net24),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(net24),
    .X(net23));
 sg13g2_buf_1 fanout24 (.A(\iro.enable ),
    .X(net24));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_tielo \iro.ro0/_6__8  (.L_LO(net8));
 sg13g2_tielo \iro.ro0/_7__9  (.L_LO(net9));
 sg13g2_tielo \iro.ro10/_7__14  (.L_LO(net14));
 sg13g2_tielo \iro.ro11/_7__17  (.L_LO(net25));
 sg13g2_tielo \iro.ro12/_7__20  (.L_LO(net28));
 sg13g2_tielo \iro.ro13/_7__23  (.L_LO(net31));
 sg13g2_tielo \iro.ro2/_7__32  (.L_LO(net40));
 sg13g2_tielo \iro.ro3/_7__40  (.L_LO(net48));
 sg13g2_tielo \iro.ro4/_7__43  (.L_LO(net51));
 sg13g2_tielo \iro.ro5/_7__46  (.L_LO(net54));
 sg13g2_tielo \iro.ro6/_7__49  (.L_LO(net57));
 sg13g2_tielo \iro.ro7/_7__52  (.L_LO(net60));
 sg13g2_tielo \iro.ro8/_7__55  (.L_LO(net63));
 sg13g2_tielo \iro.ro9/_7__58  (.L_LO(net66));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_127 ();
 sg13g2_fill_2 FILLER_28_134 ();
 sg13g2_decap_8 FILLER_28_159 ();
 sg13g2_decap_8 FILLER_28_166 ();
 sg13g2_decap_8 FILLER_28_173 ();
 sg13g2_decap_8 FILLER_28_180 ();
 sg13g2_decap_8 FILLER_28_187 ();
 sg13g2_decap_8 FILLER_28_194 ();
 sg13g2_decap_8 FILLER_28_201 ();
 sg13g2_decap_8 FILLER_28_208 ();
 sg13g2_decap_8 FILLER_28_215 ();
 sg13g2_decap_8 FILLER_28_222 ();
 sg13g2_decap_8 FILLER_28_229 ();
 sg13g2_decap_8 FILLER_28_236 ();
 sg13g2_decap_8 FILLER_28_243 ();
 sg13g2_decap_8 FILLER_28_250 ();
 sg13g2_decap_8 FILLER_28_257 ();
 sg13g2_decap_8 FILLER_28_264 ();
 sg13g2_decap_8 FILLER_28_271 ();
 sg13g2_decap_8 FILLER_28_278 ();
 sg13g2_decap_8 FILLER_28_285 ();
 sg13g2_decap_8 FILLER_28_292 ();
 sg13g2_decap_8 FILLER_28_299 ();
 sg13g2_decap_8 FILLER_28_306 ();
 sg13g2_decap_8 FILLER_28_313 ();
 sg13g2_decap_8 FILLER_28_320 ();
 sg13g2_decap_8 FILLER_28_327 ();
 sg13g2_decap_8 FILLER_28_334 ();
 sg13g2_decap_8 FILLER_28_341 ();
 sg13g2_decap_8 FILLER_28_348 ();
 sg13g2_decap_8 FILLER_28_355 ();
 sg13g2_decap_8 FILLER_28_362 ();
 sg13g2_decap_8 FILLER_28_369 ();
 sg13g2_decap_8 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_28_383 ();
 sg13g2_decap_8 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_fill_2 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_107 ();
 sg13g2_decap_4 FILLER_29_132 ();
 sg13g2_decap_4 FILLER_29_140 ();
 sg13g2_fill_2 FILLER_29_144 ();
 sg13g2_decap_4 FILLER_29_159 ();
 sg13g2_fill_1 FILLER_29_163 ();
 sg13g2_decap_8 FILLER_29_181 ();
 sg13g2_decap_8 FILLER_29_188 ();
 sg13g2_decap_8 FILLER_29_195 ();
 sg13g2_decap_8 FILLER_29_202 ();
 sg13g2_decap_8 FILLER_29_209 ();
 sg13g2_decap_8 FILLER_29_216 ();
 sg13g2_decap_8 FILLER_29_223 ();
 sg13g2_decap_8 FILLER_29_230 ();
 sg13g2_decap_8 FILLER_29_237 ();
 sg13g2_decap_8 FILLER_29_244 ();
 sg13g2_decap_8 FILLER_29_251 ();
 sg13g2_decap_8 FILLER_29_258 ();
 sg13g2_decap_8 FILLER_29_265 ();
 sg13g2_decap_8 FILLER_29_272 ();
 sg13g2_decap_8 FILLER_29_279 ();
 sg13g2_decap_8 FILLER_29_286 ();
 sg13g2_decap_8 FILLER_29_293 ();
 sg13g2_decap_8 FILLER_29_300 ();
 sg13g2_decap_8 FILLER_29_307 ();
 sg13g2_decap_8 FILLER_29_314 ();
 sg13g2_decap_8 FILLER_29_321 ();
 sg13g2_decap_8 FILLER_29_328 ();
 sg13g2_decap_8 FILLER_29_335 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_decap_8 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_decap_8 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_29_370 ();
 sg13g2_decap_8 FILLER_29_377 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_4 FILLER_30_91 ();
 sg13g2_fill_2 FILLER_30_95 ();
 sg13g2_decap_8 FILLER_30_101 ();
 sg13g2_fill_2 FILLER_30_108 ();
 sg13g2_fill_1 FILLER_30_110 ();
 sg13g2_decap_4 FILLER_30_115 ();
 sg13g2_fill_2 FILLER_30_127 ();
 sg13g2_fill_2 FILLER_30_143 ();
 sg13g2_fill_2 FILLER_30_162 ();
 sg13g2_fill_1 FILLER_30_164 ();
 sg13g2_fill_2 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_109 ();
 sg13g2_fill_2 FILLER_31_134 ();
 sg13g2_fill_1 FILLER_31_136 ();
 sg13g2_fill_2 FILLER_31_148 ();
 sg13g2_fill_1 FILLER_31_150 ();
 sg13g2_fill_2 FILLER_31_172 ();
 sg13g2_fill_1 FILLER_31_174 ();
 sg13g2_decap_8 FILLER_31_179 ();
 sg13g2_fill_1 FILLER_31_186 ();
 sg13g2_decap_8 FILLER_31_197 ();
 sg13g2_decap_8 FILLER_31_204 ();
 sg13g2_decap_8 FILLER_31_211 ();
 sg13g2_decap_8 FILLER_31_218 ();
 sg13g2_decap_8 FILLER_31_225 ();
 sg13g2_decap_8 FILLER_31_232 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_decap_8 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_decap_8 FILLER_31_260 ();
 sg13g2_decap_8 FILLER_31_267 ();
 sg13g2_decap_8 FILLER_31_274 ();
 sg13g2_decap_8 FILLER_31_281 ();
 sg13g2_decap_8 FILLER_31_288 ();
 sg13g2_decap_8 FILLER_31_295 ();
 sg13g2_decap_8 FILLER_31_302 ();
 sg13g2_decap_8 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_316 ();
 sg13g2_decap_8 FILLER_31_323 ();
 sg13g2_decap_8 FILLER_31_330 ();
 sg13g2_decap_8 FILLER_31_337 ();
 sg13g2_decap_8 FILLER_31_344 ();
 sg13g2_decap_8 FILLER_31_351 ();
 sg13g2_decap_8 FILLER_31_358 ();
 sg13g2_decap_8 FILLER_31_365 ();
 sg13g2_decap_8 FILLER_31_372 ();
 sg13g2_decap_8 FILLER_31_379 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_decap_8 FILLER_31_393 ();
 sg13g2_decap_8 FILLER_31_400 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_96 ();
 sg13g2_fill_2 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_108 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_135 ();
 sg13g2_fill_2 FILLER_32_150 ();
 sg13g2_fill_1 FILLER_32_152 ();
 sg13g2_fill_2 FILLER_32_157 ();
 sg13g2_fill_1 FILLER_32_159 ();
 sg13g2_fill_2 FILLER_32_163 ();
 sg13g2_fill_1 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_204 ();
 sg13g2_decap_8 FILLER_32_211 ();
 sg13g2_decap_8 FILLER_32_218 ();
 sg13g2_decap_8 FILLER_32_225 ();
 sg13g2_decap_8 FILLER_32_232 ();
 sg13g2_decap_8 FILLER_32_239 ();
 sg13g2_decap_8 FILLER_32_246 ();
 sg13g2_decap_8 FILLER_32_253 ();
 sg13g2_decap_8 FILLER_32_260 ();
 sg13g2_decap_8 FILLER_32_267 ();
 sg13g2_decap_8 FILLER_32_274 ();
 sg13g2_decap_8 FILLER_32_281 ();
 sg13g2_decap_8 FILLER_32_288 ();
 sg13g2_decap_8 FILLER_32_295 ();
 sg13g2_decap_8 FILLER_32_302 ();
 sg13g2_decap_8 FILLER_32_309 ();
 sg13g2_decap_8 FILLER_32_316 ();
 sg13g2_decap_8 FILLER_32_323 ();
 sg13g2_decap_8 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_decap_8 FILLER_32_351 ();
 sg13g2_decap_8 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_91 ();
 sg13g2_fill_1 FILLER_33_106 ();
 sg13g2_fill_1 FILLER_33_112 ();
 sg13g2_decap_4 FILLER_33_121 ();
 sg13g2_fill_2 FILLER_33_125 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_fill_1 FILLER_33_150 ();
 sg13g2_fill_2 FILLER_33_156 ();
 sg13g2_fill_1 FILLER_33_158 ();
 sg13g2_decap_8 FILLER_33_179 ();
 sg13g2_fill_2 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_199 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_decap_4 FILLER_33_213 ();
 sg13g2_fill_1 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_221 ();
 sg13g2_decap_8 FILLER_33_228 ();
 sg13g2_decap_8 FILLER_33_235 ();
 sg13g2_decap_8 FILLER_33_242 ();
 sg13g2_decap_8 FILLER_33_249 ();
 sg13g2_decap_8 FILLER_33_256 ();
 sg13g2_decap_8 FILLER_33_263 ();
 sg13g2_decap_8 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_decap_8 FILLER_33_284 ();
 sg13g2_decap_8 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_decap_8 FILLER_33_305 ();
 sg13g2_decap_8 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_319 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_4 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_88 ();
 sg13g2_fill_2 FILLER_34_101 ();
 sg13g2_fill_1 FILLER_34_103 ();
 sg13g2_fill_2 FILLER_34_129 ();
 sg13g2_fill_1 FILLER_34_131 ();
 sg13g2_decap_4 FILLER_34_153 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_fill_2 FILLER_34_174 ();
 sg13g2_fill_1 FILLER_34_176 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_decap_8 FILLER_34_232 ();
 sg13g2_decap_8 FILLER_34_239 ();
 sg13g2_decap_8 FILLER_34_246 ();
 sg13g2_decap_8 FILLER_34_253 ();
 sg13g2_decap_8 FILLER_34_260 ();
 sg13g2_decap_8 FILLER_34_267 ();
 sg13g2_decap_8 FILLER_34_274 ();
 sg13g2_decap_8 FILLER_34_281 ();
 sg13g2_decap_8 FILLER_34_288 ();
 sg13g2_decap_8 FILLER_34_295 ();
 sg13g2_decap_8 FILLER_34_302 ();
 sg13g2_decap_8 FILLER_34_309 ();
 sg13g2_decap_8 FILLER_34_316 ();
 sg13g2_decap_8 FILLER_34_323 ();
 sg13g2_decap_8 FILLER_34_330 ();
 sg13g2_decap_8 FILLER_34_337 ();
 sg13g2_decap_8 FILLER_34_344 ();
 sg13g2_decap_8 FILLER_34_351 ();
 sg13g2_decap_8 FILLER_34_358 ();
 sg13g2_decap_8 FILLER_34_365 ();
 sg13g2_decap_8 FILLER_34_372 ();
 sg13g2_decap_8 FILLER_34_379 ();
 sg13g2_decap_8 FILLER_34_386 ();
 sg13g2_decap_8 FILLER_34_393 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_4 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_88 ();
 sg13g2_fill_1 FILLER_35_102 ();
 sg13g2_decap_4 FILLER_35_115 ();
 sg13g2_fill_1 FILLER_35_119 ();
 sg13g2_fill_2 FILLER_35_124 ();
 sg13g2_fill_1 FILLER_35_134 ();
 sg13g2_decap_8 FILLER_35_143 ();
 sg13g2_decap_4 FILLER_35_150 ();
 sg13g2_fill_1 FILLER_35_162 ();
 sg13g2_decap_4 FILLER_35_181 ();
 sg13g2_fill_1 FILLER_35_185 ();
 sg13g2_decap_8 FILLER_35_198 ();
 sg13g2_fill_2 FILLER_35_205 ();
 sg13g2_fill_1 FILLER_35_212 ();
 sg13g2_decap_8 FILLER_35_234 ();
 sg13g2_decap_8 FILLER_35_241 ();
 sg13g2_decap_8 FILLER_35_248 ();
 sg13g2_decap_8 FILLER_35_255 ();
 sg13g2_decap_8 FILLER_35_262 ();
 sg13g2_decap_8 FILLER_35_269 ();
 sg13g2_decap_8 FILLER_35_276 ();
 sg13g2_decap_8 FILLER_35_283 ();
 sg13g2_decap_8 FILLER_35_290 ();
 sg13g2_decap_8 FILLER_35_297 ();
 sg13g2_decap_8 FILLER_35_304 ();
 sg13g2_decap_8 FILLER_35_311 ();
 sg13g2_decap_8 FILLER_35_318 ();
 sg13g2_decap_8 FILLER_35_325 ();
 sg13g2_decap_8 FILLER_35_332 ();
 sg13g2_decap_8 FILLER_35_339 ();
 sg13g2_decap_8 FILLER_35_346 ();
 sg13g2_decap_8 FILLER_35_353 ();
 sg13g2_decap_8 FILLER_35_360 ();
 sg13g2_decap_8 FILLER_35_367 ();
 sg13g2_decap_8 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_4 FILLER_36_91 ();
 sg13g2_fill_2 FILLER_36_95 ();
 sg13g2_fill_2 FILLER_36_118 ();
 sg13g2_fill_1 FILLER_36_120 ();
 sg13g2_decap_4 FILLER_36_125 ();
 sg13g2_fill_1 FILLER_36_145 ();
 sg13g2_decap_8 FILLER_36_150 ();
 sg13g2_fill_1 FILLER_36_157 ();
 sg13g2_decap_4 FILLER_36_202 ();
 sg13g2_decap_4 FILLER_36_210 ();
 sg13g2_fill_2 FILLER_36_214 ();
 sg13g2_decap_8 FILLER_36_232 ();
 sg13g2_decap_8 FILLER_36_239 ();
 sg13g2_decap_8 FILLER_36_246 ();
 sg13g2_decap_8 FILLER_36_253 ();
 sg13g2_decap_8 FILLER_36_260 ();
 sg13g2_decap_8 FILLER_36_267 ();
 sg13g2_decap_8 FILLER_36_274 ();
 sg13g2_decap_8 FILLER_36_281 ();
 sg13g2_decap_8 FILLER_36_288 ();
 sg13g2_decap_8 FILLER_36_295 ();
 sg13g2_decap_8 FILLER_36_302 ();
 sg13g2_decap_8 FILLER_36_309 ();
 sg13g2_decap_8 FILLER_36_316 ();
 sg13g2_decap_8 FILLER_36_323 ();
 sg13g2_decap_8 FILLER_36_330 ();
 sg13g2_decap_8 FILLER_36_337 ();
 sg13g2_decap_8 FILLER_36_344 ();
 sg13g2_decap_8 FILLER_36_351 ();
 sg13g2_decap_8 FILLER_36_358 ();
 sg13g2_decap_8 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_4 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_102 ();
 sg13g2_decap_8 FILLER_37_108 ();
 sg13g2_fill_1 FILLER_37_115 ();
 sg13g2_fill_2 FILLER_37_120 ();
 sg13g2_decap_8 FILLER_37_157 ();
 sg13g2_decap_4 FILLER_37_164 ();
 sg13g2_fill_2 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_174 ();
 sg13g2_fill_1 FILLER_37_181 ();
 sg13g2_fill_1 FILLER_37_206 ();
 sg13g2_fill_2 FILLER_37_211 ();
 sg13g2_decap_8 FILLER_37_234 ();
 sg13g2_decap_8 FILLER_37_241 ();
 sg13g2_decap_8 FILLER_37_248 ();
 sg13g2_decap_8 FILLER_37_255 ();
 sg13g2_decap_8 FILLER_37_262 ();
 sg13g2_decap_8 FILLER_37_269 ();
 sg13g2_decap_8 FILLER_37_276 ();
 sg13g2_decap_8 FILLER_37_283 ();
 sg13g2_decap_8 FILLER_37_290 ();
 sg13g2_decap_8 FILLER_37_297 ();
 sg13g2_decap_8 FILLER_37_304 ();
 sg13g2_decap_8 FILLER_37_311 ();
 sg13g2_decap_8 FILLER_37_318 ();
 sg13g2_decap_8 FILLER_37_325 ();
 sg13g2_decap_8 FILLER_37_332 ();
 sg13g2_decap_8 FILLER_37_339 ();
 sg13g2_decap_8 FILLER_37_346 ();
 sg13g2_decap_8 FILLER_37_353 ();
 sg13g2_decap_8 FILLER_37_360 ();
 sg13g2_decap_8 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_374 ();
 sg13g2_decap_8 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_123 ();
 sg13g2_fill_2 FILLER_38_130 ();
 sg13g2_fill_2 FILLER_38_136 ();
 sg13g2_fill_1 FILLER_38_138 ();
 sg13g2_decap_8 FILLER_38_151 ();
 sg13g2_decap_8 FILLER_38_158 ();
 sg13g2_decap_8 FILLER_38_165 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_decap_4 FILLER_38_186 ();
 sg13g2_fill_1 FILLER_38_190 ();
 sg13g2_decap_8 FILLER_38_211 ();
 sg13g2_decap_8 FILLER_38_234 ();
 sg13g2_decap_8 FILLER_38_241 ();
 sg13g2_decap_8 FILLER_38_248 ();
 sg13g2_decap_8 FILLER_38_255 ();
 sg13g2_decap_8 FILLER_38_262 ();
 sg13g2_decap_8 FILLER_38_269 ();
 sg13g2_decap_8 FILLER_38_276 ();
 sg13g2_decap_8 FILLER_38_283 ();
 sg13g2_decap_8 FILLER_38_290 ();
 sg13g2_decap_8 FILLER_38_297 ();
 sg13g2_decap_8 FILLER_38_304 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_decap_8 FILLER_38_341 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_decap_4 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_4 FILLER_38_386 ();
 sg13g2_fill_2 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net68;
 assign uio_oe[1] = net69;
 assign uio_oe[2] = net70;
 assign uio_oe[3] = net71;
 assign uio_oe[4] = net72;
 assign uio_oe[5] = net73;
 assign uio_oe[6] = net74;
 assign uio_oe[7] = net75;
endmodule

module tt_um_faramire_stopwatch (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \SPI_driver1.Cs ;
 wire \SPI_driver1.Mosi ;
 wire \SPI_driver1.SPI_Master1.count_bit[0] ;
 wire \SPI_driver1.SPI_Master1.count_bit[1] ;
 wire \SPI_driver1.SPI_Master1.count_bit[2] ;
 wire \SPI_driver1.SPI_Master1.count_bit[3] ;
 wire \SPI_driver1.SPI_Master1.count_word[0] ;
 wire \SPI_driver1.SPI_Master1.count_word[1] ;
 wire \SPI_driver1.SPI_Master1.count_word[2] ;
 wire \SPI_driver1.SPI_Master1.count_word[3] ;
 wire \SPI_driver1.SPI_Master1.report_ready ;
 wire \SPI_driver1.SPI_Master1.res ;
 wire \SPI_driver1.SPI_Master1.sclk ;
 wire \SPI_driver1.SPI_Master1.send_order ;
 wire \SPI_driver1.SPI_Master1.state[0] ;
 wire \SPI_driver1.SPI_Master1.state[1] ;
 wire \SPI_driver1.SPI_Master1.state[2] ;
 wire \SPI_driver1.SPI_Master1.word_in[0] ;
 wire \SPI_driver1.SPI_Master1.word_in[10] ;
 wire \SPI_driver1.SPI_Master1.word_in[11] ;
 wire \SPI_driver1.SPI_Master1.word_in[12] ;
 wire \SPI_driver1.SPI_Master1.word_in[13] ;
 wire \SPI_driver1.SPI_Master1.word_in[14] ;
 wire \SPI_driver1.SPI_Master1.word_in[15] ;
 wire \SPI_driver1.SPI_Master1.word_in[1] ;
 wire \SPI_driver1.SPI_Master1.word_in[2] ;
 wire \SPI_driver1.SPI_Master1.word_in[3] ;
 wire \SPI_driver1.SPI_Master1.word_in[4] ;
 wire \SPI_driver1.SPI_Master1.word_in[5] ;
 wire \SPI_driver1.SPI_Master1.word_in[6] ;
 wire \SPI_driver1.SPI_Master1.word_in[7] ;
 wire \SPI_driver1.SPI_Master1.word_in[8] ;
 wire \SPI_driver1.SPI_Master1.word_in[9] ;
 wire \SPI_driver1.SPI_Master1.word_out[0] ;
 wire \SPI_driver1.SPI_Master1.word_out[10] ;
 wire \SPI_driver1.SPI_Master1.word_out[11] ;
 wire \SPI_driver1.SPI_Master1.word_out[12] ;
 wire \SPI_driver1.SPI_Master1.word_out[13] ;
 wire \SPI_driver1.SPI_Master1.word_out[14] ;
 wire \SPI_driver1.SPI_Master1.word_out[15] ;
 wire \SPI_driver1.SPI_Master1.word_out[1] ;
 wire \SPI_driver1.SPI_Master1.word_out[2] ;
 wire \SPI_driver1.SPI_Master1.word_out[3] ;
 wire \SPI_driver1.SPI_Master1.word_out[4] ;
 wire \SPI_driver1.SPI_Master1.word_out[5] ;
 wire \SPI_driver1.SPI_Master1.word_out[6] ;
 wire \SPI_driver1.SPI_Master1.word_out[7] ;
 wire \SPI_driver1.SPI_Master1.word_out[8] ;
 wire \SPI_driver1.SPI_Master1.word_out[9] ;
 wire \SPI_driver1.ces_0X[0] ;
 wire \SPI_driver1.ces_0X[1] ;
 wire \SPI_driver1.ces_0X[2] ;
 wire \SPI_driver1.ces_0X[3] ;
 wire \SPI_driver1.ces_X0[0] ;
 wire \SPI_driver1.ces_X0[1] ;
 wire \SPI_driver1.ces_X0[2] ;
 wire \SPI_driver1.ces_X0[3] ;
 wire \SPI_driver1.clk_div ;
 wire \SPI_driver1.digit_count[0] ;
 wire \SPI_driver1.digit_count[1] ;
 wire \SPI_driver1.digit_count[2] ;
 wire \SPI_driver1.digit_count[3] ;
 wire \SPI_driver1.digit_count[4] ;
 wire \SPI_driver1.digit_count[5] ;
 wire \SPI_driver1.digit_count[6] ;
 wire \SPI_driver1.ena ;
 wire \SPI_driver1.min_0X[0] ;
 wire \SPI_driver1.min_0X[1] ;
 wire \SPI_driver1.min_0X[2] ;
 wire \SPI_driver1.min_0X[3] ;
 wire \SPI_driver1.min_X0[0] ;
 wire \SPI_driver1.min_X0[1] ;
 wire \SPI_driver1.min_X0[2] ;
 wire \SPI_driver1.sec_0X[0] ;
 wire \SPI_driver1.sec_0X[1] ;
 wire \SPI_driver1.sec_0X[2] ;
 wire \SPI_driver1.sec_0X[3] ;
 wire \SPI_driver1.sec_X0[0] ;
 wire \SPI_driver1.sec_X0[1] ;
 wire \SPI_driver1.sec_X0[2] ;
 wire \SPI_driver1.sent_BCD ;
 wire \SPI_driver1.sent_LUX ;
 wire \SPI_driver1.sent_PWR ;
 wire \SPI_driver1.sent_SCN ;
 wire \SPI_driver1.sent_TST ;
 wire \SPI_driver1.state[0] ;
 wire \SPI_driver1.state[1] ;
 wire \SPI_driver1.state[2] ;
 wire \SPI_driver1.state[3] ;
 wire \SPI_driver1.wait_count[0] ;
 wire \SPI_driver1.wait_count[1] ;
 wire \SPI_driver1.wait_count[2] ;
 wire \SPI_driver1.wait_count[3] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire clknet_0_clk;
 wire _0769_;
 wire \clockDivider1.counter[0] ;
 wire \clockDivider1.counter[10] ;
 wire \clockDivider1.counter[11] ;
 wire \clockDivider1.counter[12] ;
 wire \clockDivider1.counter[13] ;
 wire \clockDivider1.counter[1] ;
 wire \clockDivider1.counter[2] ;
 wire \clockDivider1.counter[3] ;
 wire \clockDivider1.counter[4] ;
 wire \clockDivider1.counter[5] ;
 wire \clockDivider1.counter[6] ;
 wire \clockDivider1.counter[7] ;
 wire \clockDivider1.counter[8] ;
 wire \clockDivider1.counter[9] ;
 wire \clockDivider1.ena ;
 wire \counter_chain1.ces_X0_ena ;
 wire \counter_chain1.inst_ces_X0.max ;
 wire \counter_chain1.inst_min_0X.max ;
 wire \counter_chain1.inst_sec_0X.max ;
 wire \counter_chain1.inst_sec_X0.max ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;

 sg13g2_inv_1 _0770_ (.Y(_0127_),
    .A(net135));
 sg13g2_inv_1 _0771_ (.Y(_0128_),
    .A(net326));
 sg13g2_inv_1 _0772_ (.Y(_0129_),
    .A(net177));
 sg13g2_inv_1 _0773_ (.Y(_0130_),
    .A(net140));
 sg13g2_inv_1 _0774_ (.Y(_0131_),
    .A(net318));
 sg13g2_inv_1 _0775_ (.Y(_0132_),
    .A(net285));
 sg13g2_inv_1 _0776_ (.Y(_0133_),
    .A(\SPI_driver1.SPI_Master1.report_ready ));
 sg13g2_inv_1 _0777_ (.Y(_0134_),
    .A(net181));
 sg13g2_inv_1 _0778_ (.Y(_0135_),
    .A(net200));
 sg13g2_inv_1 _0779_ (.Y(_0136_),
    .A(\SPI_driver1.SPI_Master1.send_order ));
 sg13g2_inv_1 _0780_ (.Y(_0137_),
    .A(\SPI_driver1.wait_count[0] ));
 sg13g2_inv_1 _0781_ (.Y(_0138_),
    .A(net198));
 sg13g2_inv_1 _0782_ (.Y(_0139_),
    .A(_0025_));
 sg13g2_inv_1 _0783_ (.Y(_0140_),
    .A(net300));
 sg13g2_inv_2 _0784_ (.Y(_0141_),
    .A(net1));
 sg13g2_inv_1 _0785_ (.Y(_0142_),
    .A(\SPI_driver1.digit_count[2] ));
 sg13g2_inv_1 _0786_ (.Y(_0143_),
    .A(\SPI_driver1.digit_count[1] ));
 sg13g2_inv_1 _0787_ (.Y(_0144_),
    .A(net291));
 sg13g2_inv_1 _0788_ (.Y(_0145_),
    .A(\SPI_driver1.digit_count[5] ));
 sg13g2_inv_1 _0789_ (.Y(_0146_),
    .A(net314));
 sg13g2_inv_1 _0790_ (.Y(_0147_),
    .A(net268));
 sg13g2_inv_1 _0791_ (.Y(_0148_),
    .A(net202));
 sg13g2_inv_2 _0792_ (.Y(_0149_),
    .A(net142));
 sg13g2_inv_1 _0793_ (.Y(_0150_),
    .A(\SPI_driver1.sent_TST ));
 sg13g2_inv_1 _0794_ (.Y(_0151_),
    .A(\SPI_driver1.SPI_Master1.word_out[0] ));
 sg13g2_and2_1 _0795_ (.A(net150),
    .B(net141),
    .X(_0152_));
 sg13g2_nand2_1 _0796_ (.Y(_0153_),
    .A(net150),
    .B(net141));
 sg13g2_nor2_1 _0797_ (.A(\SPI_driver1.SPI_Master1.state[0] ),
    .B(_0153_),
    .Y(_0154_));
 sg13g2_o21ai_1 _0798_ (.B1(net303),
    .Y(_0155_),
    .A1(net200),
    .A2(_0153_));
 sg13g2_nand3_1 _0799_ (.B(net297),
    .C(net141),
    .A(net200),
    .Y(_0156_));
 sg13g2_nand2_1 _0800_ (.Y(_0157_),
    .A(net150),
    .B(\SPI_driver1.SPI_Master1.count_bit[3] ));
 sg13g2_nand2_1 _0801_ (.Y(_0158_),
    .A(net249),
    .B(_0152_));
 sg13g2_nand3_1 _0802_ (.B(_0156_),
    .C(_0158_),
    .A(_0155_),
    .Y(_0001_));
 sg13g2_nor2_1 _0803_ (.A(net307),
    .B(\SPI_driver1.SPI_Master1.count_word[0] ),
    .Y(_0159_));
 sg13g2_nor3_2 _0804_ (.A(\SPI_driver1.SPI_Master1.count_word[1] ),
    .B(\SPI_driver1.SPI_Master1.count_word[0] ),
    .C(net266),
    .Y(_0160_));
 sg13g2_nand2b_1 _0805_ (.Y(_0161_),
    .B(_0160_),
    .A_N(net238));
 sg13g2_nor2_1 _0806_ (.A(net204),
    .B(_0157_),
    .Y(_0162_));
 sg13g2_nand2b_1 _0807_ (.Y(_0163_),
    .B(net150),
    .A_N(\SPI_driver1.SPI_Master1.count_bit[3] ));
 sg13g2_inv_1 _0808_ (.Y(_0164_),
    .A(_0163_));
 sg13g2_a22oi_1 _0809_ (.Y(_0165_),
    .B1(_0164_),
    .B2(net141),
    .A2(net205),
    .A1(_0161_));
 sg13g2_nand2_1 _0810_ (.Y(_0006_),
    .A(_0156_),
    .B(net312));
 sg13g2_and3_1 _0811_ (.X(_0166_),
    .A(\SPI_driver1.SPI_Master1.state[0] ),
    .B(_0136_),
    .C(net141));
 sg13g2_or3_1 _0812_ (.A(net215),
    .B(net204),
    .C(_0166_),
    .X(_0005_));
 sg13g2_nor2b_2 _0813_ (.A(net201),
    .B_N(_0156_),
    .Y(_0167_));
 sg13g2_o21ai_1 _0814_ (.B1(_0156_),
    .Y(_0168_),
    .A1(\SPI_driver1.SPI_Master1.state[0] ),
    .A2(_0153_));
 sg13g2_a22oi_1 _0815_ (.Y(_0169_),
    .B1(_0167_),
    .B2(net249),
    .A2(_0152_),
    .A1(net198));
 sg13g2_inv_1 _0816_ (.Y(_0004_),
    .A(_0169_));
 sg13g2_a22oi_1 _0817_ (.Y(_0170_),
    .B1(_0167_),
    .B2(net194),
    .A2(_0152_),
    .A1(\SPI_driver1.SPI_Master1.count_bit[0] ));
 sg13g2_inv_1 _0818_ (.Y(_0003_),
    .A(net195));
 sg13g2_nor2b_2 _0819_ (.A(net133),
    .B_N(net131),
    .Y(_0171_));
 sg13g2_nand2b_2 _0820_ (.Y(_0172_),
    .B(net131),
    .A_N(net132));
 sg13g2_nor2b_2 _0821_ (.A(net126),
    .B_N(net129),
    .Y(_0173_));
 sg13g2_nand2b_2 _0822_ (.Y(_0174_),
    .B(net129),
    .A_N(net126));
 sg13g2_nor2_1 _0823_ (.A(_0172_),
    .B(_0174_),
    .Y(_0175_));
 sg13g2_nand2_1 _0824_ (.Y(_0176_),
    .A(_0171_),
    .B(_0173_));
 sg13g2_nor3_2 _0825_ (.A(_0133_),
    .B(_0172_),
    .C(_0174_),
    .Y(_0177_));
 sg13g2_nand3_1 _0826_ (.B(_0171_),
    .C(_0173_),
    .A(net270),
    .Y(_0178_));
 sg13g2_nand2_1 _0827_ (.Y(_0179_),
    .A(net300),
    .B(_0177_));
 sg13g2_nand3b_1 _0828_ (.B(net131),
    .C(net127),
    .Y(_0180_),
    .A_N(net133));
 sg13g2_nor2_1 _0829_ (.A(net130),
    .B(_0180_),
    .Y(_0181_));
 sg13g2_nor2_1 _0830_ (.A(_0128_),
    .B(_0130_),
    .Y(_0182_));
 sg13g2_nand2_1 _0831_ (.Y(_0183_),
    .A(\SPI_driver1.ena ),
    .B(net140));
 sg13g2_nor3_2 _0832_ (.A(net129),
    .B(_0180_),
    .C(_0182_),
    .Y(_0184_));
 sg13g2_and2_2 _0833_ (.A(net130),
    .B(net126),
    .X(_0185_));
 sg13g2_nand2_2 _0834_ (.Y(_0186_),
    .A(net129),
    .B(net127));
 sg13g2_nor2_1 _0835_ (.A(net129),
    .B(net126),
    .Y(_0187_));
 sg13g2_or2_1 _0836_ (.X(_0188_),
    .B(net126),
    .A(net130));
 sg13g2_nor3_1 _0837_ (.A(_0172_),
    .B(_0185_),
    .C(_0187_),
    .Y(_0189_));
 sg13g2_o21ai_1 _0838_ (.B1(_0189_),
    .Y(_0190_),
    .A1(net145),
    .A2(_0176_));
 sg13g2_o21ai_1 _0839_ (.B1(net156),
    .Y(_0191_),
    .A1(_0184_),
    .A2(_0190_));
 sg13g2_o21ai_1 _0840_ (.B1(net301),
    .Y(_0009_),
    .A1(_0142_),
    .A2(_0191_));
 sg13g2_nand2_1 _0841_ (.Y(_0192_),
    .A(net291),
    .B(_0177_));
 sg13g2_o21ai_1 _0842_ (.B1(net292),
    .Y(_0008_),
    .A1(_0143_),
    .A2(_0191_));
 sg13g2_nand2_2 _0843_ (.Y(_0193_),
    .A(_0181_),
    .B(_0182_));
 sg13g2_nand3_1 _0844_ (.B(net207),
    .C(_0193_),
    .A(net156),
    .Y(_0194_));
 sg13g2_o21ai_1 _0845_ (.B1(_0194_),
    .Y(_0010_),
    .A1(_0145_),
    .A2(_0178_));
 sg13g2_a22oi_1 _0846_ (.Y(_0195_),
    .B1(_0167_),
    .B2(net198),
    .A2(_0152_),
    .A1(net194));
 sg13g2_inv_1 _0847_ (.Y(_0002_),
    .A(_0195_));
 sg13g2_nand2_1 _0848_ (.Y(_0196_),
    .A(net304),
    .B(_0177_));
 sg13g2_o21ai_1 _0849_ (.B1(net305),
    .Y(_0011_),
    .A1(_0140_),
    .A2(_0191_));
 sg13g2_nand2_1 _0850_ (.Y(_0197_),
    .A(net294),
    .B(_0177_));
 sg13g2_o21ai_1 _0851_ (.B1(net295),
    .Y(_0012_),
    .A1(_0145_),
    .A2(_0191_));
 sg13g2_nand2_1 _0852_ (.Y(_0198_),
    .A(net313),
    .B(_0177_));
 sg13g2_o21ai_1 _0853_ (.B1(_0198_),
    .Y(_0013_),
    .A1(_0144_),
    .A2(_0191_));
 sg13g2_nand3b_1 _0854_ (.B(net144),
    .C(net130),
    .Y(_0199_),
    .A_N(net126));
 sg13g2_nand3_1 _0855_ (.B(_0188_),
    .C(_0199_),
    .A(_0171_),
    .Y(_0200_));
 sg13g2_o21ai_1 _0856_ (.B1(net304),
    .Y(_0201_),
    .A1(_0185_),
    .A2(_0200_));
 sg13g2_nand2b_1 _0857_ (.Y(_0202_),
    .B(_0181_),
    .A_N(net306));
 sg13g2_nand3_1 _0858_ (.B(_0193_),
    .C(_0202_),
    .A(net156),
    .Y(_0203_));
 sg13g2_o21ai_1 _0859_ (.B1(_0203_),
    .Y(_0204_),
    .A1(net207),
    .A2(_0178_));
 sg13g2_nand2_1 _0860_ (.Y(_0007_),
    .A(_0201_),
    .B(_0204_));
 sg13g2_nor2_2 _0861_ (.A(net132),
    .B(net131),
    .Y(_0205_));
 sg13g2_or2_2 _0862_ (.X(_0206_),
    .B(\SPI_driver1.state[2] ),
    .A(net132));
 sg13g2_nor3_2 _0863_ (.A(net129),
    .B(net132),
    .C(net131),
    .Y(_0207_));
 sg13g2_inv_1 _0864_ (.Y(_0208_),
    .A(_0207_));
 sg13g2_nor4_2 _0865_ (.A(net129),
    .B(net127),
    .C(net132),
    .Y(_0209_),
    .D(net131));
 sg13g2_and2_2 _0866_ (.A(net154),
    .B(_0209_),
    .X(_0210_));
 sg13g2_a21o_1 _0867_ (.A2(net154),
    .A1(net141),
    .B1(_0210_),
    .X(_0015_));
 sg13g2_a22oi_1 _0868_ (.Y(_0211_),
    .B1(_0210_),
    .B2(net145),
    .A2(net288),
    .A1(net154));
 sg13g2_inv_1 _0869_ (.Y(_0020_),
    .A(_0211_));
 sg13g2_nand2_1 _0870_ (.Y(_0212_),
    .A(net128),
    .B(_0207_));
 sg13g2_nor2_1 _0871_ (.A(net284),
    .B(_0212_),
    .Y(_0213_));
 sg13g2_nand3b_1 _0872_ (.B(_0207_),
    .C(net128),
    .Y(_0214_),
    .A_N(\SPI_driver1.sent_SCN ));
 sg13g2_a22oi_1 _0873_ (.Y(_0215_),
    .B1(_0213_),
    .B2(net145),
    .A2(net284),
    .A1(net152));
 sg13g2_inv_1 _0874_ (.Y(_0019_),
    .A(_0215_));
 sg13g2_nand2_2 _0875_ (.Y(_0216_),
    .A(_0173_),
    .B(_0205_));
 sg13g2_nor3_2 _0876_ (.A(net310),
    .B(_0174_),
    .C(_0206_),
    .Y(_0217_));
 sg13g2_nand3b_1 _0877_ (.B(_0173_),
    .C(_0205_),
    .Y(_0218_),
    .A_N(\SPI_driver1.sent_LUX ));
 sg13g2_a22oi_1 _0878_ (.Y(_0219_),
    .B1(_0217_),
    .B2(net145),
    .A2(net310),
    .A1(net155));
 sg13g2_inv_1 _0879_ (.Y(_0017_),
    .A(_0219_));
 sg13g2_nand2_1 _0880_ (.Y(_0220_),
    .A(net128),
    .B(_0205_));
 sg13g2_nor2_2 _0881_ (.A(_0186_),
    .B(_0206_),
    .Y(_0221_));
 sg13g2_nor3_2 _0882_ (.A(net299),
    .B(_0186_),
    .C(_0206_),
    .Y(_0222_));
 sg13g2_a22oi_1 _0883_ (.Y(_0223_),
    .B1(_0222_),
    .B2(net145),
    .A2(net299),
    .A1(net154));
 sg13g2_inv_1 _0884_ (.Y(_0016_),
    .A(_0223_));
 sg13g2_nor2_2 _0885_ (.A(_0172_),
    .B(_0188_),
    .Y(_0224_));
 sg13g2_nand2_1 _0886_ (.Y(_0225_),
    .A(_0171_),
    .B(_0187_));
 sg13g2_nor3_2 _0887_ (.A(\SPI_driver1.sent_PWR ),
    .B(_0172_),
    .C(_0188_),
    .Y(_0226_));
 sg13g2_a22oi_1 _0888_ (.Y(_0227_),
    .B1(_0226_),
    .B2(net270),
    .A2(\SPI_driver1.sent_PWR ),
    .A1(net153));
 sg13g2_inv_1 _0889_ (.Y(_0018_),
    .A(net271));
 sg13g2_nand2_1 _0890_ (.Y(_0228_),
    .A(net229),
    .B(net153));
 sg13g2_nor2_2 _0891_ (.A(net142),
    .B(net288),
    .Y(_0229_));
 sg13g2_inv_1 _0892_ (.Y(_0230_),
    .A(_0229_));
 sg13g2_a21oi_1 _0893_ (.A1(_0209_),
    .A2(_0230_),
    .Y(_0231_),
    .B1(_0221_));
 sg13g2_nand3_1 _0894_ (.B(_0216_),
    .C(_0231_),
    .A(_0212_),
    .Y(_0232_));
 sg13g2_or3_1 _0895_ (.A(\SPI_driver1.digit_count[1] ),
    .B(\SPI_driver1.digit_count[6] ),
    .C(\SPI_driver1.digit_count[5] ),
    .X(_0233_));
 sg13g2_nand2_1 _0896_ (.Y(_0234_),
    .A(_0140_),
    .B(_0142_));
 sg13g2_or3_1 _0897_ (.A(\SPI_driver1.digit_count[4] ),
    .B(\SPI_driver1.digit_count[2] ),
    .C(\SPI_driver1.digit_count[0] ),
    .X(_0235_));
 sg13g2_nor2_1 _0898_ (.A(_0233_),
    .B(_0235_),
    .Y(_0236_));
 sg13g2_o21ai_1 _0899_ (.B1(net145),
    .Y(_0237_),
    .A1(_0233_),
    .A2(_0235_));
 sg13g2_nand2_1 _0900_ (.Y(_0238_),
    .A(_0175_),
    .B(_0237_));
 sg13g2_a21oi_1 _0901_ (.A1(net126),
    .A2(net131),
    .Y(_0239_),
    .B1(net132));
 sg13g2_a221oi_1 _0902_ (.B2(_0237_),
    .C1(net132),
    .B1(_0175_),
    .A1(net126),
    .Y(_0240_),
    .A2(net131));
 sg13g2_nand2_1 _0903_ (.Y(_0241_),
    .A(_0238_),
    .B(_0239_));
 sg13g2_nor2_1 _0904_ (.A(_0232_),
    .B(_0241_),
    .Y(_0242_));
 sg13g2_and2_2 _0905_ (.A(_0149_),
    .B(_0222_),
    .X(_0243_));
 sg13g2_a21oi_1 _0906_ (.A1(_0214_),
    .A2(_0218_),
    .Y(_0244_),
    .B1(net142));
 sg13g2_or2_1 _0907_ (.X(_0245_),
    .B(_0244_),
    .A(_0243_));
 sg13g2_nor2_1 _0908_ (.A(_0178_),
    .B(_0236_),
    .Y(_0246_));
 sg13g2_a22oi_1 _0909_ (.Y(_0247_),
    .B1(\SPI_driver1.digit_count[0] ),
    .B2(\SPI_driver1.ces_0X[0] ),
    .A2(\SPI_driver1.digit_count[6] ),
    .A1(\SPI_driver1.sec_X0[0] ));
 sg13g2_a22oi_1 _0910_ (.Y(_0248_),
    .B1(\SPI_driver1.digit_count[5] ),
    .B2(\SPI_driver1.min_X0[0] ),
    .A2(\SPI_driver1.digit_count[4] ),
    .A1(\SPI_driver1.ces_X0[0] ));
 sg13g2_a22oi_1 _0911_ (.Y(_0249_),
    .B1(\SPI_driver1.digit_count[1] ),
    .B2(\SPI_driver1.min_0X[0] ),
    .A2(\SPI_driver1.digit_count[2] ),
    .A1(\SPI_driver1.sec_0X[0] ));
 sg13g2_nand3_1 _0912_ (.B(_0248_),
    .C(_0249_),
    .A(_0247_),
    .Y(_0250_));
 sg13g2_nor2_1 _0913_ (.A(net142),
    .B(\SPI_driver1.sent_PWR ),
    .Y(_0251_));
 sg13g2_o21ai_1 _0914_ (.B1(_0228_),
    .Y(_0252_),
    .A1(net142),
    .A2(net283));
 sg13g2_a221oi_1 _0915_ (.B2(_0224_),
    .C1(_0245_),
    .B1(_0252_),
    .A1(net123),
    .Y(_0253_),
    .A2(_0250_));
 sg13g2_o21ai_1 _0916_ (.B1(_0253_),
    .Y(_0111_),
    .A1(_0228_),
    .A2(_0242_));
 sg13g2_nand2_1 _0917_ (.Y(_0254_),
    .A(net152),
    .B(net253));
 sg13g2_o21ai_1 _0918_ (.B1(_0240_),
    .Y(_0255_),
    .A1(_0225_),
    .A2(_0251_));
 sg13g2_nand3_1 _0919_ (.B(\SPI_driver1.sent_SCN ),
    .C(_0207_),
    .A(net128),
    .Y(_0256_));
 sg13g2_nand3_1 _0920_ (.B(_0173_),
    .C(_0205_),
    .A(\SPI_driver1.sent_LUX ),
    .Y(_0257_));
 sg13g2_nand3_1 _0921_ (.B(net142),
    .C(_0207_),
    .A(net128),
    .Y(_0258_));
 sg13g2_nand3_1 _0922_ (.B(_0173_),
    .C(_0205_),
    .A(net142),
    .Y(_0259_));
 sg13g2_and4_1 _0923_ (.A(_0256_),
    .B(_0257_),
    .C(_0258_),
    .D(_0259_),
    .X(_0260_));
 sg13g2_nand2_1 _0924_ (.Y(_0261_),
    .A(_0231_),
    .B(_0260_));
 sg13g2_nor2_2 _0925_ (.A(_0255_),
    .B(_0261_),
    .Y(_0262_));
 sg13g2_a22oi_1 _0926_ (.Y(_0263_),
    .B1(\SPI_driver1.digit_count[0] ),
    .B2(\SPI_driver1.ces_0X[1] ),
    .A2(\SPI_driver1.digit_count[1] ),
    .A1(\SPI_driver1.min_0X[1] ));
 sg13g2_a22oi_1 _0927_ (.Y(_0264_),
    .B1(\SPI_driver1.digit_count[6] ),
    .B2(\SPI_driver1.sec_X0[1] ),
    .A2(\SPI_driver1.digit_count[2] ),
    .A1(\SPI_driver1.sec_0X[1] ));
 sg13g2_a22oi_1 _0928_ (.Y(_0265_),
    .B1(\SPI_driver1.digit_count[5] ),
    .B2(\SPI_driver1.min_X0[1] ),
    .A2(\SPI_driver1.digit_count[4] ),
    .A1(\SPI_driver1.ces_X0[1] ));
 sg13g2_nand3_1 _0929_ (.B(_0264_),
    .C(_0265_),
    .A(_0263_),
    .Y(_0266_));
 sg13g2_a21oi_1 _0930_ (.A1(net123),
    .A2(_0266_),
    .Y(_0267_),
    .B1(_0243_));
 sg13g2_o21ai_1 _0931_ (.B1(_0267_),
    .Y(_0118_),
    .A1(_0254_),
    .A2(_0262_));
 sg13g2_and2_1 _0932_ (.A(net152),
    .B(net325),
    .X(_0268_));
 sg13g2_o21ai_1 _0933_ (.B1(_0232_),
    .Y(_0269_),
    .A1(_0245_),
    .A2(_0268_));
 sg13g2_a22oi_1 _0934_ (.Y(_0270_),
    .B1(\SPI_driver1.digit_count[0] ),
    .B2(\SPI_driver1.ces_0X[2] ),
    .A2(\SPI_driver1.digit_count[5] ),
    .A1(\SPI_driver1.min_X0[2] ));
 sg13g2_a22oi_1 _0935_ (.Y(_0271_),
    .B1(\SPI_driver1.digit_count[1] ),
    .B2(\SPI_driver1.min_0X[2] ),
    .A2(\SPI_driver1.digit_count[4] ),
    .A1(\SPI_driver1.ces_X0[2] ));
 sg13g2_a22oi_1 _0936_ (.Y(_0272_),
    .B1(\SPI_driver1.digit_count[6] ),
    .B2(\SPI_driver1.sec_X0[2] ),
    .A2(\SPI_driver1.digit_count[2] ),
    .A1(\SPI_driver1.sec_0X[2] ));
 sg13g2_nand3_1 _0937_ (.B(_0271_),
    .C(_0272_),
    .A(_0270_),
    .Y(_0273_));
 sg13g2_a22oi_1 _0938_ (.Y(_0274_),
    .B1(_0273_),
    .B2(net123),
    .A2(_0268_),
    .A1(_0255_));
 sg13g2_nand2_1 _0939_ (.Y(_0119_),
    .A(_0269_),
    .B(_0274_));
 sg13g2_a22oi_1 _0940_ (.Y(_0275_),
    .B1(\SPI_driver1.digit_count[0] ),
    .B2(\SPI_driver1.ces_0X[3] ),
    .A2(\SPI_driver1.digit_count[1] ),
    .A1(\SPI_driver1.min_0X[3] ));
 sg13g2_a22oi_1 _0941_ (.Y(_0276_),
    .B1(\SPI_driver1.digit_count[2] ),
    .B2(\SPI_driver1.sec_0X[3] ),
    .A2(\SPI_driver1.digit_count[4] ),
    .A1(\SPI_driver1.ces_X0[3] ));
 sg13g2_nand2_1 _0942_ (.Y(_0277_),
    .A(_0275_),
    .B(_0276_));
 sg13g2_nand2_1 _0943_ (.Y(_0278_),
    .A(net123),
    .B(_0277_));
 sg13g2_a21oi_1 _0944_ (.A1(net152),
    .A2(net290),
    .Y(_0279_),
    .B1(_0243_));
 sg13g2_o21ai_1 _0945_ (.B1(_0278_),
    .Y(_0120_),
    .A1(_0262_),
    .A2(_0279_));
 sg13g2_a21oi_1 _0946_ (.A1(net152),
    .A2(net259),
    .Y(_0280_),
    .B1(_0243_));
 sg13g2_nor2_1 _0947_ (.A(_0262_),
    .B(_0280_),
    .Y(_0121_));
 sg13g2_a21oi_1 _0948_ (.A1(net152),
    .A2(net262),
    .Y(_0281_),
    .B1(_0243_));
 sg13g2_nor2_1 _0949_ (.A(_0262_),
    .B(_0281_),
    .Y(_0122_));
 sg13g2_nand2_1 _0950_ (.Y(_0282_),
    .A(\SPI_driver1.sent_PWR ),
    .B(_0224_));
 sg13g2_and3_1 _0951_ (.X(_0283_),
    .A(_0240_),
    .B(_0257_),
    .C(_0282_));
 sg13g2_or4_1 _0952_ (.A(_0207_),
    .B(_0217_),
    .C(_0222_),
    .D(_0224_),
    .X(_0284_));
 sg13g2_nand3_1 _0953_ (.B(_0185_),
    .C(_0205_),
    .A(\SPI_driver1.sent_BCD ),
    .Y(_0285_));
 sg13g2_nand2_1 _0954_ (.Y(_0286_),
    .A(_0256_),
    .B(_0285_));
 sg13g2_a221oi_1 _0955_ (.B2(_0133_),
    .C1(_0286_),
    .B1(_0284_),
    .A1(\SPI_driver1.sent_TST ),
    .Y(_0287_),
    .A2(_0209_));
 sg13g2_a21oi_2 _0956_ (.B1(_0141_),
    .Y(_0288_),
    .A2(_0287_),
    .A1(_0283_));
 sg13g2_and2_1 _0957_ (.A(net187),
    .B(_0288_),
    .X(_0123_));
 sg13g2_o21ai_1 _0958_ (.B1(_0177_),
    .Y(_0289_),
    .A1(\SPI_driver1.digit_count[2] ),
    .A2(\SPI_driver1.digit_count[1] ));
 sg13g2_inv_1 _0959_ (.Y(_0290_),
    .A(_0289_));
 sg13g2_a21o_1 _0960_ (.A2(_0288_),
    .A1(net231),
    .B1(_0290_),
    .X(_0124_));
 sg13g2_nand3_1 _0961_ (.B(_0257_),
    .C(_0259_),
    .A(_0220_),
    .Y(_0291_));
 sg13g2_and2_1 _0962_ (.A(net153),
    .B(net322),
    .X(_0292_));
 sg13g2_o21ai_1 _0963_ (.B1(_0292_),
    .Y(_0293_),
    .A1(_0255_),
    .A2(_0291_));
 sg13g2_or2_1 _0964_ (.X(_0294_),
    .B(_0229_),
    .A(net322));
 sg13g2_a221oi_1 _0965_ (.B2(_0210_),
    .C1(_0243_),
    .B1(_0294_),
    .A1(_0149_),
    .Y(_0295_),
    .A2(_0213_));
 sg13g2_nand2b_2 _0966_ (.Y(_0296_),
    .B(_0246_),
    .A_N(net306));
 sg13g2_nand4_1 _0967_ (.B(_0293_),
    .C(_0295_),
    .A(_0289_),
    .Y(_0125_),
    .D(_0296_));
 sg13g2_and2_1 _0968_ (.A(net152),
    .B(net320),
    .X(_0297_));
 sg13g2_nand2_1 _0969_ (.Y(_0298_),
    .A(_0255_),
    .B(_0297_));
 sg13g2_o21ai_1 _0970_ (.B1(_0221_),
    .Y(_0299_),
    .A1(net143),
    .A2(\SPI_driver1.sent_BCD ));
 sg13g2_nand3_1 _0971_ (.B(_0216_),
    .C(_0299_),
    .A(_0212_),
    .Y(_0300_));
 sg13g2_o21ai_1 _0972_ (.B1(_0300_),
    .Y(_0301_),
    .A1(_0244_),
    .A2(_0297_));
 sg13g2_o21ai_1 _0973_ (.B1(net123),
    .Y(_0302_),
    .A1(\SPI_driver1.digit_count[5] ),
    .A2(_0234_));
 sg13g2_o21ai_1 _0974_ (.B1(_0210_),
    .Y(_0303_),
    .A1(net320),
    .A2(_0229_));
 sg13g2_nand4_1 _0975_ (.B(_0301_),
    .C(_0302_),
    .A(_0298_),
    .Y(_0126_),
    .D(_0303_));
 sg13g2_o21ai_1 _0976_ (.B1(_0210_),
    .Y(_0304_),
    .A1(net289),
    .A2(_0229_));
 sg13g2_nand4_1 _0977_ (.B(_0240_),
    .C(_0260_),
    .A(_0225_),
    .Y(_0305_),
    .D(_0299_));
 sg13g2_nand3_1 _0978_ (.B(net289),
    .C(_0305_),
    .A(net152),
    .Y(_0306_));
 sg13g2_a22oi_1 _0979_ (.Y(_0307_),
    .B1(_0233_),
    .B2(_0177_),
    .A2(_0226_),
    .A1(_0149_));
 sg13g2_nand3_1 _0980_ (.B(_0306_),
    .C(_0307_),
    .A(_0304_),
    .Y(_0112_));
 sg13g2_nand2_1 _0981_ (.Y(_0308_),
    .A(net154),
    .B(net317));
 sg13g2_a21oi_1 _0982_ (.A1(_0208_),
    .A2(_0283_),
    .Y(_0309_),
    .B1(_0308_));
 sg13g2_nand2_1 _0983_ (.Y(_0310_),
    .A(_0150_),
    .B(_0210_));
 sg13g2_nor2_1 _0984_ (.A(_0217_),
    .B(_0226_),
    .Y(_0311_));
 sg13g2_nand3_1 _0985_ (.B(_0310_),
    .C(_0311_),
    .A(_0214_),
    .Y(_0312_));
 sg13g2_nand2b_1 _0986_ (.Y(_0313_),
    .B(_0311_),
    .A_N(_0221_));
 sg13g2_nand2b_1 _0987_ (.Y(_0314_),
    .B(_0308_),
    .A_N(_0243_));
 sg13g2_a22oi_1 _0988_ (.Y(_0315_),
    .B1(_0313_),
    .B2(_0314_),
    .A2(_0312_),
    .A1(_0149_));
 sg13g2_nand2b_1 _0989_ (.Y(_0113_),
    .B(_0315_),
    .A_N(_0309_));
 sg13g2_and2_1 _0990_ (.A(net184),
    .B(_0288_),
    .X(_0114_));
 sg13g2_and2_1 _0991_ (.A(net186),
    .B(_0288_),
    .X(_0115_));
 sg13g2_and2_1 _0992_ (.A(net185),
    .B(_0288_),
    .X(_0116_));
 sg13g2_and2_1 _0993_ (.A(net183),
    .B(_0288_),
    .X(_0117_));
 sg13g2_o21ai_1 _0994_ (.B1(net143),
    .Y(_0316_),
    .A1(_0136_),
    .A2(_0141_));
 sg13g2_o21ai_1 _0995_ (.B1(_0316_),
    .Y(_0317_),
    .A1(_0222_),
    .A2(_0312_));
 sg13g2_nor2_2 _0996_ (.A(_0172_),
    .B(_0186_),
    .Y(_0318_));
 sg13g2_nand2_2 _0997_ (.Y(_0319_),
    .A(_0171_),
    .B(_0185_));
 sg13g2_nand4_1 _0998_ (.B(net154),
    .C(_0241_),
    .A(net297),
    .Y(_0320_),
    .D(_0319_));
 sg13g2_nand3_1 _0999_ (.B(_0317_),
    .C(_0320_),
    .A(_0296_),
    .Y(_0769_));
 sg13g2_nor2b_1 _1000_ (.A(_0161_),
    .B_N(net205),
    .Y(_0000_));
 sg13g2_a221oi_1 _1001_ (.B2(_0177_),
    .C1(_0200_),
    .B1(_0236_),
    .A1(_0181_),
    .Y(_0321_),
    .A2(_0183_));
 sg13g2_nand2_1 _1002_ (.Y(_0322_),
    .A(\SPI_driver1.wait_count[0] ),
    .B(net314));
 sg13g2_nand3_1 _1003_ (.B(\SPI_driver1.wait_count[1] ),
    .C(\SPI_driver1.wait_count[2] ),
    .A(\SPI_driver1.wait_count[0] ),
    .Y(_0323_));
 sg13g2_nor2_1 _1004_ (.A(_0148_),
    .B(_0323_),
    .Y(_0324_));
 sg13g2_o21ai_1 _1005_ (.B1(_0318_),
    .Y(_0325_),
    .A1(net144),
    .A2(_0324_));
 sg13g2_nand2_2 _1006_ (.Y(_0326_),
    .A(_0321_),
    .B(_0325_));
 sg13g2_nand2_1 _1007_ (.Y(_0327_),
    .A(net179),
    .B(_0318_));
 sg13g2_nand2_1 _1008_ (.Y(_0328_),
    .A(\SPI_driver1.wait_count[0] ),
    .B(_0326_));
 sg13g2_o21ai_1 _1009_ (.B1(_0328_),
    .Y(_0035_),
    .A1(_0326_),
    .A2(_0327_));
 sg13g2_a21oi_1 _1010_ (.A1(_0318_),
    .A2(_0322_),
    .Y(_0329_),
    .B1(_0326_));
 sg13g2_o21ai_1 _1011_ (.B1(_0146_),
    .Y(_0330_),
    .A1(_0137_),
    .A2(_0326_));
 sg13g2_nor2b_1 _1012_ (.A(_0329_),
    .B_N(net315),
    .Y(_0036_));
 sg13g2_or4_1 _1013_ (.A(net268),
    .B(_0319_),
    .C(_0322_),
    .D(_0326_),
    .X(_0331_));
 sg13g2_o21ai_1 _1014_ (.B1(_0331_),
    .Y(_0037_),
    .A1(_0147_),
    .A2(_0329_));
 sg13g2_or2_1 _1015_ (.X(_0332_),
    .B(_0326_),
    .A(_0323_));
 sg13g2_a22oi_1 _1016_ (.Y(_0038_),
    .B1(_0332_),
    .B2(_0148_),
    .A2(_0321_),
    .A1(_0319_));
 sg13g2_nor2b_1 _1017_ (.A(\SPI_driver1.SPI_Master1.count_bit[0] ),
    .B_N(net151),
    .Y(_0333_));
 sg13g2_nor2_1 _1018_ (.A(_0167_),
    .B(_0333_),
    .Y(_0334_));
 sg13g2_nor2b_1 _1019_ (.A(net148),
    .B_N(\SPI_driver1.SPI_Master1.word_in[1] ),
    .Y(_0335_));
 sg13g2_a21oi_1 _1020_ (.A1(net147),
    .A2(\SPI_driver1.SPI_Master1.word_out[0] ),
    .Y(_0336_),
    .B1(_0335_));
 sg13g2_nor2_1 _1021_ (.A(net224),
    .B(net118),
    .Y(_0337_));
 sg13g2_a21oi_1 _1022_ (.A1(net118),
    .A2(_0336_),
    .Y(_0039_),
    .B1(_0337_));
 sg13g2_nor2b_1 _1023_ (.A(net148),
    .B_N(\SPI_driver1.SPI_Master1.word_in[2] ),
    .Y(_0338_));
 sg13g2_a21oi_1 _1024_ (.A1(net147),
    .A2(\SPI_driver1.SPI_Master1.word_out[1] ),
    .Y(_0339_),
    .B1(_0338_));
 sg13g2_nor2_1 _1025_ (.A(net213),
    .B(net118),
    .Y(_0340_));
 sg13g2_a21oi_1 _1026_ (.A1(net118),
    .A2(_0339_),
    .Y(_0040_),
    .B1(_0340_));
 sg13g2_nor2b_1 _1027_ (.A(net147),
    .B_N(\SPI_driver1.SPI_Master1.word_in[3] ),
    .Y(_0341_));
 sg13g2_a21oi_1 _1028_ (.A1(net147),
    .A2(net213),
    .Y(_0342_),
    .B1(_0341_));
 sg13g2_nor2_1 _1029_ (.A(net236),
    .B(net118),
    .Y(_0343_));
 sg13g2_a21oi_1 _1030_ (.A1(net118),
    .A2(_0342_),
    .Y(_0041_),
    .B1(_0343_));
 sg13g2_nor2b_1 _1031_ (.A(net147),
    .B_N(\SPI_driver1.SPI_Master1.word_in[4] ),
    .Y(_0344_));
 sg13g2_a21oi_1 _1032_ (.A1(net148),
    .A2(\SPI_driver1.SPI_Master1.word_out[3] ),
    .Y(_0345_),
    .B1(_0344_));
 sg13g2_nor2_1 _1033_ (.A(net217),
    .B(net118),
    .Y(_0346_));
 sg13g2_a21oi_1 _1034_ (.A1(net118),
    .A2(_0345_),
    .Y(_0042_),
    .B1(_0346_));
 sg13g2_nor2b_1 _1035_ (.A(net147),
    .B_N(\SPI_driver1.SPI_Master1.word_in[5] ),
    .Y(_0347_));
 sg13g2_a21oi_1 _1036_ (.A1(net147),
    .A2(net217),
    .Y(_0348_),
    .B1(_0347_));
 sg13g2_nor2_1 _1037_ (.A(net222),
    .B(net120),
    .Y(_0349_));
 sg13g2_a21oi_1 _1038_ (.A1(net120),
    .A2(_0348_),
    .Y(_0043_),
    .B1(_0349_));
 sg13g2_nor2b_1 _1039_ (.A(net146),
    .B_N(net187),
    .Y(_0350_));
 sg13g2_a21oi_1 _1040_ (.A1(net146),
    .A2(net222),
    .Y(_0351_),
    .B1(_0350_));
 sg13g2_nor2_1 _1041_ (.A(net243),
    .B(net120),
    .Y(_0352_));
 sg13g2_a21oi_1 _1042_ (.A1(net120),
    .A2(_0351_),
    .Y(_0044_),
    .B1(_0352_));
 sg13g2_nor2b_1 _1043_ (.A(net147),
    .B_N(\SPI_driver1.SPI_Master1.word_in[7] ),
    .Y(_0353_));
 sg13g2_a21oi_1 _1044_ (.A1(net146),
    .A2(\SPI_driver1.SPI_Master1.word_out[6] ),
    .Y(_0354_),
    .B1(_0353_));
 sg13g2_nor2_1 _1045_ (.A(net226),
    .B(net119),
    .Y(_0355_));
 sg13g2_a21oi_1 _1046_ (.A1(net119),
    .A2(_0354_),
    .Y(_0045_),
    .B1(_0355_));
 sg13g2_nor2b_1 _1047_ (.A(net149),
    .B_N(\SPI_driver1.SPI_Master1.word_in[8] ),
    .Y(_0356_));
 sg13g2_a21oi_1 _1048_ (.A1(net149),
    .A2(net226),
    .Y(_0357_),
    .B1(_0356_));
 sg13g2_nor2_1 _1049_ (.A(net234),
    .B(net122),
    .Y(_0358_));
 sg13g2_a21oi_1 _1050_ (.A1(net119),
    .A2(_0357_),
    .Y(_0046_),
    .B1(_0358_));
 sg13g2_nor2b_1 _1051_ (.A(net148),
    .B_N(\SPI_driver1.SPI_Master1.word_in[9] ),
    .Y(_0359_));
 sg13g2_a21oi_1 _1052_ (.A1(net148),
    .A2(\SPI_driver1.SPI_Master1.word_out[8] ),
    .Y(_0360_),
    .B1(_0359_));
 sg13g2_nor2_1 _1053_ (.A(net209),
    .B(net122),
    .Y(_0361_));
 sg13g2_a21oi_1 _1054_ (.A1(net122),
    .A2(_0360_),
    .Y(_0047_),
    .B1(_0361_));
 sg13g2_nor2b_1 _1055_ (.A(net148),
    .B_N(\SPI_driver1.SPI_Master1.word_in[10] ),
    .Y(_0362_));
 sg13g2_a21oi_1 _1056_ (.A1(net148),
    .A2(net209),
    .Y(_0363_),
    .B1(_0362_));
 sg13g2_nor2_1 _1057_ (.A(net232),
    .B(net122),
    .Y(_0364_));
 sg13g2_a21oi_1 _1058_ (.A1(net122),
    .A2(_0363_),
    .Y(_0048_),
    .B1(_0364_));
 sg13g2_nor2b_1 _1059_ (.A(net150),
    .B_N(\SPI_driver1.SPI_Master1.word_in[11] ),
    .Y(_0365_));
 sg13g2_a21oi_1 _1060_ (.A1(net151),
    .A2(net232),
    .Y(_0366_),
    .B1(_0365_));
 sg13g2_nor2_1 _1061_ (.A(net244),
    .B(net121),
    .Y(_0367_));
 sg13g2_a21oi_1 _1062_ (.A1(net121),
    .A2(_0366_),
    .Y(_0049_),
    .B1(_0367_));
 sg13g2_nor2b_1 _1063_ (.A(net146),
    .B_N(net184),
    .Y(_0368_));
 sg13g2_a21oi_1 _1064_ (.A1(net146),
    .A2(net244),
    .Y(_0369_),
    .B1(_0368_));
 sg13g2_nor2_1 _1065_ (.A(net246),
    .B(net120),
    .Y(_0370_));
 sg13g2_a21oi_1 _1066_ (.A1(net121),
    .A2(_0369_),
    .Y(_0050_),
    .B1(_0370_));
 sg13g2_nor2b_1 _1067_ (.A(net146),
    .B_N(net186),
    .Y(_0371_));
 sg13g2_a21oi_1 _1068_ (.A1(net149),
    .A2(\SPI_driver1.SPI_Master1.word_out[12] ),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_nor2_1 _1069_ (.A(net211),
    .B(net121),
    .Y(_0373_));
 sg13g2_a21oi_1 _1070_ (.A1(net121),
    .A2(_0372_),
    .Y(_0051_),
    .B1(_0373_));
 sg13g2_nor2b_1 _1071_ (.A(net146),
    .B_N(net185),
    .Y(_0374_));
 sg13g2_a21oi_1 _1072_ (.A1(net146),
    .A2(net211),
    .Y(_0375_),
    .B1(_0374_));
 sg13g2_nor2_1 _1073_ (.A(net228),
    .B(net121),
    .Y(_0376_));
 sg13g2_a21oi_1 _1074_ (.A1(net121),
    .A2(_0375_),
    .Y(_0052_),
    .B1(_0376_));
 sg13g2_nor2b_1 _1075_ (.A(net150),
    .B_N(net183),
    .Y(_0377_));
 sg13g2_a21oi_1 _1076_ (.A1(net150),
    .A2(net228),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_nor2_1 _1077_ (.A(net247),
    .B(net122),
    .Y(_0379_));
 sg13g2_a21oi_1 _1078_ (.A1(net121),
    .A2(_0378_),
    .Y(_0053_),
    .B1(_0379_));
 sg13g2_nor2_2 _1079_ (.A(net150),
    .B(_0156_),
    .Y(_0380_));
 sg13g2_and3_1 _1080_ (.X(_0381_),
    .A(_0161_),
    .B(_0163_),
    .C(_0168_));
 sg13g2_nor2_1 _1081_ (.A(_0380_),
    .B(_0381_),
    .Y(_0382_));
 sg13g2_nand2_1 _1082_ (.Y(_0383_),
    .A(\SPI_driver1.SPI_Master1.count_word[0] ),
    .B(_0382_));
 sg13g2_a21oi_1 _1083_ (.A1(net189),
    .A2(_0381_),
    .Y(_0384_),
    .B1(_0380_));
 sg13g2_nand2_1 _1084_ (.Y(_0054_),
    .A(_0383_),
    .B(_0384_));
 sg13g2_o21ai_1 _1085_ (.B1(net307),
    .Y(_0385_),
    .A1(\SPI_driver1.SPI_Master1.count_word[0] ),
    .A2(_0382_));
 sg13g2_o21ai_1 _1086_ (.B1(_0159_),
    .Y(_0386_),
    .A1(_0380_),
    .A2(_0381_));
 sg13g2_nand3b_1 _1087_ (.B(net308),
    .C(_0386_),
    .Y(_0055_),
    .A_N(_0380_));
 sg13g2_nand3_1 _1088_ (.B(_0163_),
    .C(_0168_),
    .A(_0160_),
    .Y(_0387_));
 sg13g2_a22oi_1 _1089_ (.Y(_0388_),
    .B1(_0386_),
    .B2(net266),
    .A2(_0381_),
    .A1(_0160_));
 sg13g2_nand2b_1 _1090_ (.Y(_0056_),
    .B(net267),
    .A_N(_0380_));
 sg13g2_a21o_1 _1091_ (.A2(_0387_),
    .A1(net238),
    .B1(_0380_),
    .X(_0057_));
 sg13g2_o21ai_1 _1092_ (.B1(net219),
    .Y(_0389_),
    .A1(_0135_),
    .A2(_0136_));
 sg13g2_nor2b_2 _1093_ (.A(net215),
    .B_N(\SPI_driver1.SPI_Master1.res ),
    .Y(_0390_));
 sg13g2_o21ai_1 _1094_ (.B1(net220),
    .Y(_0058_),
    .A1(_0166_),
    .A2(_0390_));
 sg13g2_o21ai_1 _1095_ (.B1(_0390_),
    .Y(_0391_),
    .A1(net151),
    .A2(\SPI_driver1.SPI_Master1.sclk ));
 sg13g2_a21oi_1 _1096_ (.A1(_0138_),
    .A2(_0164_),
    .Y(_0059_),
    .B1(_0391_));
 sg13g2_a21oi_1 _1097_ (.A1(net151),
    .A2(\SPI_driver1.SPI_Master1.count_bit[0] ),
    .Y(_0392_),
    .B1(net191));
 sg13g2_nand2b_1 _1098_ (.Y(_0393_),
    .B(net151),
    .A_N(\SPI_driver1.SPI_Master1.word_out[15] ));
 sg13g2_a22oi_1 _1099_ (.Y(_0394_),
    .B1(_0390_),
    .B2(_0393_),
    .A2(_0333_),
    .A1(net141));
 sg13g2_nor2_1 _1100_ (.A(net192),
    .B(_0394_),
    .Y(_0060_));
 sg13g2_o21ai_1 _1101_ (.B1(net141),
    .Y(_0395_),
    .A1(net145),
    .A2(\SPI_driver1.SPI_Master1.state[0] ));
 sg13g2_a21oi_1 _1102_ (.A1(_0134_),
    .A2(\SPI_driver1.SPI_Master1.state[0] ),
    .Y(_0061_),
    .B1(_0395_));
 sg13g2_nand2_1 _1103_ (.Y(_0396_),
    .A(net229),
    .B(_0380_));
 sg13g2_o21ai_1 _1104_ (.B1(_0396_),
    .Y(_0062_),
    .A1(_0151_),
    .A2(net119));
 sg13g2_nand2_1 _1105_ (.Y(_0397_),
    .A(net254),
    .B(net250));
 sg13g2_nand3_1 _1106_ (.B(\clockDivider1.counter[8] ),
    .C(\clockDivider1.counter[7] ),
    .A(\clockDivider1.counter[9] ),
    .Y(_0398_));
 sg13g2_nor2b_1 _1107_ (.A(\clockDivider1.counter[10] ),
    .B_N(_0398_),
    .Y(_0399_));
 sg13g2_or3_1 _1108_ (.A(\clockDivider1.counter[5] ),
    .B(\clockDivider1.counter[4] ),
    .C(\clockDivider1.counter[3] ),
    .X(_0400_));
 sg13g2_nor4_1 _1109_ (.A(\clockDivider1.counter[10] ),
    .B(\clockDivider1.counter[6] ),
    .C(_0398_),
    .D(_0400_),
    .Y(_0401_));
 sg13g2_o21ai_1 _1110_ (.B1(_0132_),
    .Y(_0402_),
    .A1(_0399_),
    .A2(_0401_));
 sg13g2_a21oi_1 _1111_ (.A1(\clockDivider1.counter[12] ),
    .A2(_0402_),
    .Y(_0403_),
    .B1(_0139_));
 sg13g2_a21oi_1 _1112_ (.A1(\clockDivider1.ena ),
    .A2(_0403_),
    .Y(_0404_),
    .B1(net256));
 sg13g2_nor2b_2 _1113_ (.A(net156),
    .B_N(net4),
    .Y(_0405_));
 sg13g2_nand2_1 _1114_ (.Y(_0406_),
    .A(_0141_),
    .B(net4));
 sg13g2_and2_1 _1115_ (.A(\clockDivider1.ena ),
    .B(net256),
    .X(_0407_));
 sg13g2_nor3_1 _1116_ (.A(net257),
    .B(_0405_),
    .C(_0407_),
    .Y(_0063_));
 sg13g2_nor2_2 _1117_ (.A(net135),
    .B(_0405_),
    .Y(_0408_));
 sg13g2_nand3_1 _1118_ (.B(\clockDivider1.counter[1] ),
    .C(\clockDivider1.counter[0] ),
    .A(\clockDivider1.counter[2] ),
    .Y(_0409_));
 sg13g2_nor4_1 _1119_ (.A(\clockDivider1.counter[13] ),
    .B(_0131_),
    .C(\clockDivider1.counter[11] ),
    .D(_0409_),
    .Y(_0410_));
 sg13g2_a221oi_1 _1120_ (.B2(_0401_),
    .C1(_0139_),
    .B1(_0410_),
    .A1(\clockDivider1.counter[12] ),
    .Y(_0411_),
    .A2(_0402_));
 sg13g2_nand2_2 _1121_ (.Y(_0412_),
    .A(net125),
    .B(_0411_));
 sg13g2_nand2b_1 _1122_ (.Y(_0413_),
    .B(net135),
    .A_N(_0411_));
 sg13g2_o21ai_1 _1123_ (.B1(net125),
    .Y(_0414_),
    .A1(_0127_),
    .A2(_0411_));
 sg13g2_nor2_1 _1124_ (.A(net274),
    .B(_0407_),
    .Y(_0415_));
 sg13g2_and2_1 _1125_ (.A(net274),
    .B(_0407_),
    .X(_0416_));
 sg13g2_nor3_1 _1126_ (.A(_0414_),
    .B(net275),
    .C(_0416_),
    .Y(_0064_));
 sg13g2_nor2_1 _1127_ (.A(net263),
    .B(_0416_),
    .Y(_0417_));
 sg13g2_and4_1 _1128_ (.A(net135),
    .B(net263),
    .C(net274),
    .D(net256),
    .X(_0418_));
 sg13g2_nor3_1 _1129_ (.A(_0414_),
    .B(net264),
    .C(_0418_),
    .Y(_0065_));
 sg13g2_nor2_1 _1130_ (.A(net277),
    .B(_0418_),
    .Y(_0419_));
 sg13g2_and2_1 _1131_ (.A(net277),
    .B(_0418_),
    .X(_0420_));
 sg13g2_nor3_1 _1132_ (.A(_0414_),
    .B(_0419_),
    .C(_0420_),
    .Y(_0066_));
 sg13g2_nor2_1 _1133_ (.A(net287),
    .B(_0420_),
    .Y(_0421_));
 sg13g2_and2_1 _1134_ (.A(net287),
    .B(_0420_),
    .X(_0422_));
 sg13g2_nor3_1 _1135_ (.A(_0414_),
    .B(_0421_),
    .C(_0422_),
    .Y(_0067_));
 sg13g2_nand2_1 _1136_ (.Y(_0423_),
    .A(net272),
    .B(_0408_));
 sg13g2_nand3_1 _1137_ (.B(\clockDivider1.counter[4] ),
    .C(\clockDivider1.counter[3] ),
    .A(\clockDivider1.counter[5] ),
    .Y(_0424_));
 sg13g2_or2_1 _1138_ (.X(_0425_),
    .B(_0424_),
    .A(_0409_));
 sg13g2_o21ai_1 _1139_ (.B1(_0425_),
    .Y(_0426_),
    .A1(net272),
    .A2(_0422_));
 sg13g2_o21ai_1 _1140_ (.B1(_0423_),
    .Y(_0068_),
    .A1(_0412_),
    .A2(_0426_));
 sg13g2_a21oi_1 _1141_ (.A1(\clockDivider1.counter[5] ),
    .A2(_0422_),
    .Y(_0427_),
    .B1(net260));
 sg13g2_and4_1 _1142_ (.A(net260),
    .B(\clockDivider1.counter[5] ),
    .C(net327),
    .D(_0420_),
    .X(_0428_));
 sg13g2_nor3_1 _1143_ (.A(_0414_),
    .B(net261),
    .C(net328),
    .Y(_0069_));
 sg13g2_nand2_1 _1144_ (.Y(_0429_),
    .A(net278),
    .B(_0408_));
 sg13g2_nand2_1 _1145_ (.Y(_0430_),
    .A(\clockDivider1.counter[7] ),
    .B(\clockDivider1.counter[6] ));
 sg13g2_or2_1 _1146_ (.X(_0431_),
    .B(_0430_),
    .A(_0425_));
 sg13g2_o21ai_1 _1147_ (.B1(_0431_),
    .Y(_0432_),
    .A1(net278),
    .A2(_0428_));
 sg13g2_o21ai_1 _1148_ (.B1(_0429_),
    .Y(_0070_),
    .A1(_0412_),
    .A2(_0432_));
 sg13g2_a21oi_1 _1149_ (.A1(\clockDivider1.counter[7] ),
    .A2(_0428_),
    .Y(_0433_),
    .B1(net250));
 sg13g2_and3_1 _1150_ (.X(_0434_),
    .A(net250),
    .B(\clockDivider1.counter[7] ),
    .C(_0428_));
 sg13g2_nor3_1 _1151_ (.A(_0414_),
    .B(net251),
    .C(_0434_),
    .Y(_0071_));
 sg13g2_nand2_1 _1152_ (.Y(_0435_),
    .A(net254),
    .B(_0408_));
 sg13g2_nor3_2 _1153_ (.A(_0397_),
    .B(_0425_),
    .C(_0430_),
    .Y(_0436_));
 sg13g2_inv_1 _1154_ (.Y(_0437_),
    .A(_0436_));
 sg13g2_o21ai_1 _1155_ (.B1(_0437_),
    .Y(_0438_),
    .A1(net254),
    .A2(_0434_));
 sg13g2_o21ai_1 _1156_ (.B1(_0435_),
    .Y(_0072_),
    .A1(_0412_),
    .A2(_0438_));
 sg13g2_a21o_1 _1157_ (.A2(_0436_),
    .A1(net135),
    .B1(net323),
    .X(_0439_));
 sg13g2_nand3_1 _1158_ (.B(\clockDivider1.counter[10] ),
    .C(_0436_),
    .A(net134),
    .Y(_0440_));
 sg13g2_and4_1 _1159_ (.A(net125),
    .B(_0413_),
    .C(_0439_),
    .D(_0440_),
    .X(_0073_));
 sg13g2_nand2_1 _1160_ (.Y(_0441_),
    .A(net285),
    .B(_0408_));
 sg13g2_nand3_1 _1161_ (.B(\clockDivider1.counter[10] ),
    .C(_0436_),
    .A(net285),
    .Y(_0442_));
 sg13g2_nand3_1 _1162_ (.B(_0411_),
    .C(_0442_),
    .A(net125),
    .Y(_0443_));
 sg13g2_a22oi_1 _1163_ (.Y(_0074_),
    .B1(_0441_),
    .B2(_0443_),
    .A2(_0440_),
    .A1(_0132_));
 sg13g2_nand4_1 _1164_ (.B(net285),
    .C(\clockDivider1.counter[10] ),
    .A(net134),
    .Y(_0444_),
    .D(_0436_));
 sg13g2_xnor2_1 _1165_ (.Y(_0445_),
    .A(_0131_),
    .B(_0444_));
 sg13g2_nor2_1 _1166_ (.A(_0414_),
    .B(net319),
    .Y(_0075_));
 sg13g2_and2_1 _1167_ (.A(net188),
    .B(_0408_),
    .X(_0076_));
 sg13g2_nor3_1 _1168_ (.A(_0127_),
    .B(net240),
    .C(_0411_),
    .Y(_0446_));
 sg13g2_a221oi_1 _1169_ (.B2(_0130_),
    .C1(net241),
    .B1(_0413_),
    .A1(_0141_),
    .Y(_0077_),
    .A2(net4));
 sg13g2_o21ai_1 _1170_ (.B1(net156),
    .Y(_0447_),
    .A1(net135),
    .A2(net2));
 sg13g2_a21oi_1 _1171_ (.A1(_0129_),
    .A2(net2),
    .Y(_0078_),
    .B1(_0447_));
 sg13g2_a21oi_1 _1172_ (.A1(net196),
    .A2(net3),
    .Y(_0448_),
    .B1(_0141_));
 sg13g2_o21ai_1 _1173_ (.B1(_0448_),
    .Y(_0079_),
    .A1(_0128_),
    .A2(net3));
 sg13g2_and2_2 _1174_ (.A(net134),
    .B(\counter_chain1.ces_X0_ena ),
    .X(_0449_));
 sg13g2_and2_1 _1175_ (.A(\counter_chain1.inst_ces_X0.max ),
    .B(_0449_),
    .X(_0450_));
 sg13g2_and4_2 _1176_ (.A(net134),
    .B(\counter_chain1.ces_X0_ena ),
    .C(\counter_chain1.inst_ces_X0.max ),
    .D(\counter_chain1.inst_sec_0X.max ),
    .X(_0451_));
 sg13g2_nand2_1 _1177_ (.Y(_0452_),
    .A(\counter_chain1.inst_sec_0X.max ),
    .B(_0450_));
 sg13g2_and2_2 _1178_ (.A(\counter_chain1.inst_sec_X0.max ),
    .B(_0451_),
    .X(_0453_));
 sg13g2_nand2_1 _1179_ (.Y(_0454_),
    .A(\counter_chain1.inst_min_0X.max ),
    .B(_0453_));
 sg13g2_nor2b_1 _1180_ (.A(\SPI_driver1.min_X0[1] ),
    .B_N(\SPI_driver1.min_X0[2] ),
    .Y(_0455_));
 sg13g2_mux2_1 _1181_ (.A0(_0030_),
    .A1(_0029_),
    .S(_0455_),
    .X(_0456_));
 sg13g2_nand3_1 _1182_ (.B(_0453_),
    .C(_0456_),
    .A(\counter_chain1.inst_min_0X.max ),
    .Y(_0457_));
 sg13g2_inv_1 _1183_ (.Y(_0458_),
    .A(_0457_));
 sg13g2_mux2_1 _1184_ (.A0(_0458_),
    .A1(_0454_),
    .S(\SPI_driver1.min_X0[0] ),
    .X(_0459_));
 sg13g2_and2_1 _1185_ (.A(net124),
    .B(_0459_),
    .X(_0080_));
 sg13g2_nand2_1 _1186_ (.Y(_0460_),
    .A(\SPI_driver1.min_X0[1] ),
    .B(\SPI_driver1.min_X0[0] ));
 sg13g2_a22oi_1 _1187_ (.Y(_0461_),
    .B1(_0458_),
    .B2(_0460_),
    .A2(_0454_),
    .A1(\SPI_driver1.min_X0[1] ));
 sg13g2_o21ai_1 _1188_ (.B1(net124),
    .Y(_0462_),
    .A1(\SPI_driver1.min_X0[1] ),
    .A2(\SPI_driver1.min_X0[0] ));
 sg13g2_nor2_1 _1189_ (.A(_0461_),
    .B(_0462_),
    .Y(_0081_));
 sg13g2_xor2_1 _1190_ (.B(_0460_),
    .A(_0030_),
    .X(_0463_));
 sg13g2_a22oi_1 _1191_ (.Y(_0464_),
    .B1(_0458_),
    .B2(_0463_),
    .A2(_0454_),
    .A1(\SPI_driver1.min_X0[2] ));
 sg13g2_nor2_1 _1192_ (.A(_0405_),
    .B(_0464_),
    .Y(_0082_));
 sg13g2_nor3_1 _1193_ (.A(\SPI_driver1.min_0X[2] ),
    .B(\SPI_driver1.min_0X[1] ),
    .C(\SPI_driver1.min_0X[0] ),
    .Y(_0465_));
 sg13g2_nand2_1 _1194_ (.Y(_0466_),
    .A(\SPI_driver1.min_0X[3] ),
    .B(_0465_));
 sg13g2_o21ai_1 _1195_ (.B1(net124),
    .Y(_0467_),
    .A1(\counter_chain1.inst_min_0X.max ),
    .A2(_0453_));
 sg13g2_a21oi_1 _1196_ (.A1(_0453_),
    .A2(_0466_),
    .Y(_0083_),
    .B1(_0467_));
 sg13g2_nand3b_1 _1197_ (.B(_0453_),
    .C(\SPI_driver1.min_0X[3] ),
    .Y(_0468_),
    .A_N(_0465_));
 sg13g2_nand2_2 _1198_ (.Y(_0469_),
    .A(net124),
    .B(_0468_));
 sg13g2_and2_1 _1199_ (.A(\SPI_driver1.min_0X[0] ),
    .B(_0453_),
    .X(_0470_));
 sg13g2_nor2_1 _1200_ (.A(\SPI_driver1.min_0X[0] ),
    .B(_0453_),
    .Y(_0471_));
 sg13g2_nor3_1 _1201_ (.A(_0469_),
    .B(_0470_),
    .C(_0471_),
    .Y(_0084_));
 sg13g2_and2_1 _1202_ (.A(\SPI_driver1.min_0X[1] ),
    .B(_0470_),
    .X(_0472_));
 sg13g2_nor2_1 _1203_ (.A(\SPI_driver1.min_0X[1] ),
    .B(_0470_),
    .Y(_0473_));
 sg13g2_nor3_1 _1204_ (.A(_0469_),
    .B(_0472_),
    .C(_0473_),
    .Y(_0085_));
 sg13g2_xnor2_1 _1205_ (.Y(_0474_),
    .A(\SPI_driver1.min_0X[2] ),
    .B(_0472_));
 sg13g2_nor2_1 _1206_ (.A(_0469_),
    .B(_0474_),
    .Y(_0086_));
 sg13g2_a21oi_1 _1207_ (.A1(\SPI_driver1.min_0X[2] ),
    .A2(_0472_),
    .Y(_0475_),
    .B1(\SPI_driver1.min_0X[3] ));
 sg13g2_nor2_1 _1208_ (.A(_0469_),
    .B(_0475_),
    .Y(_0087_));
 sg13g2_nor2_1 _1209_ (.A(\SPI_driver1.sec_X0[1] ),
    .B(\SPI_driver1.sec_X0[0] ),
    .Y(_0476_));
 sg13g2_nand2_1 _1210_ (.Y(_0477_),
    .A(\SPI_driver1.sec_X0[2] ),
    .B(_0476_));
 sg13g2_o21ai_1 _1211_ (.B1(net124),
    .Y(_0478_),
    .A1(\counter_chain1.inst_sec_X0.max ),
    .A2(_0451_));
 sg13g2_a21oi_1 _1212_ (.A1(_0451_),
    .A2(_0477_),
    .Y(_0088_),
    .B1(_0478_));
 sg13g2_nor2b_1 _1213_ (.A(\SPI_driver1.sec_X0[1] ),
    .B_N(\SPI_driver1.sec_X0[2] ),
    .Y(_0479_));
 sg13g2_mux2_1 _1214_ (.A0(_0032_),
    .A1(_0031_),
    .S(_0479_),
    .X(_0480_));
 sg13g2_nand2_1 _1215_ (.Y(_0481_),
    .A(_0451_),
    .B(_0480_));
 sg13g2_inv_1 _1216_ (.Y(_0482_),
    .A(_0481_));
 sg13g2_o21ai_1 _1217_ (.B1(net124),
    .Y(_0483_),
    .A1(\SPI_driver1.sec_X0[0] ),
    .A2(_0482_));
 sg13g2_a21oi_1 _1218_ (.A1(\SPI_driver1.sec_X0[0] ),
    .A2(_0451_),
    .Y(_0089_),
    .B1(_0483_));
 sg13g2_nand2_1 _1219_ (.Y(_0484_),
    .A(\SPI_driver1.sec_X0[1] ),
    .B(\SPI_driver1.sec_X0[0] ));
 sg13g2_a22oi_1 _1220_ (.Y(_0485_),
    .B1(_0482_),
    .B2(_0484_),
    .A2(_0452_),
    .A1(\SPI_driver1.sec_X0[1] ));
 sg13g2_nor3_1 _1221_ (.A(_0405_),
    .B(_0476_),
    .C(_0485_),
    .Y(_0090_));
 sg13g2_xor2_1 _1222_ (.B(_0484_),
    .A(_0032_),
    .X(_0486_));
 sg13g2_a22oi_1 _1223_ (.Y(_0487_),
    .B1(_0482_),
    .B2(_0486_),
    .A2(_0452_),
    .A1(\SPI_driver1.sec_X0[2] ));
 sg13g2_nor2_1 _1224_ (.A(_0405_),
    .B(_0487_),
    .Y(_0091_));
 sg13g2_nand2b_1 _1225_ (.Y(_0488_),
    .B(\counter_chain1.inst_sec_0X.max ),
    .A_N(_0450_));
 sg13g2_nor3_1 _1226_ (.A(\SPI_driver1.sec_0X[2] ),
    .B(\SPI_driver1.sec_0X[1] ),
    .C(\SPI_driver1.sec_0X[0] ),
    .Y(_0489_));
 sg13g2_nand2_1 _1227_ (.Y(_0490_),
    .A(\SPI_driver1.sec_0X[3] ),
    .B(_0450_));
 sg13g2_nand3_1 _1228_ (.B(_0450_),
    .C(_0489_),
    .A(\SPI_driver1.sec_0X[3] ),
    .Y(_0491_));
 sg13g2_a21oi_1 _1229_ (.A1(_0488_),
    .A2(_0491_),
    .Y(_0092_),
    .B1(_0405_));
 sg13g2_o21ai_1 _1230_ (.B1(net125),
    .Y(_0492_),
    .A1(_0489_),
    .A2(_0490_));
 sg13g2_nor2_1 _1231_ (.A(\SPI_driver1.sec_0X[0] ),
    .B(_0450_),
    .Y(_0493_));
 sg13g2_and2_1 _1232_ (.A(\SPI_driver1.sec_0X[0] ),
    .B(_0450_),
    .X(_0494_));
 sg13g2_nor3_1 _1233_ (.A(_0492_),
    .B(_0493_),
    .C(_0494_),
    .Y(_0093_));
 sg13g2_and2_1 _1234_ (.A(\SPI_driver1.sec_0X[1] ),
    .B(_0494_),
    .X(_0495_));
 sg13g2_nor2_1 _1235_ (.A(\SPI_driver1.sec_0X[1] ),
    .B(_0494_),
    .Y(_0496_));
 sg13g2_nor3_1 _1236_ (.A(_0492_),
    .B(_0495_),
    .C(_0496_),
    .Y(_0094_));
 sg13g2_xnor2_1 _1237_ (.Y(_0497_),
    .A(\SPI_driver1.sec_0X[2] ),
    .B(_0495_));
 sg13g2_nor2_1 _1238_ (.A(_0492_),
    .B(_0497_),
    .Y(_0095_));
 sg13g2_a21oi_1 _1239_ (.A1(\SPI_driver1.sec_0X[2] ),
    .A2(_0495_),
    .Y(_0498_),
    .B1(\SPI_driver1.sec_0X[3] ));
 sg13g2_nor2_1 _1240_ (.A(_0492_),
    .B(_0498_),
    .Y(_0096_));
 sg13g2_nor3_1 _1241_ (.A(\SPI_driver1.ces_X0[2] ),
    .B(\SPI_driver1.ces_X0[1] ),
    .C(\SPI_driver1.ces_X0[0] ),
    .Y(_0499_));
 sg13g2_nand2_1 _1242_ (.Y(_0500_),
    .A(\SPI_driver1.ces_X0[3] ),
    .B(_0449_));
 sg13g2_nand3_1 _1243_ (.B(_0449_),
    .C(_0499_),
    .A(\SPI_driver1.ces_X0[3] ),
    .Y(_0501_));
 sg13g2_nand2b_1 _1244_ (.Y(_0502_),
    .B(\counter_chain1.inst_ces_X0.max ),
    .A_N(_0449_));
 sg13g2_a21oi_1 _1245_ (.A1(_0501_),
    .A2(_0502_),
    .Y(_0097_),
    .B1(_0405_));
 sg13g2_o21ai_1 _1246_ (.B1(net124),
    .Y(_0503_),
    .A1(_0499_),
    .A2(_0500_));
 sg13g2_and2_1 _1247_ (.A(\SPI_driver1.ces_X0[0] ),
    .B(_0449_),
    .X(_0504_));
 sg13g2_nor2_1 _1248_ (.A(\SPI_driver1.ces_X0[0] ),
    .B(_0449_),
    .Y(_0505_));
 sg13g2_nor3_1 _1249_ (.A(_0503_),
    .B(_0504_),
    .C(_0505_),
    .Y(_0098_));
 sg13g2_and2_1 _1250_ (.A(\SPI_driver1.ces_X0[1] ),
    .B(_0504_),
    .X(_0506_));
 sg13g2_nor2_1 _1251_ (.A(\SPI_driver1.ces_X0[1] ),
    .B(_0504_),
    .Y(_0507_));
 sg13g2_nor3_1 _1252_ (.A(_0503_),
    .B(_0506_),
    .C(_0507_),
    .Y(_0099_));
 sg13g2_xnor2_1 _1253_ (.Y(_0508_),
    .A(\SPI_driver1.ces_X0[2] ),
    .B(_0506_));
 sg13g2_nor2_1 _1254_ (.A(_0503_),
    .B(_0508_),
    .Y(_0100_));
 sg13g2_a21oi_1 _1255_ (.A1(\SPI_driver1.ces_X0[2] ),
    .A2(_0506_),
    .Y(_0509_),
    .B1(\SPI_driver1.ces_X0[3] ));
 sg13g2_nor2_1 _1256_ (.A(_0503_),
    .B(_0509_),
    .Y(_0101_));
 sg13g2_nand2_1 _1257_ (.Y(_0510_),
    .A(\counter_chain1.ces_X0_ena ),
    .B(_0408_));
 sg13g2_nor3_1 _1258_ (.A(\SPI_driver1.ces_0X[2] ),
    .B(\SPI_driver1.ces_0X[1] ),
    .C(\SPI_driver1.ces_0X[0] ),
    .Y(_0511_));
 sg13g2_nand2_1 _1259_ (.Y(_0512_),
    .A(\SPI_driver1.ces_0X[3] ),
    .B(net134));
 sg13g2_nand4_1 _1260_ (.B(net134),
    .C(net124),
    .A(\SPI_driver1.ces_0X[3] ),
    .Y(_0513_),
    .D(_0511_));
 sg13g2_nand2_1 _1261_ (.Y(_0102_),
    .A(_0510_),
    .B(_0513_));
 sg13g2_o21ai_1 _1262_ (.B1(\SPI_driver1.ces_0X[3] ),
    .Y(_0514_),
    .A1(\SPI_driver1.ces_0X[2] ),
    .A2(\SPI_driver1.ces_0X[1] ));
 sg13g2_a21oi_1 _1263_ (.A1(net134),
    .A2(_0514_),
    .Y(_0515_),
    .B1(\SPI_driver1.ces_0X[0] ));
 sg13g2_and2_1 _1264_ (.A(net134),
    .B(\SPI_driver1.ces_0X[0] ),
    .X(_0516_));
 sg13g2_nor3_1 _1265_ (.A(_0405_),
    .B(_0515_),
    .C(_0516_),
    .Y(_0103_));
 sg13g2_o21ai_1 _1266_ (.B1(net125),
    .Y(_0517_),
    .A1(_0511_),
    .A2(_0512_));
 sg13g2_xnor2_1 _1267_ (.Y(_0518_),
    .A(\SPI_driver1.ces_0X[1] ),
    .B(_0516_));
 sg13g2_nor2_1 _1268_ (.A(_0517_),
    .B(_0518_),
    .Y(_0104_));
 sg13g2_a21oi_1 _1269_ (.A1(\SPI_driver1.ces_0X[1] ),
    .A2(_0516_),
    .Y(_0519_),
    .B1(\SPI_driver1.ces_0X[2] ));
 sg13g2_and3_1 _1270_ (.X(_0520_),
    .A(\SPI_driver1.ces_0X[2] ),
    .B(\SPI_driver1.ces_0X[1] ),
    .C(_0516_));
 sg13g2_nor3_1 _1271_ (.A(_0517_),
    .B(_0519_),
    .C(_0520_),
    .Y(_0105_));
 sg13g2_nor2_1 _1272_ (.A(\SPI_driver1.ces_0X[3] ),
    .B(_0520_),
    .Y(_0521_));
 sg13g2_nor2_1 _1273_ (.A(_0517_),
    .B(_0521_),
    .Y(_0106_));
 sg13g2_nand3b_1 _1274_ (.B(_0187_),
    .C(net133),
    .Y(_0522_),
    .A_N(\SPI_driver1.state[2] ));
 sg13g2_nand2_1 _1275_ (.Y(_0523_),
    .A(_0130_),
    .B(net145));
 sg13g2_nand3_1 _1276_ (.B(net1),
    .C(_0523_),
    .A(net133),
    .Y(_0524_));
 sg13g2_nor2_1 _1277_ (.A(_0133_),
    .B(net280),
    .Y(_0525_));
 sg13g2_nand2_1 _1278_ (.Y(_0526_),
    .A(_0175_),
    .B(net281));
 sg13g2_a22oi_1 _1279_ (.Y(_0107_),
    .B1(_0524_),
    .B2(_0526_),
    .A2(_0522_),
    .A1(net133));
 sg13g2_nor2b_1 _1280_ (.A(net154),
    .B_N(net5),
    .Y(_0527_));
 sg13g2_a21oi_1 _1281_ (.A1(\SPI_driver1.state[2] ),
    .A2(net155),
    .Y(_0528_),
    .B1(_0527_));
 sg13g2_a21o_1 _1282_ (.A2(_0285_),
    .A1(_0282_),
    .B1(net143),
    .X(_0529_));
 sg13g2_nand3_1 _1283_ (.B(_0216_),
    .C(_0258_),
    .A(_0214_),
    .Y(_0530_));
 sg13g2_nand3_1 _1284_ (.B(\SPI_driver1.sent_LUX ),
    .C(_0214_),
    .A(_0149_),
    .Y(_0531_));
 sg13g2_a221oi_1 _1285_ (.B2(_0531_),
    .C1(_0224_),
    .B1(_0530_),
    .A1(_0185_),
    .Y(_0532_),
    .A2(_0205_));
 sg13g2_a21oi_1 _1286_ (.A1(_0528_),
    .A2(_0529_),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_a21oi_1 _1287_ (.A1(_0236_),
    .A2(_0525_),
    .Y(_0534_),
    .B1(_0176_));
 sg13g2_nor2b_1 _1288_ (.A(_0534_),
    .B_N(_0180_),
    .Y(_0535_));
 sg13g2_nor2_1 _1289_ (.A(_0528_),
    .B(_0535_),
    .Y(_0536_));
 sg13g2_a22oi_1 _1290_ (.Y(_0537_),
    .B1(_0527_),
    .B2(_0209_),
    .A2(_0522_),
    .A1(net132));
 sg13g2_a21oi_1 _1291_ (.A1(_0523_),
    .A2(_0528_),
    .Y(_0538_),
    .B1(_0522_));
 sg13g2_and2_1 _1292_ (.A(_0318_),
    .B(_0324_),
    .X(_0539_));
 sg13g2_nor3_1 _1293_ (.A(net123),
    .B(_0538_),
    .C(_0539_),
    .Y(_0540_));
 sg13g2_nand3_1 _1294_ (.B(_0537_),
    .C(_0540_),
    .A(_0193_),
    .Y(_0541_));
 sg13g2_or3_1 _1295_ (.A(_0533_),
    .B(_0536_),
    .C(_0541_),
    .X(_0108_));
 sg13g2_a21oi_1 _1296_ (.A1(_0256_),
    .A2(_0257_),
    .Y(_0542_),
    .B1(net143));
 sg13g2_and2_1 _1297_ (.A(net129),
    .B(net155),
    .X(_0543_));
 sg13g2_nor4_1 _1298_ (.A(net123),
    .B(_0539_),
    .C(_0542_),
    .D(_0543_),
    .Y(_0544_));
 sg13g2_a21oi_1 _1299_ (.A1(net143),
    .A2(_0221_),
    .Y(_0545_),
    .B1(_0222_));
 sg13g2_nand3_1 _1300_ (.B(_0256_),
    .C(_0319_),
    .A(_0216_),
    .Y(_0546_));
 sg13g2_nor2_1 _1301_ (.A(_0534_),
    .B(_0546_),
    .Y(_0547_));
 sg13g2_and2_1 _1302_ (.A(_0545_),
    .B(_0547_),
    .X(_0548_));
 sg13g2_o21ai_1 _1303_ (.B1(_0193_),
    .Y(_0109_),
    .A1(_0544_),
    .A2(_0548_));
 sg13g2_a21oi_1 _1304_ (.A1(net127),
    .A2(net155),
    .Y(_0549_),
    .B1(_0527_));
 sg13g2_o21ai_1 _1305_ (.B1(_0225_),
    .Y(_0550_),
    .A1(_0176_),
    .A2(_0525_));
 sg13g2_o21ai_1 _1306_ (.B1(_0545_),
    .Y(_0551_),
    .A1(_0319_),
    .A2(_0324_));
 sg13g2_nor4_2 _1307_ (.A(_0184_),
    .B(_0530_),
    .C(_0550_),
    .Y(_0552_),
    .D(_0551_));
 sg13g2_a21o_1 _1308_ (.A2(_0549_),
    .A1(net144),
    .B1(_0150_),
    .X(_0553_));
 sg13g2_o21ai_1 _1309_ (.B1(_0209_),
    .Y(_0554_),
    .A1(net155),
    .A2(net5));
 sg13g2_a21oi_1 _1310_ (.A1(net154),
    .A2(_0553_),
    .Y(_0555_),
    .B1(_0554_));
 sg13g2_a21oi_1 _1311_ (.A1(_0257_),
    .A2(_0282_),
    .Y(_0556_),
    .B1(net142));
 sg13g2_nor4_1 _1312_ (.A(net123),
    .B(_0538_),
    .C(_0555_),
    .D(_0556_),
    .Y(_0557_));
 sg13g2_o21ai_1 _1313_ (.B1(_0557_),
    .Y(_0110_),
    .A1(_0549_),
    .A2(_0552_));
 sg13g2_dfrbp_1 _1314_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net27),
    .D(_0007_),
    .Q_N(_0027_),
    .Q(\SPI_driver1.digit_count[0] ));
 sg13g2_dfrbp_1 _1315_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net28),
    .D(net293),
    .Q_N(_0625_),
    .Q(\SPI_driver1.digit_count[1] ));
 sg13g2_dfrbp_1 _1316_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net29),
    .D(net302),
    .Q_N(_0626_),
    .Q(\SPI_driver1.digit_count[2] ));
 sg13g2_dfrbp_1 _1317_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net30),
    .D(net208),
    .Q_N(_0028_),
    .Q(\SPI_driver1.digit_count[3] ));
 sg13g2_dfrbp_1 _1318_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net31),
    .D(_0011_),
    .Q_N(_0627_),
    .Q(\SPI_driver1.digit_count[4] ));
 sg13g2_dfrbp_1 _1319_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net32),
    .D(net296),
    .Q_N(_0628_),
    .Q(\SPI_driver1.digit_count[5] ));
 sg13g2_dfrbp_1 _1320_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net33),
    .D(_0013_),
    .Q_N(_0629_),
    .Q(\SPI_driver1.digit_count[6] ));
 sg13g2_dfrbp_1 _1321_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net34),
    .D(net216),
    .Q_N(_0630_),
    .Q(\SPI_driver1.SPI_Master1.state[0] ));
 sg13g2_dfrbp_1 _1322_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net35),
    .D(net206),
    .Q_N(_0631_),
    .Q(\SPI_driver1.SPI_Master1.state[1] ));
 sg13g2_dfrbp_1 _1323_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net36),
    .D(_0006_),
    .Q_N(_0632_),
    .Q(\SPI_driver1.SPI_Master1.state[2] ));
 sg13g2_dfrbp_1 _1324_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net37),
    .D(_0001_),
    .Q_N(_0633_),
    .Q(\SPI_driver1.SPI_Master1.count_bit[0] ));
 sg13g2_dfrbp_1 _1325_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net38),
    .D(_0002_),
    .Q_N(_0634_),
    .Q(\SPI_driver1.SPI_Master1.count_bit[1] ));
 sg13g2_dfrbp_1 _1326_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net66),
    .D(_0003_),
    .Q_N(_0635_),
    .Q(\SPI_driver1.SPI_Master1.count_bit[2] ));
 sg13g2_dfrbp_1 _1327_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net26),
    .D(_0004_),
    .Q_N(_0624_),
    .Q(\SPI_driver1.SPI_Master1.count_bit[3] ));
 sg13g2_dfrbp_1 _1328_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net47),
    .D(net180),
    .Q_N(_0034_),
    .Q(\SPI_driver1.wait_count[0] ));
 sg13g2_dfrbp_1 _1329_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net45),
    .D(net316),
    .Q_N(_0623_),
    .Q(\SPI_driver1.wait_count[1] ));
 sg13g2_dfrbp_1 _1330_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net43),
    .D(net269),
    .Q_N(_0622_),
    .Q(\SPI_driver1.wait_count[2] ));
 sg13g2_dfrbp_1 _1331_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net41),
    .D(net203),
    .Q_N(_0621_),
    .Q(\SPI_driver1.wait_count[3] ));
 sg13g2_dfrbp_1 _1332_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net39),
    .D(net225),
    .Q_N(_0620_),
    .Q(\SPI_driver1.SPI_Master1.word_out[1] ));
 sg13g2_dfrbp_1 _1333_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net25),
    .D(net214),
    .Q_N(_0619_),
    .Q(\SPI_driver1.SPI_Master1.word_out[2] ));
 sg13g2_dfrbp_1 _1334_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net176),
    .D(net237),
    .Q_N(_0618_),
    .Q(\SPI_driver1.SPI_Master1.word_out[3] ));
 sg13g2_dfrbp_1 _1335_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net175),
    .D(net218),
    .Q_N(_0617_),
    .Q(\SPI_driver1.SPI_Master1.word_out[4] ));
 sg13g2_dfrbp_1 _1336_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net174),
    .D(net223),
    .Q_N(_0616_),
    .Q(\SPI_driver1.SPI_Master1.word_out[5] ));
 sg13g2_dfrbp_1 _1337_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net173),
    .D(_0044_),
    .Q_N(_0615_),
    .Q(\SPI_driver1.SPI_Master1.word_out[6] ));
 sg13g2_dfrbp_1 _1338_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net172),
    .D(net227),
    .Q_N(_0614_),
    .Q(\SPI_driver1.SPI_Master1.word_out[7] ));
 sg13g2_dfrbp_1 _1339_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net171),
    .D(net235),
    .Q_N(_0613_),
    .Q(\SPI_driver1.SPI_Master1.word_out[8] ));
 sg13g2_dfrbp_1 _1340_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net170),
    .D(net210),
    .Q_N(_0612_),
    .Q(\SPI_driver1.SPI_Master1.word_out[9] ));
 sg13g2_dfrbp_1 _1341_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net169),
    .D(net233),
    .Q_N(_0611_),
    .Q(\SPI_driver1.SPI_Master1.word_out[10] ));
 sg13g2_dfrbp_1 _1342_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net168),
    .D(net245),
    .Q_N(_0610_),
    .Q(\SPI_driver1.SPI_Master1.word_out[11] ));
 sg13g2_dfrbp_1 _1343_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net167),
    .D(_0050_),
    .Q_N(_0609_),
    .Q(\SPI_driver1.SPI_Master1.word_out[12] ));
 sg13g2_dfrbp_1 _1344_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net166),
    .D(net212),
    .Q_N(_0608_),
    .Q(\SPI_driver1.SPI_Master1.word_out[13] ));
 sg13g2_dfrbp_1 _1345_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net165),
    .D(_0052_),
    .Q_N(_0607_),
    .Q(\SPI_driver1.SPI_Master1.word_out[14] ));
 sg13g2_dfrbp_1 _1346_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net164),
    .D(net248),
    .Q_N(_0606_),
    .Q(\SPI_driver1.SPI_Master1.word_out[15] ));
 sg13g2_dfrbp_1 _1347_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net163),
    .D(net190),
    .Q_N(_0033_),
    .Q(\SPI_driver1.SPI_Master1.count_word[0] ));
 sg13g2_dfrbp_1 _1348_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net161),
    .D(net309),
    .Q_N(_0605_),
    .Q(\SPI_driver1.SPI_Master1.count_word[1] ));
 sg13g2_dfrbp_1 _1349_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net159),
    .D(_0056_),
    .Q_N(_0604_),
    .Q(\SPI_driver1.SPI_Master1.count_word[2] ));
 sg13g2_dfrbp_1 _1350_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net157),
    .D(net239),
    .Q_N(_0603_),
    .Q(\SPI_driver1.SPI_Master1.count_word[3] ));
 sg13g2_dfrbp_1 _1351_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net116),
    .D(net221),
    .Q_N(_0602_),
    .Q(\SPI_driver1.Cs ));
 sg13g2_dfrbp_1 _1352_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net114),
    .D(net199),
    .Q_N(_0601_),
    .Q(\SPI_driver1.SPI_Master1.sclk ));
 sg13g2_dfrbp_1 _1353_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net112),
    .D(net193),
    .Q_N(_0600_),
    .Q(\SPI_driver1.Mosi ));
 sg13g2_dfrbp_1 _1354_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net67),
    .D(net182),
    .Q_N(_0026_),
    .Q(\SPI_driver1.SPI_Master1.report_ready ));
 sg13g2_dfrbp_1 _1355_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net68),
    .D(_0111_),
    .Q_N(_0636_),
    .Q(\SPI_driver1.SPI_Master1.word_in[0] ));
 sg13g2_dfrbp_1 _1356_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net69),
    .D(_0118_),
    .Q_N(_0637_),
    .Q(\SPI_driver1.SPI_Master1.word_in[1] ));
 sg13g2_dfrbp_1 _1357_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net70),
    .D(_0119_),
    .Q_N(_0638_),
    .Q(\SPI_driver1.SPI_Master1.word_in[2] ));
 sg13g2_dfrbp_1 _1358_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net71),
    .D(_0120_),
    .Q_N(_0639_),
    .Q(\SPI_driver1.SPI_Master1.word_in[3] ));
 sg13g2_dfrbp_1 _1359_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net72),
    .D(_0121_),
    .Q_N(_0640_),
    .Q(\SPI_driver1.SPI_Master1.word_in[4] ));
 sg13g2_dfrbp_1 _1360_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net73),
    .D(_0122_),
    .Q_N(_0641_),
    .Q(\SPI_driver1.SPI_Master1.word_in[5] ));
 sg13g2_dfrbp_1 _1361_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net74),
    .D(_0123_),
    .Q_N(_0642_),
    .Q(\SPI_driver1.SPI_Master1.word_in[6] ));
 sg13g2_dfrbp_1 _1362_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net75),
    .D(_0124_),
    .Q_N(_0643_),
    .Q(\SPI_driver1.SPI_Master1.word_in[7] ));
 sg13g2_dfrbp_1 _1363_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net76),
    .D(_0125_),
    .Q_N(_0644_),
    .Q(\SPI_driver1.SPI_Master1.word_in[8] ));
 sg13g2_dfrbp_1 _1364_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net77),
    .D(net321),
    .Q_N(_0645_),
    .Q(\SPI_driver1.SPI_Master1.word_in[9] ));
 sg13g2_dfrbp_1 _1365_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net78),
    .D(_0112_),
    .Q_N(_0646_),
    .Q(\SPI_driver1.SPI_Master1.word_in[10] ));
 sg13g2_dfrbp_1 _1366_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net79),
    .D(_0113_),
    .Q_N(_0647_),
    .Q(\SPI_driver1.SPI_Master1.word_in[11] ));
 sg13g2_dfrbp_1 _1367_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net80),
    .D(_0114_),
    .Q_N(_0648_),
    .Q(\SPI_driver1.SPI_Master1.word_in[12] ));
 sg13g2_dfrbp_1 _1368_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net81),
    .D(_0115_),
    .Q_N(_0649_),
    .Q(\SPI_driver1.SPI_Master1.word_in[13] ));
 sg13g2_dfrbp_1 _1369_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net83),
    .D(_0116_),
    .Q_N(_0650_),
    .Q(\SPI_driver1.SPI_Master1.word_in[14] ));
 sg13g2_dfrbp_1 _1370_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net110),
    .D(_0117_),
    .Q_N(_0599_),
    .Q(\SPI_driver1.SPI_Master1.word_in[15] ));
 sg13g2_dfrbp_1 _1371_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net84),
    .D(net230),
    .Q_N(_0651_),
    .Q(\SPI_driver1.SPI_Master1.word_out[0] ));
 sg13g2_dfrbp_1 _1372_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net85),
    .D(_0015_),
    .Q_N(_0024_),
    .Q(\SPI_driver1.SPI_Master1.res ));
 sg13g2_dfrbp_1 _1373_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net86),
    .D(net298),
    .Q_N(_0014_),
    .Q(\SPI_driver1.SPI_Master1.send_order ));
 sg13g2_dfrbp_1 _1374_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net87),
    .D(_0020_),
    .Q_N(_0652_),
    .Q(\SPI_driver1.sent_TST ));
 sg13g2_dfrbp_1 _1375_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net88),
    .D(_0019_),
    .Q_N(_0653_),
    .Q(\SPI_driver1.sent_SCN ));
 sg13g2_dfrbp_1 _1376_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net89),
    .D(_0017_),
    .Q_N(_0654_),
    .Q(\SPI_driver1.sent_LUX ));
 sg13g2_dfrbp_1 _1377_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net82),
    .D(_0016_),
    .Q_N(_0655_),
    .Q(\SPI_driver1.sent_BCD ));
 sg13g2_dfrbp_1 _1378_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net108),
    .D(_0018_),
    .Q_N(_0598_),
    .Q(\SPI_driver1.sent_PWR ));
 sg13g2_dfrbp_1 _1379_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net106),
    .D(net258),
    .Q_N(_0597_),
    .Q(\clockDivider1.counter[0] ));
 sg13g2_dfrbp_1 _1380_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net104),
    .D(net276),
    .Q_N(_0596_),
    .Q(\clockDivider1.counter[1] ));
 sg13g2_dfrbp_1 _1381_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net102),
    .D(net265),
    .Q_N(_0595_),
    .Q(\clockDivider1.counter[2] ));
 sg13g2_dfrbp_1 _1382_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net100),
    .D(_0066_),
    .Q_N(_0594_),
    .Q(\clockDivider1.counter[3] ));
 sg13g2_dfrbp_1 _1383_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net98),
    .D(_0067_),
    .Q_N(_0593_),
    .Q(\clockDivider1.counter[4] ));
 sg13g2_dfrbp_1 _1384_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net96),
    .D(net273),
    .Q_N(_0592_),
    .Q(\clockDivider1.counter[5] ));
 sg13g2_dfrbp_1 _1385_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net94),
    .D(_0069_),
    .Q_N(_0591_),
    .Q(\clockDivider1.counter[6] ));
 sg13g2_dfrbp_1 _1386_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net92),
    .D(net279),
    .Q_N(_0590_),
    .Q(\clockDivider1.counter[7] ));
 sg13g2_dfrbp_1 _1387_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net90),
    .D(net252),
    .Q_N(_0589_),
    .Q(\clockDivider1.counter[8] ));
 sg13g2_dfrbp_1 _1388_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net65),
    .D(net255),
    .Q_N(_0588_),
    .Q(\clockDivider1.counter[9] ));
 sg13g2_dfrbp_1 _1389_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net63),
    .D(net324),
    .Q_N(_0587_),
    .Q(\clockDivider1.counter[10] ));
 sg13g2_dfrbp_1 _1390_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net61),
    .D(net286),
    .Q_N(_0586_),
    .Q(\clockDivider1.counter[11] ));
 sg13g2_dfrbp_1 _1391_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net59),
    .D(_0075_),
    .Q_N(_0585_),
    .Q(\clockDivider1.counter[12] ));
 sg13g2_dfrbp_1 _1392_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net57),
    .D(_0076_),
    .Q_N(_0025_),
    .Q(\clockDivider1.counter[13] ));
 sg13g2_dfrbp_1 _1393_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net55),
    .D(net242),
    .Q_N(_0021_),
    .Q(\SPI_driver1.clk_div ));
 sg13g2_dfrbp_1 _1394_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net53),
    .D(net178),
    .Q_N(_0022_),
    .Q(\clockDivider1.ena ));
 sg13g2_dfrbp_1 _1395_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net51),
    .D(net197),
    .Q_N(_0023_),
    .Q(\SPI_driver1.ena ));
 sg13g2_dfrbp_1 _1396_ (.CLK(net136),
    .RESET_B(net49),
    .D(_0080_),
    .Q_N(_0029_),
    .Q(\SPI_driver1.min_X0[0] ));
 sg13g2_dfrbp_1 _1397_ (.CLK(net136),
    .RESET_B(net46),
    .D(_0081_),
    .Q_N(_0584_),
    .Q(\SPI_driver1.min_X0[1] ));
 sg13g2_dfrbp_1 _1398_ (.CLK(net137),
    .RESET_B(net42),
    .D(_0082_),
    .Q_N(_0030_),
    .Q(\SPI_driver1.min_X0[2] ));
 sg13g2_dfrbp_1 _1399_ (.CLK(net136),
    .RESET_B(net162),
    .D(_0083_),
    .Q_N(_0583_),
    .Q(\counter_chain1.inst_min_0X.max ));
 sg13g2_dfrbp_1 _1400_ (.CLK(net136),
    .RESET_B(net158),
    .D(_0084_),
    .Q_N(_0582_),
    .Q(\SPI_driver1.min_0X[0] ));
 sg13g2_dfrbp_1 _1401_ (.CLK(net137),
    .RESET_B(net115),
    .D(_0085_),
    .Q_N(_0581_),
    .Q(\SPI_driver1.min_0X[1] ));
 sg13g2_dfrbp_1 _1402_ (.CLK(net137),
    .RESET_B(net111),
    .D(_0086_),
    .Q_N(_0580_),
    .Q(\SPI_driver1.min_0X[2] ));
 sg13g2_dfrbp_1 _1403_ (.CLK(net137),
    .RESET_B(net107),
    .D(_0087_),
    .Q_N(_0579_),
    .Q(\SPI_driver1.min_0X[3] ));
 sg13g2_dfrbp_1 _1404_ (.CLK(net139),
    .RESET_B(net103),
    .D(_0088_),
    .Q_N(_0578_),
    .Q(\counter_chain1.inst_sec_X0.max ));
 sg13g2_dfrbp_1 _1405_ (.CLK(net139),
    .RESET_B(net99),
    .D(_0089_),
    .Q_N(_0031_),
    .Q(\SPI_driver1.sec_X0[0] ));
 sg13g2_dfrbp_1 _1406_ (.CLK(net138),
    .RESET_B(net95),
    .D(_0090_),
    .Q_N(_0577_),
    .Q(\SPI_driver1.sec_X0[1] ));
 sg13g2_dfrbp_1 _1407_ (.CLK(net138),
    .RESET_B(net91),
    .D(_0091_),
    .Q_N(_0032_),
    .Q(\SPI_driver1.sec_X0[2] ));
 sg13g2_dfrbp_1 _1408_ (.CLK(net138),
    .RESET_B(net64),
    .D(_0092_),
    .Q_N(_0576_),
    .Q(\counter_chain1.inst_sec_0X.max ));
 sg13g2_dfrbp_1 _1409_ (.CLK(net138),
    .RESET_B(net60),
    .D(_0093_),
    .Q_N(_0575_),
    .Q(\SPI_driver1.sec_0X[0] ));
 sg13g2_dfrbp_1 _1410_ (.CLK(net138),
    .RESET_B(net56),
    .D(_0094_),
    .Q_N(_0574_),
    .Q(\SPI_driver1.sec_0X[1] ));
 sg13g2_dfrbp_1 _1411_ (.CLK(net138),
    .RESET_B(net52),
    .D(_0095_),
    .Q_N(_0573_),
    .Q(\SPI_driver1.sec_0X[2] ));
 sg13g2_dfrbp_1 _1412_ (.CLK(net138),
    .RESET_B(net48),
    .D(_0096_),
    .Q_N(_0572_),
    .Q(\SPI_driver1.sec_0X[3] ));
 sg13g2_dfrbp_1 _1413_ (.CLK(net138),
    .RESET_B(net40),
    .D(_0097_),
    .Q_N(_0571_),
    .Q(\counter_chain1.inst_ces_X0.max ));
 sg13g2_dfrbp_1 _1414_ (.CLK(net136),
    .RESET_B(net117),
    .D(_0098_),
    .Q_N(_0570_),
    .Q(\SPI_driver1.ces_X0[0] ));
 sg13g2_dfrbp_1 _1415_ (.CLK(net136),
    .RESET_B(net109),
    .D(_0099_),
    .Q_N(_0569_),
    .Q(\SPI_driver1.ces_X0[1] ));
 sg13g2_dfrbp_1 _1416_ (.CLK(net136),
    .RESET_B(net101),
    .D(_0100_),
    .Q_N(_0568_),
    .Q(\SPI_driver1.ces_X0[2] ));
 sg13g2_dfrbp_1 _1417_ (.CLK(net136),
    .RESET_B(net93),
    .D(_0101_),
    .Q_N(_0567_),
    .Q(\SPI_driver1.ces_X0[3] ));
 sg13g2_dfrbp_1 _1418_ (.CLK(net139),
    .RESET_B(net62),
    .D(_0102_),
    .Q_N(_0566_),
    .Q(\counter_chain1.ces_X0_ena ));
 sg13g2_dfrbp_1 _1419_ (.CLK(net139),
    .RESET_B(net54),
    .D(_0103_),
    .Q_N(_0565_),
    .Q(\SPI_driver1.ces_0X[0] ));
 sg13g2_dfrbp_1 _1420_ (.CLK(net139),
    .RESET_B(net44),
    .D(_0104_),
    .Q_N(_0564_),
    .Q(\SPI_driver1.ces_0X[1] ));
 sg13g2_dfrbp_1 _1421_ (.CLK(net139),
    .RESET_B(net113),
    .D(_0105_),
    .Q_N(_0563_),
    .Q(\SPI_driver1.ces_0X[2] ));
 sg13g2_dfrbp_1 _1422_ (.CLK(net139),
    .RESET_B(net97),
    .D(_0106_),
    .Q_N(_0562_),
    .Q(\SPI_driver1.ces_0X[3] ));
 sg13g2_dfrbp_1 _1423_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net58),
    .D(net282),
    .Q_N(_0561_),
    .Q(\SPI_driver1.state[3] ));
 sg13g2_dfrbp_1 _1424_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net50),
    .D(_0108_),
    .Q_N(_0560_),
    .Q(\SPI_driver1.state[2] ));
 sg13g2_dfrbp_1 _1425_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net160),
    .D(_0109_),
    .Q_N(_0559_),
    .Q(\SPI_driver1.state[1] ));
 sg13g2_dfrbp_1 _1426_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net105),
    .D(_0110_),
    .Q_N(_0558_),
    .Q(\SPI_driver1.state[0] ));
 sg13g2_tiehi _1327__26 (.L_HI(net26));
 sg13g2_tiehi _1314__27 (.L_HI(net27));
 sg13g2_tiehi _1315__28 (.L_HI(net28));
 sg13g2_tiehi _1316__29 (.L_HI(net29));
 sg13g2_tiehi _1317__30 (.L_HI(net30));
 sg13g2_tiehi _1318__31 (.L_HI(net31));
 sg13g2_tiehi _1319__32 (.L_HI(net32));
 sg13g2_tiehi _1320__33 (.L_HI(net33));
 sg13g2_tiehi _1321__34 (.L_HI(net34));
 sg13g2_tiehi _1322__35 (.L_HI(net35));
 sg13g2_tiehi _1323__36 (.L_HI(net36));
 sg13g2_tiehi _1324__37 (.L_HI(net37));
 sg13g2_tiehi _1325__38 (.L_HI(net38));
 sg13g2_tiehi _1332__39 (.L_HI(net39));
 sg13g2_tiehi _1413__40 (.L_HI(net40));
 sg13g2_tiehi _1331__41 (.L_HI(net41));
 sg13g2_tiehi _1398__42 (.L_HI(net42));
 sg13g2_tiehi _1330__43 (.L_HI(net43));
 sg13g2_tiehi _1420__44 (.L_HI(net44));
 sg13g2_tiehi _1329__45 (.L_HI(net45));
 sg13g2_tiehi _1397__46 (.L_HI(net46));
 sg13g2_tiehi _1328__47 (.L_HI(net47));
 sg13g2_tiehi _1412__48 (.L_HI(net48));
 sg13g2_tiehi _1396__49 (.L_HI(net49));
 sg13g2_tiehi _1424__50 (.L_HI(net50));
 sg13g2_tiehi _1395__51 (.L_HI(net51));
 sg13g2_tiehi _1411__52 (.L_HI(net52));
 sg13g2_tiehi _1394__53 (.L_HI(net53));
 sg13g2_tiehi _1419__54 (.L_HI(net54));
 sg13g2_tiehi _1393__55 (.L_HI(net55));
 sg13g2_tiehi _1410__56 (.L_HI(net56));
 sg13g2_tiehi _1392__57 (.L_HI(net57));
 sg13g2_tiehi _1423__58 (.L_HI(net58));
 sg13g2_tiehi _1391__59 (.L_HI(net59));
 sg13g2_tiehi _1409__60 (.L_HI(net60));
 sg13g2_tiehi _1390__61 (.L_HI(net61));
 sg13g2_tiehi _1418__62 (.L_HI(net62));
 sg13g2_tiehi _1389__63 (.L_HI(net63));
 sg13g2_tiehi _1408__64 (.L_HI(net64));
 sg13g2_tiehi _1388__65 (.L_HI(net65));
 sg13g2_tiehi _1326__66 (.L_HI(net66));
 sg13g2_tiehi _1354__67 (.L_HI(net67));
 sg13g2_tiehi _1355__68 (.L_HI(net68));
 sg13g2_tiehi _1356__69 (.L_HI(net69));
 sg13g2_tiehi _1357__70 (.L_HI(net70));
 sg13g2_tiehi _1358__71 (.L_HI(net71));
 sg13g2_tiehi _1359__72 (.L_HI(net72));
 sg13g2_tiehi _1360__73 (.L_HI(net73));
 sg13g2_tiehi _1361__74 (.L_HI(net74));
 sg13g2_tiehi _1362__75 (.L_HI(net75));
 sg13g2_tiehi _1363__76 (.L_HI(net76));
 sg13g2_tiehi _1364__77 (.L_HI(net77));
 sg13g2_tiehi _1365__78 (.L_HI(net78));
 sg13g2_tiehi _1366__79 (.L_HI(net79));
 sg13g2_tiehi _1367__80 (.L_HI(net80));
 sg13g2_tiehi _1368__81 (.L_HI(net81));
 sg13g2_tiehi _1377__82 (.L_HI(net82));
 sg13g2_tiehi _1369__83 (.L_HI(net83));
 sg13g2_tiehi _1371__84 (.L_HI(net84));
 sg13g2_tiehi _1372__85 (.L_HI(net85));
 sg13g2_tiehi _1373__86 (.L_HI(net86));
 sg13g2_tiehi _1374__87 (.L_HI(net87));
 sg13g2_tiehi _1375__88 (.L_HI(net88));
 sg13g2_tiehi _1376__89 (.L_HI(net89));
 sg13g2_tiehi _1387__90 (.L_HI(net90));
 sg13g2_tiehi _1407__91 (.L_HI(net91));
 sg13g2_tiehi _1386__92 (.L_HI(net92));
 sg13g2_tiehi _1417__93 (.L_HI(net93));
 sg13g2_tiehi _1385__94 (.L_HI(net94));
 sg13g2_tiehi _1406__95 (.L_HI(net95));
 sg13g2_tiehi _1384__96 (.L_HI(net96));
 sg13g2_tiehi _1422__97 (.L_HI(net97));
 sg13g2_tiehi _1383__98 (.L_HI(net98));
 sg13g2_tiehi _1405__99 (.L_HI(net99));
 sg13g2_tiehi _1382__100 (.L_HI(net100));
 sg13g2_tiehi _1416__101 (.L_HI(net101));
 sg13g2_tiehi _1381__102 (.L_HI(net102));
 sg13g2_tiehi _1404__103 (.L_HI(net103));
 sg13g2_tiehi _1380__104 (.L_HI(net104));
 sg13g2_tiehi _1426__105 (.L_HI(net105));
 sg13g2_tiehi _1379__106 (.L_HI(net106));
 sg13g2_tiehi _1403__107 (.L_HI(net107));
 sg13g2_tiehi _1378__108 (.L_HI(net108));
 sg13g2_tiehi _1415__109 (.L_HI(net109));
 sg13g2_tiehi _1370__110 (.L_HI(net110));
 sg13g2_tiehi _1402__111 (.L_HI(net111));
 sg13g2_tiehi _1353__112 (.L_HI(net112));
 sg13g2_tiehi _1421__113 (.L_HI(net113));
 sg13g2_tiehi _1352__114 (.L_HI(net114));
 sg13g2_tiehi _1401__115 (.L_HI(net115));
 sg13g2_tiehi _1351__116 (.L_HI(net116));
 sg13g2_tiehi _1414__117 (.L_HI(net117));
 sg13g2_tiehi _1350__118 (.L_HI(net157));
 sg13g2_tiehi _1400__119 (.L_HI(net158));
 sg13g2_tiehi _1349__120 (.L_HI(net159));
 sg13g2_tiehi _1425__121 (.L_HI(net160));
 sg13g2_tiehi _1348__122 (.L_HI(net161));
 sg13g2_tiehi _1399__123 (.L_HI(net162));
 sg13g2_tiehi _1347__124 (.L_HI(net163));
 sg13g2_tiehi _1346__125 (.L_HI(net164));
 sg13g2_tiehi _1345__126 (.L_HI(net165));
 sg13g2_tiehi _1344__127 (.L_HI(net166));
 sg13g2_tiehi _1343__128 (.L_HI(net167));
 sg13g2_tiehi _1342__129 (.L_HI(net168));
 sg13g2_tiehi _1341__130 (.L_HI(net169));
 sg13g2_tiehi _1340__131 (.L_HI(net170));
 sg13g2_tiehi _1339__132 (.L_HI(net171));
 sg13g2_tiehi _1338__133 (.L_HI(net172));
 sg13g2_tiehi _1337__134 (.L_HI(net173));
 sg13g2_tiehi _1336__135 (.L_HI(net174));
 sg13g2_tiehi _1335__136 (.L_HI(net175));
 sg13g2_tiehi _1334__137 (.L_HI(net176));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_faramire_stopwatch_7 (.L_LO(net7));
 sg13g2_tielo tt_um_faramire_stopwatch_8 (.L_LO(net8));
 sg13g2_tielo tt_um_faramire_stopwatch_9 (.L_LO(net9));
 sg13g2_tielo tt_um_faramire_stopwatch_10 (.L_LO(net10));
 sg13g2_tielo tt_um_faramire_stopwatch_11 (.L_LO(net11));
 sg13g2_tielo tt_um_faramire_stopwatch_12 (.L_LO(net12));
 sg13g2_tielo tt_um_faramire_stopwatch_13 (.L_LO(net13));
 sg13g2_tielo tt_um_faramire_stopwatch_14 (.L_LO(net14));
 sg13g2_tielo tt_um_faramire_stopwatch_15 (.L_LO(net15));
 sg13g2_tielo tt_um_faramire_stopwatch_16 (.L_LO(net16));
 sg13g2_tielo tt_um_faramire_stopwatch_17 (.L_LO(net17));
 sg13g2_tielo tt_um_faramire_stopwatch_18 (.L_LO(net18));
 sg13g2_tielo tt_um_faramire_stopwatch_19 (.L_LO(net19));
 sg13g2_tielo tt_um_faramire_stopwatch_20 (.L_LO(net20));
 sg13g2_tielo tt_um_faramire_stopwatch_21 (.L_LO(net21));
 sg13g2_tielo tt_um_faramire_stopwatch_22 (.L_LO(net22));
 sg13g2_tielo tt_um_faramire_stopwatch_23 (.L_LO(net23));
 sg13g2_tielo tt_um_faramire_stopwatch_24 (.L_LO(net24));
 sg13g2_tiehi _1333__25 (.L_HI(net25));
 sg13g2_buf_1 _1559_ (.A(\SPI_driver1.Mosi ),
    .X(uo_out[0]));
 sg13g2_buf_1 _1560_ (.A(\SPI_driver1.Cs ),
    .X(uo_out[1]));
 sg13g2_buf_1 _1561_ (.A(\SPI_driver1.SPI_Master1.sclk ),
    .X(uo_out[2]));
 sg13g2_buf_1 _1562_ (.A(net135),
    .X(uo_out[3]));
 sg13g2_buf_1 _1563_ (.A(\SPI_driver1.ena ),
    .X(uo_out[4]));
 sg13g2_buf_2 fanout118 (.A(net120),
    .X(net118));
 sg13g2_buf_1 fanout119 (.A(net120),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_0334_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(net122),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_0334_),
    .X(net122));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(_0246_));
 sg13g2_buf_2 fanout124 (.A(net125),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_0406_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(net128),
    .X(net126));
 sg13g2_buf_1 fanout127 (.A(net128),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(\SPI_driver1.state[0] ),
    .X(net128));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(\SPI_driver1.state[1] ));
 sg13g2_buf_1 fanout130 (.A(\SPI_driver1.state[1] ),
    .X(net130));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(\SPI_driver1.state[2] ));
 sg13g2_buf_2 fanout132 (.A(\SPI_driver1.state[3] ),
    .X(net132));
 sg13g2_buf_1 fanout133 (.A(\SPI_driver1.state[3] ),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(net135),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(\clockDivider1.ena ),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(net140),
    .X(net136));
 sg13g2_buf_1 fanout137 (.A(net140),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(\SPI_driver1.clk_div ),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(net311),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(net144),
    .X(net142));
 sg13g2_buf_1 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_0026_),
    .X(net144));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(net270));
 sg13g2_buf_2 fanout146 (.A(net149),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(net149),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(\SPI_driver1.SPI_Master1.state[2] ),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(\SPI_driver1.SPI_Master1.state[2] ),
    .X(net150));
 sg13g2_buf_1 fanout151 (.A(\SPI_driver1.SPI_Master1.state[2] ),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(net153),
    .X(net152));
 sg13g2_buf_1 fanout153 (.A(net156),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(net156),
    .X(net154));
 sg13g2_buf_1 fanout155 (.A(net156),
    .X(net155));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(net1));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_tielo tt_um_faramire_stopwatch_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0022_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0078_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0034_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0035_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0014_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0061_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold7 (.A(\SPI_driver1.SPI_Master1.word_in[15] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold8 (.A(\SPI_driver1.SPI_Master1.word_in[12] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold9 (.A(\SPI_driver1.SPI_Master1.word_in[14] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold10 (.A(\SPI_driver1.SPI_Master1.word_in[13] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold11 (.A(\SPI_driver1.SPI_Master1.word_in[6] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold12 (.A(\clockDivider1.counter[13] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0033_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0054_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold15 (.A(\SPI_driver1.Mosi ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0392_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0060_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold18 (.A(\SPI_driver1.SPI_Master1.count_bit[2] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0170_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0023_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0079_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold22 (.A(\SPI_driver1.SPI_Master1.count_bit[1] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0059_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold24 (.A(\SPI_driver1.SPI_Master1.state[0] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0154_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold26 (.A(\SPI_driver1.wait_count[3] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0038_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0024_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0162_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0000_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold31 (.A(\SPI_driver1.digit_count[3] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0010_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold33 (.A(\SPI_driver1.SPI_Master1.word_out[9] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0047_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold35 (.A(\SPI_driver1.SPI_Master1.word_out[13] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0051_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold37 (.A(\SPI_driver1.SPI_Master1.word_out[2] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0040_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold39 (.A(\SPI_driver1.SPI_Master1.state[1] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0005_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold41 (.A(\SPI_driver1.SPI_Master1.word_out[4] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0042_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold43 (.A(\SPI_driver1.Cs ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0389_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0058_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold46 (.A(\SPI_driver1.SPI_Master1.word_out[5] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0043_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold48 (.A(\SPI_driver1.SPI_Master1.word_out[1] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0039_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold50 (.A(\SPI_driver1.SPI_Master1.word_out[7] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0045_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold52 (.A(\SPI_driver1.SPI_Master1.word_out[14] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold53 (.A(\SPI_driver1.SPI_Master1.word_in[0] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0062_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold55 (.A(\SPI_driver1.SPI_Master1.word_in[7] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold56 (.A(\SPI_driver1.SPI_Master1.word_out[10] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0048_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold58 (.A(\SPI_driver1.SPI_Master1.word_out[8] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0046_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold60 (.A(\SPI_driver1.SPI_Master1.word_out[3] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0041_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold62 (.A(\SPI_driver1.SPI_Master1.count_word[3] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0057_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0021_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0446_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0077_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold67 (.A(\SPI_driver1.SPI_Master1.word_out[6] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold68 (.A(\SPI_driver1.SPI_Master1.word_out[11] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0049_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold70 (.A(\SPI_driver1.SPI_Master1.word_out[12] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold71 (.A(\SPI_driver1.SPI_Master1.word_out[15] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0053_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold73 (.A(\SPI_driver1.SPI_Master1.count_bit[3] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold74 (.A(\clockDivider1.counter[8] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0433_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0071_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold77 (.A(\SPI_driver1.SPI_Master1.word_in[1] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold78 (.A(\clockDivider1.counter[9] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0072_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold80 (.A(\clockDivider1.counter[0] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0404_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0063_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold83 (.A(\SPI_driver1.SPI_Master1.word_in[4] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold84 (.A(\clockDivider1.counter[6] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0427_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold86 (.A(\SPI_driver1.SPI_Master1.word_in[5] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold87 (.A(\clockDivider1.counter[2] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0417_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0065_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold90 (.A(\SPI_driver1.SPI_Master1.count_word[2] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0388_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold92 (.A(\SPI_driver1.wait_count[2] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0037_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold94 (.A(\SPI_driver1.SPI_Master1.report_ready ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0227_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold96 (.A(\clockDivider1.counter[5] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0068_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold98 (.A(\clockDivider1.counter[1] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0415_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0064_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold101 (.A(\clockDivider1.counter[3] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold102 (.A(\clockDivider1.counter[7] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0070_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0028_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0525_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0107_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold107 (.A(\SPI_driver1.sent_PWR ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold108 (.A(\SPI_driver1.sent_SCN ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold109 (.A(\clockDivider1.counter[11] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0074_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold111 (.A(\clockDivider1.counter[4] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold112 (.A(\SPI_driver1.sent_TST ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold113 (.A(\SPI_driver1.SPI_Master1.word_in[10] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold114 (.A(\SPI_driver1.SPI_Master1.word_in[3] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold115 (.A(\SPI_driver1.digit_count[6] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0192_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0008_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold118 (.A(\SPI_driver1.digit_count[1] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0197_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0012_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold121 (.A(\SPI_driver1.SPI_Master1.send_order ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0769_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold123 (.A(\SPI_driver1.sent_BCD ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold124 (.A(\SPI_driver1.digit_count[4] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0179_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0009_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold127 (.A(\SPI_driver1.SPI_Master1.count_bit[0] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold128 (.A(\SPI_driver1.digit_count[0] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0196_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0027_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold131 (.A(\SPI_driver1.SPI_Master1.count_word[1] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0385_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0055_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold134 (.A(\SPI_driver1.sent_LUX ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold135 (.A(\SPI_driver1.SPI_Master1.res ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0165_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold137 (.A(\SPI_driver1.digit_count[2] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold138 (.A(\SPI_driver1.wait_count[1] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0330_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0036_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold141 (.A(\SPI_driver1.SPI_Master1.word_in[11] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold142 (.A(\clockDivider1.counter[12] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0445_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold144 (.A(\SPI_driver1.SPI_Master1.word_in[9] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0126_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold146 (.A(\SPI_driver1.SPI_Master1.word_in[8] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold147 (.A(\clockDivider1.counter[10] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0073_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold149 (.A(\SPI_driver1.SPI_Master1.word_in[2] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold150 (.A(\SPI_driver1.ena ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold151 (.A(\clockDivider1.counter[4] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0428_),
    .X(net328));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_fill_2 FILLER_15_119 ();
 sg13g2_fill_1 FILLER_15_121 ();
 sg13g2_decap_4 FILLER_15_126 ();
 sg13g2_fill_2 FILLER_15_130 ();
 sg13g2_decap_8 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_decap_8 FILLER_15_172 ();
 sg13g2_decap_8 FILLER_15_179 ();
 sg13g2_decap_8 FILLER_15_186 ();
 sg13g2_decap_8 FILLER_15_193 ();
 sg13g2_decap_8 FILLER_15_200 ();
 sg13g2_decap_8 FILLER_15_207 ();
 sg13g2_decap_4 FILLER_15_218 ();
 sg13g2_fill_1 FILLER_15_222 ();
 sg13g2_fill_2 FILLER_15_231 ();
 sg13g2_decap_4 FILLER_15_238 ();
 sg13g2_fill_2 FILLER_15_242 ();
 sg13g2_decap_8 FILLER_15_274 ();
 sg13g2_decap_8 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_295 ();
 sg13g2_decap_4 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_352 ();
 sg13g2_decap_8 FILLER_15_359 ();
 sg13g2_decap_8 FILLER_15_366 ();
 sg13g2_decap_8 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_4 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_125 ();
 sg13g2_fill_2 FILLER_16_131 ();
 sg13g2_decap_8 FILLER_16_146 ();
 sg13g2_decap_8 FILLER_16_153 ();
 sg13g2_decap_8 FILLER_16_160 ();
 sg13g2_decap_8 FILLER_16_167 ();
 sg13g2_decap_8 FILLER_16_174 ();
 sg13g2_decap_8 FILLER_16_181 ();
 sg13g2_decap_8 FILLER_16_188 ();
 sg13g2_decap_8 FILLER_16_195 ();
 sg13g2_fill_1 FILLER_16_202 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_4 FILLER_16_266 ();
 sg13g2_fill_2 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_298 ();
 sg13g2_fill_2 FILLER_16_305 ();
 sg13g2_fill_1 FILLER_16_311 ();
 sg13g2_decap_4 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_fill_1 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_4 FILLER_17_49 ();
 sg13g2_fill_2 FILLER_17_79 ();
 sg13g2_fill_2 FILLER_17_94 ();
 sg13g2_fill_2 FILLER_17_118 ();
 sg13g2_fill_2 FILLER_17_129 ();
 sg13g2_fill_2 FILLER_17_161 ();
 sg13g2_fill_1 FILLER_17_163 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_4 FILLER_17_203 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_decap_8 FILLER_17_213 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_4 FILLER_17_231 ();
 sg13g2_fill_2 FILLER_17_244 ();
 sg13g2_fill_1 FILLER_17_246 ();
 sg13g2_decap_8 FILLER_17_265 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_292 ();
 sg13g2_fill_1 FILLER_17_299 ();
 sg13g2_fill_1 FILLER_17_336 ();
 sg13g2_fill_1 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_18 ();
 sg13g2_decap_8 FILLER_18_23 ();
 sg13g2_fill_1 FILLER_18_30 ();
 sg13g2_decap_8 FILLER_18_57 ();
 sg13g2_fill_2 FILLER_18_68 ();
 sg13g2_fill_1 FILLER_18_70 ();
 sg13g2_fill_1 FILLER_18_97 ();
 sg13g2_fill_1 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_230 ();
 sg13g2_decap_8 FILLER_18_237 ();
 sg13g2_fill_1 FILLER_18_244 ();
 sg13g2_decap_4 FILLER_18_259 ();
 sg13g2_fill_2 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_300 ();
 sg13g2_decap_4 FILLER_18_307 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_4 FILLER_18_333 ();
 sg13g2_fill_2 FILLER_18_337 ();
 sg13g2_decap_4 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_62 ();
 sg13g2_fill_1 FILLER_19_78 ();
 sg13g2_fill_1 FILLER_19_133 ();
 sg13g2_fill_2 FILLER_19_139 ();
 sg13g2_fill_2 FILLER_19_184 ();
 sg13g2_decap_8 FILLER_19_190 ();
 sg13g2_decap_8 FILLER_19_197 ();
 sg13g2_decap_8 FILLER_19_204 ();
 sg13g2_fill_2 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_213 ();
 sg13g2_decap_8 FILLER_19_240 ();
 sg13g2_fill_2 FILLER_19_247 ();
 sg13g2_fill_2 FILLER_19_258 ();
 sg13g2_decap_4 FILLER_19_265 ();
 sg13g2_fill_2 FILLER_19_285 ();
 sg13g2_decap_8 FILLER_19_297 ();
 sg13g2_decap_4 FILLER_19_304 ();
 sg13g2_fill_1 FILLER_19_313 ();
 sg13g2_decap_4 FILLER_19_320 ();
 sg13g2_fill_2 FILLER_19_329 ();
 sg13g2_fill_1 FILLER_19_340 ();
 sg13g2_fill_2 FILLER_19_356 ();
 sg13g2_decap_4 FILLER_19_362 ();
 sg13g2_fill_1 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_fill_2 FILLER_19_379 ();
 sg13g2_fill_1 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_fill_2 FILLER_20_35 ();
 sg13g2_decap_4 FILLER_20_42 ();
 sg13g2_fill_1 FILLER_20_46 ();
 sg13g2_fill_2 FILLER_20_52 ();
 sg13g2_fill_1 FILLER_20_54 ();
 sg13g2_decap_4 FILLER_20_60 ();
 sg13g2_fill_1 FILLER_20_68 ();
 sg13g2_fill_2 FILLER_20_100 ();
 sg13g2_fill_1 FILLER_20_102 ();
 sg13g2_decap_8 FILLER_20_107 ();
 sg13g2_fill_1 FILLER_20_114 ();
 sg13g2_fill_2 FILLER_20_164 ();
 sg13g2_fill_1 FILLER_20_166 ();
 sg13g2_fill_1 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_229 ();
 sg13g2_fill_2 FILLER_20_236 ();
 sg13g2_fill_2 FILLER_20_248 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_decap_8 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_fill_1 FILLER_20_339 ();
 sg13g2_fill_2 FILLER_20_350 ();
 sg13g2_fill_2 FILLER_20_356 ();
 sg13g2_fill_1 FILLER_20_358 ();
 sg13g2_fill_1 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_23 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_fill_2 FILLER_21_175 ();
 sg13g2_fill_2 FILLER_21_181 ();
 sg13g2_decap_8 FILLER_21_192 ();
 sg13g2_decap_4 FILLER_21_199 ();
 sg13g2_fill_1 FILLER_21_203 ();
 sg13g2_fill_1 FILLER_21_208 ();
 sg13g2_decap_8 FILLER_21_213 ();
 sg13g2_fill_2 FILLER_21_220 ();
 sg13g2_fill_2 FILLER_21_236 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_decap_4 FILLER_21_256 ();
 sg13g2_fill_2 FILLER_21_260 ();
 sg13g2_decap_8 FILLER_21_268 ();
 sg13g2_decap_4 FILLER_21_280 ();
 sg13g2_fill_2 FILLER_21_288 ();
 sg13g2_decap_8 FILLER_21_299 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_fill_2 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_fill_2 FILLER_21_361 ();
 sg13g2_fill_1 FILLER_21_383 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_4 ();
 sg13g2_fill_2 FILLER_22_32 ();
 sg13g2_fill_2 FILLER_22_43 ();
 sg13g2_fill_1 FILLER_22_45 ();
 sg13g2_fill_2 FILLER_22_51 ();
 sg13g2_fill_1 FILLER_22_53 ();
 sg13g2_decap_4 FILLER_22_71 ();
 sg13g2_fill_2 FILLER_22_75 ();
 sg13g2_fill_1 FILLER_22_103 ();
 sg13g2_fill_2 FILLER_22_123 ();
 sg13g2_fill_2 FILLER_22_135 ();
 sg13g2_fill_1 FILLER_22_177 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_4 FILLER_22_189 ();
 sg13g2_fill_2 FILLER_22_219 ();
 sg13g2_fill_1 FILLER_22_230 ();
 sg13g2_decap_4 FILLER_22_257 ();
 sg13g2_fill_1 FILLER_22_261 ();
 sg13g2_fill_1 FILLER_22_273 ();
 sg13g2_decap_4 FILLER_22_312 ();
 sg13g2_fill_2 FILLER_22_342 ();
 sg13g2_decap_4 FILLER_22_349 ();
 sg13g2_fill_2 FILLER_22_353 ();
 sg13g2_fill_2 FILLER_22_376 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_14 ();
 sg13g2_fill_1 FILLER_23_137 ();
 sg13g2_fill_1 FILLER_23_154 ();
 sg13g2_fill_2 FILLER_23_159 ();
 sg13g2_fill_2 FILLER_23_193 ();
 sg13g2_fill_1 FILLER_23_195 ();
 sg13g2_fill_2 FILLER_23_230 ();
 sg13g2_fill_2 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_fill_2 FILLER_23_273 ();
 sg13g2_fill_1 FILLER_23_275 ();
 sg13g2_fill_2 FILLER_23_284 ();
 sg13g2_fill_1 FILLER_23_286 ();
 sg13g2_decap_8 FILLER_23_292 ();
 sg13g2_fill_2 FILLER_23_299 ();
 sg13g2_decap_4 FILLER_23_330 ();
 sg13g2_fill_1 FILLER_23_334 ();
 sg13g2_fill_2 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_8 FILLER_23_360 ();
 sg13g2_fill_2 FILLER_23_379 ();
 sg13g2_fill_2 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_4 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_35 ();
 sg13g2_fill_2 FILLER_24_45 ();
 sg13g2_fill_2 FILLER_24_92 ();
 sg13g2_fill_2 FILLER_24_117 ();
 sg13g2_decap_4 FILLER_24_127 ();
 sg13g2_fill_1 FILLER_24_131 ();
 sg13g2_decap_4 FILLER_24_193 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_decap_4 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_206 ();
 sg13g2_decap_8 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_222 ();
 sg13g2_decap_8 FILLER_24_229 ();
 sg13g2_decap_4 FILLER_24_236 ();
 sg13g2_fill_2 FILLER_24_240 ();
 sg13g2_fill_2 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_304 ();
 sg13g2_fill_2 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_331 ();
 sg13g2_fill_2 FILLER_24_336 ();
 sg13g2_fill_1 FILLER_24_338 ();
 sg13g2_fill_1 FILLER_24_347 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_46 ();
 sg13g2_fill_1 FILLER_25_48 ();
 sg13g2_fill_2 FILLER_25_53 ();
 sg13g2_fill_1 FILLER_25_55 ();
 sg13g2_fill_2 FILLER_25_74 ();
 sg13g2_fill_2 FILLER_25_104 ();
 sg13g2_fill_2 FILLER_25_111 ();
 sg13g2_fill_2 FILLER_25_147 ();
 sg13g2_fill_1 FILLER_25_149 ();
 sg13g2_fill_2 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_172 ();
 sg13g2_fill_1 FILLER_25_178 ();
 sg13g2_fill_2 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_256 ();
 sg13g2_fill_2 FILLER_25_309 ();
 sg13g2_fill_1 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_317 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_fill_1 FILLER_25_354 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_9 ();
 sg13g2_fill_1 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_90 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_fill_1 FILLER_26_106 ();
 sg13g2_fill_2 FILLER_26_111 ();
 sg13g2_fill_2 FILLER_26_121 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_fill_2 FILLER_26_128 ();
 sg13g2_fill_1 FILLER_26_130 ();
 sg13g2_fill_1 FILLER_26_160 ();
 sg13g2_fill_1 FILLER_26_225 ();
 sg13g2_fill_2 FILLER_26_230 ();
 sg13g2_fill_1 FILLER_26_232 ();
 sg13g2_fill_2 FILLER_26_310 ();
 sg13g2_fill_1 FILLER_26_312 ();
 sg13g2_fill_1 FILLER_26_343 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_59 ();
 sg13g2_fill_1 FILLER_27_61 ();
 sg13g2_fill_1 FILLER_27_95 ();
 sg13g2_fill_1 FILLER_27_101 ();
 sg13g2_decap_8 FILLER_27_128 ();
 sg13g2_fill_1 FILLER_27_135 ();
 sg13g2_fill_2 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_149 ();
 sg13g2_fill_2 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_fill_2 FILLER_27_179 ();
 sg13g2_fill_1 FILLER_27_181 ();
 sg13g2_decap_4 FILLER_27_228 ();
 sg13g2_fill_1 FILLER_27_232 ();
 sg13g2_fill_2 FILLER_27_327 ();
 sg13g2_fill_2 FILLER_27_355 ();
 sg13g2_fill_1 FILLER_28_59 ();
 sg13g2_fill_1 FILLER_28_110 ();
 sg13g2_fill_2 FILLER_28_137 ();
 sg13g2_fill_1 FILLER_28_153 ();
 sg13g2_fill_1 FILLER_28_159 ();
 sg13g2_fill_2 FILLER_28_170 ();
 sg13g2_fill_1 FILLER_28_172 ();
 sg13g2_fill_1 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_209 ();
 sg13g2_decap_8 FILLER_28_216 ();
 sg13g2_fill_2 FILLER_28_223 ();
 sg13g2_fill_1 FILLER_28_228 ();
 sg13g2_fill_1 FILLER_28_234 ();
 sg13g2_fill_1 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_307 ();
 sg13g2_fill_2 FILLER_28_326 ();
 sg13g2_fill_2 FILLER_28_370 ();
 sg13g2_fill_2 FILLER_28_381 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_44 ();
 sg13g2_fill_2 FILLER_29_71 ();
 sg13g2_fill_1 FILLER_29_73 ();
 sg13g2_fill_1 FILLER_29_93 ();
 sg13g2_fill_2 FILLER_29_114 ();
 sg13g2_fill_2 FILLER_29_146 ();
 sg13g2_fill_2 FILLER_29_166 ();
 sg13g2_decap_8 FILLER_29_193 ();
 sg13g2_fill_2 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_29_226 ();
 sg13g2_fill_2 FILLER_29_244 ();
 sg13g2_fill_1 FILLER_29_269 ();
 sg13g2_fill_2 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_333 ();
 sg13g2_fill_2 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_368 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_2 FILLER_30_26 ();
 sg13g2_fill_1 FILLER_30_43 ();
 sg13g2_fill_2 FILLER_30_83 ();
 sg13g2_fill_2 FILLER_30_94 ();
 sg13g2_fill_2 FILLER_30_122 ();
 sg13g2_fill_2 FILLER_30_155 ();
 sg13g2_decap_4 FILLER_30_198 ();
 sg13g2_fill_1 FILLER_30_202 ();
 sg13g2_fill_2 FILLER_30_219 ();
 sg13g2_fill_2 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_fill_1 FILLER_30_263 ();
 sg13g2_fill_2 FILLER_30_272 ();
 sg13g2_fill_2 FILLER_30_302 ();
 sg13g2_fill_2 FILLER_30_311 ();
 sg13g2_fill_1 FILLER_30_330 ();
 sg13g2_fill_1 FILLER_30_373 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_40 ();
 sg13g2_fill_1 FILLER_31_119 ();
 sg13g2_fill_2 FILLER_31_134 ();
 sg13g2_decap_4 FILLER_31_150 ();
 sg13g2_fill_2 FILLER_31_164 ();
 sg13g2_decap_8 FILLER_31_174 ();
 sg13g2_fill_2 FILLER_31_191 ();
 sg13g2_fill_1 FILLER_31_208 ();
 sg13g2_decap_4 FILLER_31_214 ();
 sg13g2_fill_1 FILLER_31_218 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_fill_1 FILLER_32_95 ();
 sg13g2_fill_2 FILLER_32_101 ();
 sg13g2_fill_1 FILLER_32_133 ();
 sg13g2_fill_2 FILLER_32_154 ();
 sg13g2_fill_2 FILLER_32_165 ();
 sg13g2_fill_1 FILLER_32_188 ();
 sg13g2_decap_8 FILLER_32_194 ();
 sg13g2_fill_2 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_203 ();
 sg13g2_fill_2 FILLER_32_217 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_226 ();
 sg13g2_fill_1 FILLER_32_228 ();
 sg13g2_decap_4 FILLER_32_245 ();
 sg13g2_fill_2 FILLER_32_249 ();
 sg13g2_fill_2 FILLER_32_274 ();
 sg13g2_fill_1 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_334 ();
 sg13g2_fill_1 FILLER_32_366 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_fill_2 FILLER_33_161 ();
 sg13g2_decap_4 FILLER_33_169 ();
 sg13g2_fill_2 FILLER_33_182 ();
 sg13g2_fill_2 FILLER_33_194 ();
 sg13g2_decap_4 FILLER_33_218 ();
 sg13g2_fill_1 FILLER_33_222 ();
 sg13g2_fill_2 FILLER_33_230 ();
 sg13g2_decap_4 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_fill_1 FILLER_33_360 ();
 sg13g2_fill_2 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_40 ();
 sg13g2_fill_1 FILLER_34_57 ();
 sg13g2_fill_2 FILLER_34_80 ();
 sg13g2_fill_1 FILLER_34_115 ();
 sg13g2_fill_2 FILLER_34_125 ();
 sg13g2_decap_8 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_160 ();
 sg13g2_fill_2 FILLER_34_195 ();
 sg13g2_fill_1 FILLER_34_202 ();
 sg13g2_decap_8 FILLER_34_213 ();
 sg13g2_decap_8 FILLER_34_220 ();
 sg13g2_fill_1 FILLER_34_234 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_122 ();
 sg13g2_fill_2 FILLER_35_176 ();
 sg13g2_fill_1 FILLER_35_178 ();
 sg13g2_fill_1 FILLER_35_189 ();
 sg13g2_fill_2 FILLER_35_305 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_55 ();
 sg13g2_fill_2 FILLER_36_100 ();
 sg13g2_fill_1 FILLER_36_111 ();
 sg13g2_fill_2 FILLER_36_117 ();
 sg13g2_fill_1 FILLER_36_124 ();
 sg13g2_decap_4 FILLER_36_156 ();
 sg13g2_fill_2 FILLER_36_160 ();
 sg13g2_fill_1 FILLER_36_202 ();
 sg13g2_decap_4 FILLER_36_214 ();
 sg13g2_fill_1 FILLER_36_218 ();
 sg13g2_fill_1 FILLER_36_301 ();
 sg13g2_fill_1 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_fill_2 FILLER_37_28 ();
 sg13g2_fill_1 FILLER_37_64 ();
 sg13g2_fill_1 FILLER_37_70 ();
 sg13g2_fill_2 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_135 ();
 sg13g2_fill_2 FILLER_37_140 ();
 sg13g2_fill_2 FILLER_37_174 ();
 sg13g2_fill_1 FILLER_37_176 ();
 sg13g2_fill_2 FILLER_37_349 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_111 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_148 ();
 sg13g2_fill_2 FILLER_38_174 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_fill_2 FILLER_38_200 ();
 sg13g2_fill_2 FILLER_38_211 ();
 sg13g2_fill_1 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_218 ();
 sg13g2_fill_1 FILLER_38_225 ();
 sg13g2_fill_1 FILLER_38_284 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net8;
 assign uio_oe[3] = net9;
 assign uio_oe[4] = net10;
 assign uio_oe[5] = net11;
 assign uio_oe[6] = net12;
 assign uio_oe[7] = net13;
 assign uio_out[0] = net14;
 assign uio_out[1] = net15;
 assign uio_out[2] = net16;
 assign uio_out[3] = net17;
 assign uio_out[4] = net18;
 assign uio_out[5] = net19;
 assign uio_out[6] = net20;
 assign uio_out[7] = net21;
 assign uo_out[5] = net22;
 assign uo_out[6] = net23;
 assign uo_out[7] = net24;
endmodule

module tt_um_dlfloatmac (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \MAC.a[0] ;
 wire \MAC.a[10] ;
 wire \MAC.a[11] ;
 wire \MAC.a[12] ;
 wire \MAC.a[13] ;
 wire \MAC.a[14] ;
 wire \MAC.a[15] ;
 wire \MAC.a[1] ;
 wire \MAC.a[2] ;
 wire \MAC.a[3] ;
 wire \MAC.a[4] ;
 wire \MAC.a[5] ;
 wire \MAC.a[6] ;
 wire \MAC.a[7] ;
 wire \MAC.a[8] ;
 wire \MAC.a[9] ;
 wire \MAC.add.a1[0] ;
 wire \MAC.add.a1[10] ;
 wire \MAC.add.a1[11] ;
 wire \MAC.add.a1[12] ;
 wire \MAC.add.a1[13] ;
 wire \MAC.add.a1[14] ;
 wire \MAC.add.a1[15] ;
 wire \MAC.add.a1[1] ;
 wire \MAC.add.a1[2] ;
 wire \MAC.add.a1[3] ;
 wire \MAC.add.a1[4] ;
 wire \MAC.add.a1[5] ;
 wire \MAC.add.a1[6] ;
 wire \MAC.add.a1[7] ;
 wire \MAC.add.a1[8] ;
 wire \MAC.add.a1[9] ;
 wire \MAC.add.b1[0] ;
 wire \MAC.add.b1[10] ;
 wire \MAC.add.b1[11] ;
 wire \MAC.add.b1[12] ;
 wire \MAC.add.b1[13] ;
 wire \MAC.add.b1[14] ;
 wire \MAC.add.b1[15] ;
 wire \MAC.add.b1[1] ;
 wire \MAC.add.b1[2] ;
 wire \MAC.add.b1[3] ;
 wire \MAC.add.b1[4] ;
 wire \MAC.add.b1[5] ;
 wire \MAC.add.b1[6] ;
 wire \MAC.add.b1[7] ;
 wire \MAC.add.b1[8] ;
 wire \MAC.add.b1[9] ;
 wire \MAC.add.c_add[0] ;
 wire \MAC.add.c_add[10] ;
 wire \MAC.add.c_add[11] ;
 wire \MAC.add.c_add[12] ;
 wire \MAC.add.c_add[13] ;
 wire \MAC.add.c_add[14] ;
 wire \MAC.add.c_add[15] ;
 wire \MAC.add.c_add[1] ;
 wire \MAC.add.c_add[2] ;
 wire \MAC.add.c_add[3] ;
 wire \MAC.add.c_add[4] ;
 wire \MAC.add.c_add[5] ;
 wire \MAC.add.c_add[6] ;
 wire \MAC.add.c_add[7] ;
 wire \MAC.add.c_add[8] ;
 wire \MAC.add.c_add[9] ;
 wire \MAC.b[0] ;
 wire \MAC.b[10] ;
 wire \MAC.b[11] ;
 wire \MAC.b[12] ;
 wire \MAC.b[13] ;
 wire \MAC.b[14] ;
 wire \MAC.b[15] ;
 wire \MAC.b[1] ;
 wire \MAC.b[2] ;
 wire \MAC.b[3] ;
 wire \MAC.b[4] ;
 wire \MAC.b[5] ;
 wire \MAC.b[6] ;
 wire \MAC.b[7] ;
 wire \MAC.b[8] ;
 wire \MAC.b[9] ;
 wire \MAC.mul.c_mul1[0] ;
 wire \MAC.mul.c_mul1[10] ;
 wire \MAC.mul.c_mul1[11] ;
 wire \MAC.mul.c_mul1[12] ;
 wire \MAC.mul.c_mul1[13] ;
 wire \MAC.mul.c_mul1[14] ;
 wire \MAC.mul.c_mul1[15] ;
 wire \MAC.mul.c_mul1[1] ;
 wire \MAC.mul.c_mul1[2] ;
 wire \MAC.mul.c_mul1[3] ;
 wire \MAC.mul.c_mul1[4] ;
 wire \MAC.mul.c_mul1[5] ;
 wire \MAC.mul.c_mul1[6] ;
 wire \MAC.mul.c_mul1[7] ;
 wire \MAC.mul.c_mul1[8] ;
 wire \MAC.mul.c_mul1[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire clknet_0_clk;
 wire \wrap.state[0] ;
 wire \wrap.temp_data[0] ;
 wire \wrap.temp_data[10] ;
 wire \wrap.temp_data[11] ;
 wire \wrap.temp_data[12] ;
 wire \wrap.temp_data[13] ;
 wire \wrap.temp_data[14] ;
 wire \wrap.temp_data[15] ;
 wire \wrap.temp_data[1] ;
 wire \wrap.temp_data[2] ;
 wire \wrap.temp_data[3] ;
 wire \wrap.temp_data[4] ;
 wire \wrap.temp_data[5] ;
 wire \wrap.temp_data[6] ;
 wire \wrap.temp_data[7] ;
 wire \wrap.temp_data[8] ;
 wire \wrap.temp_data[9] ;
 wire \wrap2.state[0] ;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;

 sg13g2_inv_1 _1271_ (.Y(_0458_),
    .A(\MAC.add.a1[12] ));
 sg13g2_inv_1 _1272_ (.Y(_0459_),
    .A(\MAC.add.a1[11] ));
 sg13g2_inv_1 _1273_ (.Y(_0460_),
    .A(_0046_));
 sg13g2_inv_1 _1274_ (.Y(_0461_),
    .A(\MAC.add.a1[2] ));
 sg13g2_inv_1 _1275_ (.Y(_0462_),
    .A(_0048_));
 sg13g2_inv_1 _1276_ (.Y(_0463_),
    .A(\MAC.add.b1[3] ));
 sg13g2_inv_1 _1277_ (.Y(_0464_),
    .A(_0052_));
 sg13g2_inv_1 _1278_ (.Y(_0465_),
    .A(_0054_));
 sg13g2_inv_1 _1279_ (.Y(_0466_),
    .A(net66));
 sg13g2_inv_1 _1280_ (.Y(_0467_),
    .A(_0056_));
 sg13g2_inv_1 _1281_ (.Y(_0468_),
    .A(\MAC.add.b1[7] ));
 sg13g2_inv_1 _1282_ (.Y(_0469_),
    .A(\MAC.add.a1[7] ));
 sg13g2_inv_2 _1283_ (.Y(_0470_),
    .A(_0058_));
 sg13g2_inv_1 _1284_ (.Y(_0471_),
    .A(\MAC.add.b1[8] ));
 sg13g2_inv_1 _1285_ (.Y(_0472_),
    .A(_0060_));
 sg13g2_inv_1 _1286_ (.Y(_0473_),
    .A(net389));
 sg13g2_inv_2 _1287_ (.Y(_0474_),
    .A(net386));
 sg13g2_inv_1 _1288_ (.Y(_0475_),
    .A(net374));
 sg13g2_inv_1 _1289_ (.Y(_0476_),
    .A(net369));
 sg13g2_and2_1 _1290_ (.A(net43),
    .B(net353),
    .X(_0002_));
 sg13g2_and2_1 _1291_ (.A(net352),
    .B(net53),
    .X(_0009_));
 sg13g2_and2_1 _1292_ (.A(net353),
    .B(net35),
    .X(_0010_));
 sg13g2_and2_1 _1293_ (.A(net353),
    .B(net54),
    .X(_0011_));
 sg13g2_and2_1 _1294_ (.A(net353),
    .B(net37),
    .X(_0012_));
 sg13g2_and2_1 _1295_ (.A(net350),
    .B(net40),
    .X(_0013_));
 sg13g2_and2_1 _1296_ (.A(net350),
    .B(net52),
    .X(_0014_));
 sg13g2_and2_1 _1297_ (.A(net351),
    .B(net49),
    .X(_0015_));
 sg13g2_and2_1 _1298_ (.A(net350),
    .B(net51),
    .X(_0016_));
 sg13g2_and2_1 _1299_ (.A(net349),
    .B(net56),
    .X(_0017_));
 sg13g2_and2_1 _1300_ (.A(net349),
    .B(net46),
    .X(_0003_));
 sg13g2_and2_1 _1301_ (.A(net347),
    .B(net42),
    .X(_0004_));
 sg13g2_and2_1 _1302_ (.A(net347),
    .B(net48),
    .X(_0005_));
 sg13g2_and2_1 _1303_ (.A(net347),
    .B(net44),
    .X(_0006_));
 sg13g2_and2_1 _1304_ (.A(net348),
    .B(net39),
    .X(_0007_));
 sg13g2_and2_1 _1305_ (.A(net348),
    .B(net45),
    .X(_0008_));
 sg13g2_and2_1 _1306_ (.A(net352),
    .B(net1),
    .X(_0018_));
 sg13g2_and2_1 _1307_ (.A(net352),
    .B(net2),
    .X(_0025_));
 sg13g2_and2_1 _1308_ (.A(net350),
    .B(net3),
    .X(_0026_));
 sg13g2_and2_1 _1309_ (.A(net353),
    .B(net4),
    .X(_0027_));
 sg13g2_and2_1 _1310_ (.A(net352),
    .B(net5),
    .X(_0028_));
 sg13g2_and2_1 _1311_ (.A(net350),
    .B(net6),
    .X(_0029_));
 sg13g2_and2_1 _1312_ (.A(net351),
    .B(net7),
    .X(_0030_));
 sg13g2_and2_1 _1313_ (.A(net351),
    .B(net8),
    .X(_0031_));
 sg13g2_and2_1 _1314_ (.A(net350),
    .B(net9),
    .X(_0032_));
 sg13g2_and2_1 _1315_ (.A(net349),
    .B(net10),
    .X(_0033_));
 sg13g2_and2_1 _1316_ (.A(net349),
    .B(net11),
    .X(_0019_));
 sg13g2_and2_1 _1317_ (.A(net347),
    .B(net12),
    .X(_0020_));
 sg13g2_and2_1 _1318_ (.A(net348),
    .B(net13),
    .X(_0021_));
 sg13g2_and2_1 _1319_ (.A(net348),
    .B(net14),
    .X(_0022_));
 sg13g2_and2_1 _1320_ (.A(net348),
    .B(net15),
    .X(_0023_));
 sg13g2_and2_1 _1321_ (.A(net348),
    .B(net16),
    .X(_0024_));
 sg13g2_nor4_1 _1322_ (.A(\MAC.add.b1[7] ),
    .B(\MAC.add.a1[7] ),
    .C(\MAC.add.b1[8] ),
    .D(\MAC.add.a1[8] ),
    .Y(_0477_));
 sg13g2_nor4_1 _1323_ (.A(\MAC.add.b1[5] ),
    .B(\MAC.add.a1[5] ),
    .C(\MAC.add.b1[6] ),
    .D(\MAC.add.a1[6] ),
    .Y(_0478_));
 sg13g2_nor4_1 _1324_ (.A(\MAC.add.b1[3] ),
    .B(\MAC.add.a1[3] ),
    .C(\MAC.add.b1[4] ),
    .D(\MAC.add.a1[4] ),
    .Y(_0479_));
 sg13g2_nand3_1 _1325_ (.B(_0478_),
    .C(_0479_),
    .A(_0477_),
    .Y(_0480_));
 sg13g2_nor2_1 _1326_ (.A(\MAC.add.b1[12] ),
    .B(\MAC.add.b1[11] ),
    .Y(_0481_));
 sg13g2_nor4_1 _1327_ (.A(\MAC.add.b1[10] ),
    .B(\MAC.add.b1[9] ),
    .C(\MAC.add.b1[14] ),
    .D(\MAC.add.b1[13] ),
    .Y(_0482_));
 sg13g2_nand2_2 _1328_ (.Y(_0483_),
    .A(_0481_),
    .B(_0482_));
 sg13g2_nor4_1 _1329_ (.A(\MAC.add.a1[10] ),
    .B(\MAC.add.a1[9] ),
    .C(\MAC.add.a1[14] ),
    .D(\MAC.add.a1[13] ),
    .Y(_0484_));
 sg13g2_nand3_1 _1330_ (.B(_0459_),
    .C(_0484_),
    .A(_0458_),
    .Y(_0485_));
 sg13g2_nor4_1 _1331_ (.A(\MAC.add.a1[15] ),
    .B(\MAC.add.b1[15] ),
    .C(\MAC.add.b1[0] ),
    .D(\MAC.add.a1[0] ),
    .Y(_0486_));
 sg13g2_nor3_1 _1332_ (.A(\MAC.add.b1[1] ),
    .B(\MAC.add.a1[1] ),
    .C(\MAC.add.b1[2] ),
    .Y(_0487_));
 sg13g2_nand3_1 _1333_ (.B(_0486_),
    .C(_0487_),
    .A(_0461_),
    .Y(_0488_));
 sg13g2_nor4_2 _1334_ (.A(_0480_),
    .B(_0483_),
    .C(_0485_),
    .Y(_0489_),
    .D(_0488_));
 sg13g2_xor2_1 _1335_ (.B(\MAC.add.b1[15] ),
    .A(\MAC.add.a1[15] ),
    .X(_0490_));
 sg13g2_xnor2_1 _1336_ (.Y(_0491_),
    .A(\MAC.add.a1[15] ),
    .B(\MAC.add.b1[15] ));
 sg13g2_nand2b_1 _1337_ (.Y(_0492_),
    .B(\MAC.add.b1[14] ),
    .A_N(\MAC.add.a1[14] ));
 sg13g2_nand2b_1 _1338_ (.Y(_0493_),
    .B(\MAC.add.a1[14] ),
    .A_N(\MAC.add.b1[14] ));
 sg13g2_nand2b_1 _1339_ (.Y(_0494_),
    .B(\MAC.add.a1[13] ),
    .A_N(\MAC.add.b1[13] ));
 sg13g2_nand2b_1 _1340_ (.Y(_0495_),
    .B(\MAC.add.b1[13] ),
    .A_N(\MAC.add.a1[13] ));
 sg13g2_nand2b_1 _1341_ (.Y(_0496_),
    .B(\MAC.add.a1[12] ),
    .A_N(\MAC.add.b1[12] ));
 sg13g2_nor2b_1 _1342_ (.A(\MAC.add.a1[11] ),
    .B_N(\MAC.add.b1[11] ),
    .Y(_0497_));
 sg13g2_nand2b_1 _1343_ (.Y(_0498_),
    .B(\MAC.add.a1[11] ),
    .A_N(\MAC.add.b1[11] ));
 sg13g2_nand2b_2 _1344_ (.Y(_0499_),
    .B(_0498_),
    .A_N(_0497_));
 sg13g2_nor2b_1 _1345_ (.A(\MAC.add.a1[10] ),
    .B_N(\MAC.add.b1[10] ),
    .Y(_0500_));
 sg13g2_nor2b_1 _1346_ (.A(\MAC.add.b1[10] ),
    .B_N(\MAC.add.a1[10] ),
    .Y(_0501_));
 sg13g2_nand2b_1 _1347_ (.Y(_0502_),
    .B(\MAC.add.a1[10] ),
    .A_N(\MAC.add.b1[10] ));
 sg13g2_nand2b_1 _1348_ (.Y(_0503_),
    .B(\MAC.add.a1[9] ),
    .A_N(\MAC.add.b1[9] ));
 sg13g2_o21ai_1 _1349_ (.B1(_0502_),
    .Y(_0504_),
    .A1(_0500_),
    .A2(_0503_));
 sg13g2_nor2_1 _1350_ (.A(_0499_),
    .B(_0504_),
    .Y(_0505_));
 sg13g2_a21oi_1 _1351_ (.A1(_0458_),
    .A2(\MAC.add.b1[12] ),
    .Y(_0506_),
    .B1(_0497_));
 sg13g2_o21ai_1 _1352_ (.B1(_0506_),
    .Y(_0507_),
    .A1(_0499_),
    .A2(_0504_));
 sg13g2_nand3_1 _1353_ (.B(_0496_),
    .C(_0507_),
    .A(_0494_),
    .Y(_0508_));
 sg13g2_nand3_1 _1354_ (.B(_0495_),
    .C(_0508_),
    .A(_0492_),
    .Y(_0509_));
 sg13g2_nand2_1 _1355_ (.Y(_0510_),
    .A(net344),
    .B(_0509_));
 sg13g2_and2_1 _1356_ (.A(net344),
    .B(_0509_),
    .X(_0511_));
 sg13g2_nand2_1 _1357_ (.Y(_0512_),
    .A(_0059_),
    .B(net334));
 sg13g2_o21ai_1 _1358_ (.B1(_0512_),
    .Y(_0513_),
    .A1(_0470_),
    .A2(net333));
 sg13g2_nor2_1 _1359_ (.A(_0472_),
    .B(net335),
    .Y(_0514_));
 sg13g2_a21oi_2 _1360_ (.B1(_0514_),
    .Y(_0515_),
    .A2(net334),
    .A1(_0061_));
 sg13g2_xnor2_1 _1361_ (.Y(_0516_),
    .A(\MAC.add.a1[12] ),
    .B(\MAC.add.b1[12] ));
 sg13g2_nor2_1 _1362_ (.A(_0497_),
    .B(_0505_),
    .Y(_0517_));
 sg13g2_nor2_1 _1363_ (.A(_0500_),
    .B(_0501_),
    .Y(_0518_));
 sg13g2_nor2b_1 _1364_ (.A(\MAC.add.a1[9] ),
    .B_N(\MAC.add.b1[9] ),
    .Y(_0519_));
 sg13g2_xor2_1 _1365_ (.B(\MAC.add.b1[9] ),
    .A(\MAC.add.a1[9] ),
    .X(_0520_));
 sg13g2_nor3_2 _1366_ (.A(_0500_),
    .B(_0501_),
    .C(_0520_),
    .Y(_0521_));
 sg13g2_nor2_1 _1367_ (.A(_0504_),
    .B(_0521_),
    .Y(_0522_));
 sg13g2_o21ai_1 _1368_ (.B1(_0498_),
    .Y(_0523_),
    .A1(_0499_),
    .A2(_0522_));
 sg13g2_and2_1 _1369_ (.A(_0483_),
    .B(_0485_),
    .X(_0524_));
 sg13g2_nand2_2 _1370_ (.Y(_0525_),
    .A(_0483_),
    .B(_0485_));
 sg13g2_xor2_1 _1371_ (.B(_0517_),
    .A(_0516_),
    .X(_0526_));
 sg13g2_and3_1 _1372_ (.X(_0527_),
    .A(net345),
    .B(net338),
    .C(_0526_));
 sg13g2_xor2_1 _1373_ (.B(_0523_),
    .A(_0516_),
    .X(_0528_));
 sg13g2_a21oi_1 _1374_ (.A1(net345),
    .A2(net338),
    .Y(_0529_),
    .B1(_0528_));
 sg13g2_nor3_2 _1375_ (.A(_0525_),
    .B(_0527_),
    .C(_0529_),
    .Y(_0530_));
 sg13g2_nand2_1 _1376_ (.Y(_0531_),
    .A(_0494_),
    .B(_0495_));
 sg13g2_inv_1 _1377_ (.Y(_0532_),
    .A(_0531_));
 sg13g2_nand3b_1 _1378_ (.B(_0516_),
    .C(_0521_),
    .Y(_0533_),
    .A_N(_0499_));
 sg13g2_nand3_1 _1379_ (.B(_0507_),
    .C(_0533_),
    .A(_0496_),
    .Y(_0534_));
 sg13g2_xnor2_1 _1380_ (.Y(_0535_),
    .A(_0532_),
    .B(_0534_));
 sg13g2_nand3_1 _1381_ (.B(net338),
    .C(_0533_),
    .A(net345),
    .Y(_0536_));
 sg13g2_or2_1 _1382_ (.X(_0537_),
    .B(_0536_),
    .A(_0535_));
 sg13g2_a21oi_2 _1383_ (.B1(_0525_),
    .Y(_0538_),
    .A2(_0536_),
    .A1(_0535_));
 sg13g2_nand2_1 _1384_ (.Y(_0539_),
    .A(_0537_),
    .B(_0538_));
 sg13g2_xnor2_1 _1385_ (.Y(_0540_),
    .A(_0499_),
    .B(_0522_));
 sg13g2_o21ai_1 _1386_ (.B1(_0540_),
    .Y(_0541_),
    .A1(net335),
    .A2(_0521_));
 sg13g2_or3_1 _1387_ (.A(net335),
    .B(_0521_),
    .C(_0540_),
    .X(_0542_));
 sg13g2_and3_2 _1388_ (.X(_0543_),
    .A(net341),
    .B(_0541_),
    .C(_0542_));
 sg13g2_nand3_1 _1389_ (.B(_0541_),
    .C(_0542_),
    .A(net341),
    .Y(_0544_));
 sg13g2_a21oi_2 _1390_ (.B1(_0530_),
    .Y(_0545_),
    .A2(_0538_),
    .A1(_0537_));
 sg13g2_a21o_2 _1391_ (.A2(_0538_),
    .A1(_0537_),
    .B1(_0530_),
    .X(_0546_));
 sg13g2_xnor2_1 _1392_ (.Y(_0547_),
    .A(_0518_),
    .B(_0519_));
 sg13g2_nand4_1 _1393_ (.B(net338),
    .C(_0520_),
    .A(net343),
    .Y(_0548_),
    .D(_0547_));
 sg13g2_a21o_1 _1394_ (.A2(_0520_),
    .A1(net331),
    .B1(_0547_),
    .X(_0549_));
 sg13g2_and2_1 _1395_ (.A(net341),
    .B(_0548_),
    .X(_0550_));
 sg13g2_and2_2 _1396_ (.A(net330),
    .B(net329),
    .X(_0551_));
 sg13g2_nand2_2 _1397_ (.Y(_0552_),
    .A(net330),
    .B(net329));
 sg13g2_a22oi_1 _1398_ (.Y(_0553_),
    .B1(_0532_),
    .B2(_0534_),
    .A2(_0508_),
    .A1(_0495_));
 sg13g2_a21o_1 _1399_ (.A2(_0508_),
    .A1(_0495_),
    .B1(_0492_),
    .X(_0554_));
 sg13g2_or2_2 _1400_ (.X(_0555_),
    .B(\MAC.add.b1[14] ),
    .A(\MAC.add.a1[14] ));
 sg13g2_nand2_1 _1401_ (.Y(_0556_),
    .A(_0492_),
    .B(net345));
 sg13g2_o21ai_1 _1402_ (.B1(_0554_),
    .Y(_0557_),
    .A1(net345),
    .A2(_0553_));
 sg13g2_nand2_2 _1403_ (.Y(_0558_),
    .A(_0520_),
    .B(net341));
 sg13g2_inv_1 _1404_ (.Y(_0559_),
    .A(_0558_));
 sg13g2_a21o_1 _1405_ (.A2(_0557_),
    .A1(net341),
    .B1(_0559_),
    .X(_0560_));
 sg13g2_a21oi_2 _1406_ (.B1(_0560_),
    .Y(_0561_),
    .A2(net329),
    .A1(net330));
 sg13g2_nand3_1 _1407_ (.B(net324),
    .C(_0561_),
    .A(_0539_),
    .Y(_0562_));
 sg13g2_nand3_1 _1408_ (.B(_0545_),
    .C(_0561_),
    .A(net323),
    .Y(_0563_));
 sg13g2_nor2_1 _1409_ (.A(_0515_),
    .B(_0563_),
    .Y(_0564_));
 sg13g2_nor2_2 _1410_ (.A(_0557_),
    .B(_0558_),
    .Y(_0565_));
 sg13g2_nand2b_1 _1411_ (.Y(_0566_),
    .B(_0559_),
    .A_N(_0557_));
 sg13g2_a21oi_1 _1412_ (.A1(net344),
    .A2(net338),
    .Y(_0567_),
    .B1(_0472_));
 sg13g2_and3_1 _1413_ (.X(_0568_),
    .A(_0061_),
    .B(net344),
    .C(net337));
 sg13g2_or4_1 _1414_ (.A(_0525_),
    .B(_0557_),
    .C(_0567_),
    .D(_0568_),
    .X(_0569_));
 sg13g2_a22oi_1 _1415_ (.Y(_0570_),
    .B1(_0566_),
    .B2(_0569_),
    .A2(_0550_),
    .A1(_0549_));
 sg13g2_nand3_1 _1416_ (.B(net323),
    .C(_0570_),
    .A(_0539_),
    .Y(_0571_));
 sg13g2_nand3_1 _1417_ (.B(_0545_),
    .C(_0570_),
    .A(net323),
    .Y(_0572_));
 sg13g2_a21o_2 _1418_ (.A2(_0572_),
    .A1(_0515_),
    .B1(_0563_),
    .X(_0573_));
 sg13g2_a21oi_2 _1419_ (.B1(_0563_),
    .Y(_0574_),
    .A2(_0572_),
    .A1(_0515_));
 sg13g2_and2_1 _1420_ (.A(_0546_),
    .B(_0562_),
    .X(_0575_));
 sg13g2_nor3_1 _1421_ (.A(_0520_),
    .B(_0525_),
    .C(_0557_),
    .Y(_0576_));
 sg13g2_a21oi_1 _1422_ (.A1(net343),
    .A2(net337),
    .Y(_0577_),
    .B1(_0470_));
 sg13g2_and3_1 _1423_ (.X(_0578_),
    .A(_0059_),
    .B(net343),
    .C(net337));
 sg13g2_nor2_1 _1424_ (.A(_0577_),
    .B(_0578_),
    .Y(_0579_));
 sg13g2_nor4_1 _1425_ (.A(_0557_),
    .B(_0558_),
    .C(_0567_),
    .D(_0568_),
    .Y(_0580_));
 sg13g2_a21oi_1 _1426_ (.A1(net327),
    .A2(_0579_),
    .Y(_0581_),
    .B1(_0580_));
 sg13g2_a21oi_1 _1427_ (.A1(net343),
    .A2(net337),
    .Y(_0582_),
    .B1(_0465_));
 sg13g2_a21oi_2 _1428_ (.B1(_0582_),
    .Y(_0583_),
    .A2(net331),
    .A1(_0055_));
 sg13g2_a21oi_1 _1429_ (.A1(net343),
    .A2(net337),
    .Y(_0584_),
    .B1(_0467_));
 sg13g2_and3_1 _1430_ (.X(_0585_),
    .A(_0057_),
    .B(net343),
    .C(net337));
 sg13g2_nor2_1 _1431_ (.A(_0584_),
    .B(_0585_),
    .Y(_0586_));
 sg13g2_nor4_1 _1432_ (.A(_0557_),
    .B(_0558_),
    .C(_0584_),
    .D(_0585_),
    .Y(_0587_));
 sg13g2_a21oi_1 _1433_ (.A1(net327),
    .A2(_0583_),
    .Y(_0588_),
    .B1(_0587_));
 sg13g2_a221oi_1 _1434_ (.B2(_0583_),
    .C1(_0587_),
    .B1(net327),
    .A1(net330),
    .Y(_0589_),
    .A2(net329));
 sg13g2_a21oi_1 _1435_ (.A1(_0551_),
    .A2(_0581_),
    .Y(_0590_),
    .B1(_0589_));
 sg13g2_a21o_1 _1436_ (.A2(_0581_),
    .A1(_0551_),
    .B1(_0589_),
    .X(_0591_));
 sg13g2_nand3b_1 _1437_ (.B(net343),
    .C(net337),
    .Y(_0592_),
    .A_N(_0051_));
 sg13g2_o21ai_1 _1438_ (.B1(_0592_),
    .Y(_0593_),
    .A1(_0050_),
    .A2(net331));
 sg13g2_a21oi_1 _1439_ (.A1(net343),
    .A2(net337),
    .Y(_0594_),
    .B1(_0464_));
 sg13g2_a21oi_1 _1440_ (.A1(_0053_),
    .A2(net331),
    .Y(_0595_),
    .B1(_0594_));
 sg13g2_a22oi_1 _1441_ (.Y(_0596_),
    .B1(_0595_),
    .B2(_0565_),
    .A2(_0593_),
    .A1(net327));
 sg13g2_nand2_1 _1442_ (.Y(_0597_),
    .A(_0551_),
    .B(_0596_));
 sg13g2_a21oi_1 _1443_ (.A1(net344),
    .A2(net338),
    .Y(_0598_),
    .B1(_0462_));
 sg13g2_a21oi_1 _1444_ (.A1(_0049_),
    .A2(net331),
    .Y(_0599_),
    .B1(_0598_));
 sg13g2_a21oi_1 _1445_ (.A1(net344),
    .A2(net338),
    .Y(_0600_),
    .B1(_0460_));
 sg13g2_a21oi_1 _1446_ (.A1(_0047_),
    .A2(net331),
    .Y(_0601_),
    .B1(_0600_));
 sg13g2_a22oi_1 _1447_ (.Y(_0602_),
    .B1(_0601_),
    .B2(net328),
    .A2(_0599_),
    .A1(_0565_));
 sg13g2_a21oi_1 _1448_ (.A1(_0552_),
    .A2(_0602_),
    .Y(_0603_),
    .B1(_0543_));
 sg13g2_a221oi_1 _1449_ (.B2(_0603_),
    .C1(_0530_),
    .B1(_0597_),
    .A1(_0543_),
    .Y(_0604_),
    .A2(_0590_));
 sg13g2_or2_1 _1450_ (.X(_0605_),
    .B(_0604_),
    .A(_0575_));
 sg13g2_nor2_1 _1451_ (.A(_0460_),
    .B(net334),
    .Y(_0606_));
 sg13g2_a21oi_2 _1452_ (.B1(_0606_),
    .Y(_0607_),
    .A2(net333),
    .A1(_0047_));
 sg13g2_nor3_1 _1453_ (.A(_0575_),
    .B(_0604_),
    .C(_0607_),
    .Y(_0608_));
 sg13g2_a22oi_1 _1454_ (.Y(_0609_),
    .B1(_0595_),
    .B2(net327),
    .A2(_0583_),
    .A1(_0565_));
 sg13g2_nor4_1 _1455_ (.A(_0557_),
    .B(_0558_),
    .C(_0577_),
    .D(_0578_),
    .Y(_0610_));
 sg13g2_a21oi_1 _1456_ (.A1(net327),
    .A2(_0586_),
    .Y(_0611_),
    .B1(_0610_));
 sg13g2_mux2_1 _1457_ (.A0(_0609_),
    .A1(_0611_),
    .S(_0551_),
    .X(_0612_));
 sg13g2_or2_1 _1458_ (.X(_0613_),
    .B(_0612_),
    .A(net324));
 sg13g2_a22oi_1 _1459_ (.Y(_0614_),
    .B1(_0599_),
    .B2(net328),
    .A2(_0593_),
    .A1(_0565_));
 sg13g2_nand2_1 _1460_ (.Y(_0615_),
    .A(_0565_),
    .B(_0601_));
 sg13g2_nor2_1 _1461_ (.A(_0045_),
    .B(net335),
    .Y(_0616_));
 sg13g2_nor2_1 _1462_ (.A(_0044_),
    .B(net332),
    .Y(_0617_));
 sg13g2_o21ai_1 _1463_ (.B1(net328),
    .Y(_0618_),
    .A1(_0616_),
    .A2(_0617_));
 sg13g2_nand3_1 _1464_ (.B(_0615_),
    .C(_0618_),
    .A(_0552_),
    .Y(_0619_));
 sg13g2_a21oi_1 _1465_ (.A1(_0551_),
    .A2(_0614_),
    .Y(_0620_),
    .B1(_0543_));
 sg13g2_a21oi_1 _1466_ (.A1(_0619_),
    .A2(_0620_),
    .Y(_0621_),
    .B1(_0530_));
 sg13g2_a22oi_1 _1467_ (.Y(_0622_),
    .B1(_0613_),
    .B2(_0621_),
    .A2(_0571_),
    .A1(_0546_));
 sg13g2_inv_1 _1468_ (.Y(_0623_),
    .A(_0622_));
 sg13g2_mux2_2 _1469_ (.A0(_0045_),
    .A1(_0044_),
    .S(net331),
    .X(_0624_));
 sg13g2_or3_1 _1470_ (.A(_0608_),
    .B(_0622_),
    .C(_0624_),
    .X(_0625_));
 sg13g2_a21o_1 _1471_ (.A2(_0609_),
    .A1(_0551_),
    .B1(_0543_),
    .X(_0626_));
 sg13g2_a21oi_1 _1472_ (.A1(_0552_),
    .A2(_0614_),
    .Y(_0627_),
    .B1(_0626_));
 sg13g2_a221oi_1 _1473_ (.B2(_0586_),
    .C1(_0610_),
    .B1(net327),
    .A1(net330),
    .Y(_0628_),
    .A2(net329));
 sg13g2_and4_1 _1474_ (.A(net330),
    .B(net329),
    .C(_0566_),
    .D(_0569_),
    .X(_0629_));
 sg13g2_nor3_1 _1475_ (.A(net323),
    .B(_0628_),
    .C(_0629_),
    .Y(_0630_));
 sg13g2_o21ai_1 _1476_ (.B1(_0545_),
    .Y(_0631_),
    .A1(_0627_),
    .A2(_0630_));
 sg13g2_nor2_1 _1477_ (.A(_0462_),
    .B(net334),
    .Y(_0632_));
 sg13g2_a21oi_2 _1478_ (.B1(_0632_),
    .Y(_0633_),
    .A2(net333),
    .A1(_0049_));
 sg13g2_a22oi_1 _1479_ (.Y(_0634_),
    .B1(_0631_),
    .B2(_0633_),
    .A2(_0607_),
    .A1(_0605_));
 sg13g2_a221oi_1 _1480_ (.B2(_0579_),
    .C1(_0580_),
    .B1(net327),
    .A1(net330),
    .Y(_0635_),
    .A2(net329));
 sg13g2_and3_1 _1481_ (.X(_0636_),
    .A(net330),
    .B(net329),
    .C(_0560_));
 sg13g2_mux4_1 _1482_ (.S0(_0552_),
    .A0(_0560_),
    .A1(_0581_),
    .A2(_0588_),
    .A3(_0596_),
    .S1(net324),
    .X(_0637_));
 sg13g2_nand2b_2 _1483_ (.Y(_0638_),
    .B(_0545_),
    .A_N(_0637_));
 sg13g2_mux2_2 _1484_ (.A0(_0051_),
    .A1(_0050_),
    .S(net331),
    .X(_0639_));
 sg13g2_nand2b_1 _1485_ (.Y(_0640_),
    .B(_0639_),
    .A_N(_0638_));
 sg13g2_o21ai_1 _1486_ (.B1(_0640_),
    .Y(_0641_),
    .A1(_0631_),
    .A2(_0633_));
 sg13g2_a21o_1 _1487_ (.A2(_0634_),
    .A1(_0625_),
    .B1(_0641_),
    .X(_0642_));
 sg13g2_nor4_2 _1488_ (.A(_0543_),
    .B(_0546_),
    .C(_0635_),
    .Y(_0643_),
    .D(_0636_));
 sg13g2_nor4_2 _1489_ (.A(_0543_),
    .B(_0546_),
    .C(_0628_),
    .Y(_0644_),
    .D(_0629_));
 sg13g2_nand2_1 _1490_ (.Y(_0645_),
    .A(_0057_),
    .B(net334));
 sg13g2_o21ai_1 _1491_ (.B1(_0645_),
    .Y(_0646_),
    .A1(_0467_),
    .A2(net333));
 sg13g2_a22oi_1 _1492_ (.Y(_0647_),
    .B1(_0644_),
    .B2(_0646_),
    .A2(_0643_),
    .A1(_0513_));
 sg13g2_o21ai_1 _1493_ (.B1(_0545_),
    .Y(_0648_),
    .A1(net323),
    .A2(_0561_));
 sg13g2_a21oi_2 _1494_ (.B1(_0648_),
    .Y(_0649_),
    .A2(_0591_),
    .A1(net323));
 sg13g2_nand2_1 _1495_ (.Y(_0650_),
    .A(_0055_),
    .B(net333));
 sg13g2_o21ai_1 _1496_ (.B1(_0650_),
    .Y(_0651_),
    .A1(_0465_),
    .A2(net333));
 sg13g2_nor2_1 _1497_ (.A(_0649_),
    .B(_0651_),
    .Y(_0652_));
 sg13g2_or2_1 _1498_ (.X(_0653_),
    .B(_0643_),
    .A(_0513_));
 sg13g2_or2_1 _1499_ (.X(_0654_),
    .B(_0646_),
    .A(_0644_));
 sg13g2_nand3_1 _1500_ (.B(_0653_),
    .C(_0654_),
    .A(_0647_),
    .Y(_0655_));
 sg13g2_nand2b_1 _1501_ (.Y(_0656_),
    .B(_0638_),
    .A_N(_0639_));
 sg13g2_o21ai_1 _1502_ (.B1(_0545_),
    .Y(_0657_),
    .A1(net323),
    .A2(_0570_));
 sg13g2_a21oi_2 _1503_ (.B1(_0657_),
    .Y(_0658_),
    .A2(_0612_),
    .A1(net323));
 sg13g2_inv_1 _1504_ (.Y(_0659_),
    .A(_0658_));
 sg13g2_nand2_1 _1505_ (.Y(_0660_),
    .A(_0053_),
    .B(net333));
 sg13g2_o21ai_1 _1506_ (.B1(_0660_),
    .Y(_0661_),
    .A1(_0464_),
    .A2(net333));
 sg13g2_inv_1 _1507_ (.Y(_0662_),
    .A(_0661_));
 sg13g2_nor2_1 _1508_ (.A(_0658_),
    .B(_0661_),
    .Y(_0663_));
 sg13g2_a22oi_1 _1509_ (.Y(_0664_),
    .B1(_0658_),
    .B2(_0661_),
    .A2(_0651_),
    .A1(_0649_));
 sg13g2_nand2_1 _1510_ (.Y(_0665_),
    .A(_0656_),
    .B(_0664_));
 sg13g2_nor4_2 _1511_ (.A(_0652_),
    .B(_0655_),
    .C(_0663_),
    .Y(_0666_),
    .D(_0665_));
 sg13g2_nor3_1 _1512_ (.A(_0652_),
    .B(_0655_),
    .C(_0664_),
    .Y(_0667_));
 sg13g2_nor3_1 _1513_ (.A(_0515_),
    .B(_0562_),
    .C(_0572_),
    .Y(_0668_));
 sg13g2_nor2b_1 _1514_ (.A(_0647_),
    .B_N(_0653_),
    .Y(_0669_));
 sg13g2_or3_1 _1515_ (.A(_0667_),
    .B(_0668_),
    .C(_0669_),
    .X(_0670_));
 sg13g2_a21oi_2 _1516_ (.B1(_0670_),
    .Y(_0671_),
    .A2(_0666_),
    .A1(_0642_));
 sg13g2_a21o_2 _1517_ (.A2(_0666_),
    .A1(_0642_),
    .B1(_0670_),
    .X(_0672_));
 sg13g2_nor2_1 _1518_ (.A(_0573_),
    .B(_0671_),
    .Y(_0673_));
 sg13g2_nand2_2 _1519_ (.Y(_0674_),
    .A(_0574_),
    .B(_0672_));
 sg13g2_nor2_1 _1520_ (.A(_0643_),
    .B(net320),
    .Y(_0675_));
 sg13g2_a21oi_2 _1521_ (.B1(_0675_),
    .Y(_0676_),
    .A2(net319),
    .A1(_0513_));
 sg13g2_nor2_1 _1522_ (.A(_0644_),
    .B(net320),
    .Y(_0677_));
 sg13g2_a21oi_2 _1523_ (.B1(_0677_),
    .Y(_0678_),
    .A2(net319),
    .A1(_0646_));
 sg13g2_a21o_1 _1524_ (.A2(_0672_),
    .A1(_0574_),
    .B1(_0649_),
    .X(_0679_));
 sg13g2_nand3_1 _1525_ (.B(_0651_),
    .C(_0672_),
    .A(_0574_),
    .Y(_0680_));
 sg13g2_nand2_1 _1526_ (.Y(_0681_),
    .A(_0679_),
    .B(_0680_));
 sg13g2_a21oi_1 _1527_ (.A1(_0574_),
    .A2(_0672_),
    .Y(_0682_),
    .B1(_0659_));
 sg13g2_a21oi_2 _1528_ (.B1(_0682_),
    .Y(_0683_),
    .A2(net319),
    .A1(_0662_));
 sg13g2_nor3_2 _1529_ (.A(_0573_),
    .B(_0639_),
    .C(_0671_),
    .Y(_0684_));
 sg13g2_a21oi_1 _1530_ (.A1(_0574_),
    .A2(_0672_),
    .Y(_0685_),
    .B1(_0638_));
 sg13g2_nor2_2 _1531_ (.A(_0684_),
    .B(_0685_),
    .Y(_0686_));
 sg13g2_o21ai_1 _1532_ (.B1(net346),
    .Y(_0687_),
    .A1(_0684_),
    .A2(_0685_));
 sg13g2_or3_1 _1533_ (.A(_0573_),
    .B(_0633_),
    .C(_0671_),
    .X(_0688_));
 sg13g2_o21ai_1 _1534_ (.B1(_0631_),
    .Y(_0689_),
    .A1(_0573_),
    .A2(_0671_));
 sg13g2_nand2_2 _1535_ (.Y(_0690_),
    .A(_0688_),
    .B(_0689_));
 sg13g2_nand3_1 _1536_ (.B(_0688_),
    .C(_0689_),
    .A(net346),
    .Y(_0691_));
 sg13g2_nand3_1 _1537_ (.B(_0624_),
    .C(_0672_),
    .A(_0574_),
    .Y(_0692_));
 sg13g2_o21ai_1 _1538_ (.B1(_0623_),
    .Y(_0693_),
    .A1(_0573_),
    .A2(_0671_));
 sg13g2_nand3_1 _1539_ (.B(_0692_),
    .C(_0693_),
    .A(net346),
    .Y(_0694_));
 sg13g2_a21oi_1 _1540_ (.A1(_0574_),
    .A2(_0672_),
    .Y(_0695_),
    .B1(_0605_));
 sg13g2_and3_1 _1541_ (.X(_0696_),
    .A(_0574_),
    .B(_0607_),
    .C(_0672_));
 sg13g2_nor2_1 _1542_ (.A(_0695_),
    .B(_0696_),
    .Y(_0697_));
 sg13g2_o21ai_1 _1543_ (.B1(net346),
    .Y(_0698_),
    .A1(_0695_),
    .A2(_0696_));
 sg13g2_a221oi_1 _1544_ (.B2(_0693_),
    .C1(_0695_),
    .B1(_0692_),
    .A1(_0607_),
    .Y(_0699_),
    .A2(net320));
 sg13g2_nor2_1 _1545_ (.A(_0491_),
    .B(_0699_),
    .Y(_0700_));
 sg13g2_a21oi_1 _1546_ (.A1(_0690_),
    .A2(_0699_),
    .Y(_0701_),
    .B1(_0491_));
 sg13g2_nand4_1 _1547_ (.B(_0691_),
    .C(_0694_),
    .A(_0687_),
    .Y(_0702_),
    .D(_0698_));
 sg13g2_nand4_1 _1548_ (.B(_0686_),
    .C(_0690_),
    .A(_0683_),
    .Y(_0703_),
    .D(_0699_));
 sg13g2_a221oi_1 _1549_ (.B2(_0680_),
    .C1(_0682_),
    .B1(_0679_),
    .A1(_0662_),
    .Y(_0704_),
    .A2(net319));
 sg13g2_nand4_1 _1550_ (.B(_0690_),
    .C(_0699_),
    .A(_0686_),
    .Y(_0705_),
    .D(_0704_));
 sg13g2_nand2_1 _1551_ (.Y(_0706_),
    .A(net346),
    .B(_0705_));
 sg13g2_o21ai_1 _1552_ (.B1(net346),
    .Y(_0707_),
    .A1(_0678_),
    .A2(_0705_));
 sg13g2_nor3_2 _1553_ (.A(_0676_),
    .B(_0678_),
    .C(_0705_),
    .Y(_0708_));
 sg13g2_nor2_1 _1554_ (.A(_0491_),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_nand3_1 _1555_ (.B(_0572_),
    .C(_0708_),
    .A(_0563_),
    .Y(_0710_));
 sg13g2_and2_1 _1556_ (.A(_0490_),
    .B(_0710_),
    .X(_0711_));
 sg13g2_nor2_1 _1557_ (.A(_0572_),
    .B(_0674_),
    .Y(_0712_));
 sg13g2_a21oi_1 _1558_ (.A1(_0515_),
    .A2(_0674_),
    .Y(_0713_),
    .B1(_0712_));
 sg13g2_nor2_1 _1559_ (.A(_0564_),
    .B(_0572_),
    .Y(_0714_));
 sg13g2_xnor2_1 _1560_ (.Y(_0715_),
    .A(_0709_),
    .B(_0714_));
 sg13g2_nor2_1 _1561_ (.A(_0713_),
    .B(_0715_),
    .Y(_0716_));
 sg13g2_nand3_1 _1562_ (.B(_0681_),
    .C(_0703_),
    .A(net346),
    .Y(_0717_));
 sg13g2_a21o_1 _1563_ (.A2(_0703_),
    .A1(net346),
    .B1(_0681_),
    .X(_0718_));
 sg13g2_nor2_1 _1564_ (.A(_0651_),
    .B(net320),
    .Y(_0719_));
 sg13g2_a21oi_2 _1565_ (.B1(_0719_),
    .Y(_0720_),
    .A2(net319),
    .A1(_0649_));
 sg13g2_nand3_1 _1566_ (.B(_0718_),
    .C(_0720_),
    .A(_0717_),
    .Y(_0721_));
 sg13g2_a21oi_1 _1567_ (.A1(_0717_),
    .A2(_0718_),
    .Y(_0722_),
    .B1(_0720_));
 sg13g2_a21o_1 _1568_ (.A2(_0718_),
    .A1(_0717_),
    .B1(_0720_),
    .X(_0723_));
 sg13g2_and2_1 _1569_ (.A(_0721_),
    .B(_0723_),
    .X(_0724_));
 sg13g2_xnor2_1 _1570_ (.Y(_0725_),
    .A(_0686_),
    .B(_0701_));
 sg13g2_mux2_1 _1571_ (.A0(_0638_),
    .A1(_0639_),
    .S(_0674_),
    .X(_0726_));
 sg13g2_inv_1 _1572_ (.Y(_0727_),
    .A(_0726_));
 sg13g2_nor2_2 _1573_ (.A(_0725_),
    .B(_0727_),
    .Y(_0728_));
 sg13g2_xor2_1 _1574_ (.B(_0700_),
    .A(_0690_),
    .X(_0729_));
 sg13g2_nor2_1 _1575_ (.A(_0631_),
    .B(_0674_),
    .Y(_0730_));
 sg13g2_a21oi_2 _1576_ (.B1(_0730_),
    .Y(_0731_),
    .A2(_0674_),
    .A1(_0633_));
 sg13g2_nor2_1 _1577_ (.A(_0729_),
    .B(_0731_),
    .Y(_0732_));
 sg13g2_xor2_1 _1578_ (.B(_0697_),
    .A(_0694_),
    .X(_0733_));
 sg13g2_nor2_1 _1579_ (.A(_0607_),
    .B(net320),
    .Y(_0734_));
 sg13g2_a21oi_2 _1580_ (.B1(_0734_),
    .Y(_0735_),
    .A2(net320),
    .A1(_0605_));
 sg13g2_nand2_1 _1581_ (.Y(_0736_),
    .A(_0733_),
    .B(_0735_));
 sg13g2_nor2_1 _1582_ (.A(_0623_),
    .B(_0624_),
    .Y(_0737_));
 sg13g2_inv_1 _1583_ (.Y(_0738_),
    .A(_0737_));
 sg13g2_xnor2_1 _1584_ (.Y(_0739_),
    .A(_0733_),
    .B(_0735_));
 sg13g2_o21ai_1 _1585_ (.B1(_0736_),
    .Y(_0740_),
    .A1(_0738_),
    .A2(_0739_));
 sg13g2_xor2_1 _1586_ (.B(_0731_),
    .A(_0729_),
    .X(_0741_));
 sg13g2_a21o_1 _1587_ (.A2(_0741_),
    .A1(_0740_),
    .B1(_0732_),
    .X(_0742_));
 sg13g2_a221oi_1 _1588_ (.B2(_0741_),
    .C1(_0732_),
    .B1(_0740_),
    .A1(_0725_),
    .Y(_0743_),
    .A2(_0727_));
 sg13g2_xor2_1 _1589_ (.B(_0702_),
    .A(_0683_),
    .X(_0744_));
 sg13g2_nor2_1 _1590_ (.A(_0659_),
    .B(_0674_),
    .Y(_0745_));
 sg13g2_a21oi_2 _1591_ (.B1(_0745_),
    .Y(_0746_),
    .A2(_0674_),
    .A1(_0662_));
 sg13g2_nor2_1 _1592_ (.A(_0744_),
    .B(_0746_),
    .Y(_0747_));
 sg13g2_xnor2_1 _1593_ (.Y(_0748_),
    .A(_0744_),
    .B(_0746_));
 sg13g2_nor3_1 _1594_ (.A(_0728_),
    .B(_0743_),
    .C(_0748_),
    .Y(_0749_));
 sg13g2_or3_1 _1595_ (.A(_0728_),
    .B(_0743_),
    .C(_0748_),
    .X(_0750_));
 sg13g2_nand3b_1 _1596_ (.B(_0723_),
    .C(_0721_),
    .Y(_0751_),
    .A_N(_0748_));
 sg13g2_nor3_1 _1597_ (.A(_0728_),
    .B(_0743_),
    .C(_0751_),
    .Y(_0752_));
 sg13g2_or3_1 _1598_ (.A(_0728_),
    .B(_0743_),
    .C(_0751_),
    .X(_0753_));
 sg13g2_xnor2_1 _1599_ (.Y(_0754_),
    .A(_0676_),
    .B(_0707_));
 sg13g2_xor2_1 _1600_ (.B(_0707_),
    .A(_0676_),
    .X(_0755_));
 sg13g2_nor2_1 _1601_ (.A(_0513_),
    .B(net319),
    .Y(_0756_));
 sg13g2_nand2_1 _1602_ (.Y(_0757_),
    .A(_0643_),
    .B(net319));
 sg13g2_nor2b_1 _1603_ (.A(_0756_),
    .B_N(_0757_),
    .Y(_0758_));
 sg13g2_nand2b_1 _1604_ (.Y(_0759_),
    .B(_0757_),
    .A_N(_0756_));
 sg13g2_nor2_1 _1605_ (.A(_0754_),
    .B(_0759_),
    .Y(_0760_));
 sg13g2_xor2_1 _1606_ (.B(_0706_),
    .A(_0678_),
    .X(_0761_));
 sg13g2_xnor2_1 _1607_ (.Y(_0762_),
    .A(_0678_),
    .B(_0706_));
 sg13g2_nand2b_1 _1608_ (.Y(_0763_),
    .B(_0674_),
    .A_N(_0646_));
 sg13g2_nand2_1 _1609_ (.Y(_0764_),
    .A(_0644_),
    .B(net319));
 sg13g2_nand2_2 _1610_ (.Y(_0765_),
    .A(_0763_),
    .B(_0764_));
 sg13g2_nand2_2 _1611_ (.Y(_0766_),
    .A(_0762_),
    .B(_0765_));
 sg13g2_a221oi_1 _1612_ (.B2(_0764_),
    .C1(_0761_),
    .B1(_0763_),
    .A1(_0755_),
    .Y(_0767_),
    .A2(_0758_));
 sg13g2_and2_1 _1613_ (.A(_0721_),
    .B(_0747_),
    .X(_0768_));
 sg13g2_or2_1 _1614_ (.X(_0769_),
    .B(_0768_),
    .A(_0722_));
 sg13g2_nor2_1 _1615_ (.A(_0755_),
    .B(_0758_),
    .Y(_0770_));
 sg13g2_nand2_1 _1616_ (.Y(_0771_),
    .A(_0754_),
    .B(_0759_));
 sg13g2_nor4_1 _1617_ (.A(_0722_),
    .B(_0767_),
    .C(_0768_),
    .D(_0770_),
    .Y(_0772_));
 sg13g2_nor2_1 _1618_ (.A(_0762_),
    .B(_0765_),
    .Y(_0773_));
 sg13g2_a21o_1 _1619_ (.A2(_0773_),
    .A1(_0771_),
    .B1(_0760_),
    .X(_0774_));
 sg13g2_a21o_1 _1620_ (.A2(_0772_),
    .A1(_0753_),
    .B1(_0774_),
    .X(_0775_));
 sg13g2_nand2b_1 _1621_ (.Y(_0776_),
    .B(_0713_),
    .A_N(_0715_));
 sg13g2_nand2b_1 _1622_ (.Y(_0777_),
    .B(_0715_),
    .A_N(_0713_));
 sg13g2_and2_1 _1623_ (.A(_0776_),
    .B(_0777_),
    .X(_0778_));
 sg13g2_a221oi_1 _1624_ (.B2(_0777_),
    .C1(_0774_),
    .B1(_0776_),
    .A1(_0753_),
    .Y(_0779_),
    .A2(_0772_));
 sg13g2_a21oi_1 _1625_ (.A1(_0490_),
    .A2(_0714_),
    .Y(_0780_),
    .B1(_0709_));
 sg13g2_xor2_1 _1626_ (.B(_0780_),
    .A(_0563_),
    .X(_0781_));
 sg13g2_or3_1 _1627_ (.A(_0716_),
    .B(_0779_),
    .C(_0781_),
    .X(_0782_));
 sg13g2_nand2_1 _1628_ (.Y(_0783_),
    .A(_0524_),
    .B(_0782_));
 sg13g2_nor2_1 _1629_ (.A(_0711_),
    .B(_0783_),
    .Y(_0784_));
 sg13g2_or2_2 _1630_ (.X(_0785_),
    .B(_0783_),
    .A(_0711_));
 sg13g2_xnor2_1 _1631_ (.Y(_0786_),
    .A(_0737_),
    .B(_0739_));
 sg13g2_xnor2_1 _1632_ (.Y(_0787_),
    .A(_0738_),
    .B(_0739_));
 sg13g2_xor2_1 _1633_ (.B(_0624_),
    .A(_0622_),
    .X(_0788_));
 sg13g2_o21ai_1 _1634_ (.B1(_0781_),
    .Y(_0789_),
    .A1(_0716_),
    .A2(_0779_));
 sg13g2_and3_2 _1635_ (.X(_0790_),
    .A(net341),
    .B(_0782_),
    .C(_0789_));
 sg13g2_nand3_1 _1636_ (.B(_0782_),
    .C(_0789_),
    .A(net341),
    .Y(_0791_));
 sg13g2_o21ai_1 _1637_ (.B1(_0724_),
    .Y(_0792_),
    .A1(_0747_),
    .A2(_0749_));
 sg13g2_or3_1 _1638_ (.A(_0724_),
    .B(_0747_),
    .C(_0749_),
    .X(_0793_));
 sg13g2_nand2_2 _1639_ (.Y(_0794_),
    .A(_0792_),
    .B(_0793_));
 sg13g2_inv_1 _1640_ (.Y(_0795_),
    .A(_0794_));
 sg13g2_o21ai_1 _1641_ (.B1(_0748_),
    .Y(_0796_),
    .A1(_0728_),
    .A2(_0743_));
 sg13g2_and2_2 _1642_ (.A(_0750_),
    .B(_0796_),
    .X(_0797_));
 sg13g2_xnor2_1 _1643_ (.Y(_0798_),
    .A(_0725_),
    .B(_0726_));
 sg13g2_xor2_1 _1644_ (.B(_0798_),
    .A(_0742_),
    .X(_0799_));
 sg13g2_xnor2_1 _1645_ (.Y(_0800_),
    .A(_0742_),
    .B(_0798_));
 sg13g2_xor2_1 _1646_ (.B(_0741_),
    .A(_0740_),
    .X(_0801_));
 sg13g2_or2_1 _1647_ (.X(_0802_),
    .B(_0788_),
    .A(_0786_));
 sg13g2_nand2b_1 _1648_ (.Y(_0803_),
    .B(_0802_),
    .A_N(_0801_));
 sg13g2_a22oi_1 _1649_ (.Y(_0804_),
    .B1(_0800_),
    .B2(_0803_),
    .A2(_0796_),
    .A1(_0750_));
 sg13g2_a21o_1 _1650_ (.A2(_0793_),
    .A1(_0792_),
    .B1(_0804_),
    .X(_0805_));
 sg13g2_xor2_1 _1651_ (.B(_0778_),
    .A(_0775_),
    .X(_0806_));
 sg13g2_xnor2_1 _1652_ (.Y(_0807_),
    .A(_0775_),
    .B(_0778_));
 sg13g2_xnor2_1 _1653_ (.Y(_0808_),
    .A(_0761_),
    .B(_0765_));
 sg13g2_nor2_1 _1654_ (.A(_0752_),
    .B(_0769_),
    .Y(_0809_));
 sg13g2_o21ai_1 _1655_ (.B1(_0808_),
    .Y(_0810_),
    .A1(_0752_),
    .A2(_0769_));
 sg13g2_xor2_1 _1656_ (.B(_0809_),
    .A(_0808_),
    .X(_0811_));
 sg13g2_inv_1 _1657_ (.Y(_0812_),
    .A(_0811_));
 sg13g2_nand3_1 _1658_ (.B(_0807_),
    .C(_0811_),
    .A(_0805_),
    .Y(_0813_));
 sg13g2_nand2_1 _1659_ (.Y(_0814_),
    .A(_0790_),
    .B(_0813_));
 sg13g2_nand2b_1 _1660_ (.Y(_0815_),
    .B(_0771_),
    .A_N(_0760_));
 sg13g2_inv_1 _1661_ (.Y(_0816_),
    .A(_0815_));
 sg13g2_a21oi_2 _1662_ (.B1(_0816_),
    .Y(_0817_),
    .A2(_0810_),
    .A1(_0766_));
 sg13g2_and3_1 _1663_ (.X(_0818_),
    .A(_0766_),
    .B(_0810_),
    .C(_0816_));
 sg13g2_or2_2 _1664_ (.X(_0819_),
    .B(_0818_),
    .A(_0817_));
 sg13g2_nor2_1 _1665_ (.A(_0817_),
    .B(_0818_),
    .Y(_0820_));
 sg13g2_o21ai_1 _1666_ (.B1(_0807_),
    .Y(_0821_),
    .A1(_0817_),
    .A2(_0818_));
 sg13g2_and3_1 _1667_ (.X(_0822_),
    .A(_0790_),
    .B(_0813_),
    .C(_0821_));
 sg13g2_nand3_1 _1668_ (.B(_0813_),
    .C(_0821_),
    .A(_0790_),
    .Y(_0823_));
 sg13g2_nor2_1 _1669_ (.A(_0788_),
    .B(net315),
    .Y(_0824_));
 sg13g2_nor2_1 _1670_ (.A(_0799_),
    .B(_0801_),
    .Y(_0825_));
 sg13g2_or3_1 _1671_ (.A(_0795_),
    .B(_0797_),
    .C(_0825_),
    .X(_0826_));
 sg13g2_and3_1 _1672_ (.X(_0827_),
    .A(_0811_),
    .B(_0820_),
    .C(_0826_));
 sg13g2_nand2_1 _1673_ (.Y(_0828_),
    .A(_0790_),
    .B(_0807_));
 sg13g2_nor2_1 _1674_ (.A(_0827_),
    .B(_0828_),
    .Y(_0829_));
 sg13g2_nor2b_2 _1675_ (.A(net310),
    .B_N(_0824_),
    .Y(_0830_));
 sg13g2_nor2_1 _1676_ (.A(_0791_),
    .B(_0819_),
    .Y(_0831_));
 sg13g2_nand2b_1 _1677_ (.Y(_0832_),
    .B(_0825_),
    .A_N(_0797_));
 sg13g2_or2_1 _1678_ (.X(_0833_),
    .B(_0832_),
    .A(_0795_));
 sg13g2_nand4_1 _1679_ (.B(_0811_),
    .C(_0831_),
    .A(_0807_),
    .Y(_0834_),
    .D(_0833_));
 sg13g2_nor3_1 _1680_ (.A(_0806_),
    .B(_0817_),
    .C(_0818_),
    .Y(_0835_));
 sg13g2_nand2_1 _1681_ (.Y(_0836_),
    .A(_0794_),
    .B(_0811_));
 sg13g2_nor4_2 _1682_ (.A(_0806_),
    .B(_0819_),
    .C(_0832_),
    .Y(_0837_),
    .D(_0836_));
 sg13g2_and2_1 _1683_ (.A(_0787_),
    .B(_0788_),
    .X(_0838_));
 sg13g2_nor2_1 _1684_ (.A(_0791_),
    .B(_0838_),
    .Y(_0839_));
 sg13g2_nand2_1 _1685_ (.Y(_0840_),
    .A(_0837_),
    .B(_0839_));
 sg13g2_and2_1 _1686_ (.A(_0834_),
    .B(_0840_),
    .X(_0841_));
 sg13g2_a21oi_1 _1687_ (.A1(_0837_),
    .A2(_0839_),
    .Y(_0842_),
    .B1(net317));
 sg13g2_and2_2 _1688_ (.A(_0834_),
    .B(_0842_),
    .X(_0843_));
 sg13g2_nand2_1 _1689_ (.Y(_0844_),
    .A(_0834_),
    .B(_0842_));
 sg13g2_a22oi_1 _1690_ (.Y(_0845_),
    .B1(_0830_),
    .B2(_0843_),
    .A2(_0786_),
    .A1(net316));
 sg13g2_or2_1 _1691_ (.X(_0846_),
    .B(_0845_),
    .A(net342));
 sg13g2_mux2_2 _1692_ (.A0(\MAC.add.a1[9] ),
    .A1(\MAC.add.b1[9] ),
    .S(net332),
    .X(_0847_));
 sg13g2_inv_1 _1693_ (.Y(_0848_),
    .A(_0847_));
 sg13g2_nor2_1 _1694_ (.A(\MAC.add.b1[11] ),
    .B(net336),
    .Y(_0849_));
 sg13g2_a21oi_2 _1695_ (.B1(_0849_),
    .Y(_0850_),
    .A2(net336),
    .A1(_0459_));
 sg13g2_inv_1 _1696_ (.Y(_0851_),
    .A(_0850_));
 sg13g2_mux2_2 _1697_ (.A0(\MAC.add.a1[10] ),
    .A1(\MAC.add.b1[10] ),
    .S(net332),
    .X(_0852_));
 sg13g2_inv_1 _1698_ (.Y(_0853_),
    .A(_0852_));
 sg13g2_nor3_2 _1699_ (.A(_0847_),
    .B(_0850_),
    .C(_0852_),
    .Y(_0854_));
 sg13g2_inv_1 _1700_ (.Y(_0855_),
    .A(_0854_));
 sg13g2_nand4_1 _1701_ (.B(_0711_),
    .C(_0782_),
    .A(net341),
    .Y(_0856_),
    .D(_0789_));
 sg13g2_nor2_1 _1702_ (.A(_0802_),
    .B(_0832_),
    .Y(_0857_));
 sg13g2_nor4_2 _1703_ (.A(_0806_),
    .B(_0819_),
    .C(_0836_),
    .Y(_0858_),
    .D(_0857_));
 sg13g2_o21ai_1 _1704_ (.B1(_0851_),
    .Y(_0859_),
    .A1(_0856_),
    .A2(_0858_));
 sg13g2_nor2_1 _1705_ (.A(_0801_),
    .B(_0802_),
    .Y(_0860_));
 sg13g2_or3_1 _1706_ (.A(_0797_),
    .B(_0799_),
    .C(_0860_),
    .X(_0861_));
 sg13g2_nand3_1 _1707_ (.B(_0811_),
    .C(_0861_),
    .A(_0794_),
    .Y(_0862_));
 sg13g2_a21o_1 _1708_ (.A2(_0862_),
    .A1(_0835_),
    .B1(_0856_),
    .X(_0863_));
 sg13g2_nor2_1 _1709_ (.A(_0853_),
    .B(_0863_),
    .Y(_0864_));
 sg13g2_a21oi_1 _1710_ (.A1(_0785_),
    .A2(_0823_),
    .Y(_0865_),
    .B1(_0848_));
 sg13g2_a221oi_1 _1711_ (.B2(_0863_),
    .C1(_0848_),
    .B1(_0853_),
    .A1(_0785_),
    .Y(_0866_),
    .A2(_0823_));
 sg13g2_nor2_1 _1712_ (.A(_0864_),
    .B(_0866_),
    .Y(_0867_));
 sg13g2_or3_1 _1713_ (.A(_0851_),
    .B(_0856_),
    .C(_0858_),
    .X(_0868_));
 sg13g2_o21ai_1 _1714_ (.B1(_0859_),
    .Y(_0869_),
    .A1(_0864_),
    .A2(_0866_));
 sg13g2_and2_1 _1715_ (.A(_0868_),
    .B(_0869_),
    .X(_0870_));
 sg13g2_a21oi_2 _1716_ (.B1(_0856_),
    .Y(_0871_),
    .A2(_0838_),
    .A1(_0837_));
 sg13g2_mux2_2 _1717_ (.A0(\MAC.add.a1[13] ),
    .A1(\MAC.add.b1[13] ),
    .S(net332),
    .X(_0872_));
 sg13g2_nor2_1 _1718_ (.A(\MAC.add.b1[12] ),
    .B(net336),
    .Y(_0873_));
 sg13g2_a21oi_2 _1719_ (.B1(_0873_),
    .Y(_0874_),
    .A2(net336),
    .A1(_0458_));
 sg13g2_nor2_1 _1720_ (.A(_0855_),
    .B(_0874_),
    .Y(_0875_));
 sg13g2_nand2b_1 _1721_ (.Y(_0876_),
    .B(_0875_),
    .A_N(_0872_));
 sg13g2_xnor2_1 _1722_ (.Y(_0877_),
    .A(_0872_),
    .B(_0875_));
 sg13g2_xnor2_1 _1723_ (.Y(_0878_),
    .A(_0555_),
    .B(_0876_));
 sg13g2_o21ai_1 _1724_ (.B1(_0878_),
    .Y(_0879_),
    .A1(_0871_),
    .A2(_0877_));
 sg13g2_xor2_1 _1725_ (.B(_0874_),
    .A(_0854_),
    .X(_0880_));
 sg13g2_a21oi_2 _1726_ (.B1(_0856_),
    .Y(_0881_),
    .A2(_0837_),
    .A1(_0787_));
 sg13g2_o21ai_1 _1727_ (.B1(_0879_),
    .Y(_0882_),
    .A1(_0880_),
    .A2(_0881_));
 sg13g2_a21oi_1 _1728_ (.A1(_0855_),
    .A2(_0870_),
    .Y(_0883_),
    .B1(_0882_));
 sg13g2_a21oi_1 _1729_ (.A1(_0871_),
    .A2(_0877_),
    .Y(_0884_),
    .B1(_0878_));
 sg13g2_nor4_1 _1730_ (.A(_0555_),
    .B(_0872_),
    .C(_0880_),
    .D(_0884_),
    .Y(_0885_));
 sg13g2_nor2b_1 _1731_ (.A(_0883_),
    .B_N(_0885_),
    .Y(_0886_));
 sg13g2_nand4_1 _1732_ (.B(\MAC.add.b1[13] ),
    .C(\MAC.add.b1[15] ),
    .A(\MAC.add.b1[14] ),
    .Y(_0887_),
    .D(\MAC.add.b1[0] ));
 sg13g2_nand4_1 _1733_ (.B(\MAC.add.b1[11] ),
    .C(\MAC.add.b1[10] ),
    .A(\MAC.add.b1[12] ),
    .Y(_0888_),
    .D(\MAC.add.b1[9] ));
 sg13g2_or2_1 _1734_ (.X(_0889_),
    .B(_0888_),
    .A(_0887_));
 sg13g2_nand4_1 _1735_ (.B(\MAC.add.b1[2] ),
    .C(\MAC.add.b1[3] ),
    .A(\MAC.add.b1[1] ),
    .Y(_0890_),
    .D(\MAC.add.b1[4] ));
 sg13g2_nand4_1 _1736_ (.B(net66),
    .C(\MAC.add.b1[7] ),
    .A(\MAC.add.b1[5] ),
    .Y(_0891_),
    .D(\MAC.add.b1[8] ));
 sg13g2_nor3_1 _1737_ (.A(_0889_),
    .B(_0890_),
    .C(_0891_),
    .Y(_0892_));
 sg13g2_nand4_1 _1738_ (.B(\MAC.add.a1[13] ),
    .C(\MAC.add.a1[15] ),
    .A(\MAC.add.a1[14] ),
    .Y(_0893_),
    .D(\MAC.add.a1[0] ));
 sg13g2_nand4_1 _1739_ (.B(\MAC.add.a1[11] ),
    .C(\MAC.add.a1[10] ),
    .A(\MAC.add.a1[12] ),
    .Y(_0894_),
    .D(\MAC.add.a1[9] ));
 sg13g2_nand4_1 _1740_ (.B(\MAC.add.a1[2] ),
    .C(\MAC.add.a1[3] ),
    .A(\MAC.add.a1[1] ),
    .Y(_0895_),
    .D(\MAC.add.a1[4] ));
 sg13g2_nand4_1 _1741_ (.B(\MAC.add.a1[6] ),
    .C(\MAC.add.a1[7] ),
    .A(\MAC.add.a1[5] ),
    .Y(_0896_),
    .D(\MAC.add.a1[8] ));
 sg13g2_nor4_2 _1742_ (.A(_0893_),
    .B(_0894_),
    .C(_0895_),
    .Y(_0897_),
    .D(_0896_));
 sg13g2_nor2_1 _1743_ (.A(_0892_),
    .B(_0897_),
    .Y(_0898_));
 sg13g2_nor3_1 _1744_ (.A(_0889_),
    .B(_0890_),
    .C(_0891_),
    .Y(_0899_));
 sg13g2_nor4_2 _1745_ (.A(_0893_),
    .B(_0894_),
    .C(_0895_),
    .Y(_0900_),
    .D(_0896_));
 sg13g2_nor2_1 _1746_ (.A(_0899_),
    .B(_0900_),
    .Y(_0901_));
 sg13g2_nor2b_1 _1747_ (.A(net307),
    .B_N(_0901_),
    .Y(_0902_));
 sg13g2_and4_1 _1748_ (.A(_0847_),
    .B(_0850_),
    .C(_0852_),
    .D(_0874_),
    .X(_0903_));
 sg13g2_and4_1 _1749_ (.A(_0555_),
    .B(net318),
    .C(_0872_),
    .D(_0903_),
    .X(_0904_));
 sg13g2_and4_1 _1750_ (.A(_0555_),
    .B(net318),
    .C(_0872_),
    .D(_0903_),
    .X(_0905_));
 sg13g2_nand4_1 _1751_ (.B(net318),
    .C(_0872_),
    .A(_0555_),
    .Y(_0906_),
    .D(_0903_));
 sg13g2_a21oi_1 _1752_ (.A1(_0846_),
    .A2(_0902_),
    .Y(\MAC.add.c_add[0] ),
    .B1(_0905_));
 sg13g2_nor2_1 _1753_ (.A(_0788_),
    .B(_0823_),
    .Y(_0907_));
 sg13g2_a21oi_1 _1754_ (.A1(_0786_),
    .A2(_0823_),
    .Y(_0908_),
    .B1(_0907_));
 sg13g2_nor2_1 _1755_ (.A(net310),
    .B(_0908_),
    .Y(_0909_));
 sg13g2_a21oi_1 _1756_ (.A1(_0841_),
    .A2(_0909_),
    .Y(_0910_),
    .B1(net317));
 sg13g2_nor2_1 _1757_ (.A(_0785_),
    .B(_0801_),
    .Y(_0911_));
 sg13g2_or2_1 _1758_ (.X(_0912_),
    .B(_0911_),
    .A(net342));
 sg13g2_nor2b_2 _1759_ (.A(_0904_),
    .B_N(_0898_),
    .Y(_0913_));
 sg13g2_o21ai_1 _1760_ (.B1(net308),
    .Y(\MAC.add.c_add[1] ),
    .A1(_0910_),
    .A2(_0912_));
 sg13g2_nor2_1 _1761_ (.A(_0801_),
    .B(_0822_),
    .Y(_0914_));
 sg13g2_a21oi_1 _1762_ (.A1(_0787_),
    .A2(_0822_),
    .Y(_0915_),
    .B1(_0914_));
 sg13g2_mux2_1 _1763_ (.A0(_0915_),
    .A1(_0824_),
    .S(net309),
    .X(_0916_));
 sg13g2_a22oi_1 _1764_ (.Y(_0917_),
    .B1(_0843_),
    .B2(_0916_),
    .A2(_0799_),
    .A1(net316));
 sg13g2_o21ai_1 _1765_ (.B1(net308),
    .Y(_0918_),
    .A1(net342),
    .A2(_0917_));
 sg13g2_nor2b_1 _1766_ (.A(net306),
    .B_N(_0918_),
    .Y(\MAC.add.c_add[2] ));
 sg13g2_nand2_1 _1767_ (.Y(_0919_),
    .A(_0801_),
    .B(net315));
 sg13g2_o21ai_1 _1768_ (.B1(_0919_),
    .Y(_0920_),
    .A1(_0800_),
    .A2(net315));
 sg13g2_nor2_1 _1769_ (.A(net309),
    .B(_0920_),
    .Y(_0921_));
 sg13g2_a21oi_2 _1770_ (.B1(_0921_),
    .Y(_0922_),
    .A2(_0908_),
    .A1(net310));
 sg13g2_a22oi_1 _1771_ (.Y(_0923_),
    .B1(_0843_),
    .B2(_0922_),
    .A2(_0797_),
    .A1(net316));
 sg13g2_o21ai_1 _1772_ (.B1(net308),
    .Y(_0924_),
    .A1(net342),
    .A2(_0923_));
 sg13g2_nor2b_1 _1773_ (.A(net306),
    .B_N(_0924_),
    .Y(\MAC.add.c_add[3] ));
 sg13g2_nor2_1 _1774_ (.A(_0800_),
    .B(_0823_),
    .Y(_0925_));
 sg13g2_a21oi_1 _1775_ (.A1(_0797_),
    .A2(_0823_),
    .Y(_0926_),
    .B1(_0925_));
 sg13g2_nor2_1 _1776_ (.A(net309),
    .B(_0926_),
    .Y(_0927_));
 sg13g2_a21oi_2 _1777_ (.B1(_0927_),
    .Y(_0928_),
    .A2(_0915_),
    .A1(net310));
 sg13g2_nor2b_2 _1778_ (.A(_0834_),
    .B_N(_0842_),
    .Y(_0929_));
 sg13g2_a22oi_1 _1779_ (.Y(_0930_),
    .B1(_0830_),
    .B2(_0929_),
    .A2(_0795_),
    .A1(net316));
 sg13g2_o21ai_1 _1780_ (.B1(_0930_),
    .Y(_0931_),
    .A1(_0844_),
    .A2(_0928_));
 sg13g2_nand2b_1 _1781_ (.Y(_0932_),
    .B(_0931_),
    .A_N(net342));
 sg13g2_a21oi_1 _1782_ (.A1(net308),
    .A2(_0932_),
    .Y(\MAC.add.c_add[4] ),
    .B1(net306));
 sg13g2_nor2_1 _1783_ (.A(_0794_),
    .B(net315),
    .Y(_0933_));
 sg13g2_a21oi_1 _1784_ (.A1(_0797_),
    .A2(net315),
    .Y(_0934_),
    .B1(_0933_));
 sg13g2_nand2b_1 _1785_ (.Y(_0935_),
    .B(_0934_),
    .A_N(net309));
 sg13g2_or3_1 _1786_ (.A(_0827_),
    .B(_0828_),
    .C(_0920_),
    .X(_0936_));
 sg13g2_nand3_1 _1787_ (.B(_0935_),
    .C(_0936_),
    .A(_0843_),
    .Y(_0937_));
 sg13g2_a22oi_1 _1788_ (.Y(_0938_),
    .B1(_0909_),
    .B2(_0929_),
    .A2(_0812_),
    .A1(net316));
 sg13g2_a21o_1 _1789_ (.A2(_0938_),
    .A1(_0937_),
    .B1(_0489_),
    .X(_0939_));
 sg13g2_a21oi_1 _1790_ (.A1(net308),
    .A2(_0939_),
    .Y(\MAC.add.c_add[5] ),
    .B1(net306));
 sg13g2_nor2_1 _1791_ (.A(_0811_),
    .B(net315),
    .Y(_0940_));
 sg13g2_a21oi_1 _1792_ (.A1(_0795_),
    .A2(net315),
    .Y(_0941_),
    .B1(_0940_));
 sg13g2_nand2b_1 _1793_ (.Y(_0942_),
    .B(_0941_),
    .A_N(net309));
 sg13g2_nand2_1 _1794_ (.Y(_0943_),
    .A(net310),
    .B(_0926_));
 sg13g2_nand3_1 _1795_ (.B(_0942_),
    .C(_0943_),
    .A(_0843_),
    .Y(_0944_));
 sg13g2_a22oi_1 _1796_ (.Y(_0945_),
    .B1(_0916_),
    .B2(_0929_),
    .A2(_0819_),
    .A1(net316));
 sg13g2_a21o_1 _1797_ (.A2(_0945_),
    .A1(_0944_),
    .B1(net342),
    .X(_0946_));
 sg13g2_a21oi_1 _1798_ (.A1(net308),
    .A2(_0946_),
    .Y(\MAC.add.c_add[6] ),
    .B1(net306));
 sg13g2_a22oi_1 _1799_ (.Y(_0947_),
    .B1(net315),
    .B2(_0811_),
    .A2(_0820_),
    .A1(_0814_));
 sg13g2_or2_1 _1800_ (.X(_0948_),
    .B(_0947_),
    .A(net309));
 sg13g2_nand2_1 _1801_ (.Y(_0949_),
    .A(net309),
    .B(_0934_));
 sg13g2_nand3_1 _1802_ (.B(_0948_),
    .C(_0949_),
    .A(_0843_),
    .Y(_0950_));
 sg13g2_a22oi_1 _1803_ (.Y(_0951_),
    .B1(_0922_),
    .B2(_0929_),
    .A2(_0806_),
    .A1(net316));
 sg13g2_a21o_1 _1804_ (.A2(_0951_),
    .A1(_0950_),
    .B1(net342),
    .X(_0952_));
 sg13g2_a21oi_1 _1805_ (.A1(net308),
    .A2(_0952_),
    .Y(\MAC.add.c_add[7] ),
    .B1(net306));
 sg13g2_nand2b_1 _1806_ (.Y(_0953_),
    .B(net309),
    .A_N(_0941_));
 sg13g2_o21ai_1 _1807_ (.B1(_0953_),
    .Y(_0954_),
    .A1(_0807_),
    .A2(_0831_));
 sg13g2_a21oi_1 _1808_ (.A1(_0830_),
    .A2(_0834_),
    .Y(_0955_),
    .B1(net317));
 sg13g2_a21oi_1 _1809_ (.A1(_0928_),
    .A2(_0955_),
    .Y(_0956_),
    .B1(_0843_));
 sg13g2_a21oi_1 _1810_ (.A1(net316),
    .A2(_0790_),
    .Y(_0957_),
    .B1(net342));
 sg13g2_o21ai_1 _1811_ (.B1(_0957_),
    .Y(_0958_),
    .A1(_0954_),
    .A2(_0956_));
 sg13g2_a21oi_1 _1812_ (.A1(net308),
    .A2(_0958_),
    .Y(\MAC.add.c_add[8] ),
    .B1(net306));
 sg13g2_nand3_1 _1813_ (.B(_0823_),
    .C(_0848_),
    .A(_0785_),
    .Y(_0959_));
 sg13g2_nand2b_1 _1814_ (.Y(_0960_),
    .B(_0959_),
    .A_N(_0865_));
 sg13g2_a21oi_1 _1815_ (.A1(_0902_),
    .A2(_0960_),
    .Y(\MAC.add.c_add[9] ),
    .B1(_0905_));
 sg13g2_xnor2_1 _1816_ (.Y(_0961_),
    .A(_0852_),
    .B(_0863_));
 sg13g2_xnor2_1 _1817_ (.Y(_0962_),
    .A(_0865_),
    .B(_0961_));
 sg13g2_nand3_1 _1818_ (.B(_0906_),
    .C(_0962_),
    .A(_0901_),
    .Y(_0963_));
 sg13g2_nor2b_1 _1819_ (.A(net306),
    .B_N(_0963_),
    .Y(\MAC.add.c_add[10] ));
 sg13g2_nand2_1 _1820_ (.Y(_0964_),
    .A(_0859_),
    .B(_0868_));
 sg13g2_xnor2_1 _1821_ (.Y(_0965_),
    .A(_0867_),
    .B(_0964_));
 sg13g2_nand3_1 _1822_ (.B(_0906_),
    .C(_0965_),
    .A(_0901_),
    .Y(_0966_));
 sg13g2_nor2b_1 _1823_ (.A(net307),
    .B_N(_0966_),
    .Y(\MAC.add.c_add[11] ));
 sg13g2_nand2_1 _1824_ (.Y(_0967_),
    .A(_0874_),
    .B(_0881_));
 sg13g2_xnor2_1 _1825_ (.Y(_0968_),
    .A(_0874_),
    .B(_0881_));
 sg13g2_a21o_1 _1826_ (.A2(_0869_),
    .A1(_0868_),
    .B1(_0968_),
    .X(_0969_));
 sg13g2_xnor2_1 _1827_ (.Y(_0970_),
    .A(_0870_),
    .B(_0968_));
 sg13g2_a21oi_1 _1828_ (.A1(_0913_),
    .A2(_0970_),
    .Y(\MAC.add.c_add[12] ),
    .B1(net307));
 sg13g2_and2_1 _1829_ (.A(_0871_),
    .B(_0872_),
    .X(_0971_));
 sg13g2_xnor2_1 _1830_ (.Y(_0972_),
    .A(_0871_),
    .B(_0872_));
 sg13g2_a21oi_1 _1831_ (.A1(_0967_),
    .A2(_0969_),
    .Y(_0973_),
    .B1(_0972_));
 sg13g2_nand3_1 _1832_ (.B(_0969_),
    .C(_0972_),
    .A(_0967_),
    .Y(_0974_));
 sg13g2_nand2b_1 _1833_ (.Y(_0975_),
    .B(_0974_),
    .A_N(_0973_));
 sg13g2_a21oi_1 _1834_ (.A1(_0913_),
    .A2(_0975_),
    .Y(\MAC.add.c_add[13] ),
    .B1(net307));
 sg13g2_xnor2_1 _1835_ (.Y(_0976_),
    .A(_0555_),
    .B(_0871_));
 sg13g2_o21ai_1 _1836_ (.B1(_0976_),
    .Y(_0977_),
    .A1(_0971_),
    .A2(_0973_));
 sg13g2_nor3_1 _1837_ (.A(_0971_),
    .B(_0973_),
    .C(_0976_),
    .Y(_0978_));
 sg13g2_nor2b_1 _1838_ (.A(_0978_),
    .B_N(_0913_),
    .Y(_0979_));
 sg13g2_a21oi_1 _1839_ (.A1(_0977_),
    .A2(_0979_),
    .Y(\MAC.add.c_add[14] ),
    .B1(net307));
 sg13g2_nor3_2 _1840_ (.A(_0531_),
    .B(_0533_),
    .C(_0556_),
    .Y(_0980_));
 sg13g2_nand2_1 _1841_ (.Y(_0981_),
    .A(_0471_),
    .B(\MAC.add.a1[8] ));
 sg13g2_nand2_1 _1842_ (.Y(_0982_),
    .A(\MAC.add.b1[7] ),
    .B(_0469_));
 sg13g2_o21ai_1 _1843_ (.B1(_0982_),
    .Y(_0983_),
    .A1(_0466_),
    .A2(\MAC.add.a1[6] ));
 sg13g2_a22oi_1 _1844_ (.Y(_0984_),
    .B1(_0468_),
    .B2(\MAC.add.a1[7] ),
    .A2(\MAC.add.a1[6] ),
    .A1(_0466_));
 sg13g2_nor2b_1 _1845_ (.A(_0983_),
    .B_N(_0984_),
    .Y(_0985_));
 sg13g2_nand2b_1 _1846_ (.Y(_0986_),
    .B(\MAC.add.a1[5] ),
    .A_N(\MAC.add.b1[5] ));
 sg13g2_nand2b_1 _1847_ (.Y(_0987_),
    .B(\MAC.add.a1[4] ),
    .A_N(\MAC.add.b1[4] ));
 sg13g2_nand3_1 _1848_ (.B(_0986_),
    .C(_0987_),
    .A(_0985_),
    .Y(_0988_));
 sg13g2_nand2_1 _1849_ (.Y(_0989_),
    .A(\MAC.add.b1[2] ),
    .B(_0461_));
 sg13g2_o21ai_1 _1850_ (.B1(_0989_),
    .Y(_0990_),
    .A1(_0463_),
    .A2(\MAC.add.a1[3] ));
 sg13g2_nand2_1 _1851_ (.Y(_0991_),
    .A(_0463_),
    .B(\MAC.add.a1[3] ));
 sg13g2_o21ai_1 _1852_ (.B1(_0991_),
    .Y(_0992_),
    .A1(\MAC.add.b1[2] ),
    .A2(_0461_));
 sg13g2_nor2_1 _1853_ (.A(_0990_),
    .B(_0992_),
    .Y(_0993_));
 sg13g2_nor2b_1 _1854_ (.A(\MAC.add.b1[0] ),
    .B_N(\MAC.add.a1[0] ),
    .Y(_0994_));
 sg13g2_nand2b_1 _1855_ (.Y(_0995_),
    .B(\MAC.add.b1[1] ),
    .A_N(\MAC.add.a1[1] ));
 sg13g2_nor2b_1 _1856_ (.A(\MAC.add.b1[1] ),
    .B_N(\MAC.add.a1[1] ),
    .Y(_0996_));
 sg13g2_nor2_1 _1857_ (.A(_0994_),
    .B(_0996_),
    .Y(_0997_));
 sg13g2_nor2b_1 _1858_ (.A(\MAC.add.a1[4] ),
    .B_N(\MAC.add.b1[4] ),
    .Y(_0998_));
 sg13g2_o21ai_1 _1859_ (.B1(_0995_),
    .Y(_0999_),
    .A1(_0994_),
    .A2(_0996_));
 sg13g2_a221oi_1 _1860_ (.B2(_0999_),
    .C1(_0998_),
    .B1(_0993_),
    .A1(_0990_),
    .Y(_1000_),
    .A2(_0991_));
 sg13g2_nor2_1 _1861_ (.A(_0988_),
    .B(_1000_),
    .Y(_1001_));
 sg13g2_nand2b_1 _1862_ (.Y(_1002_),
    .B(\MAC.add.b1[5] ),
    .A_N(\MAC.add.a1[5] ));
 sg13g2_nand3b_1 _1863_ (.B(_0985_),
    .C(\MAC.add.b1[5] ),
    .Y(_1003_),
    .A_N(\MAC.add.a1[5] ));
 sg13g2_o21ai_1 _1864_ (.B1(_0983_),
    .Y(_1004_),
    .A1(\MAC.add.b1[7] ),
    .A2(_0469_));
 sg13g2_nand2b_1 _1865_ (.Y(_1005_),
    .B(\MAC.add.b1[8] ),
    .A_N(\MAC.add.a1[8] ));
 sg13g2_nand3_1 _1866_ (.B(_1004_),
    .C(_1005_),
    .A(_1003_),
    .Y(_1006_));
 sg13g2_o21ai_1 _1867_ (.B1(_0981_),
    .Y(_1007_),
    .A1(_1001_),
    .A2(_1006_));
 sg13g2_nand2b_1 _1868_ (.Y(_1008_),
    .B(\MAC.add.b1[0] ),
    .A_N(\MAC.add.a1[0] ));
 sg13g2_nand3_1 _1869_ (.B(_1005_),
    .C(_1008_),
    .A(_1002_),
    .Y(_1009_));
 sg13g2_a21oi_1 _1870_ (.A1(_0471_),
    .A2(\MAC.add.a1[8] ),
    .Y(_1010_),
    .B1(_0998_));
 sg13g2_nand4_1 _1871_ (.B(_0995_),
    .C(_0997_),
    .A(_0993_),
    .Y(_1011_),
    .D(_1010_));
 sg13g2_nor3_1 _1872_ (.A(_0988_),
    .B(_1009_),
    .C(_1011_),
    .Y(_1012_));
 sg13g2_o21ai_1 _1873_ (.B1(_0980_),
    .Y(_1013_),
    .A1(_1007_),
    .A2(_1012_));
 sg13g2_and2_1 _1874_ (.A(\MAC.add.a1[15] ),
    .B(_0980_),
    .X(_1014_));
 sg13g2_a22oi_1 _1875_ (.Y(_1015_),
    .B1(_1014_),
    .B2(_1007_),
    .A2(_1013_),
    .A1(\MAC.add.b1[15] ));
 sg13g2_xnor2_1 _1876_ (.Y(_1016_),
    .A(net336),
    .B(_1015_));
 sg13g2_a21o_1 _1877_ (.A2(\MAC.add.b1[15] ),
    .A1(\MAC.add.a1[15] ),
    .B1(_1016_),
    .X(_1017_));
 sg13g2_o21ai_1 _1878_ (.B1(_1017_),
    .Y(_1018_),
    .A1(net78),
    .A2(\MAC.add.b1[15] ));
 sg13g2_o21ai_1 _1879_ (.B1(net79),
    .Y(\MAC.add.c_add[15] ),
    .A1(_0898_),
    .A2(_0904_));
 sg13g2_nor2_1 _1880_ (.A(\MAC.b[14] ),
    .B(\MAC.a[14] ),
    .Y(_1019_));
 sg13g2_xnor2_1 _1881_ (.Y(_1020_),
    .A(\MAC.b[14] ),
    .B(\MAC.a[14] ));
 sg13g2_and2_1 _1882_ (.A(\MAC.b[13] ),
    .B(\MAC.a[13] ),
    .X(_1021_));
 sg13g2_nand2_1 _1883_ (.Y(_1022_),
    .A(\MAC.b[12] ),
    .B(\MAC.a[12] ));
 sg13g2_xnor2_1 _1884_ (.Y(_1023_),
    .A(\MAC.b[12] ),
    .B(\MAC.a[12] ));
 sg13g2_nand2_1 _1885_ (.Y(_1024_),
    .A(\MAC.b[10] ),
    .B(\MAC.a[10] ));
 sg13g2_nand2_1 _1886_ (.Y(_1025_),
    .A(\MAC.b[9] ),
    .B(\MAC.a[9] ));
 sg13g2_xor2_1 _1887_ (.B(\MAC.a[10] ),
    .A(\MAC.b[10] ),
    .X(_1026_));
 sg13g2_nand2b_1 _1888_ (.Y(_1027_),
    .B(_1026_),
    .A_N(_1025_));
 sg13g2_xnor2_1 _1889_ (.Y(_1028_),
    .A(\MAC.b[11] ),
    .B(\MAC.a[11] ));
 sg13g2_a21oi_1 _1890_ (.A1(_1024_),
    .A2(_1027_),
    .Y(_1029_),
    .B1(_1028_));
 sg13g2_a21oi_1 _1891_ (.A1(\MAC.b[11] ),
    .A2(\MAC.a[11] ),
    .Y(_1030_),
    .B1(_1029_));
 sg13g2_o21ai_1 _1892_ (.B1(_1022_),
    .Y(_1031_),
    .A1(_1023_),
    .A2(_1030_));
 sg13g2_xor2_1 _1893_ (.B(\MAC.a[13] ),
    .A(\MAC.b[13] ),
    .X(_1032_));
 sg13g2_a21oi_2 _1894_ (.B1(_1021_),
    .Y(_1033_),
    .A2(_1032_),
    .A1(_1031_));
 sg13g2_nor2_1 _1895_ (.A(_1020_),
    .B(_1033_),
    .Y(_1034_));
 sg13g2_a21oi_1 _1896_ (.A1(\MAC.b[14] ),
    .A2(\MAC.a[14] ),
    .Y(_1035_),
    .B1(_1034_));
 sg13g2_xor2_1 _1897_ (.B(\MAC.a[9] ),
    .A(\MAC.b[9] ),
    .X(_1036_));
 sg13g2_nand2_1 _1898_ (.Y(_1037_),
    .A(_1026_),
    .B(_1036_));
 sg13g2_nor3_1 _1899_ (.A(_1023_),
    .B(_1028_),
    .C(_1037_),
    .Y(_1038_));
 sg13g2_nand2_1 _1900_ (.Y(_1039_),
    .A(_1032_),
    .B(_1038_));
 sg13g2_xor2_1 _1901_ (.B(_1033_),
    .A(_1020_),
    .X(_1040_));
 sg13g2_xnor2_1 _1902_ (.Y(_1041_),
    .A(_1039_),
    .B(_1040_));
 sg13g2_nand2b_1 _1903_ (.Y(_1042_),
    .B(_1041_),
    .A_N(_1035_));
 sg13g2_and2_1 _1904_ (.A(_1019_),
    .B(_1033_),
    .X(_1043_));
 sg13g2_inv_1 _1905_ (.Y(_1044_),
    .A(net326));
 sg13g2_nand2_1 _1906_ (.Y(_1045_),
    .A(_1042_),
    .B(_1044_));
 sg13g2_nor4_1 _1907_ (.A(\MAC.b[14] ),
    .B(\MAC.b[13] ),
    .C(net374),
    .D(net372),
    .Y(_1046_));
 sg13g2_nor4_1 _1908_ (.A(\MAC.b[10] ),
    .B(\MAC.b[9] ),
    .C(\MAC.b[12] ),
    .D(\MAC.b[11] ),
    .Y(_1047_));
 sg13g2_nor4_1 _1909_ (.A(net370),
    .B(net368),
    .C(net366),
    .D(net364),
    .Y(_1048_));
 sg13g2_nor4_1 _1910_ (.A(net362),
    .B(net359),
    .C(net357),
    .D(\MAC.b[15] ),
    .Y(_1049_));
 sg13g2_and3_1 _1911_ (.X(_1050_),
    .A(_1046_),
    .B(_1047_),
    .C(_1049_));
 sg13g2_nor4_1 _1912_ (.A(\MAC.a[14] ),
    .B(\MAC.a[13] ),
    .C(net392),
    .D(net391),
    .Y(_1051_));
 sg13g2_nor4_1 _1913_ (.A(\MAC.a[10] ),
    .B(\MAC.a[9] ),
    .C(\MAC.a[12] ),
    .D(\MAC.a[11] ),
    .Y(_1052_));
 sg13g2_nor4_1 _1914_ (.A(net389),
    .B(net387),
    .C(net385),
    .D(net382),
    .Y(_1053_));
 sg13g2_nor4_1 _1915_ (.A(net381),
    .B(net379),
    .C(net377),
    .D(\MAC.a[15] ),
    .Y(_1054_));
 sg13g2_and3_1 _1916_ (.X(_1055_),
    .A(_1051_),
    .B(_1052_),
    .C(_1054_));
 sg13g2_a22oi_1 _1917_ (.Y(_1056_),
    .B1(_1053_),
    .B2(_1055_),
    .A2(_1050_),
    .A1(_1048_));
 sg13g2_nand2_1 _1918_ (.Y(_1057_),
    .A(net376),
    .B(net356));
 sg13g2_nand2_2 _1919_ (.Y(_1058_),
    .A(net379),
    .B(net358));
 sg13g2_nor2_1 _1920_ (.A(net376),
    .B(net357),
    .Y(_1059_));
 sg13g2_o21ai_1 _1921_ (.B1(_1057_),
    .Y(_1060_),
    .A1(_1058_),
    .A2(_1059_));
 sg13g2_and2_2 _1922_ (.A(net380),
    .B(net378),
    .X(_1061_));
 sg13g2_nand2_1 _1923_ (.Y(_1062_),
    .A(net356),
    .B(_1061_));
 sg13g2_nand2_1 _1924_ (.Y(_1063_),
    .A(net376),
    .B(net358));
 sg13g2_a21oi_1 _1925_ (.A1(net378),
    .A2(net356),
    .Y(_1064_),
    .B1(net380));
 sg13g2_a21oi_1 _1926_ (.A1(net356),
    .A2(_1061_),
    .Y(_1065_),
    .B1(_1064_));
 sg13g2_o21ai_1 _1927_ (.B1(_1062_),
    .Y(_1066_),
    .A1(_1063_),
    .A2(_1064_));
 sg13g2_nor2_1 _1928_ (.A(net378),
    .B(_1057_),
    .Y(_1067_));
 sg13g2_xor2_1 _1929_ (.B(_1057_),
    .A(net378),
    .X(_1068_));
 sg13g2_nand2b_1 _1930_ (.Y(_1069_),
    .B(net358),
    .A_N(_1068_));
 sg13g2_xnor2_1 _1931_ (.Y(_1070_),
    .A(net358),
    .B(_1068_));
 sg13g2_nand2_1 _1932_ (.Y(_1071_),
    .A(_1066_),
    .B(_1070_));
 sg13g2_xnor2_1 _1933_ (.Y(_1072_),
    .A(_1066_),
    .B(_1070_));
 sg13g2_nand3_1 _1934_ (.B(net381),
    .C(\MAC.b[8] ),
    .A(net383),
    .Y(_1073_));
 sg13g2_a21o_1 _1935_ (.A2(net357),
    .A1(net381),
    .B1(net383),
    .X(_1074_));
 sg13g2_nand2_1 _1936_ (.Y(_1075_),
    .A(_1073_),
    .B(_1074_));
 sg13g2_o21ai_1 _1937_ (.B1(_1073_),
    .Y(_1076_),
    .A1(_1058_),
    .A2(_1075_));
 sg13g2_xnor2_1 _1938_ (.Y(_1077_),
    .A(_1063_),
    .B(_1065_));
 sg13g2_nand2_1 _1939_ (.Y(_1078_),
    .A(_1076_),
    .B(_1077_));
 sg13g2_xnor2_1 _1940_ (.Y(_1079_),
    .A(_1076_),
    .B(_1077_));
 sg13g2_inv_1 _1941_ (.Y(_1080_),
    .A(_1079_));
 sg13g2_nand2_1 _1942_ (.Y(_1081_),
    .A(net360),
    .B(_1080_));
 sg13g2_a21oi_1 _1943_ (.A1(_1078_),
    .A2(_1081_),
    .Y(_1082_),
    .B1(_1072_));
 sg13g2_nor2_1 _1944_ (.A(_1059_),
    .B(_1067_),
    .Y(_1083_));
 sg13g2_xnor2_1 _1945_ (.Y(_1084_),
    .A(_1069_),
    .B(_1083_));
 sg13g2_a22oi_1 _1946_ (.Y(_1085_),
    .B1(_1082_),
    .B2(_1084_),
    .A2(_1070_),
    .A1(_1066_));
 sg13g2_nand2b_1 _1947_ (.Y(_1086_),
    .B(_1085_),
    .A_N(_1060_));
 sg13g2_nand3_1 _1948_ (.B(_1078_),
    .C(_1081_),
    .A(_1072_),
    .Y(_1087_));
 sg13g2_nand2b_1 _1949_ (.Y(_1088_),
    .B(_1087_),
    .A_N(_1082_));
 sg13g2_and2_1 _1950_ (.A(net385),
    .B(net382),
    .X(_1089_));
 sg13g2_nand2_1 _1951_ (.Y(_1090_),
    .A(net357),
    .B(_1089_));
 sg13g2_nand2_1 _1952_ (.Y(_1091_),
    .A(net381),
    .B(net359));
 sg13g2_a21oi_1 _1953_ (.A1(net383),
    .A2(net357),
    .Y(_1092_),
    .B1(net385));
 sg13g2_a21oi_1 _1954_ (.A1(net357),
    .A2(_1089_),
    .Y(_1093_),
    .B1(_1092_));
 sg13g2_o21ai_1 _1955_ (.B1(_1090_),
    .Y(_1094_),
    .A1(_1091_),
    .A2(_1092_));
 sg13g2_xor2_1 _1956_ (.B(_1075_),
    .A(_1058_),
    .X(_1095_));
 sg13g2_nand2_1 _1957_ (.Y(_1096_),
    .A(_1094_),
    .B(_1095_));
 sg13g2_nand2_1 _1958_ (.Y(_1097_),
    .A(net377),
    .B(net362));
 sg13g2_nor2_1 _1959_ (.A(_0042_),
    .B(_1097_),
    .Y(_1098_));
 sg13g2_xnor2_1 _1960_ (.Y(_1099_),
    .A(_0042_),
    .B(_1097_));
 sg13g2_xnor2_1 _1961_ (.Y(_1100_),
    .A(_1094_),
    .B(_1095_));
 sg13g2_o21ai_1 _1962_ (.B1(_1096_),
    .Y(_1101_),
    .A1(_1099_),
    .A2(_1100_));
 sg13g2_xor2_1 _1963_ (.B(_1079_),
    .A(net360),
    .X(_1102_));
 sg13g2_nor2b_1 _1964_ (.A(_1102_),
    .B_N(_1101_),
    .Y(_1103_));
 sg13g2_xnor2_1 _1965_ (.Y(_1104_),
    .A(_1101_),
    .B(_1102_));
 sg13g2_a21o_1 _1966_ (.A2(_1104_),
    .A1(_1098_),
    .B1(_1103_),
    .X(_1105_));
 sg13g2_nor2b_1 _1967_ (.A(_1088_),
    .B_N(_1105_),
    .Y(_1106_));
 sg13g2_nand2_1 _1968_ (.Y(_1107_),
    .A(_1071_),
    .B(_1084_));
 sg13g2_and3_1 _1969_ (.X(_1108_),
    .A(_1071_),
    .B(_1084_),
    .C(_1106_));
 sg13g2_xnor2_1 _1970_ (.Y(_1109_),
    .A(_1098_),
    .B(_1104_));
 sg13g2_nand3_1 _1971_ (.B(net385),
    .C(net356),
    .A(net387),
    .Y(_1110_));
 sg13g2_nand2_1 _1972_ (.Y(_1111_),
    .A(net383),
    .B(net359));
 sg13g2_a21o_1 _1973_ (.A2(net356),
    .A1(net385),
    .B1(net387),
    .X(_1112_));
 sg13g2_nand2_1 _1974_ (.Y(_1113_),
    .A(_1110_),
    .B(_1112_));
 sg13g2_o21ai_1 _1975_ (.B1(_1110_),
    .Y(_1114_),
    .A1(_1111_),
    .A2(_1113_));
 sg13g2_xnor2_1 _1976_ (.Y(_1115_),
    .A(_1091_),
    .B(_1093_));
 sg13g2_nand2_1 _1977_ (.Y(_1116_),
    .A(_1114_),
    .B(_1115_));
 sg13g2_xnor2_1 _1978_ (.Y(_1117_),
    .A(_1114_),
    .B(_1115_));
 sg13g2_nand2_1 _1979_ (.Y(_1118_),
    .A(net378),
    .B(net360));
 sg13g2_nand2_1 _1980_ (.Y(_1119_),
    .A(net376),
    .B(net363));
 sg13g2_xor2_1 _1981_ (.B(_1119_),
    .A(_1118_),
    .X(_1120_));
 sg13g2_nand2_1 _1982_ (.Y(_1121_),
    .A(net365),
    .B(_1120_));
 sg13g2_xnor2_1 _1983_ (.Y(_1122_),
    .A(net365),
    .B(_1120_));
 sg13g2_o21ai_1 _1984_ (.B1(_1116_),
    .Y(_1123_),
    .A1(_1117_),
    .A2(_1122_));
 sg13g2_xnor2_1 _1985_ (.Y(_1124_),
    .A(_1099_),
    .B(_1100_));
 sg13g2_nand2b_1 _1986_ (.Y(_1125_),
    .B(_1123_),
    .A_N(_1124_));
 sg13g2_o21ai_1 _1987_ (.B1(_1121_),
    .Y(_1126_),
    .A1(_1118_),
    .A2(_1119_));
 sg13g2_inv_1 _1988_ (.Y(_1127_),
    .A(_1126_));
 sg13g2_xor2_1 _1989_ (.B(_1124_),
    .A(_1123_),
    .X(_1128_));
 sg13g2_o21ai_1 _1990_ (.B1(_1125_),
    .Y(_1129_),
    .A1(_1127_),
    .A2(_1128_));
 sg13g2_nand2b_1 _1991_ (.Y(_1130_),
    .B(_1129_),
    .A_N(_1109_));
 sg13g2_xor2_1 _1992_ (.B(_1105_),
    .A(_1088_),
    .X(_1131_));
 sg13g2_or2_1 _1993_ (.X(_1132_),
    .B(_1131_),
    .A(_1130_));
 sg13g2_nor2_1 _1994_ (.A(_1082_),
    .B(_1106_),
    .Y(_1133_));
 sg13g2_xnor2_1 _1995_ (.Y(_1134_),
    .A(_1107_),
    .B(_1133_));
 sg13g2_xor2_1 _1996_ (.B(_1134_),
    .A(_1132_),
    .X(_1135_));
 sg13g2_xor2_1 _1997_ (.B(_1129_),
    .A(_1109_),
    .X(_1136_));
 sg13g2_xnor2_1 _1998_ (.Y(_1137_),
    .A(_1127_),
    .B(_1128_));
 sg13g2_nor2_2 _1999_ (.A(_0473_),
    .B(_0474_),
    .Y(_1138_));
 sg13g2_nand2_1 _2000_ (.Y(_1139_),
    .A(net356),
    .B(_1138_));
 sg13g2_nand2_1 _2001_ (.Y(_1140_),
    .A(net384),
    .B(net359));
 sg13g2_a21oi_1 _2002_ (.A1(net386),
    .A2(net355),
    .Y(_1141_),
    .B1(net388));
 sg13g2_a21oi_1 _2003_ (.A1(net355),
    .A2(_1138_),
    .Y(_1142_),
    .B1(_1141_));
 sg13g2_o21ai_1 _2004_ (.B1(_1139_),
    .Y(_1143_),
    .A1(_1140_),
    .A2(_1141_));
 sg13g2_xor2_1 _2005_ (.B(_1113_),
    .A(_1111_),
    .X(_1144_));
 sg13g2_nand2_1 _2006_ (.Y(_1145_),
    .A(_1143_),
    .B(_1144_));
 sg13g2_and2_1 _2007_ (.A(net377),
    .B(net365),
    .X(_1146_));
 sg13g2_and2_2 _2008_ (.A(net363),
    .B(net361),
    .X(_1147_));
 sg13g2_nand2_1 _2009_ (.Y(_1148_),
    .A(net380),
    .B(net360));
 sg13g2_a22oi_1 _2010_ (.Y(_1149_),
    .B1(net361),
    .B2(net380),
    .A2(net363),
    .A1(net378));
 sg13g2_a21oi_1 _2011_ (.A1(_1061_),
    .A2(_1147_),
    .Y(_1150_),
    .B1(_1149_));
 sg13g2_xor2_1 _2012_ (.B(_1150_),
    .A(_1146_),
    .X(_1151_));
 sg13g2_inv_1 _2013_ (.Y(_1152_),
    .A(_1151_));
 sg13g2_xnor2_1 _2014_ (.Y(_1153_),
    .A(_1143_),
    .B(_1144_));
 sg13g2_o21ai_1 _2015_ (.B1(_1145_),
    .Y(_1154_),
    .A1(_1152_),
    .A2(_1153_));
 sg13g2_xor2_1 _2016_ (.B(_1122_),
    .A(_1117_),
    .X(_1155_));
 sg13g2_nand2_1 _2017_ (.Y(_1156_),
    .A(_1154_),
    .B(_1155_));
 sg13g2_a22oi_1 _2018_ (.Y(_1157_),
    .B1(_1150_),
    .B2(_1146_),
    .A2(_1147_),
    .A1(_1061_));
 sg13g2_xnor2_1 _2019_ (.Y(_1158_),
    .A(_1154_),
    .B(_1155_));
 sg13g2_o21ai_1 _2020_ (.B1(_1156_),
    .Y(_1159_),
    .A1(_1157_),
    .A2(_1158_));
 sg13g2_nand2b_2 _2021_ (.Y(_1160_),
    .B(_1159_),
    .A_N(_1137_));
 sg13g2_nor2_1 _2022_ (.A(_1136_),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_nor3_1 _2023_ (.A(_1131_),
    .B(_1136_),
    .C(_1160_),
    .Y(_1162_));
 sg13g2_xnor2_1 _2024_ (.Y(_1163_),
    .A(_1137_),
    .B(_1159_));
 sg13g2_and2_1 _2025_ (.A(net390),
    .B(net355),
    .X(_1164_));
 sg13g2_nand2_1 _2026_ (.Y(_1165_),
    .A(net388),
    .B(_1164_));
 sg13g2_a21oi_1 _2027_ (.A1(net389),
    .A2(net355),
    .Y(_1166_),
    .B1(net390));
 sg13g2_a21oi_1 _2028_ (.A1(net388),
    .A2(_1164_),
    .Y(_1167_),
    .B1(_1166_));
 sg13g2_nand2_1 _2029_ (.Y(_1168_),
    .A(net386),
    .B(net359));
 sg13g2_o21ai_1 _2030_ (.B1(_1165_),
    .Y(_1169_),
    .A1(_1166_),
    .A2(_1168_));
 sg13g2_xnor2_1 _2031_ (.Y(_1170_),
    .A(_1140_),
    .B(_1142_));
 sg13g2_nand2_1 _2032_ (.Y(_1171_),
    .A(_1169_),
    .B(_1170_));
 sg13g2_nand2_1 _2033_ (.Y(_1172_),
    .A(net378),
    .B(net365));
 sg13g2_nand2_2 _2034_ (.Y(_1173_),
    .A(net382),
    .B(net363));
 sg13g2_nor2_1 _2035_ (.A(_1148_),
    .B(_1173_),
    .Y(_1174_));
 sg13g2_or2_1 _2036_ (.X(_1175_),
    .B(_1173_),
    .A(_1148_));
 sg13g2_a22oi_1 _2037_ (.Y(_1176_),
    .B1(net360),
    .B2(net382),
    .A2(net363),
    .A1(net380));
 sg13g2_nor2_1 _2038_ (.A(_1174_),
    .B(_1176_),
    .Y(_1177_));
 sg13g2_xnor2_1 _2039_ (.Y(_1178_),
    .A(_1172_),
    .B(_1177_));
 sg13g2_inv_1 _2040_ (.Y(_1179_),
    .A(_1178_));
 sg13g2_xnor2_1 _2041_ (.Y(_1180_),
    .A(_1169_),
    .B(_1170_));
 sg13g2_o21ai_1 _2042_ (.B1(_1171_),
    .Y(_1181_),
    .A1(_1179_),
    .A2(_1180_));
 sg13g2_xnor2_1 _2043_ (.Y(_1182_),
    .A(_1151_),
    .B(_1153_));
 sg13g2_nand2_1 _2044_ (.Y(_1183_),
    .A(_1181_),
    .B(_1182_));
 sg13g2_xnor2_1 _2045_ (.Y(_1184_),
    .A(_1181_),
    .B(_1182_));
 sg13g2_o21ai_1 _2046_ (.B1(_1175_),
    .Y(_1185_),
    .A1(_1172_),
    .A2(_1176_));
 sg13g2_nand2_1 _2047_ (.Y(_1186_),
    .A(net376),
    .B(net367));
 sg13g2_nor2_1 _2048_ (.A(_0043_),
    .B(_1186_),
    .Y(_1187_));
 sg13g2_o21ai_1 _2049_ (.B1(net367),
    .Y(_1188_),
    .A1(_0043_),
    .A2(_1186_));
 sg13g2_xnor2_1 _2050_ (.Y(_1189_),
    .A(_1185_),
    .B(_1188_));
 sg13g2_inv_1 _2051_ (.Y(_1190_),
    .A(_1189_));
 sg13g2_o21ai_1 _2052_ (.B1(_1183_),
    .Y(_1191_),
    .A1(_1184_),
    .A2(_1190_));
 sg13g2_xnor2_1 _2053_ (.Y(_1192_),
    .A(_1157_),
    .B(_1158_));
 sg13g2_nor2b_1 _2054_ (.A(_1192_),
    .B_N(_1191_),
    .Y(_1193_));
 sg13g2_a21oi_1 _2055_ (.A1(net367),
    .A2(_1185_),
    .Y(_1194_),
    .B1(_1187_));
 sg13g2_xor2_1 _2056_ (.B(_1192_),
    .A(_1191_),
    .X(_1195_));
 sg13g2_nor2_1 _2057_ (.A(_1194_),
    .B(_1195_),
    .Y(_1196_));
 sg13g2_o21ai_1 _2058_ (.B1(_1163_),
    .Y(_1197_),
    .A1(_1193_),
    .A2(_1196_));
 sg13g2_or2_1 _2059_ (.X(_1198_),
    .B(_1197_),
    .A(_1136_));
 sg13g2_xnor2_1 _2060_ (.Y(_1199_),
    .A(_1136_),
    .B(_1197_));
 sg13g2_a21oi_1 _2061_ (.A1(_1160_),
    .A2(_1199_),
    .Y(_1200_),
    .B1(_1161_));
 sg13g2_xor2_1 _2062_ (.B(_1195_),
    .A(_1194_),
    .X(_1201_));
 sg13g2_and2_2 _2063_ (.A(net392),
    .B(net390),
    .X(_1202_));
 sg13g2_nand2_1 _2064_ (.Y(_0078_),
    .A(net355),
    .B(_1202_));
 sg13g2_nor2_1 _2065_ (.A(net392),
    .B(_1164_),
    .Y(_0079_));
 sg13g2_a21oi_1 _2066_ (.A1(net355),
    .A2(_1202_),
    .Y(_0080_),
    .B1(_0079_));
 sg13g2_nand2_1 _2067_ (.Y(_0081_),
    .A(net388),
    .B(net358));
 sg13g2_o21ai_1 _2068_ (.B1(_0078_),
    .Y(_0082_),
    .A1(_0079_),
    .A2(_0081_));
 sg13g2_xnor2_1 _2069_ (.Y(_0083_),
    .A(_1167_),
    .B(_1168_));
 sg13g2_xnor2_1 _2070_ (.Y(_0084_),
    .A(_0082_),
    .B(_0083_));
 sg13g2_nand2_1 _2071_ (.Y(_0085_),
    .A(net380),
    .B(net365));
 sg13g2_nand2_1 _2072_ (.Y(_0086_),
    .A(net384),
    .B(net360));
 sg13g2_xor2_1 _2073_ (.B(_0086_),
    .A(_1173_),
    .X(_0087_));
 sg13g2_nand2b_1 _2074_ (.Y(_0088_),
    .B(_0087_),
    .A_N(_0085_));
 sg13g2_xnor2_1 _2075_ (.Y(_0089_),
    .A(_0085_),
    .B(_0087_));
 sg13g2_nor2b_1 _2076_ (.A(_0084_),
    .B_N(_0089_),
    .Y(_0090_));
 sg13g2_a21o_1 _2077_ (.A2(_0083_),
    .A1(_0082_),
    .B1(_0090_),
    .X(_0091_));
 sg13g2_xnor2_1 _2078_ (.Y(_0092_),
    .A(_1178_),
    .B(_1180_));
 sg13g2_nand2_1 _2079_ (.Y(_0093_),
    .A(_0091_),
    .B(_0092_));
 sg13g2_nand2_1 _2080_ (.Y(_0094_),
    .A(net379),
    .B(net369));
 sg13g2_nand2_1 _2081_ (.Y(_0095_),
    .A(net378),
    .B(net367));
 sg13g2_nand2_1 _2082_ (.Y(_0096_),
    .A(net376),
    .B(net369));
 sg13g2_xor2_1 _2083_ (.B(_0096_),
    .A(_0095_),
    .X(_0097_));
 sg13g2_nand2_1 _2084_ (.Y(_0098_),
    .A(net371),
    .B(_0097_));
 sg13g2_o21ai_1 _2085_ (.B1(_0098_),
    .Y(_0099_),
    .A1(_0095_),
    .A2(_0096_));
 sg13g2_o21ai_1 _2086_ (.B1(_0088_),
    .Y(_0100_),
    .A1(_1173_),
    .A2(_0086_));
 sg13g2_xor2_1 _2087_ (.B(_1186_),
    .A(_0043_),
    .X(_0101_));
 sg13g2_nand2_1 _2088_ (.Y(_0102_),
    .A(_0100_),
    .B(_0101_));
 sg13g2_xnor2_1 _2089_ (.Y(_0103_),
    .A(_0100_),
    .B(_0101_));
 sg13g2_nand2b_1 _2090_ (.Y(_0104_),
    .B(_0099_),
    .A_N(_0103_));
 sg13g2_xor2_1 _2091_ (.B(_0103_),
    .A(_0099_),
    .X(_0105_));
 sg13g2_xnor2_1 _2092_ (.Y(_0106_),
    .A(_0091_),
    .B(_0092_));
 sg13g2_o21ai_1 _2093_ (.B1(_0093_),
    .Y(_0107_),
    .A1(_0105_),
    .A2(_0106_));
 sg13g2_xnor2_1 _2094_ (.Y(_0108_),
    .A(_1184_),
    .B(_1189_));
 sg13g2_and2_1 _2095_ (.A(_0107_),
    .B(_0108_),
    .X(_0109_));
 sg13g2_nand2_1 _2096_ (.Y(_0110_),
    .A(_0102_),
    .B(_0104_));
 sg13g2_xnor2_1 _2097_ (.Y(_0111_),
    .A(_0107_),
    .B(_0108_));
 sg13g2_nor2b_1 _2098_ (.A(_0111_),
    .B_N(_0110_),
    .Y(_0112_));
 sg13g2_o21ai_1 _2099_ (.B1(_1201_),
    .Y(_0113_),
    .A1(_0109_),
    .A2(_0112_));
 sg13g2_or3_1 _2100_ (.A(_1163_),
    .B(_1193_),
    .C(_1196_),
    .X(_0114_));
 sg13g2_nand2_1 _2101_ (.Y(_0115_),
    .A(_1197_),
    .B(_0114_));
 sg13g2_nor2_1 _2102_ (.A(_0113_),
    .B(_0115_),
    .Y(_0116_));
 sg13g2_xor2_1 _2103_ (.B(_0111_),
    .A(_0110_),
    .X(_0117_));
 sg13g2_nand2_1 _2104_ (.Y(_0118_),
    .A(net392),
    .B(net358));
 sg13g2_and3_1 _2105_ (.X(_0119_),
    .A(net358),
    .B(net355),
    .C(_1202_));
 sg13g2_nor2_1 _2106_ (.A(_0080_),
    .B(_0119_),
    .Y(_0120_));
 sg13g2_xnor2_1 _2107_ (.Y(_0121_),
    .A(_0081_),
    .B(_0120_));
 sg13g2_nand2_1 _2108_ (.Y(_0122_),
    .A(net382),
    .B(net365));
 sg13g2_nand2_1 _2109_ (.Y(_0123_),
    .A(net384),
    .B(net364));
 sg13g2_nand2_1 _2110_ (.Y(_0124_),
    .A(net386),
    .B(net361));
 sg13g2_or2_1 _2111_ (.X(_0125_),
    .B(_0124_),
    .A(_0123_));
 sg13g2_xnor2_1 _2112_ (.Y(_0126_),
    .A(_0123_),
    .B(_0124_));
 sg13g2_xor2_1 _2113_ (.B(_0126_),
    .A(_0122_),
    .X(_0127_));
 sg13g2_nor2b_1 _2114_ (.A(_0121_),
    .B_N(_0127_),
    .Y(_0128_));
 sg13g2_a21o_1 _2115_ (.A2(_0119_),
    .A1(net388),
    .B1(_0128_),
    .X(_0129_));
 sg13g2_xnor2_1 _2116_ (.Y(_0130_),
    .A(_0084_),
    .B(_0089_));
 sg13g2_nand2_1 _2117_ (.Y(_0131_),
    .A(_0129_),
    .B(_0130_));
 sg13g2_xnor2_1 _2118_ (.Y(_0132_),
    .A(_0129_),
    .B(_0130_));
 sg13g2_nand2_1 _2119_ (.Y(_0133_),
    .A(net370),
    .B(net368));
 sg13g2_inv_2 _2120_ (.Y(_0134_),
    .A(_0133_));
 sg13g2_nand2_1 _2121_ (.Y(_0135_),
    .A(net381),
    .B(net367));
 sg13g2_xnor2_1 _2122_ (.Y(_0136_),
    .A(_0094_),
    .B(_0135_));
 sg13g2_nand2_1 _2123_ (.Y(_0137_),
    .A(net376),
    .B(net371));
 sg13g2_nor2_1 _2124_ (.A(_0136_),
    .B(_0137_),
    .Y(_0138_));
 sg13g2_a21oi_2 _2125_ (.B1(_0138_),
    .Y(_0139_),
    .A2(_0134_),
    .A1(_1061_));
 sg13g2_o21ai_1 _2126_ (.B1(_0125_),
    .Y(_0140_),
    .A1(_0122_),
    .A2(_0126_));
 sg13g2_xnor2_1 _2127_ (.Y(_0141_),
    .A(net371),
    .B(_0097_));
 sg13g2_nand2b_1 _2128_ (.Y(_0142_),
    .B(_0140_),
    .A_N(_0141_));
 sg13g2_xor2_1 _2129_ (.B(_0141_),
    .A(_0140_),
    .X(_0143_));
 sg13g2_xnor2_1 _2130_ (.Y(_0144_),
    .A(_0139_),
    .B(_0143_));
 sg13g2_o21ai_1 _2131_ (.B1(_0131_),
    .Y(_0145_),
    .A1(_0132_),
    .A2(_0144_));
 sg13g2_xor2_1 _2132_ (.B(_0106_),
    .A(_0105_),
    .X(_0146_));
 sg13g2_nand2_1 _2133_ (.Y(_0147_),
    .A(_0145_),
    .B(_0146_));
 sg13g2_o21ai_1 _2134_ (.B1(_0142_),
    .Y(_0148_),
    .A1(_0139_),
    .A2(_0143_));
 sg13g2_xor2_1 _2135_ (.B(_0146_),
    .A(_0145_),
    .X(_0149_));
 sg13g2_nand2_1 _2136_ (.Y(_0150_),
    .A(_0148_),
    .B(_0149_));
 sg13g2_a21oi_2 _2137_ (.B1(_0117_),
    .Y(_0151_),
    .A2(_0150_),
    .A1(_0147_));
 sg13g2_or3_1 _2138_ (.A(_1201_),
    .B(_0109_),
    .C(_0112_),
    .X(_0152_));
 sg13g2_and2_1 _2139_ (.A(_0113_),
    .B(_0152_),
    .X(_0153_));
 sg13g2_nand2_1 _2140_ (.Y(_0154_),
    .A(_0151_),
    .B(_0153_));
 sg13g2_xnor2_1 _2141_ (.Y(_0155_),
    .A(_0148_),
    .B(_0149_));
 sg13g2_and2_1 _2142_ (.A(net384),
    .B(net366),
    .X(_0156_));
 sg13g2_a22oi_1 _2143_ (.Y(_0157_),
    .B1(net361),
    .B2(net388),
    .A2(net364),
    .A1(net386));
 sg13g2_a21oi_1 _2144_ (.A1(_1138_),
    .A2(_1147_),
    .Y(_0158_),
    .B1(_0157_));
 sg13g2_xor2_1 _2145_ (.B(_0158_),
    .A(_0156_),
    .X(_0159_));
 sg13g2_a22oi_1 _2146_ (.Y(_0160_),
    .B1(net355),
    .B2(net392),
    .A2(net358),
    .A1(net390));
 sg13g2_nor2_1 _2147_ (.A(_0119_),
    .B(_0160_),
    .Y(_0161_));
 sg13g2_nand2_1 _2148_ (.Y(_0162_),
    .A(_0159_),
    .B(_0161_));
 sg13g2_xnor2_1 _2149_ (.Y(_0163_),
    .A(_0121_),
    .B(_0127_));
 sg13g2_nor2b_1 _2150_ (.A(_0162_),
    .B_N(_0163_),
    .Y(_0164_));
 sg13g2_xnor2_1 _2151_ (.Y(_0165_),
    .A(_0162_),
    .B(_0163_));
 sg13g2_nand2_1 _2152_ (.Y(_0166_),
    .A(net382),
    .B(net369));
 sg13g2_nor2_1 _2153_ (.A(_0135_),
    .B(_0166_),
    .Y(_0167_));
 sg13g2_nand2_1 _2154_ (.Y(_0168_),
    .A(net379),
    .B(net371));
 sg13g2_a22oi_1 _2155_ (.Y(_0169_),
    .B1(net367),
    .B2(net382),
    .A2(net369),
    .A1(net381));
 sg13g2_nor3_1 _2156_ (.A(_0167_),
    .B(_0168_),
    .C(_0169_),
    .Y(_0170_));
 sg13g2_or2_1 _2157_ (.X(_0171_),
    .B(_0170_),
    .A(_0167_));
 sg13g2_a22oi_1 _2158_ (.Y(_0172_),
    .B1(_0156_),
    .B2(_0158_),
    .A2(_1147_),
    .A1(_1138_));
 sg13g2_xnor2_1 _2159_ (.Y(_0173_),
    .A(_0136_),
    .B(_0137_));
 sg13g2_xor2_1 _2160_ (.B(_0173_),
    .A(_0172_),
    .X(_0174_));
 sg13g2_nand2_1 _2161_ (.Y(_0175_),
    .A(_0171_),
    .B(_0174_));
 sg13g2_xnor2_1 _2162_ (.Y(_0176_),
    .A(_0171_),
    .B(_0174_));
 sg13g2_inv_1 _2163_ (.Y(_0177_),
    .A(_0176_));
 sg13g2_a21oi_1 _2164_ (.A1(_0165_),
    .A2(_0177_),
    .Y(_0178_),
    .B1(_0164_));
 sg13g2_xor2_1 _2165_ (.B(_0144_),
    .A(_0132_),
    .X(_0179_));
 sg13g2_nand2b_1 _2166_ (.Y(_0180_),
    .B(_0179_),
    .A_N(_0178_));
 sg13g2_o21ai_1 _2167_ (.B1(_0175_),
    .Y(_0181_),
    .A1(_0172_),
    .A2(_0173_));
 sg13g2_xnor2_1 _2168_ (.Y(_0182_),
    .A(_0178_),
    .B(_0179_));
 sg13g2_nand2_1 _2169_ (.Y(_0183_),
    .A(_0181_),
    .B(_0182_));
 sg13g2_a21o_1 _2170_ (.A2(_0183_),
    .A1(_0180_),
    .B1(_0155_),
    .X(_0184_));
 sg13g2_nand3_1 _2171_ (.B(_0147_),
    .C(_0150_),
    .A(_0117_),
    .Y(_0185_));
 sg13g2_nand2b_1 _2172_ (.Y(_0186_),
    .B(_0185_),
    .A_N(_0151_));
 sg13g2_nor2_1 _2173_ (.A(_0184_),
    .B(_0186_),
    .Y(_0187_));
 sg13g2_xnor2_1 _2174_ (.Y(_0188_),
    .A(_0181_),
    .B(_0182_));
 sg13g2_nand2_1 _2175_ (.Y(_0189_),
    .A(net386),
    .B(net366));
 sg13g2_nand2_1 _2176_ (.Y(_0190_),
    .A(net388),
    .B(net363));
 sg13g2_nand2_1 _2177_ (.Y(_0191_),
    .A(net390),
    .B(net360));
 sg13g2_or2_1 _2178_ (.X(_0192_),
    .B(_0191_),
    .A(_0190_));
 sg13g2_xor2_1 _2179_ (.B(_0191_),
    .A(_0190_),
    .X(_0193_));
 sg13g2_nand2b_1 _2180_ (.Y(_0194_),
    .B(_0193_),
    .A_N(_0189_));
 sg13g2_xnor2_1 _2181_ (.Y(_0195_),
    .A(_0189_),
    .B(_0193_));
 sg13g2_nand2b_1 _2182_ (.Y(_0196_),
    .B(_0195_),
    .A_N(_0118_));
 sg13g2_inv_1 _2183_ (.Y(_0197_),
    .A(_0196_));
 sg13g2_xor2_1 _2184_ (.B(_0161_),
    .A(_0159_),
    .X(_0198_));
 sg13g2_xnor2_1 _2185_ (.Y(_0199_),
    .A(_0196_),
    .B(_0198_));
 sg13g2_inv_1 _2186_ (.Y(_0200_),
    .A(_0199_));
 sg13g2_nand2_2 _2187_ (.Y(_0201_),
    .A(net384),
    .B(net367));
 sg13g2_nand2_1 _2188_ (.Y(_0202_),
    .A(net380),
    .B(net371));
 sg13g2_xor2_1 _2189_ (.B(_0201_),
    .A(_0166_),
    .X(_0203_));
 sg13g2_nand2b_1 _2190_ (.Y(_0204_),
    .B(_0203_),
    .A_N(_0202_));
 sg13g2_o21ai_1 _2191_ (.B1(_0204_),
    .Y(_0205_),
    .A1(_0166_),
    .A2(_0201_));
 sg13g2_and2_1 _2192_ (.A(_0192_),
    .B(_0194_),
    .X(_0206_));
 sg13g2_o21ai_1 _2193_ (.B1(_0168_),
    .Y(_0207_),
    .A1(_0167_),
    .A2(_0169_));
 sg13g2_nor2b_1 _2194_ (.A(_0170_),
    .B_N(_0207_),
    .Y(_0208_));
 sg13g2_nor2b_1 _2195_ (.A(_0206_),
    .B_N(_0208_),
    .Y(_0209_));
 sg13g2_xnor2_1 _2196_ (.Y(_0210_),
    .A(_0206_),
    .B(_0208_));
 sg13g2_xnor2_1 _2197_ (.Y(_0211_),
    .A(_0205_),
    .B(_0210_));
 sg13g2_nor2_1 _2198_ (.A(_0200_),
    .B(_0211_),
    .Y(_0212_));
 sg13g2_a21oi_1 _2199_ (.A1(_0197_),
    .A2(_0198_),
    .Y(_0213_),
    .B1(_0212_));
 sg13g2_xor2_1 _2200_ (.B(_0176_),
    .A(_0165_),
    .X(_0214_));
 sg13g2_nor2_1 _2201_ (.A(_0213_),
    .B(_0214_),
    .Y(_0215_));
 sg13g2_a21o_1 _2202_ (.A2(_0210_),
    .A1(_0205_),
    .B1(_0209_),
    .X(_0216_));
 sg13g2_xor2_1 _2203_ (.B(_0214_),
    .A(_0213_),
    .X(_0217_));
 sg13g2_a21oi_2 _2204_ (.B1(_0215_),
    .Y(_0218_),
    .A2(_0217_),
    .A1(_0216_));
 sg13g2_nor2_1 _2205_ (.A(_0188_),
    .B(_0218_),
    .Y(_0219_));
 sg13g2_nand3_1 _2206_ (.B(_0180_),
    .C(_0183_),
    .A(_0155_),
    .Y(_0220_));
 sg13g2_nand2_1 _2207_ (.Y(_0221_),
    .A(_0184_),
    .B(_0220_));
 sg13g2_nand3_1 _2208_ (.B(_0219_),
    .C(_0220_),
    .A(_0184_),
    .Y(_0222_));
 sg13g2_xnor2_1 _2209_ (.Y(_0223_),
    .A(_0188_),
    .B(_0218_));
 sg13g2_nor3_1 _2210_ (.A(_0474_),
    .B(_0476_),
    .C(_0201_),
    .Y(_0224_));
 sg13g2_nand2_1 _2211_ (.Y(_0225_),
    .A(net382),
    .B(net371));
 sg13g2_a22oi_1 _2212_ (.Y(_0226_),
    .B1(net367),
    .B2(net386),
    .A2(net369),
    .A1(net384));
 sg13g2_nor3_1 _2213_ (.A(_0224_),
    .B(_0225_),
    .C(_0226_),
    .Y(_0227_));
 sg13g2_or2_1 _2214_ (.X(_0228_),
    .B(_0227_),
    .A(_0224_));
 sg13g2_and2_1 _2215_ (.A(net388),
    .B(net366),
    .X(_0229_));
 sg13g2_a22oi_1 _2216_ (.Y(_0230_),
    .B1(net360),
    .B2(net392),
    .A2(net363),
    .A1(net390));
 sg13g2_a21oi_1 _2217_ (.A1(_1147_),
    .A2(_1202_),
    .Y(_0231_),
    .B1(_0230_));
 sg13g2_a22oi_1 _2218_ (.Y(_0232_),
    .B1(_0229_),
    .B2(_0231_),
    .A2(_1202_),
    .A1(_1147_));
 sg13g2_xnor2_1 _2219_ (.Y(_0233_),
    .A(_0202_),
    .B(_0203_));
 sg13g2_nor2b_1 _2220_ (.A(_0232_),
    .B_N(_0233_),
    .Y(_0234_));
 sg13g2_xnor2_1 _2221_ (.Y(_0235_),
    .A(_0232_),
    .B(_0233_));
 sg13g2_xnor2_1 _2222_ (.Y(_0236_),
    .A(_0228_),
    .B(_0235_));
 sg13g2_xnor2_1 _2223_ (.Y(_0237_),
    .A(_0118_),
    .B(_0195_));
 sg13g2_nand2b_1 _2224_ (.Y(_0238_),
    .B(_0237_),
    .A_N(_0236_));
 sg13g2_xor2_1 _2225_ (.B(_0211_),
    .A(_0199_),
    .X(_0239_));
 sg13g2_nor2_1 _2226_ (.A(_0238_),
    .B(_0239_),
    .Y(_0240_));
 sg13g2_a21o_1 _2227_ (.A2(_0235_),
    .A1(_0228_),
    .B1(_0234_),
    .X(_0241_));
 sg13g2_xor2_1 _2228_ (.B(_0239_),
    .A(_0238_),
    .X(_0242_));
 sg13g2_a21oi_1 _2229_ (.A1(_0241_),
    .A2(_0242_),
    .Y(_0243_),
    .B1(_0240_));
 sg13g2_xnor2_1 _2230_ (.Y(_0244_),
    .A(_0216_),
    .B(_0217_));
 sg13g2_nor2_1 _2231_ (.A(_0243_),
    .B(_0244_),
    .Y(_0245_));
 sg13g2_xor2_1 _2232_ (.B(_0244_),
    .A(_0243_),
    .X(_0246_));
 sg13g2_a21oi_2 _2233_ (.B1(_0245_),
    .Y(_0247_),
    .A2(_0246_),
    .A1(net373));
 sg13g2_nor2_1 _2234_ (.A(_0223_),
    .B(_0247_),
    .Y(_0248_));
 sg13g2_nor3_1 _2235_ (.A(_0473_),
    .B(_0474_),
    .C(_0133_),
    .Y(_0249_));
 sg13g2_nand2_1 _2236_ (.Y(_0250_),
    .A(net385),
    .B(net372));
 sg13g2_a22oi_1 _2237_ (.Y(_0251_),
    .B1(net368),
    .B2(net389),
    .A2(net370),
    .A1(net386));
 sg13g2_or3_1 _2238_ (.A(_0249_),
    .B(_0250_),
    .C(_0251_),
    .X(_0252_));
 sg13g2_nand2b_1 _2239_ (.Y(_0253_),
    .B(_0252_),
    .A_N(_0249_));
 sg13g2_nand2_1 _2240_ (.Y(_0254_),
    .A(\MAC.a[0] ),
    .B(net366));
 sg13g2_and4_1 _2241_ (.A(net392),
    .B(net390),
    .C(net365),
    .D(net363),
    .X(_0255_));
 sg13g2_o21ai_1 _2242_ (.B1(_0225_),
    .Y(_0256_),
    .A1(_0224_),
    .A2(_0226_));
 sg13g2_nor2b_1 _2243_ (.A(_0227_),
    .B_N(_0256_),
    .Y(_0257_));
 sg13g2_and2_1 _2244_ (.A(_0255_),
    .B(_0257_),
    .X(_0258_));
 sg13g2_xor2_1 _2245_ (.B(_0257_),
    .A(_0255_),
    .X(_0259_));
 sg13g2_xor2_1 _2246_ (.B(_0259_),
    .A(_0253_),
    .X(_0260_));
 sg13g2_xor2_1 _2247_ (.B(_0231_),
    .A(_0229_),
    .X(_0261_));
 sg13g2_nand2_1 _2248_ (.Y(_0262_),
    .A(_0260_),
    .B(_0261_));
 sg13g2_xor2_1 _2249_ (.B(_0237_),
    .A(_0236_),
    .X(_0263_));
 sg13g2_nor2_1 _2250_ (.A(_0262_),
    .B(_0263_),
    .Y(_0264_));
 sg13g2_a21o_1 _2251_ (.A2(_0259_),
    .A1(_0253_),
    .B1(_0258_),
    .X(_0265_));
 sg13g2_xor2_1 _2252_ (.B(_0263_),
    .A(_0262_),
    .X(_0266_));
 sg13g2_a21oi_1 _2253_ (.A1(_0265_),
    .A2(_0266_),
    .Y(_0267_),
    .B1(_0264_));
 sg13g2_xnor2_1 _2254_ (.Y(_0268_),
    .A(_0241_),
    .B(_0242_));
 sg13g2_nor2_1 _2255_ (.A(_0267_),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_and2_1 _2256_ (.A(net376),
    .B(net373),
    .X(_0270_));
 sg13g2_xor2_1 _2257_ (.B(_0268_),
    .A(_0267_),
    .X(_0271_));
 sg13g2_a21oi_1 _2258_ (.A1(_0270_),
    .A2(_0271_),
    .Y(_0272_),
    .B1(_0269_));
 sg13g2_xnor2_1 _2259_ (.Y(_0273_),
    .A(net373),
    .B(_0246_));
 sg13g2_or2_1 _2260_ (.X(_0274_),
    .B(_0273_),
    .A(_0272_));
 sg13g2_xnor2_1 _2261_ (.Y(_0275_),
    .A(_0272_),
    .B(_0273_));
 sg13g2_xor2_1 _2262_ (.B(_0271_),
    .A(_0270_),
    .X(_0276_));
 sg13g2_xor2_1 _2263_ (.B(_0261_),
    .A(_0260_),
    .X(_0277_));
 sg13g2_and4_1 _2264_ (.A(net391),
    .B(net389),
    .C(net370),
    .D(net368),
    .X(_0278_));
 sg13g2_nand2_1 _2265_ (.Y(_0279_),
    .A(net387),
    .B(net372));
 sg13g2_a22oi_1 _2266_ (.Y(_0280_),
    .B1(net368),
    .B2(net391),
    .A2(net370),
    .A1(net389));
 sg13g2_or3_1 _2267_ (.A(_0278_),
    .B(_0279_),
    .C(_0280_),
    .X(_0281_));
 sg13g2_nand2b_1 _2268_ (.Y(_0282_),
    .B(_0281_),
    .A_N(_0278_));
 sg13g2_o21ai_1 _2269_ (.B1(_0250_),
    .Y(_0283_),
    .A1(_0249_),
    .A2(_0251_));
 sg13g2_nand2_1 _2270_ (.Y(_0284_),
    .A(_0252_),
    .B(_0283_));
 sg13g2_nor2b_1 _2271_ (.A(_0284_),
    .B_N(_0282_),
    .Y(_0285_));
 sg13g2_a22oi_1 _2272_ (.Y(_0286_),
    .B1(net364),
    .B2(net392),
    .A2(net365),
    .A1(net390));
 sg13g2_nor2_1 _2273_ (.A(_0255_),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_xnor2_1 _2274_ (.Y(_0288_),
    .A(_0282_),
    .B(_0284_));
 sg13g2_a21o_1 _2275_ (.A2(_0288_),
    .A1(_0287_),
    .B1(_0285_),
    .X(_0289_));
 sg13g2_nand2_1 _2276_ (.Y(_0290_),
    .A(_0277_),
    .B(_0289_));
 sg13g2_xnor2_1 _2277_ (.Y(_0291_),
    .A(_0265_),
    .B(_0266_));
 sg13g2_nand2_1 _2278_ (.Y(_0292_),
    .A(net379),
    .B(net373));
 sg13g2_xor2_1 _2279_ (.B(_0291_),
    .A(_0290_),
    .X(_0293_));
 sg13g2_nand2b_1 _2280_ (.Y(_0294_),
    .B(_0293_),
    .A_N(_0292_));
 sg13g2_o21ai_1 _2281_ (.B1(_0294_),
    .Y(_0295_),
    .A1(_0290_),
    .A2(_0291_));
 sg13g2_nor2_1 _2282_ (.A(_0276_),
    .B(_0295_),
    .Y(_0296_));
 sg13g2_nand2_1 _2283_ (.Y(_0297_),
    .A(_0276_),
    .B(_0295_));
 sg13g2_xor2_1 _2284_ (.B(_0289_),
    .A(_0277_),
    .X(_0298_));
 sg13g2_xor2_1 _2285_ (.B(_0288_),
    .A(_0287_),
    .X(_0299_));
 sg13g2_and3_1 _2286_ (.X(_0300_),
    .A(net370),
    .B(net368),
    .C(_1202_));
 sg13g2_nand2_1 _2287_ (.Y(_0301_),
    .A(net389),
    .B(net372));
 sg13g2_a22oi_1 _2288_ (.Y(_0302_),
    .B1(net368),
    .B2(\MAC.a[0] ),
    .A2(net369),
    .A1(net391));
 sg13g2_nor3_1 _2289_ (.A(_0300_),
    .B(_0301_),
    .C(_0302_),
    .Y(_0303_));
 sg13g2_or2_1 _2290_ (.X(_0304_),
    .B(_0303_),
    .A(_0300_));
 sg13g2_o21ai_1 _2291_ (.B1(_0279_),
    .Y(_0305_),
    .A1(_0278_),
    .A2(_0280_));
 sg13g2_nand2_1 _2292_ (.Y(_0306_),
    .A(_0281_),
    .B(_0305_));
 sg13g2_nand2b_1 _2293_ (.Y(_0307_),
    .B(_0304_),
    .A_N(_0306_));
 sg13g2_xnor2_1 _2294_ (.Y(_0308_),
    .A(_0304_),
    .B(_0306_));
 sg13g2_nand2b_1 _2295_ (.Y(_0309_),
    .B(_0308_),
    .A_N(_0254_));
 sg13g2_nand2_1 _2296_ (.Y(_0310_),
    .A(_0307_),
    .B(_0309_));
 sg13g2_nand2_1 _2297_ (.Y(_0311_),
    .A(_0299_),
    .B(_0310_));
 sg13g2_inv_1 _2298_ (.Y(_0312_),
    .A(_0311_));
 sg13g2_nand2_1 _2299_ (.Y(_0313_),
    .A(_0298_),
    .B(_0312_));
 sg13g2_nand2_1 _2300_ (.Y(_0314_),
    .A(net380),
    .B(net373));
 sg13g2_xnor2_1 _2301_ (.Y(_0315_),
    .A(_0298_),
    .B(_0312_));
 sg13g2_o21ai_1 _2302_ (.B1(_0313_),
    .Y(_0316_),
    .A1(_0314_),
    .A2(_0315_));
 sg13g2_xnor2_1 _2303_ (.Y(_0317_),
    .A(_0292_),
    .B(_0293_));
 sg13g2_nor2_1 _2304_ (.A(_0316_),
    .B(_0317_),
    .Y(_0318_));
 sg13g2_and2_1 _2305_ (.A(\MAC.a[0] ),
    .B(net369),
    .X(_0319_));
 sg13g2_nand3_1 _2306_ (.B(net372),
    .C(_0319_),
    .A(net391),
    .Y(_0320_));
 sg13g2_o21ai_1 _2307_ (.B1(_0301_),
    .Y(_0321_),
    .A1(_0300_),
    .A2(_0302_));
 sg13g2_nor2b_1 _2308_ (.A(_0303_),
    .B_N(_0321_),
    .Y(_0322_));
 sg13g2_nand2b_1 _2309_ (.Y(_0323_),
    .B(_0322_),
    .A_N(_0320_));
 sg13g2_xnor2_1 _2310_ (.Y(_0324_),
    .A(_0254_),
    .B(_0308_));
 sg13g2_nand2b_1 _2311_ (.Y(_0325_),
    .B(_0324_),
    .A_N(_0323_));
 sg13g2_xnor2_1 _2312_ (.Y(_0326_),
    .A(_0299_),
    .B(_0310_));
 sg13g2_nor2_1 _2313_ (.A(_0325_),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_and2_1 _2314_ (.A(net383),
    .B(net374),
    .X(_0328_));
 sg13g2_xor2_1 _2315_ (.B(_0326_),
    .A(_0325_),
    .X(_0329_));
 sg13g2_a21oi_1 _2316_ (.A1(_0328_),
    .A2(_0329_),
    .Y(_0330_),
    .B1(_0327_));
 sg13g2_xnor2_1 _2317_ (.Y(_0331_),
    .A(_0323_),
    .B(_0324_));
 sg13g2_a21o_1 _2318_ (.A2(net371),
    .A1(net391),
    .B1(_0319_),
    .X(_0332_));
 sg13g2_nand2_1 _2319_ (.Y(_0333_),
    .A(_0320_),
    .B(_0332_));
 sg13g2_xor2_1 _2320_ (.B(_0322_),
    .A(_0320_),
    .X(_0334_));
 sg13g2_and2_1 _2321_ (.A(_0474_),
    .B(_0334_),
    .X(_0335_));
 sg13g2_nor4_1 _2322_ (.A(_0473_),
    .B(_0475_),
    .C(_0333_),
    .D(_0335_),
    .Y(_0336_));
 sg13g2_nor3_1 _2323_ (.A(_0474_),
    .B(_0475_),
    .C(_0334_),
    .Y(_0337_));
 sg13g2_nand3_1 _2324_ (.B(net371),
    .C(_1202_),
    .A(net374),
    .Y(_0338_));
 sg13g2_xnor2_1 _2325_ (.Y(_0339_),
    .A(_0473_),
    .B(_0333_));
 sg13g2_nor3_1 _2326_ (.A(_0306_),
    .B(_0338_),
    .C(_0339_),
    .Y(_0340_));
 sg13g2_nor3_1 _2327_ (.A(_0336_),
    .B(_0337_),
    .C(_0340_),
    .Y(_0341_));
 sg13g2_nand3_1 _2328_ (.B(net373),
    .C(_0331_),
    .A(net384),
    .Y(_0342_));
 sg13g2_a21oi_1 _2329_ (.A1(net384),
    .A2(net373),
    .Y(_0343_),
    .B1(_0331_));
 sg13g2_a221oi_1 _2330_ (.B2(_0342_),
    .C1(_0343_),
    .B1(_0341_),
    .A1(_0328_),
    .Y(_0344_),
    .A2(_0329_));
 sg13g2_o21ai_1 _2331_ (.B1(_0344_),
    .Y(_0345_),
    .A1(_0328_),
    .A2(_0329_));
 sg13g2_xnor2_1 _2332_ (.Y(_0346_),
    .A(_0314_),
    .B(_0315_));
 sg13g2_nand2_1 _2333_ (.Y(_0347_),
    .A(_0330_),
    .B(_0346_));
 sg13g2_o21ai_1 _2334_ (.B1(_0345_),
    .Y(_0348_),
    .A1(_0330_),
    .A2(_0346_));
 sg13g2_a22oi_1 _2335_ (.Y(_0349_),
    .B1(_0347_),
    .B2(_0348_),
    .A2(_0317_),
    .A1(_0316_));
 sg13g2_or3_1 _2336_ (.A(_0296_),
    .B(_0318_),
    .C(_0349_),
    .X(_0350_));
 sg13g2_a21o_1 _2337_ (.A2(_0350_),
    .A1(_0297_),
    .B1(_0275_),
    .X(_0351_));
 sg13g2_xnor2_1 _2338_ (.Y(_0352_),
    .A(_0223_),
    .B(_0247_));
 sg13g2_a21oi_1 _2339_ (.A1(_0274_),
    .A2(_0351_),
    .Y(_0353_),
    .B1(_0352_));
 sg13g2_xnor2_1 _2340_ (.Y(_0354_),
    .A(_0219_),
    .B(_0221_));
 sg13g2_o21ai_1 _2341_ (.B1(_0354_),
    .Y(_0355_),
    .A1(_0248_),
    .A2(_0353_));
 sg13g2_xnor2_1 _2342_ (.Y(_0356_),
    .A(_0184_),
    .B(_0186_));
 sg13g2_a21oi_1 _2343_ (.A1(_0222_),
    .A2(_0355_),
    .Y(_0357_),
    .B1(_0356_));
 sg13g2_nor2_1 _2344_ (.A(_0187_),
    .B(_0357_),
    .Y(_0358_));
 sg13g2_xnor2_1 _2345_ (.Y(_0359_),
    .A(_0151_),
    .B(_0153_));
 sg13g2_o21ai_1 _2346_ (.B1(_0154_),
    .Y(_0360_),
    .A1(_0358_),
    .A2(_0359_));
 sg13g2_xor2_1 _2347_ (.B(_0115_),
    .A(_0113_),
    .X(_0361_));
 sg13g2_and2_1 _2348_ (.A(_0360_),
    .B(_0361_),
    .X(_0362_));
 sg13g2_o21ai_1 _2349_ (.B1(_1200_),
    .Y(_0363_),
    .A1(_0116_),
    .A2(_0362_));
 sg13g2_o21ai_1 _2350_ (.B1(_1130_),
    .Y(_0364_),
    .A1(_1136_),
    .A2(_1160_));
 sg13g2_xor2_1 _2351_ (.B(_0364_),
    .A(_1131_),
    .X(_0365_));
 sg13g2_a21oi_1 _2352_ (.A1(_1198_),
    .A2(_0363_),
    .Y(_0366_),
    .B1(_0365_));
 sg13g2_o21ai_1 _2353_ (.B1(_1135_),
    .Y(_0367_),
    .A1(_1162_),
    .A2(_0366_));
 sg13g2_o21ai_1 _2354_ (.B1(_0367_),
    .Y(_0368_),
    .A1(_1132_),
    .A2(_1134_));
 sg13g2_nor2_1 _2355_ (.A(_1108_),
    .B(_0368_),
    .Y(_0369_));
 sg13g2_xor2_1 _2356_ (.B(_1085_),
    .A(_1060_),
    .X(_0370_));
 sg13g2_nor3_1 _2357_ (.A(_1086_),
    .B(_1108_),
    .C(_0368_),
    .Y(_0371_));
 sg13g2_nand3_1 _2358_ (.B(_0351_),
    .C(_0352_),
    .A(_0274_),
    .Y(_0372_));
 sg13g2_nand2b_1 _2359_ (.Y(_0373_),
    .B(_0372_),
    .A_N(_0353_));
 sg13g2_nor2_1 _2360_ (.A(net313),
    .B(_0373_),
    .Y(_0374_));
 sg13g2_nand3_1 _2361_ (.B(_0297_),
    .C(_0350_),
    .A(_0275_),
    .Y(_0375_));
 sg13g2_and3_1 _2362_ (.X(_0376_),
    .A(_0351_),
    .B(net313),
    .C(_0375_));
 sg13g2_o21ai_1 _2363_ (.B1(net339),
    .Y(_0377_),
    .A1(_0374_),
    .A2(_0376_));
 sg13g2_xor2_1 _2364_ (.B(_1032_),
    .A(_1031_),
    .X(_0378_));
 sg13g2_nand3_1 _2365_ (.B(_1027_),
    .C(_1028_),
    .A(_1024_),
    .Y(_0379_));
 sg13g2_nand2b_1 _2366_ (.Y(_0380_),
    .B(_0379_),
    .A_N(_1029_));
 sg13g2_xor2_1 _2367_ (.B(_0380_),
    .A(_1037_),
    .X(_0381_));
 sg13g2_xor2_1 _2368_ (.B(_1026_),
    .A(_1025_),
    .X(_0382_));
 sg13g2_xnor2_1 _2369_ (.Y(_0383_),
    .A(_1023_),
    .B(_1030_));
 sg13g2_nor3_1 _2370_ (.A(_1036_),
    .B(_0382_),
    .C(_0383_),
    .Y(_0384_));
 sg13g2_nand3_1 _2371_ (.B(_0381_),
    .C(_0384_),
    .A(_0378_),
    .Y(_0385_));
 sg13g2_nor3_1 _2372_ (.A(_1035_),
    .B(_1040_),
    .C(_0385_),
    .Y(_0386_));
 sg13g2_nand4_1 _2373_ (.B(_1089_),
    .C(_1138_),
    .A(_1061_),
    .Y(_0387_),
    .D(_1202_));
 sg13g2_nand4_1 _2374_ (.B(\MAC.a[13] ),
    .C(net377),
    .A(\MAC.a[14] ),
    .Y(_0388_),
    .D(\MAC.a[15] ));
 sg13g2_nand4_1 _2375_ (.B(\MAC.a[9] ),
    .C(\MAC.a[12] ),
    .A(\MAC.a[10] ),
    .Y(_0389_),
    .D(\MAC.a[11] ));
 sg13g2_nor3_1 _2376_ (.A(_0387_),
    .B(_0388_),
    .C(_0389_),
    .Y(_0390_));
 sg13g2_nand4_1 _2377_ (.B(\MAC.b[9] ),
    .C(net373),
    .A(\MAC.b[10] ),
    .Y(_0391_),
    .D(net372));
 sg13g2_nand2_1 _2378_ (.Y(_0392_),
    .A(_1147_),
    .B(_0134_));
 sg13g2_nand4_1 _2379_ (.B(\MAC.b[11] ),
    .C(\MAC.b[14] ),
    .A(\MAC.b[12] ),
    .Y(_0393_),
    .D(\MAC.b[13] ));
 sg13g2_nand4_1 _2380_ (.B(net359),
    .C(net357),
    .A(net366),
    .Y(_0394_),
    .D(\MAC.b[15] ));
 sg13g2_nor4_1 _2381_ (.A(_0391_),
    .B(_0392_),
    .C(_0393_),
    .D(_0394_),
    .Y(_0395_));
 sg13g2_nor3_2 _2382_ (.A(_0386_),
    .B(_0390_),
    .C(_0395_),
    .Y(_0396_));
 sg13g2_a21oi_1 _2383_ (.A1(_0377_),
    .A2(_0396_),
    .Y(\MAC.mul.c_mul1[0] ),
    .B1(_1045_));
 sg13g2_and2_1 _2384_ (.A(_1042_),
    .B(_0396_),
    .X(_0397_));
 sg13g2_or3_1 _2385_ (.A(_0248_),
    .B(_0353_),
    .C(_0354_),
    .X(_0398_));
 sg13g2_and2_1 _2386_ (.A(_0355_),
    .B(_0398_),
    .X(_0399_));
 sg13g2_o21ai_1 _2387_ (.B1(net339),
    .Y(_0400_),
    .A1(net311),
    .A2(_0399_));
 sg13g2_a21o_1 _2388_ (.A2(_0373_),
    .A1(net312),
    .B1(_0400_),
    .X(_0401_));
 sg13g2_a21oi_1 _2389_ (.A1(net321),
    .A2(_0401_),
    .Y(\MAC.mul.c_mul1[1] ),
    .B1(net325));
 sg13g2_nand2b_1 _2390_ (.Y(_0402_),
    .B(net311),
    .A_N(_0399_));
 sg13g2_nand3_1 _2391_ (.B(_0355_),
    .C(_0356_),
    .A(_0222_),
    .Y(_0403_));
 sg13g2_nand2b_1 _2392_ (.Y(_0404_),
    .B(_0403_),
    .A_N(_0357_));
 sg13g2_nand2b_1 _2393_ (.Y(_0405_),
    .B(_0404_),
    .A_N(net311));
 sg13g2_nand3_1 _2394_ (.B(_0402_),
    .C(_0405_),
    .A(net339),
    .Y(_0406_));
 sg13g2_a21oi_1 _2395_ (.A1(net321),
    .A2(_0406_),
    .Y(\MAC.mul.c_mul1[2] ),
    .B1(net325));
 sg13g2_xor2_1 _2396_ (.B(_0359_),
    .A(_0358_),
    .X(_0407_));
 sg13g2_o21ai_1 _2397_ (.B1(net339),
    .Y(_0408_),
    .A1(net311),
    .A2(_0407_));
 sg13g2_a21o_1 _2398_ (.A2(_0404_),
    .A1(net311),
    .B1(_0408_),
    .X(_0409_));
 sg13g2_a21oi_1 _2399_ (.A1(net321),
    .A2(_0409_),
    .Y(\MAC.mul.c_mul1[3] ),
    .B1(net325));
 sg13g2_nand2b_1 _2400_ (.Y(_0410_),
    .B(net311),
    .A_N(_0407_));
 sg13g2_xnor2_1 _2401_ (.Y(_0411_),
    .A(_0360_),
    .B(_0361_));
 sg13g2_nand2b_1 _2402_ (.Y(_0412_),
    .B(_0411_),
    .A_N(net311));
 sg13g2_nand3_1 _2403_ (.B(_0410_),
    .C(_0412_),
    .A(net339),
    .Y(_0413_));
 sg13g2_a21oi_1 _2404_ (.A1(net321),
    .A2(_0413_),
    .Y(\MAC.mul.c_mul1[4] ),
    .B1(net325));
 sg13g2_or3_1 _2405_ (.A(_1200_),
    .B(_0116_),
    .C(_0362_),
    .X(_0414_));
 sg13g2_nand2_1 _2406_ (.Y(_0415_),
    .A(_0363_),
    .B(_0414_));
 sg13g2_nand2b_1 _2407_ (.Y(_0416_),
    .B(_0415_),
    .A_N(net312));
 sg13g2_nand2_1 _2408_ (.Y(_0417_),
    .A(net311),
    .B(_0411_));
 sg13g2_nand3_1 _2409_ (.B(_0416_),
    .C(_0417_),
    .A(net339),
    .Y(_0418_));
 sg13g2_a21oi_1 _2410_ (.A1(net321),
    .A2(_0418_),
    .Y(\MAC.mul.c_mul1[5] ),
    .B1(net325));
 sg13g2_nand3_1 _2411_ (.B(_0363_),
    .C(_0365_),
    .A(_1198_),
    .Y(_0419_));
 sg13g2_nand2b_1 _2412_ (.Y(_0420_),
    .B(_0419_),
    .A_N(_0366_));
 sg13g2_nand2b_1 _2413_ (.Y(_0421_),
    .B(_0420_),
    .A_N(net312));
 sg13g2_nand2_1 _2414_ (.Y(_0422_),
    .A(net312),
    .B(_0415_));
 sg13g2_nand3_1 _2415_ (.B(_0421_),
    .C(_0422_),
    .A(net339),
    .Y(_0423_));
 sg13g2_a21oi_1 _2416_ (.A1(net321),
    .A2(_0423_),
    .Y(\MAC.mul.c_mul1[6] ),
    .B1(net325));
 sg13g2_or3_1 _2417_ (.A(_1135_),
    .B(_1162_),
    .C(_0366_),
    .X(_0424_));
 sg13g2_nand2_1 _2418_ (.Y(_0425_),
    .A(_0367_),
    .B(_0424_));
 sg13g2_nand2b_1 _2419_ (.Y(_0426_),
    .B(_0425_),
    .A_N(net313));
 sg13g2_nand2_1 _2420_ (.Y(_0427_),
    .A(net313),
    .B(_0420_));
 sg13g2_nand3_1 _2421_ (.B(_0426_),
    .C(_0427_),
    .A(net340),
    .Y(_0428_));
 sg13g2_a21oi_1 _2422_ (.A1(net321),
    .A2(_0428_),
    .Y(\MAC.mul.c_mul1[7] ),
    .B1(net325));
 sg13g2_xnor2_1 _2423_ (.Y(_0429_),
    .A(_0369_),
    .B(_0370_));
 sg13g2_nand2_1 _2424_ (.Y(_0430_),
    .A(net313),
    .B(_0425_));
 sg13g2_nand3_1 _2425_ (.B(_0429_),
    .C(_0430_),
    .A(net339),
    .Y(_0431_));
 sg13g2_a21oi_1 _2426_ (.A1(net321),
    .A2(_0431_),
    .Y(\MAC.mul.c_mul1[8] ),
    .B1(net325));
 sg13g2_nor2b_1 _2427_ (.A(_1036_),
    .B_N(net314),
    .Y(_0432_));
 sg13g2_nor2b_1 _2428_ (.A(net314),
    .B_N(_1036_),
    .Y(_0433_));
 sg13g2_o21ai_1 _2429_ (.B1(_1056_),
    .Y(_0434_),
    .A1(_0432_),
    .A2(_0433_));
 sg13g2_a21oi_1 _2430_ (.A1(_0396_),
    .A2(_0434_),
    .Y(\MAC.mul.c_mul1[9] ),
    .B1(_1045_));
 sg13g2_o21ai_1 _2431_ (.B1(net340),
    .Y(_0435_),
    .A1(_0382_),
    .A2(_0432_));
 sg13g2_a21o_1 _2432_ (.A2(_0432_),
    .A1(_0382_),
    .B1(_0435_),
    .X(_0436_));
 sg13g2_a21oi_1 _2433_ (.A1(net322),
    .A2(_0436_),
    .Y(\MAC.mul.c_mul1[10] ),
    .B1(net326));
 sg13g2_nor3_1 _2434_ (.A(_1036_),
    .B(net314),
    .C(_0382_),
    .Y(_0437_));
 sg13g2_nand2_2 _2435_ (.Y(_0438_),
    .A(_0381_),
    .B(_0437_));
 sg13g2_o21ai_1 _2436_ (.B1(net340),
    .Y(_0439_),
    .A1(_0381_),
    .A2(_0437_));
 sg13g2_nand2b_1 _2437_ (.Y(_0440_),
    .B(_0438_),
    .A_N(_0439_));
 sg13g2_a21oi_1 _2438_ (.A1(net322),
    .A2(_0440_),
    .Y(\MAC.mul.c_mul1[11] ),
    .B1(net326));
 sg13g2_o21ai_1 _2439_ (.B1(_0438_),
    .Y(_0441_),
    .A1(_1037_),
    .A2(_0380_));
 sg13g2_nand2b_1 _2440_ (.Y(_0442_),
    .B(_0441_),
    .A_N(_0383_));
 sg13g2_nand2b_1 _2441_ (.Y(_0443_),
    .B(_0383_),
    .A_N(_0441_));
 sg13g2_nand3_1 _2442_ (.B(_0442_),
    .C(_0443_),
    .A(net340),
    .Y(_0444_));
 sg13g2_a21oi_1 _2443_ (.A1(net322),
    .A2(_0444_),
    .Y(\MAC.mul.c_mul1[12] ),
    .B1(net326));
 sg13g2_o21ai_1 _2444_ (.B1(_1039_),
    .Y(_0445_),
    .A1(_1038_),
    .A2(_0378_));
 sg13g2_nor3_1 _2445_ (.A(_0383_),
    .B(_0438_),
    .C(_0445_),
    .Y(_0446_));
 sg13g2_o21ai_1 _2446_ (.B1(_0445_),
    .Y(_0447_),
    .A1(_0383_),
    .A2(_0438_));
 sg13g2_nand3b_1 _2447_ (.B(_0447_),
    .C(net340),
    .Y(_0448_),
    .A_N(_0446_));
 sg13g2_a21oi_1 _2448_ (.A1(net322),
    .A2(_0448_),
    .Y(\MAC.mul.c_mul1[13] ),
    .B1(net326));
 sg13g2_nand2b_1 _2449_ (.Y(_0449_),
    .B(_1041_),
    .A_N(_0446_));
 sg13g2_nand2b_1 _2450_ (.Y(_0450_),
    .B(_0446_),
    .A_N(_1040_));
 sg13g2_nand3_1 _2451_ (.B(_0449_),
    .C(_0450_),
    .A(net340),
    .Y(_0451_));
 sg13g2_a21oi_1 _2452_ (.A1(net322),
    .A2(_0451_),
    .Y(\MAC.mul.c_mul1[14] ),
    .B1(net326));
 sg13g2_xor2_1 _2453_ (.B(net76),
    .A(\MAC.a[15] ),
    .X(_0452_));
 sg13g2_nand2_1 _2454_ (.Y(_0453_),
    .A(net340),
    .B(net77));
 sg13g2_o21ai_1 _2455_ (.B1(_1044_),
    .Y(_0454_),
    .A1(_1042_),
    .A2(net77));
 sg13g2_a21oi_1 _2456_ (.A1(net322),
    .A2(_0453_),
    .Y(\MAC.mul.c_mul1[15] ),
    .B1(_0454_));
 sg13g2_nand2_1 _2457_ (.Y(_0455_),
    .A(net58),
    .B(\MAC.add.b1[0] ));
 sg13g2_o21ai_1 _2458_ (.B1(net59),
    .Y(_0034_),
    .A1(net58),
    .A2(_0471_));
 sg13g2_mux2_1 _2459_ (.A0(\MAC.add.b1[9] ),
    .A1(net62),
    .S(net58),
    .X(_0035_));
 sg13g2_mux2_1 _2460_ (.A0(net68),
    .A1(\MAC.add.b1[2] ),
    .S(net375),
    .X(_0036_));
 sg13g2_nor2_1 _2461_ (.A(net375),
    .B(net64),
    .Y(_0456_));
 sg13g2_a21oi_1 _2462_ (.A1(net375),
    .A2(_0463_),
    .Y(_0037_),
    .B1(_0456_));
 sg13g2_mux2_1 _2463_ (.A0(\MAC.add.b1[12] ),
    .A1(net70),
    .S(net375),
    .X(_0038_));
 sg13g2_mux2_1 _2464_ (.A0(net74),
    .A1(\MAC.add.b1[5] ),
    .S(net375),
    .X(_0039_));
 sg13g2_nor2_1 _2465_ (.A(net375),
    .B(\MAC.add.b1[14] ),
    .Y(_0457_));
 sg13g2_a21oi_1 _2466_ (.A1(net375),
    .A2(_0466_),
    .Y(_0040_),
    .B1(_0457_));
 sg13g2_mux2_1 _2467_ (.A0(\MAC.add.b1[15] ),
    .A1(net72),
    .S(net375),
    .X(_0041_));
 sg13g2_mux2_1 _2468_ (.A0(net1),
    .A1(net43),
    .S(net352),
    .X(_0062_));
 sg13g2_mux2_1 _2469_ (.A0(net2),
    .A1(net53),
    .S(net352),
    .X(_0063_));
 sg13g2_mux2_1 _2470_ (.A0(net3),
    .A1(net35),
    .S(net353),
    .X(_0064_));
 sg13g2_mux2_1 _2471_ (.A0(net4),
    .A1(net54),
    .S(net352),
    .X(_0065_));
 sg13g2_mux2_1 _2472_ (.A0(net5),
    .A1(net37),
    .S(net352),
    .X(_0066_));
 sg13g2_mux2_1 _2473_ (.A0(net6),
    .A1(net40),
    .S(net350),
    .X(_0067_));
 sg13g2_mux2_1 _2474_ (.A0(net7),
    .A1(net52),
    .S(net351),
    .X(_0068_));
 sg13g2_mux2_1 _2475_ (.A0(net8),
    .A1(net49),
    .S(net350),
    .X(_0069_));
 sg13g2_mux2_1 _2476_ (.A0(net9),
    .A1(net51),
    .S(net351),
    .X(_0070_));
 sg13g2_mux2_1 _2477_ (.A0(net10),
    .A1(net56),
    .S(net349),
    .X(_0071_));
 sg13g2_mux2_1 _2478_ (.A0(net11),
    .A1(net46),
    .S(net349),
    .X(_0072_));
 sg13g2_mux2_1 _2479_ (.A0(net12),
    .A1(net42),
    .S(net347),
    .X(_0073_));
 sg13g2_mux2_1 _2480_ (.A0(net13),
    .A1(net48),
    .S(net347),
    .X(_0074_));
 sg13g2_mux2_1 _2481_ (.A0(net14),
    .A1(net44),
    .S(net347),
    .X(_0075_));
 sg13g2_mux2_1 _2482_ (.A0(net15),
    .A1(net39),
    .S(net347),
    .X(_0076_));
 sg13g2_mux2_1 _2483_ (.A0(net16),
    .A1(net45),
    .S(net348),
    .X(_0077_));
 sg13g2_dfrbp_1 _2484_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net405),
    .D(_0002_),
    .Q_N(_1220_),
    .Q(\MAC.a[0] ));
 sg13g2_dfrbp_1 _2485_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net405),
    .D(_0009_),
    .Q_N(_1221_),
    .Q(\MAC.a[1] ));
 sg13g2_dfrbp_1 _2486_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net407),
    .D(net36),
    .Q_N(_1222_),
    .Q(\MAC.a[2] ));
 sg13g2_dfrbp_1 _2487_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net407),
    .D(net55),
    .Q_N(_1223_),
    .Q(\MAC.a[3] ));
 sg13g2_dfrbp_1 _2488_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net404),
    .D(net38),
    .Q_N(_1224_),
    .Q(\MAC.a[4] ));
 sg13g2_dfrbp_1 _2489_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net404),
    .D(net41),
    .Q_N(_1225_),
    .Q(\MAC.a[5] ));
 sg13g2_dfrbp_1 _2490_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net404),
    .D(_0014_),
    .Q_N(_1226_),
    .Q(\MAC.a[6] ));
 sg13g2_dfrbp_1 _2491_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net404),
    .D(net50),
    .Q_N(_1227_),
    .Q(\MAC.a[7] ));
 sg13g2_dfrbp_1 _2492_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net404),
    .D(_0016_),
    .Q_N(_1228_),
    .Q(\MAC.a[8] ));
 sg13g2_dfrbp_1 _2493_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net403),
    .D(net57),
    .Q_N(_1229_),
    .Q(\MAC.a[9] ));
 sg13g2_dfrbp_1 _2494_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net403),
    .D(net47),
    .Q_N(_1230_),
    .Q(\MAC.a[10] ));
 sg13g2_dfrbp_1 _2495_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net402),
    .D(_0004_),
    .Q_N(_1231_),
    .Q(\MAC.a[11] ));
 sg13g2_dfrbp_1 _2496_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net402),
    .D(_0005_),
    .Q_N(_1232_),
    .Q(\MAC.a[12] ));
 sg13g2_dfrbp_1 _2497_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net399),
    .D(_0006_),
    .Q_N(_1233_),
    .Q(\MAC.a[13] ));
 sg13g2_dfrbp_1 _2498_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net400),
    .D(_0007_),
    .Q_N(_1234_),
    .Q(\MAC.a[14] ));
 sg13g2_dfrbp_1 _2499_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net400),
    .D(_0008_),
    .Q_N(_1235_),
    .Q(\MAC.a[15] ));
 sg13g2_dfrbp_1 _2500_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net397),
    .D(net34),
    .Q_N(_0001_),
    .Q(\wrap2.state[0] ));
 sg13g2_dfrbp_1 _2501_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net405),
    .D(_0018_),
    .Q_N(_1236_),
    .Q(\MAC.b[0] ));
 sg13g2_dfrbp_1 _2502_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net405),
    .D(_0025_),
    .Q_N(_1237_),
    .Q(\MAC.b[1] ));
 sg13g2_dfrbp_1 _2503_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net404),
    .D(_0026_),
    .Q_N(_0043_),
    .Q(\MAC.b[2] ));
 sg13g2_dfrbp_1 _2504_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net407),
    .D(_0027_),
    .Q_N(_1238_),
    .Q(\MAC.b[3] ));
 sg13g2_dfrbp_1 _2505_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net405),
    .D(_0028_),
    .Q_N(_1239_),
    .Q(\MAC.b[4] ));
 sg13g2_dfrbp_1 _2506_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net403),
    .D(_0029_),
    .Q_N(_0042_),
    .Q(\MAC.b[5] ));
 sg13g2_dfrbp_1 _2507_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net404),
    .D(_0030_),
    .Q_N(_1240_),
    .Q(\MAC.b[6] ));
 sg13g2_dfrbp_1 _2508_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net406),
    .D(_0031_),
    .Q_N(_1241_),
    .Q(\MAC.b[7] ));
 sg13g2_dfrbp_1 _2509_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net403),
    .D(_0032_),
    .Q_N(_1242_),
    .Q(\MAC.b[8] ));
 sg13g2_dfrbp_1 _2510_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net402),
    .D(_0033_),
    .Q_N(_1243_),
    .Q(\MAC.b[9] ));
 sg13g2_dfrbp_1 _2511_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net402),
    .D(_0019_),
    .Q_N(_1244_),
    .Q(\MAC.b[10] ));
 sg13g2_dfrbp_1 _2512_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net402),
    .D(_0020_),
    .Q_N(_1245_),
    .Q(\MAC.b[11] ));
 sg13g2_dfrbp_1 _2513_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net402),
    .D(_0021_),
    .Q_N(_1246_),
    .Q(\MAC.b[12] ));
 sg13g2_dfrbp_1 _2514_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net399),
    .D(_0022_),
    .Q_N(_1247_),
    .Q(\MAC.b[13] ));
 sg13g2_dfrbp_1 _2515_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net400),
    .D(_0023_),
    .Q_N(_1248_),
    .Q(\MAC.b[14] ));
 sg13g2_dfrbp_1 _2516_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net400),
    .D(_0024_),
    .Q_N(_1249_),
    .Q(\MAC.b[15] ));
 sg13g2_dfrbp_1 _2517_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net399),
    .D(net60),
    .Q_N(_1250_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _2518_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net399),
    .D(net63),
    .Q_N(_1251_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _2519_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net399),
    .D(net69),
    .Q_N(_1252_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _2520_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net398),
    .D(net65),
    .Q_N(_1253_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _2521_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net397),
    .D(net71),
    .Q_N(_1254_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _2522_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net397),
    .D(net75),
    .Q_N(_1255_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _2523_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net397),
    .D(net67),
    .Q_N(_1256_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _2524_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net397),
    .D(net73),
    .Q_N(_1257_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _2525_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net399),
    .D(net33),
    .Q_N(_0000_),
    .Q(\wrap.state[0] ));
 sg13g2_dfrbp_1 _2526_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net395),
    .D(\MAC.mul.c_mul1[0] ),
    .Q_N(_0045_),
    .Q(\MAC.add.a1[0] ));
 sg13g2_dfrbp_1 _2527_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net394),
    .D(\MAC.mul.c_mul1[1] ),
    .Q_N(_0047_),
    .Q(\MAC.add.a1[1] ));
 sg13g2_dfrbp_1 _2528_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net394),
    .D(\MAC.mul.c_mul1[2] ),
    .Q_N(_0049_),
    .Q(\MAC.add.a1[2] ));
 sg13g2_dfrbp_1 _2529_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net394),
    .D(\MAC.mul.c_mul1[3] ),
    .Q_N(_0051_),
    .Q(\MAC.add.a1[3] ));
 sg13g2_dfrbp_1 _2530_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net394),
    .D(\MAC.mul.c_mul1[4] ),
    .Q_N(_0053_),
    .Q(\MAC.add.a1[4] ));
 sg13g2_dfrbp_1 _2531_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net394),
    .D(\MAC.mul.c_mul1[5] ),
    .Q_N(_0055_),
    .Q(\MAC.add.a1[5] ));
 sg13g2_dfrbp_1 _2532_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net393),
    .D(\MAC.mul.c_mul1[6] ),
    .Q_N(_0057_),
    .Q(\MAC.add.a1[6] ));
 sg13g2_dfrbp_1 _2533_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net394),
    .D(\MAC.mul.c_mul1[7] ),
    .Q_N(_0059_),
    .Q(\MAC.add.a1[7] ));
 sg13g2_dfrbp_1 _2534_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net394),
    .D(\MAC.mul.c_mul1[8] ),
    .Q_N(_0061_),
    .Q(\MAC.add.a1[8] ));
 sg13g2_dfrbp_1 _2535_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net395),
    .D(\MAC.mul.c_mul1[9] ),
    .Q_N(_1258_),
    .Q(\MAC.add.a1[9] ));
 sg13g2_dfrbp_1 _2536_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net395),
    .D(\MAC.mul.c_mul1[10] ),
    .Q_N(_1259_),
    .Q(\MAC.add.a1[10] ));
 sg13g2_dfrbp_1 _2537_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net395),
    .D(\MAC.mul.c_mul1[11] ),
    .Q_N(_1260_),
    .Q(\MAC.add.a1[11] ));
 sg13g2_dfrbp_1 _2538_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net395),
    .D(\MAC.mul.c_mul1[12] ),
    .Q_N(_1261_),
    .Q(\MAC.add.a1[12] ));
 sg13g2_dfrbp_1 _2539_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net394),
    .D(\MAC.mul.c_mul1[13] ),
    .Q_N(_1262_),
    .Q(\MAC.add.a1[13] ));
 sg13g2_dfrbp_1 _2540_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net400),
    .D(\MAC.mul.c_mul1[14] ),
    .Q_N(_1263_),
    .Q(\MAC.add.a1[14] ));
 sg13g2_dfrbp_1 _2541_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net395),
    .D(\MAC.mul.c_mul1[15] ),
    .Q_N(_1264_),
    .Q(\MAC.add.a1[15] ));
 sg13g2_dfrbp_1 _2542_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net398),
    .D(\MAC.add.c_add[0] ),
    .Q_N(_0044_),
    .Q(\MAC.add.b1[0] ));
 sg13g2_dfrbp_1 _2543_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net393),
    .D(\MAC.add.c_add[1] ),
    .Q_N(_0046_),
    .Q(\MAC.add.b1[1] ));
 sg13g2_dfrbp_1 _2544_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net393),
    .D(\MAC.add.c_add[2] ),
    .Q_N(_0048_),
    .Q(\MAC.add.b1[2] ));
 sg13g2_dfrbp_1 _2545_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net393),
    .D(\MAC.add.c_add[3] ),
    .Q_N(_0050_),
    .Q(\MAC.add.b1[3] ));
 sg13g2_dfrbp_1 _2546_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net393),
    .D(\MAC.add.c_add[4] ),
    .Q_N(_0052_),
    .Q(\MAC.add.b1[4] ));
 sg13g2_dfrbp_1 _2547_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net396),
    .D(\MAC.add.c_add[5] ),
    .Q_N(_0054_),
    .Q(\MAC.add.b1[5] ));
 sg13g2_dfrbp_1 _2548_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net393),
    .D(\MAC.add.c_add[6] ),
    .Q_N(_0056_),
    .Q(\MAC.add.b1[6] ));
 sg13g2_dfrbp_1 _2549_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net393),
    .D(\MAC.add.c_add[7] ),
    .Q_N(_0058_),
    .Q(\MAC.add.b1[7] ));
 sg13g2_dfrbp_1 _2550_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net393),
    .D(\MAC.add.c_add[8] ),
    .Q_N(_0060_),
    .Q(\MAC.add.b1[8] ));
 sg13g2_dfrbp_1 _2551_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net398),
    .D(\MAC.add.c_add[9] ),
    .Q_N(_1265_),
    .Q(\MAC.add.b1[9] ));
 sg13g2_dfrbp_1 _2552_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net398),
    .D(\MAC.add.c_add[10] ),
    .Q_N(_1266_),
    .Q(\MAC.add.b1[10] ));
 sg13g2_dfrbp_1 _2553_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net398),
    .D(\MAC.add.c_add[11] ),
    .Q_N(_1267_),
    .Q(\MAC.add.b1[11] ));
 sg13g2_dfrbp_1 _2554_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net397),
    .D(\MAC.add.c_add[12] ),
    .Q_N(_1268_),
    .Q(\MAC.add.b1[12] ));
 sg13g2_dfrbp_1 _2555_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net397),
    .D(\MAC.add.c_add[13] ),
    .Q_N(_1269_),
    .Q(\MAC.add.b1[13] ));
 sg13g2_dfrbp_1 _2556_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net397),
    .D(\MAC.add.c_add[14] ),
    .Q_N(_1270_),
    .Q(\MAC.add.b1[14] ));
 sg13g2_dfrbp_1 _2557_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net398),
    .D(\MAC.add.c_add[15] ),
    .Q_N(_1219_),
    .Q(\MAC.add.b1[15] ));
 sg13g2_dfrbp_1 _2558_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net406),
    .D(_0062_),
    .Q_N(_1218_),
    .Q(\wrap.temp_data[0] ));
 sg13g2_dfrbp_1 _2559_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net406),
    .D(_0063_),
    .Q_N(_1217_),
    .Q(\wrap.temp_data[1] ));
 sg13g2_dfrbp_1 _2560_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net405),
    .D(_0064_),
    .Q_N(_1216_),
    .Q(\wrap.temp_data[2] ));
 sg13g2_dfrbp_1 _2561_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net405),
    .D(_0065_),
    .Q_N(_1215_),
    .Q(\wrap.temp_data[3] ));
 sg13g2_dfrbp_1 _2562_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net405),
    .D(_0066_),
    .Q_N(_1214_),
    .Q(\wrap.temp_data[4] ));
 sg13g2_dfrbp_1 _2563_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net404),
    .D(_0067_),
    .Q_N(_1213_),
    .Q(\wrap.temp_data[5] ));
 sg13g2_dfrbp_1 _2564_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net406),
    .D(_0068_),
    .Q_N(_1212_),
    .Q(\wrap.temp_data[6] ));
 sg13g2_dfrbp_1 _2565_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net406),
    .D(_0069_),
    .Q_N(_1211_),
    .Q(\wrap.temp_data[7] ));
 sg13g2_dfrbp_1 _2566_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net403),
    .D(_0070_),
    .Q_N(_1210_),
    .Q(\wrap.temp_data[8] ));
 sg13g2_dfrbp_1 _2567_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net402),
    .D(_0071_),
    .Q_N(_1209_),
    .Q(\wrap.temp_data[9] ));
 sg13g2_dfrbp_1 _2568_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net402),
    .D(_0072_),
    .Q_N(_1208_),
    .Q(\wrap.temp_data[10] ));
 sg13g2_dfrbp_1 _2569_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net400),
    .D(_0073_),
    .Q_N(_1207_),
    .Q(\wrap.temp_data[11] ));
 sg13g2_dfrbp_1 _2570_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net401),
    .D(_0074_),
    .Q_N(_1206_),
    .Q(\wrap.temp_data[12] ));
 sg13g2_dfrbp_1 _2571_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net400),
    .D(_0075_),
    .Q_N(_1205_),
    .Q(\wrap.temp_data[13] ));
 sg13g2_dfrbp_1 _2572_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net399),
    .D(_0076_),
    .Q_N(_1204_),
    .Q(\wrap.temp_data[14] ));
 sg13g2_dfrbp_1 _2573_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net399),
    .D(_0077_),
    .Q_N(_1203_),
    .Q(\wrap.temp_data[15] ));
 sg13g2_tielo tt_um_dlfloatmac_18 (.L_LO(net18));
 sg13g2_tielo tt_um_dlfloatmac_19 (.L_LO(net19));
 sg13g2_tielo tt_um_dlfloatmac_20 (.L_LO(net20));
 sg13g2_tielo tt_um_dlfloatmac_21 (.L_LO(net21));
 sg13g2_tielo tt_um_dlfloatmac_22 (.L_LO(net22));
 sg13g2_tielo tt_um_dlfloatmac_23 (.L_LO(net23));
 sg13g2_tielo tt_um_dlfloatmac_24 (.L_LO(net24));
 sg13g2_tielo tt_um_dlfloatmac_25 (.L_LO(net25));
 sg13g2_tielo tt_um_dlfloatmac_26 (.L_LO(net26));
 sg13g2_tielo tt_um_dlfloatmac_27 (.L_LO(net27));
 sg13g2_tielo tt_um_dlfloatmac_28 (.L_LO(net28));
 sg13g2_tielo tt_um_dlfloatmac_29 (.L_LO(net29));
 sg13g2_tielo tt_um_dlfloatmac_30 (.L_LO(net30));
 sg13g2_tielo tt_um_dlfloatmac_31 (.L_LO(net31));
 sg13g2_tielo tt_um_dlfloatmac_32 (.L_LO(net32));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 fanout306 (.A(_0886_),
    .X(net306));
 sg13g2_buf_1 fanout307 (.A(_0886_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_0913_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(net310),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_0829_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(net312),
    .X(net311));
 sg13g2_buf_1 fanout312 (.A(net313),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(net314),
    .X(net313));
 sg13g2_buf_1 fanout314 (.A(_0371_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_0822_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(net317),
    .X(net316));
 sg13g2_buf_1 fanout317 (.A(net318),
    .X(net317));
 sg13g2_buf_1 fanout318 (.A(_0784_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(net320),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_0673_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_0397_),
    .X(net321));
 sg13g2_buf_1 fanout322 (.A(_0397_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_0544_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_1043_),
    .X(net325));
 sg13g2_buf_1 fanout326 (.A(_1043_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(net328),
    .X(net327));
 sg13g2_buf_1 fanout328 (.A(_0576_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_0550_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_0549_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(net332),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_0511_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(net334),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(net335),
    .X(net334));
 sg13g2_buf_1 fanout335 (.A(net336),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_0510_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(net338),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_0509_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(net340),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_1056_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_0524_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_0489_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(net345),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(net345),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_0493_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_0490_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(net348),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(net349),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(net354),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(net354),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(net354),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(net353),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(net354),
    .X(net353));
 sg13g2_buf_1 fanout354 (.A(net61),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(net356),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(net357),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(\MAC.b[8] ),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(net359),
    .X(net358));
 sg13g2_buf_4 fanout359 (.X(net359),
    .A(\MAC.b[7] ));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(net362));
 sg13g2_buf_1 fanout361 (.A(net362),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(\MAC.b[6] ),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(net364),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(\MAC.b[5] ),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(net366),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(\MAC.b[4] ),
    .X(net366));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(\MAC.b[3] ));
 sg13g2_buf_2 fanout368 (.A(\MAC.b[3] ),
    .X(net368));
 sg13g2_buf_4 fanout369 (.X(net369),
    .A(\MAC.b[2] ));
 sg13g2_buf_2 fanout370 (.A(\MAC.b[2] ),
    .X(net370));
 sg13g2_buf_4 fanout371 (.X(net371),
    .A(\MAC.b[1] ));
 sg13g2_buf_2 fanout372 (.A(\MAC.b[1] ),
    .X(net372));
 sg13g2_buf_4 fanout373 (.X(net373),
    .A(\MAC.b[0] ));
 sg13g2_buf_1 fanout374 (.A(\MAC.b[0] ),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(net58),
    .X(net375));
 sg13g2_buf_4 fanout376 (.X(net376),
    .A(net377));
 sg13g2_buf_2 fanout377 (.A(\MAC.a[8] ),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(net379),
    .X(net378));
 sg13g2_buf_4 fanout379 (.X(net379),
    .A(\MAC.a[7] ));
 sg13g2_buf_4 fanout380 (.X(net380),
    .A(net381));
 sg13g2_buf_4 fanout381 (.X(net381),
    .A(\MAC.a[6] ));
 sg13g2_buf_4 fanout382 (.X(net382),
    .A(\MAC.a[5] ));
 sg13g2_buf_1 fanout383 (.A(\MAC.a[5] ),
    .X(net383));
 sg13g2_buf_4 fanout384 (.X(net384),
    .A(\MAC.a[4] ));
 sg13g2_buf_2 fanout385 (.A(\MAC.a[4] ),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(\MAC.a[3] ),
    .X(net386));
 sg13g2_buf_1 fanout387 (.A(\MAC.a[3] ),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(net389),
    .X(net388));
 sg13g2_buf_4 fanout389 (.X(net389),
    .A(\MAC.a[2] ));
 sg13g2_buf_2 fanout390 (.A(\MAC.a[1] ),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(\MAC.a[1] ),
    .X(net391));
 sg13g2_buf_4 fanout392 (.X(net392),
    .A(\MAC.a[0] ));
 sg13g2_buf_4 fanout393 (.X(net393),
    .A(net396));
 sg13g2_buf_4 fanout394 (.X(net394),
    .A(net396));
 sg13g2_buf_4 fanout395 (.X(net395),
    .A(net396));
 sg13g2_buf_2 fanout396 (.A(net401),
    .X(net396));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(net398));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(net401));
 sg13g2_buf_4 fanout399 (.X(net399),
    .A(net400));
 sg13g2_buf_4 fanout400 (.X(net400),
    .A(net401));
 sg13g2_buf_2 fanout401 (.A(rst_n),
    .X(net401));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(net403));
 sg13g2_buf_4 fanout403 (.X(net403),
    .A(rst_n));
 sg13g2_buf_4 fanout404 (.X(net404),
    .A(net407));
 sg13g2_buf_4 fanout405 (.X(net405),
    .A(net406));
 sg13g2_buf_4 fanout406 (.X(net406),
    .A(net407));
 sg13g2_buf_2 fanout407 (.A(rst_n),
    .X(net407));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_tielo tt_um_dlfloatmac_17 (.L_LO(net17));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0000_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0001_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold3 (.A(\wrap.temp_data[2] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0010_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold5 (.A(\wrap.temp_data[4] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0012_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold7 (.A(\wrap.temp_data[14] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold8 (.A(\wrap.temp_data[5] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0013_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold10 (.A(\wrap.temp_data[11] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold11 (.A(\wrap.temp_data[0] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold12 (.A(\wrap.temp_data[13] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold13 (.A(\wrap.temp_data[15] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold14 (.A(\wrap.temp_data[10] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0003_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold16 (.A(\wrap.temp_data[12] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold17 (.A(\wrap.temp_data[7] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0015_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold19 (.A(\wrap.temp_data[8] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold20 (.A(\wrap.temp_data[6] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold21 (.A(\wrap.temp_data[1] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold22 (.A(\wrap.temp_data[3] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0011_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold24 (.A(\wrap.temp_data[9] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0017_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold26 (.A(\wrap2.state[0] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0455_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0034_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold29 (.A(\wrap.state[0] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold30 (.A(\MAC.add.b1[1] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0035_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold32 (.A(\MAC.add.b1[11] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0037_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold34 (.A(\MAC.add.b1[6] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0040_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold36 (.A(\MAC.add.b1[10] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0036_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold38 (.A(\MAC.add.b1[4] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0038_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold40 (.A(\MAC.add.b1[7] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0041_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold42 (.A(\MAC.add.b1[13] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0039_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold44 (.A(\MAC.b[15] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0452_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold46 (.A(\MAC.add.a1[15] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold47 (.A(_1018_),
    .X(net79));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_decap_8 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_fill_1 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_313 ();
 sg13g2_decap_8 FILLER_34_320 ();
 sg13g2_decap_8 FILLER_34_327 ();
 sg13g2_fill_2 FILLER_34_334 ();
 sg13g2_decap_8 FILLER_34_348 ();
 sg13g2_decap_8 FILLER_34_355 ();
 sg13g2_decap_8 FILLER_34_362 ();
 sg13g2_decap_8 FILLER_34_369 ();
 sg13g2_decap_8 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_34_383 ();
 sg13g2_decap_8 FILLER_34_390 ();
 sg13g2_decap_8 FILLER_34_397 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_fill_2 FILLER_35_301 ();
 sg13g2_fill_1 FILLER_35_303 ();
 sg13g2_decap_8 FILLER_35_321 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_fill_2 FILLER_36_294 ();
 sg13g2_fill_1 FILLER_36_296 ();
 sg13g2_fill_1 FILLER_36_302 ();
 sg13g2_fill_1 FILLER_36_347 ();
 sg13g2_fill_1 FILLER_36_366 ();
 sg13g2_fill_1 FILLER_36_377 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_fill_2 FILLER_37_287 ();
 sg13g2_fill_1 FILLER_37_289 ();
 sg13g2_decap_4 FILLER_37_330 ();
 sg13g2_fill_2 FILLER_37_334 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_4 FILLER_38_284 ();
 sg13g2_fill_2 FILLER_38_297 ();
 sg13g2_fill_2 FILLER_38_312 ();
 sg13g2_fill_1 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_fill_2 FILLER_38_347 ();
 sg13g2_fill_1 FILLER_38_370 ();
 sg13g2_fill_1 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_decap_8 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_238 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_4 FILLER_39_266 ();
 sg13g2_fill_2 FILLER_39_270 ();
 sg13g2_decap_8 FILLER_39_310 ();
 sg13g2_fill_2 FILLER_39_317 ();
 sg13g2_fill_1 FILLER_39_319 ();
 sg13g2_fill_2 FILLER_39_324 ();
 sg13g2_decap_8 FILLER_39_344 ();
 sg13g2_decap_4 FILLER_39_351 ();
 sg13g2_fill_1 FILLER_39_355 ();
 sg13g2_fill_1 FILLER_39_364 ();
 sg13g2_fill_2 FILLER_39_373 ();
 sg13g2_decap_4 FILLER_39_384 ();
 sg13g2_fill_2 FILLER_39_388 ();
 sg13g2_decap_8 FILLER_39_394 ();
 sg13g2_decap_8 FILLER_39_401 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_fill_1 FILLER_40_147 ();
 sg13g2_fill_2 FILLER_40_153 ();
 sg13g2_fill_1 FILLER_40_155 ();
 sg13g2_decap_8 FILLER_40_176 ();
 sg13g2_decap_8 FILLER_40_183 ();
 sg13g2_decap_8 FILLER_40_190 ();
 sg13g2_decap_8 FILLER_40_197 ();
 sg13g2_decap_8 FILLER_40_204 ();
 sg13g2_decap_8 FILLER_40_211 ();
 sg13g2_decap_8 FILLER_40_218 ();
 sg13g2_decap_8 FILLER_40_225 ();
 sg13g2_decap_8 FILLER_40_232 ();
 sg13g2_decap_8 FILLER_40_239 ();
 sg13g2_decap_8 FILLER_40_246 ();
 sg13g2_decap_8 FILLER_40_253 ();
 sg13g2_decap_8 FILLER_40_260 ();
 sg13g2_fill_2 FILLER_40_286 ();
 sg13g2_fill_2 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_decap_8 FILLER_40_323 ();
 sg13g2_decap_4 FILLER_40_330 ();
 sg13g2_fill_2 FILLER_40_338 ();
 sg13g2_fill_2 FILLER_40_361 ();
 sg13g2_fill_2 FILLER_40_371 ();
 sg13g2_fill_1 FILLER_40_373 ();
 sg13g2_fill_2 FILLER_40_389 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_4 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_183 ();
 sg13g2_decap_8 FILLER_41_190 ();
 sg13g2_decap_8 FILLER_41_197 ();
 sg13g2_decap_8 FILLER_41_204 ();
 sg13g2_decap_8 FILLER_41_211 ();
 sg13g2_decap_8 FILLER_41_218 ();
 sg13g2_decap_8 FILLER_41_225 ();
 sg13g2_decap_8 FILLER_41_232 ();
 sg13g2_decap_8 FILLER_41_239 ();
 sg13g2_decap_8 FILLER_41_246 ();
 sg13g2_decap_8 FILLER_41_253 ();
 sg13g2_decap_8 FILLER_41_260 ();
 sg13g2_decap_4 FILLER_41_267 ();
 sg13g2_fill_1 FILLER_41_287 ();
 sg13g2_fill_2 FILLER_41_293 ();
 sg13g2_decap_8 FILLER_41_307 ();
 sg13g2_fill_2 FILLER_41_314 ();
 sg13g2_fill_2 FILLER_41_329 ();
 sg13g2_fill_1 FILLER_41_331 ();
 sg13g2_fill_2 FILLER_41_343 ();
 sg13g2_fill_1 FILLER_41_345 ();
 sg13g2_fill_2 FILLER_41_376 ();
 sg13g2_fill_1 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_fill_2 FILLER_42_153 ();
 sg13g2_fill_1 FILLER_42_163 ();
 sg13g2_decap_8 FILLER_42_191 ();
 sg13g2_decap_8 FILLER_42_198 ();
 sg13g2_decap_8 FILLER_42_205 ();
 sg13g2_decap_8 FILLER_42_212 ();
 sg13g2_decap_8 FILLER_42_219 ();
 sg13g2_decap_8 FILLER_42_226 ();
 sg13g2_decap_8 FILLER_42_233 ();
 sg13g2_decap_8 FILLER_42_240 ();
 sg13g2_decap_8 FILLER_42_247 ();
 sg13g2_decap_8 FILLER_42_254 ();
 sg13g2_decap_8 FILLER_42_261 ();
 sg13g2_decap_8 FILLER_42_268 ();
 sg13g2_decap_8 FILLER_42_275 ();
 sg13g2_decap_8 FILLER_42_286 ();
 sg13g2_decap_8 FILLER_42_293 ();
 sg13g2_fill_2 FILLER_42_333 ();
 sg13g2_fill_2 FILLER_42_345 ();
 sg13g2_fill_1 FILLER_42_347 ();
 sg13g2_fill_2 FILLER_42_353 ();
 sg13g2_decap_4 FILLER_42_360 ();
 sg13g2_fill_2 FILLER_42_372 ();
 sg13g2_decap_4 FILLER_42_382 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_4 FILLER_43_84 ();
 sg13g2_fill_1 FILLER_43_88 ();
 sg13g2_decap_4 FILLER_43_93 ();
 sg13g2_fill_1 FILLER_43_97 ();
 sg13g2_decap_8 FILLER_43_103 ();
 sg13g2_decap_4 FILLER_43_110 ();
 sg13g2_fill_2 FILLER_43_165 ();
 sg13g2_fill_2 FILLER_43_174 ();
 sg13g2_fill_1 FILLER_43_176 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_259 ();
 sg13g2_decap_4 FILLER_43_266 ();
 sg13g2_fill_2 FILLER_43_270 ();
 sg13g2_fill_2 FILLER_43_297 ();
 sg13g2_fill_1 FILLER_43_308 ();
 sg13g2_fill_1 FILLER_43_312 ();
 sg13g2_fill_1 FILLER_43_318 ();
 sg13g2_fill_2 FILLER_43_350 ();
 sg13g2_fill_1 FILLER_43_352 ();
 sg13g2_decap_8 FILLER_43_361 ();
 sg13g2_decap_4 FILLER_43_368 ();
 sg13g2_fill_2 FILLER_43_389 ();
 sg13g2_fill_1 FILLER_43_391 ();
 sg13g2_decap_8 FILLER_43_401 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_4 FILLER_44_77 ();
 sg13g2_fill_2 FILLER_44_94 ();
 sg13g2_fill_1 FILLER_44_96 ();
 sg13g2_fill_1 FILLER_44_118 ();
 sg13g2_decap_8 FILLER_44_180 ();
 sg13g2_fill_2 FILLER_44_187 ();
 sg13g2_decap_8 FILLER_44_194 ();
 sg13g2_decap_8 FILLER_44_201 ();
 sg13g2_decap_8 FILLER_44_208 ();
 sg13g2_decap_8 FILLER_44_215 ();
 sg13g2_decap_8 FILLER_44_222 ();
 sg13g2_decap_8 FILLER_44_229 ();
 sg13g2_decap_8 FILLER_44_236 ();
 sg13g2_decap_8 FILLER_44_243 ();
 sg13g2_decap_8 FILLER_44_250 ();
 sg13g2_decap_8 FILLER_44_257 ();
 sg13g2_decap_4 FILLER_44_264 ();
 sg13g2_fill_1 FILLER_44_268 ();
 sg13g2_fill_2 FILLER_44_277 ();
 sg13g2_fill_1 FILLER_44_279 ();
 sg13g2_fill_2 FILLER_44_293 ();
 sg13g2_fill_1 FILLER_44_310 ();
 sg13g2_fill_2 FILLER_44_323 ();
 sg13g2_fill_1 FILLER_44_341 ();
 sg13g2_fill_2 FILLER_44_369 ();
 sg13g2_fill_1 FILLER_44_371 ();
 sg13g2_fill_2 FILLER_44_384 ();
 sg13g2_fill_1 FILLER_44_386 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_4 FILLER_45_77 ();
 sg13g2_fill_2 FILLER_45_145 ();
 sg13g2_fill_1 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_158 ();
 sg13g2_decap_4 FILLER_45_165 ();
 sg13g2_fill_1 FILLER_45_169 ();
 sg13g2_fill_2 FILLER_45_175 ();
 sg13g2_decap_4 FILLER_45_188 ();
 sg13g2_decap_4 FILLER_45_197 ();
 sg13g2_decap_8 FILLER_45_227 ();
 sg13g2_decap_8 FILLER_45_234 ();
 sg13g2_decap_8 FILLER_45_241 ();
 sg13g2_decap_8 FILLER_45_248 ();
 sg13g2_decap_4 FILLER_45_255 ();
 sg13g2_fill_1 FILLER_45_259 ();
 sg13g2_fill_2 FILLER_45_269 ();
 sg13g2_fill_1 FILLER_45_271 ();
 sg13g2_decap_8 FILLER_45_295 ();
 sg13g2_fill_1 FILLER_45_302 ();
 sg13g2_fill_1 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_314 ();
 sg13g2_decap_4 FILLER_45_321 ();
 sg13g2_fill_2 FILLER_45_325 ();
 sg13g2_fill_2 FILLER_45_339 ();
 sg13g2_fill_2 FILLER_45_366 ();
 sg13g2_fill_1 FILLER_45_368 ();
 sg13g2_fill_1 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_389 ();
 sg13g2_decap_4 FILLER_45_404 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_4 FILLER_46_77 ();
 sg13g2_fill_2 FILLER_46_105 ();
 sg13g2_fill_2 FILLER_46_117 ();
 sg13g2_fill_1 FILLER_46_124 ();
 sg13g2_fill_2 FILLER_46_138 ();
 sg13g2_decap_4 FILLER_46_156 ();
 sg13g2_fill_2 FILLER_46_160 ();
 sg13g2_fill_2 FILLER_46_201 ();
 sg13g2_fill_1 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_230 ();
 sg13g2_decap_8 FILLER_46_237 ();
 sg13g2_decap_4 FILLER_46_244 ();
 sg13g2_fill_2 FILLER_46_248 ();
 sg13g2_fill_2 FILLER_46_277 ();
 sg13g2_fill_1 FILLER_46_279 ();
 sg13g2_fill_2 FILLER_46_285 ();
 sg13g2_fill_1 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_4 FILLER_46_336 ();
 sg13g2_fill_2 FILLER_46_354 ();
 sg13g2_fill_1 FILLER_46_356 ();
 sg13g2_fill_1 FILLER_46_367 ();
 sg13g2_fill_2 FILLER_46_392 ();
 sg13g2_fill_1 FILLER_46_394 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_fill_2 FILLER_47_70 ();
 sg13g2_fill_1 FILLER_47_72 ();
 sg13g2_fill_2 FILLER_47_83 ();
 sg13g2_fill_1 FILLER_47_85 ();
 sg13g2_fill_2 FILLER_47_109 ();
 sg13g2_fill_1 FILLER_47_111 ();
 sg13g2_decap_8 FILLER_47_128 ();
 sg13g2_decap_4 FILLER_47_135 ();
 sg13g2_fill_1 FILLER_47_139 ();
 sg13g2_fill_1 FILLER_47_151 ();
 sg13g2_fill_1 FILLER_47_163 ();
 sg13g2_fill_2 FILLER_47_178 ();
 sg13g2_fill_2 FILLER_47_190 ();
 sg13g2_fill_1 FILLER_47_192 ();
 sg13g2_fill_2 FILLER_47_202 ();
 sg13g2_fill_1 FILLER_47_204 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_fill_1 FILLER_47_280 ();
 sg13g2_fill_2 FILLER_47_286 ();
 sg13g2_fill_2 FILLER_47_297 ();
 sg13g2_fill_1 FILLER_47_299 ();
 sg13g2_decap_4 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_337 ();
 sg13g2_decap_4 FILLER_47_344 ();
 sg13g2_fill_2 FILLER_47_348 ();
 sg13g2_fill_1 FILLER_47_360 ();
 sg13g2_decap_4 FILLER_47_369 ();
 sg13g2_fill_2 FILLER_47_373 ();
 sg13g2_decap_8 FILLER_47_380 ();
 sg13g2_fill_1 FILLER_47_387 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_4 FILLER_48_70 ();
 sg13g2_fill_2 FILLER_48_74 ();
 sg13g2_fill_1 FILLER_48_96 ();
 sg13g2_decap_4 FILLER_48_113 ();
 sg13g2_decap_8 FILLER_48_121 ();
 sg13g2_fill_2 FILLER_48_128 ();
 sg13g2_fill_1 FILLER_48_130 ();
 sg13g2_fill_1 FILLER_48_154 ();
 sg13g2_fill_1 FILLER_48_161 ();
 sg13g2_fill_1 FILLER_48_171 ();
 sg13g2_fill_1 FILLER_48_176 ();
 sg13g2_decap_8 FILLER_48_186 ();
 sg13g2_fill_1 FILLER_48_193 ();
 sg13g2_decap_8 FILLER_48_227 ();
 sg13g2_decap_8 FILLER_48_234 ();
 sg13g2_decap_4 FILLER_48_241 ();
 sg13g2_decap_8 FILLER_48_250 ();
 sg13g2_fill_1 FILLER_48_257 ();
 sg13g2_decap_4 FILLER_48_272 ();
 sg13g2_decap_4 FILLER_48_296 ();
 sg13g2_fill_1 FILLER_48_300 ();
 sg13g2_fill_2 FILLER_48_317 ();
 sg13g2_fill_2 FILLER_48_340 ();
 sg13g2_fill_1 FILLER_48_346 ();
 sg13g2_decap_4 FILLER_48_352 ();
 sg13g2_fill_2 FILLER_48_356 ();
 sg13g2_decap_4 FILLER_48_363 ();
 sg13g2_fill_2 FILLER_48_367 ();
 sg13g2_decap_4 FILLER_48_373 ();
 sg13g2_fill_1 FILLER_48_377 ();
 sg13g2_fill_2 FILLER_48_383 ();
 sg13g2_fill_1 FILLER_48_385 ();
 sg13g2_fill_1 FILLER_48_394 ();
 sg13g2_fill_2 FILLER_48_407 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_93 ();
 sg13g2_decap_4 FILLER_49_100 ();
 sg13g2_fill_2 FILLER_49_104 ();
 sg13g2_fill_2 FILLER_49_120 ();
 sg13g2_fill_2 FILLER_49_127 ();
 sg13g2_fill_2 FILLER_49_134 ();
 sg13g2_decap_4 FILLER_49_141 ();
 sg13g2_decap_4 FILLER_49_150 ();
 sg13g2_decap_4 FILLER_49_160 ();
 sg13g2_fill_1 FILLER_49_164 ();
 sg13g2_decap_8 FILLER_49_173 ();
 sg13g2_decap_8 FILLER_49_180 ();
 sg13g2_decap_4 FILLER_49_187 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_210 ();
 sg13g2_fill_2 FILLER_49_217 ();
 sg13g2_fill_1 FILLER_49_219 ();
 sg13g2_fill_1 FILLER_49_246 ();
 sg13g2_decap_4 FILLER_49_252 ();
 sg13g2_fill_2 FILLER_49_256 ();
 sg13g2_decap_4 FILLER_49_269 ();
 sg13g2_fill_2 FILLER_49_273 ();
 sg13g2_fill_2 FILLER_49_293 ();
 sg13g2_fill_1 FILLER_49_295 ();
 sg13g2_fill_2 FILLER_49_304 ();
 sg13g2_fill_1 FILLER_49_306 ();
 sg13g2_fill_2 FILLER_49_360 ();
 sg13g2_fill_2 FILLER_49_375 ();
 sg13g2_decap_4 FILLER_49_403 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_fill_2 FILLER_50_77 ();
 sg13g2_fill_1 FILLER_50_79 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_4 FILLER_50_91 ();
 sg13g2_fill_2 FILLER_50_95 ();
 sg13g2_fill_2 FILLER_50_134 ();
 sg13g2_fill_1 FILLER_50_136 ();
 sg13g2_fill_2 FILLER_50_148 ();
 sg13g2_fill_2 FILLER_50_159 ();
 sg13g2_fill_1 FILLER_50_179 ();
 sg13g2_decap_8 FILLER_50_210 ();
 sg13g2_decap_8 FILLER_50_217 ();
 sg13g2_decap_8 FILLER_50_224 ();
 sg13g2_decap_8 FILLER_50_231 ();
 sg13g2_decap_8 FILLER_50_238 ();
 sg13g2_fill_1 FILLER_50_245 ();
 sg13g2_decap_8 FILLER_50_251 ();
 sg13g2_fill_2 FILLER_50_272 ();
 sg13g2_decap_4 FILLER_50_286 ();
 sg13g2_fill_1 FILLER_50_305 ();
 sg13g2_fill_2 FILLER_50_319 ();
 sg13g2_fill_2 FILLER_50_330 ();
 sg13g2_fill_1 FILLER_50_379 ();
 sg13g2_decap_4 FILLER_50_387 ();
 sg13g2_fill_2 FILLER_50_391 ();
 sg13g2_decap_8 FILLER_50_401 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_4 FILLER_51_63 ();
 sg13g2_fill_2 FILLER_51_104 ();
 sg13g2_fill_1 FILLER_51_106 ();
 sg13g2_fill_2 FILLER_51_123 ();
 sg13g2_fill_2 FILLER_51_132 ();
 sg13g2_fill_1 FILLER_51_134 ();
 sg13g2_fill_2 FILLER_51_140 ();
 sg13g2_fill_1 FILLER_51_142 ();
 sg13g2_fill_2 FILLER_51_151 ();
 sg13g2_fill_1 FILLER_51_166 ();
 sg13g2_fill_2 FILLER_51_190 ();
 sg13g2_decap_4 FILLER_51_243 ();
 sg13g2_fill_2 FILLER_51_257 ();
 sg13g2_fill_1 FILLER_51_282 ();
 sg13g2_decap_8 FILLER_51_296 ();
 sg13g2_decap_4 FILLER_51_303 ();
 sg13g2_fill_2 FILLER_51_307 ();
 sg13g2_decap_8 FILLER_51_314 ();
 sg13g2_decap_8 FILLER_51_321 ();
 sg13g2_fill_2 FILLER_51_328 ();
 sg13g2_fill_2 FILLER_51_333 ();
 sg13g2_fill_2 FILLER_51_339 ();
 sg13g2_fill_2 FILLER_51_367 ();
 sg13g2_fill_2 FILLER_51_388 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_fill_2 FILLER_52_63 ();
 sg13g2_fill_2 FILLER_52_109 ();
 sg13g2_decap_4 FILLER_52_118 ();
 sg13g2_fill_2 FILLER_52_130 ();
 sg13g2_fill_2 FILLER_52_142 ();
 sg13g2_fill_2 FILLER_52_156 ();
 sg13g2_fill_1 FILLER_52_158 ();
 sg13g2_fill_1 FILLER_52_184 ();
 sg13g2_decap_8 FILLER_52_239 ();
 sg13g2_decap_8 FILLER_52_246 ();
 sg13g2_fill_2 FILLER_52_253 ();
 sg13g2_fill_2 FILLER_52_270 ();
 sg13g2_fill_1 FILLER_52_272 ();
 sg13g2_fill_2 FILLER_52_284 ();
 sg13g2_fill_1 FILLER_52_295 ();
 sg13g2_decap_8 FILLER_52_300 ();
 sg13g2_decap_8 FILLER_52_307 ();
 sg13g2_fill_2 FILLER_52_314 ();
 sg13g2_fill_1 FILLER_52_316 ();
 sg13g2_fill_2 FILLER_52_333 ();
 sg13g2_fill_1 FILLER_52_335 ();
 sg13g2_decap_4 FILLER_52_340 ();
 sg13g2_fill_1 FILLER_52_344 ();
 sg13g2_decap_8 FILLER_52_353 ();
 sg13g2_fill_2 FILLER_52_360 ();
 sg13g2_fill_1 FILLER_52_362 ();
 sg13g2_fill_1 FILLER_52_368 ();
 sg13g2_decap_8 FILLER_52_372 ();
 sg13g2_decap_8 FILLER_52_379 ();
 sg13g2_fill_2 FILLER_52_386 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_fill_1 FILLER_53_56 ();
 sg13g2_fill_1 FILLER_53_87 ();
 sg13g2_fill_2 FILLER_53_110 ();
 sg13g2_fill_1 FILLER_53_112 ();
 sg13g2_fill_1 FILLER_53_131 ();
 sg13g2_decap_8 FILLER_53_147 ();
 sg13g2_decap_4 FILLER_53_154 ();
 sg13g2_fill_1 FILLER_53_158 ();
 sg13g2_decap_8 FILLER_53_183 ();
 sg13g2_decap_8 FILLER_53_190 ();
 sg13g2_decap_4 FILLER_53_217 ();
 sg13g2_decap_8 FILLER_53_255 ();
 sg13g2_decap_4 FILLER_53_262 ();
 sg13g2_fill_2 FILLER_53_266 ();
 sg13g2_fill_1 FILLER_53_273 ();
 sg13g2_fill_2 FILLER_53_287 ();
 sg13g2_fill_1 FILLER_53_289 ();
 sg13g2_fill_1 FILLER_53_298 ();
 sg13g2_fill_2 FILLER_53_309 ();
 sg13g2_fill_1 FILLER_53_331 ();
 sg13g2_fill_2 FILLER_53_337 ();
 sg13g2_fill_1 FILLER_53_339 ();
 sg13g2_fill_2 FILLER_53_345 ();
 sg13g2_fill_1 FILLER_53_347 ();
 sg13g2_decap_8 FILLER_53_353 ();
 sg13g2_fill_2 FILLER_53_360 ();
 sg13g2_fill_1 FILLER_53_362 ();
 sg13g2_fill_2 FILLER_53_386 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_4 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_85 ();
 sg13g2_decap_4 FILLER_54_92 ();
 sg13g2_fill_1 FILLER_54_96 ();
 sg13g2_decap_8 FILLER_54_135 ();
 sg13g2_decap_8 FILLER_54_142 ();
 sg13g2_fill_1 FILLER_54_149 ();
 sg13g2_decap_4 FILLER_54_167 ();
 sg13g2_decap_8 FILLER_54_175 ();
 sg13g2_decap_4 FILLER_54_182 ();
 sg13g2_fill_2 FILLER_54_186 ();
 sg13g2_decap_4 FILLER_54_195 ();
 sg13g2_fill_2 FILLER_54_199 ();
 sg13g2_decap_8 FILLER_54_206 ();
 sg13g2_fill_1 FILLER_54_213 ();
 sg13g2_decap_8 FILLER_54_245 ();
 sg13g2_decap_8 FILLER_54_252 ();
 sg13g2_fill_2 FILLER_54_259 ();
 sg13g2_fill_1 FILLER_54_261 ();
 sg13g2_decap_8 FILLER_54_266 ();
 sg13g2_decap_8 FILLER_54_273 ();
 sg13g2_fill_1 FILLER_54_280 ();
 sg13g2_fill_2 FILLER_54_301 ();
 sg13g2_fill_1 FILLER_54_331 ();
 sg13g2_fill_2 FILLER_54_345 ();
 sg13g2_fill_2 FILLER_54_361 ();
 sg13g2_fill_2 FILLER_54_369 ();
 sg13g2_fill_2 FILLER_54_388 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_4 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_78 ();
 sg13g2_decap_4 FILLER_55_85 ();
 sg13g2_decap_8 FILLER_55_107 ();
 sg13g2_decap_8 FILLER_55_114 ();
 sg13g2_fill_2 FILLER_55_125 ();
 sg13g2_fill_1 FILLER_55_127 ();
 sg13g2_decap_8 FILLER_55_136 ();
 sg13g2_decap_8 FILLER_55_143 ();
 sg13g2_decap_8 FILLER_55_150 ();
 sg13g2_decap_8 FILLER_55_157 ();
 sg13g2_fill_2 FILLER_55_164 ();
 sg13g2_fill_1 FILLER_55_166 ();
 sg13g2_decap_8 FILLER_55_211 ();
 sg13g2_decap_8 FILLER_55_218 ();
 sg13g2_fill_2 FILLER_55_233 ();
 sg13g2_fill_1 FILLER_55_235 ();
 sg13g2_decap_8 FILLER_55_275 ();
 sg13g2_decap_4 FILLER_55_282 ();
 sg13g2_fill_2 FILLER_55_286 ();
 sg13g2_fill_1 FILLER_55_293 ();
 sg13g2_fill_2 FILLER_55_316 ();
 sg13g2_fill_2 FILLER_55_323 ();
 sg13g2_fill_1 FILLER_55_325 ();
 sg13g2_fill_1 FILLER_55_334 ();
 sg13g2_fill_2 FILLER_55_345 ();
 sg13g2_fill_1 FILLER_55_347 ();
 sg13g2_fill_1 FILLER_55_353 ();
 sg13g2_fill_2 FILLER_55_360 ();
 sg13g2_fill_2 FILLER_55_391 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_fill_2 FILLER_56_77 ();
 sg13g2_fill_1 FILLER_56_79 ();
 sg13g2_fill_2 FILLER_56_92 ();
 sg13g2_fill_1 FILLER_56_94 ();
 sg13g2_decap_4 FILLER_56_111 ();
 sg13g2_fill_1 FILLER_56_125 ();
 sg13g2_fill_2 FILLER_56_135 ();
 sg13g2_fill_1 FILLER_56_137 ();
 sg13g2_fill_2 FILLER_56_146 ();
 sg13g2_decap_4 FILLER_56_177 ();
 sg13g2_fill_1 FILLER_56_181 ();
 sg13g2_decap_8 FILLER_56_208 ();
 sg13g2_decap_8 FILLER_56_227 ();
 sg13g2_fill_2 FILLER_56_234 ();
 sg13g2_fill_2 FILLER_56_281 ();
 sg13g2_decap_8 FILLER_56_288 ();
 sg13g2_decap_8 FILLER_56_295 ();
 sg13g2_decap_4 FILLER_56_302 ();
 sg13g2_fill_1 FILLER_56_306 ();
 sg13g2_fill_1 FILLER_56_351 ();
 sg13g2_fill_2 FILLER_56_360 ();
 sg13g2_decap_8 FILLER_56_374 ();
 sg13g2_decap_4 FILLER_56_381 ();
 sg13g2_fill_2 FILLER_56_393 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_fill_1 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_4 FILLER_57_111 ();
 sg13g2_fill_2 FILLER_57_136 ();
 sg13g2_decap_8 FILLER_57_146 ();
 sg13g2_decap_4 FILLER_57_153 ();
 sg13g2_fill_2 FILLER_57_157 ();
 sg13g2_fill_2 FILLER_57_170 ();
 sg13g2_fill_1 FILLER_57_172 ();
 sg13g2_fill_1 FILLER_57_191 ();
 sg13g2_fill_1 FILLER_57_196 ();
 sg13g2_decap_8 FILLER_57_205 ();
 sg13g2_fill_1 FILLER_57_212 ();
 sg13g2_decap_8 FILLER_57_245 ();
 sg13g2_decap_4 FILLER_57_257 ();
 sg13g2_decap_4 FILLER_57_274 ();
 sg13g2_decap_8 FILLER_57_293 ();
 sg13g2_fill_1 FILLER_57_300 ();
 sg13g2_fill_1 FILLER_57_308 ();
 sg13g2_decap_8 FILLER_57_317 ();
 sg13g2_decap_8 FILLER_57_332 ();
 sg13g2_decap_4 FILLER_57_339 ();
 sg13g2_fill_2 FILLER_57_343 ();
 sg13g2_decap_4 FILLER_57_349 ();
 sg13g2_fill_1 FILLER_57_353 ();
 sg13g2_decap_4 FILLER_57_358 ();
 sg13g2_fill_2 FILLER_57_362 ();
 sg13g2_decap_8 FILLER_57_368 ();
 sg13g2_decap_8 FILLER_57_375 ();
 sg13g2_fill_2 FILLER_57_394 ();
 sg13g2_fill_1 FILLER_57_396 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_4 FILLER_58_63 ();
 sg13g2_fill_1 FILLER_58_92 ();
 sg13g2_fill_2 FILLER_58_103 ();
 sg13g2_fill_1 FILLER_58_105 ();
 sg13g2_fill_1 FILLER_58_118 ();
 sg13g2_decap_4 FILLER_58_123 ();
 sg13g2_decap_8 FILLER_58_132 ();
 sg13g2_fill_2 FILLER_58_139 ();
 sg13g2_fill_2 FILLER_58_167 ();
 sg13g2_fill_2 FILLER_58_190 ();
 sg13g2_fill_1 FILLER_58_192 ();
 sg13g2_decap_4 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_225 ();
 sg13g2_fill_2 FILLER_58_258 ();
 sg13g2_fill_1 FILLER_58_260 ();
 sg13g2_decap_4 FILLER_58_271 ();
 sg13g2_fill_2 FILLER_58_275 ();
 sg13g2_fill_1 FILLER_58_284 ();
 sg13g2_decap_4 FILLER_58_295 ();
 sg13g2_fill_1 FILLER_58_299 ();
 sg13g2_fill_1 FILLER_58_325 ();
 sg13g2_decap_8 FILLER_58_348 ();
 sg13g2_fill_2 FILLER_58_355 ();
 sg13g2_decap_4 FILLER_58_363 ();
 sg13g2_fill_1 FILLER_58_376 ();
 sg13g2_decap_4 FILLER_58_384 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_4 FILLER_59_63 ();
 sg13g2_fill_2 FILLER_59_67 ();
 sg13g2_decap_4 FILLER_59_96 ();
 sg13g2_fill_2 FILLER_59_100 ();
 sg13g2_fill_2 FILLER_59_115 ();
 sg13g2_fill_2 FILLER_59_139 ();
 sg13g2_decap_8 FILLER_59_146 ();
 sg13g2_decap_8 FILLER_59_153 ();
 sg13g2_fill_2 FILLER_59_160 ();
 sg13g2_fill_1 FILLER_59_162 ();
 sg13g2_decap_8 FILLER_59_166 ();
 sg13g2_decap_4 FILLER_59_193 ();
 sg13g2_fill_1 FILLER_59_197 ();
 sg13g2_decap_8 FILLER_59_201 ();
 sg13g2_decap_4 FILLER_59_208 ();
 sg13g2_fill_1 FILLER_59_212 ();
 sg13g2_fill_1 FILLER_59_225 ();
 sg13g2_decap_4 FILLER_59_229 ();
 sg13g2_fill_2 FILLER_59_233 ();
 sg13g2_fill_2 FILLER_59_266 ();
 sg13g2_fill_1 FILLER_59_268 ();
 sg13g2_fill_2 FILLER_59_276 ();
 sg13g2_fill_1 FILLER_59_278 ();
 sg13g2_fill_1 FILLER_59_284 ();
 sg13g2_fill_2 FILLER_59_301 ();
 sg13g2_fill_1 FILLER_59_328 ();
 sg13g2_fill_1 FILLER_59_389 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_4 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_86 ();
 sg13g2_fill_2 FILLER_60_93 ();
 sg13g2_fill_1 FILLER_60_95 ();
 sg13g2_fill_2 FILLER_60_142 ();
 sg13g2_fill_2 FILLER_60_173 ();
 sg13g2_decap_4 FILLER_60_186 ();
 sg13g2_fill_2 FILLER_60_190 ();
 sg13g2_fill_2 FILLER_60_209 ();
 sg13g2_fill_1 FILLER_60_211 ();
 sg13g2_decap_4 FILLER_60_227 ();
 sg13g2_fill_2 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_238 ();
 sg13g2_decap_8 FILLER_60_245 ();
 sg13g2_decap_8 FILLER_60_252 ();
 sg13g2_decap_4 FILLER_60_264 ();
 sg13g2_fill_1 FILLER_60_273 ();
 sg13g2_decap_8 FILLER_60_298 ();
 sg13g2_decap_8 FILLER_60_305 ();
 sg13g2_fill_1 FILLER_60_312 ();
 sg13g2_fill_1 FILLER_60_334 ();
 sg13g2_fill_2 FILLER_60_340 ();
 sg13g2_fill_2 FILLER_60_372 ();
 sg13g2_decap_8 FILLER_60_379 ();
 sg13g2_decap_8 FILLER_60_386 ();
 sg13g2_fill_2 FILLER_60_393 ();
 sg13g2_decap_8 FILLER_60_399 ();
 sg13g2_fill_2 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_4 FILLER_61_91 ();
 sg13g2_decap_4 FILLER_61_121 ();
 sg13g2_fill_2 FILLER_61_125 ();
 sg13g2_fill_2 FILLER_61_132 ();
 sg13g2_fill_2 FILLER_61_138 ();
 sg13g2_decap_4 FILLER_61_149 ();
 sg13g2_fill_2 FILLER_61_179 ();
 sg13g2_fill_1 FILLER_61_181 ();
 sg13g2_fill_2 FILLER_61_197 ();
 sg13g2_fill_1 FILLER_61_199 ();
 sg13g2_fill_1 FILLER_61_212 ();
 sg13g2_fill_1 FILLER_61_237 ();
 sg13g2_decap_8 FILLER_61_264 ();
 sg13g2_fill_2 FILLER_61_271 ();
 sg13g2_decap_8 FILLER_61_301 ();
 sg13g2_decap_8 FILLER_61_308 ();
 sg13g2_decap_8 FILLER_61_315 ();
 sg13g2_fill_2 FILLER_61_322 ();
 sg13g2_fill_1 FILLER_61_324 ();
 sg13g2_fill_2 FILLER_61_336 ();
 sg13g2_fill_2 FILLER_61_371 ();
 sg13g2_fill_1 FILLER_61_393 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_fill_2 FILLER_62_63 ();
 sg13g2_fill_1 FILLER_62_83 ();
 sg13g2_fill_1 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_108 ();
 sg13g2_decap_8 FILLER_62_115 ();
 sg13g2_fill_2 FILLER_62_172 ();
 sg13g2_fill_1 FILLER_62_174 ();
 sg13g2_fill_2 FILLER_62_222 ();
 sg13g2_decap_8 FILLER_62_252 ();
 sg13g2_decap_8 FILLER_62_259 ();
 sg13g2_fill_1 FILLER_62_266 ();
 sg13g2_decap_8 FILLER_62_311 ();
 sg13g2_decap_8 FILLER_62_318 ();
 sg13g2_decap_4 FILLER_62_325 ();
 sg13g2_fill_1 FILLER_62_329 ();
 sg13g2_decap_8 FILLER_62_335 ();
 sg13g2_fill_2 FILLER_62_342 ();
 sg13g2_fill_1 FILLER_62_344 ();
 sg13g2_fill_2 FILLER_62_364 ();
 sg13g2_fill_1 FILLER_62_366 ();
 sg13g2_fill_2 FILLER_62_372 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_fill_1 FILLER_63_85 ();
 sg13g2_decap_8 FILLER_63_92 ();
 sg13g2_decap_8 FILLER_63_99 ();
 sg13g2_decap_8 FILLER_63_106 ();
 sg13g2_decap_8 FILLER_63_113 ();
 sg13g2_decap_4 FILLER_63_120 ();
 sg13g2_fill_2 FILLER_63_124 ();
 sg13g2_decap_8 FILLER_63_146 ();
 sg13g2_decap_8 FILLER_63_153 ();
 sg13g2_decap_8 FILLER_63_160 ();
 sg13g2_decap_8 FILLER_63_167 ();
 sg13g2_decap_4 FILLER_63_174 ();
 sg13g2_fill_1 FILLER_63_178 ();
 sg13g2_decap_4 FILLER_63_182 ();
 sg13g2_fill_2 FILLER_63_186 ();
 sg13g2_decap_8 FILLER_63_200 ();
 sg13g2_fill_2 FILLER_63_216 ();
 sg13g2_fill_1 FILLER_63_233 ();
 sg13g2_fill_2 FILLER_63_277 ();
 sg13g2_fill_1 FILLER_63_279 ();
 sg13g2_fill_1 FILLER_63_294 ();
 sg13g2_fill_1 FILLER_63_308 ();
 sg13g2_fill_1 FILLER_63_318 ();
 sg13g2_fill_1 FILLER_63_330 ();
 sg13g2_decap_8 FILLER_63_342 ();
 sg13g2_fill_2 FILLER_63_349 ();
 sg13g2_fill_1 FILLER_63_351 ();
 sg13g2_fill_1 FILLER_63_377 ();
 sg13g2_fill_2 FILLER_63_386 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_4 FILLER_64_63 ();
 sg13g2_fill_1 FILLER_64_67 ();
 sg13g2_fill_1 FILLER_64_83 ();
 sg13g2_fill_1 FILLER_64_91 ();
 sg13g2_fill_2 FILLER_64_117 ();
 sg13g2_decap_8 FILLER_64_129 ();
 sg13g2_fill_1 FILLER_64_136 ();
 sg13g2_decap_8 FILLER_64_141 ();
 sg13g2_fill_1 FILLER_64_148 ();
 sg13g2_fill_1 FILLER_64_179 ();
 sg13g2_fill_2 FILLER_64_193 ();
 sg13g2_fill_1 FILLER_64_195 ();
 sg13g2_fill_1 FILLER_64_233 ();
 sg13g2_fill_1 FILLER_64_243 ();
 sg13g2_fill_2 FILLER_64_300 ();
 sg13g2_fill_1 FILLER_64_327 ();
 sg13g2_decap_8 FILLER_64_340 ();
 sg13g2_decap_8 FILLER_64_347 ();
 sg13g2_decap_8 FILLER_64_367 ();
 sg13g2_fill_1 FILLER_64_374 ();
 sg13g2_decap_4 FILLER_64_390 ();
 sg13g2_fill_1 FILLER_64_394 ();
 sg13g2_decap_4 FILLER_64_404 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_fill_1 FILLER_65_98 ();
 sg13g2_fill_2 FILLER_65_110 ();
 sg13g2_fill_1 FILLER_65_133 ();
 sg13g2_fill_2 FILLER_65_141 ();
 sg13g2_fill_1 FILLER_65_143 ();
 sg13g2_decap_4 FILLER_65_154 ();
 sg13g2_fill_1 FILLER_65_189 ();
 sg13g2_decap_4 FILLER_65_256 ();
 sg13g2_fill_1 FILLER_65_308 ();
 sg13g2_fill_1 FILLER_65_315 ();
 sg13g2_fill_1 FILLER_65_322 ();
 sg13g2_fill_1 FILLER_65_348 ();
 sg13g2_decap_4 FILLER_65_361 ();
 sg13g2_fill_2 FILLER_65_365 ();
 sg13g2_fill_2 FILLER_65_378 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_4 FILLER_66_84 ();
 sg13g2_fill_2 FILLER_66_88 ();
 sg13g2_fill_2 FILLER_66_120 ();
 sg13g2_fill_1 FILLER_66_128 ();
 sg13g2_fill_1 FILLER_66_139 ();
 sg13g2_decap_8 FILLER_66_176 ();
 sg13g2_fill_2 FILLER_66_183 ();
 sg13g2_fill_1 FILLER_66_201 ();
 sg13g2_fill_1 FILLER_66_207 ();
 sg13g2_decap_8 FILLER_66_248 ();
 sg13g2_decap_8 FILLER_66_255 ();
 sg13g2_decap_8 FILLER_66_262 ();
 sg13g2_fill_1 FILLER_66_269 ();
 sg13g2_fill_2 FILLER_66_274 ();
 sg13g2_fill_1 FILLER_66_276 ();
 sg13g2_fill_2 FILLER_66_303 ();
 sg13g2_decap_8 FILLER_66_323 ();
 sg13g2_fill_2 FILLER_66_330 ();
 sg13g2_decap_8 FILLER_66_338 ();
 sg13g2_decap_8 FILLER_66_345 ();
 sg13g2_fill_2 FILLER_66_352 ();
 sg13g2_fill_1 FILLER_66_354 ();
 sg13g2_fill_2 FILLER_66_389 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_fill_2 FILLER_67_70 ();
 sg13g2_fill_2 FILLER_67_110 ();
 sg13g2_fill_1 FILLER_67_142 ();
 sg13g2_decap_4 FILLER_67_169 ();
 sg13g2_fill_2 FILLER_67_173 ();
 sg13g2_fill_1 FILLER_67_203 ();
 sg13g2_fill_1 FILLER_67_218 ();
 sg13g2_decap_8 FILLER_67_232 ();
 sg13g2_fill_2 FILLER_67_239 ();
 sg13g2_fill_2 FILLER_67_246 ();
 sg13g2_decap_8 FILLER_67_274 ();
 sg13g2_decap_8 FILLER_67_281 ();
 sg13g2_decap_4 FILLER_67_288 ();
 sg13g2_fill_1 FILLER_67_292 ();
 sg13g2_fill_1 FILLER_67_314 ();
 sg13g2_decap_4 FILLER_67_351 ();
 sg13g2_fill_2 FILLER_67_355 ();
 sg13g2_fill_2 FILLER_67_365 ();
 sg13g2_fill_1 FILLER_67_367 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_fill_1 FILLER_68_84 ();
 sg13g2_fill_1 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_141 ();
 sg13g2_decap_8 FILLER_68_148 ();
 sg13g2_fill_1 FILLER_68_155 ();
 sg13g2_decap_8 FILLER_68_161 ();
 sg13g2_decap_8 FILLER_68_168 ();
 sg13g2_fill_2 FILLER_68_182 ();
 sg13g2_fill_1 FILLER_68_184 ();
 sg13g2_fill_2 FILLER_68_210 ();
 sg13g2_decap_8 FILLER_68_221 ();
 sg13g2_fill_1 FILLER_68_228 ();
 sg13g2_fill_2 FILLER_68_243 ();
 sg13g2_fill_1 FILLER_68_245 ();
 sg13g2_fill_2 FILLER_68_272 ();
 sg13g2_decap_4 FILLER_68_300 ();
 sg13g2_fill_2 FILLER_68_304 ();
 sg13g2_fill_2 FILLER_68_332 ();
 sg13g2_fill_2 FILLER_68_365 ();
 sg13g2_decap_4 FILLER_68_377 ();
 sg13g2_fill_1 FILLER_68_381 ();
 sg13g2_decap_8 FILLER_68_387 ();
 sg13g2_decap_4 FILLER_68_394 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_fill_2 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_95 ();
 sg13g2_decap_8 FILLER_69_102 ();
 sg13g2_decap_4 FILLER_69_109 ();
 sg13g2_fill_1 FILLER_69_113 ();
 sg13g2_fill_2 FILLER_69_118 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_4 FILLER_69_138 ();
 sg13g2_fill_2 FILLER_69_142 ();
 sg13g2_fill_1 FILLER_69_147 ();
 sg13g2_decap_4 FILLER_69_153 ();
 sg13g2_fill_1 FILLER_69_157 ();
 sg13g2_fill_1 FILLER_69_200 ();
 sg13g2_decap_4 FILLER_69_210 ();
 sg13g2_fill_1 FILLER_69_214 ();
 sg13g2_fill_2 FILLER_69_220 ();
 sg13g2_fill_1 FILLER_69_222 ();
 sg13g2_decap_8 FILLER_69_254 ();
 sg13g2_decap_8 FILLER_69_261 ();
 sg13g2_decap_4 FILLER_69_268 ();
 sg13g2_decap_8 FILLER_69_298 ();
 sg13g2_fill_2 FILLER_69_320 ();
 sg13g2_decap_8 FILLER_69_378 ();
 sg13g2_decap_8 FILLER_69_385 ();
 sg13g2_decap_8 FILLER_69_392 ();
 sg13g2_decap_8 FILLER_69_399 ();
 sg13g2_fill_2 FILLER_69_406 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_4 FILLER_70_77 ();
 sg13g2_fill_2 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_107 ();
 sg13g2_decap_8 FILLER_70_114 ();
 sg13g2_decap_8 FILLER_70_125 ();
 sg13g2_fill_1 FILLER_70_139 ();
 sg13g2_fill_1 FILLER_70_196 ();
 sg13g2_fill_2 FILLER_70_256 ();
 sg13g2_fill_2 FILLER_70_273 ();
 sg13g2_decap_4 FILLER_70_289 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_4 FILLER_71_77 ();
 sg13g2_fill_1 FILLER_71_89 ();
 sg13g2_fill_2 FILLER_71_118 ();
 sg13g2_fill_1 FILLER_71_120 ();
 sg13g2_fill_2 FILLER_71_126 ();
 sg13g2_fill_2 FILLER_71_201 ();
 sg13g2_decap_8 FILLER_71_238 ();
 sg13g2_fill_1 FILLER_71_271 ();
 sg13g2_decap_8 FILLER_71_298 ();
 sg13g2_fill_2 FILLER_71_305 ();
 sg13g2_fill_1 FILLER_71_312 ();
 sg13g2_fill_1 FILLER_71_377 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_4 FILLER_72_77 ();
 sg13g2_fill_2 FILLER_72_147 ();
 sg13g2_fill_1 FILLER_72_157 ();
 sg13g2_decap_8 FILLER_72_173 ();
 sg13g2_fill_1 FILLER_72_242 ();
 sg13g2_fill_1 FILLER_72_251 ();
 sg13g2_decap_4 FILLER_72_267 ();
 sg13g2_fill_1 FILLER_72_297 ();
 sg13g2_fill_2 FILLER_72_346 ();
 sg13g2_decap_4 FILLER_72_374 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_4 FILLER_73_77 ();
 sg13g2_fill_1 FILLER_73_81 ();
 sg13g2_fill_1 FILLER_73_111 ();
 sg13g2_fill_2 FILLER_73_149 ();
 sg13g2_decap_4 FILLER_73_238 ();
 sg13g2_fill_2 FILLER_73_242 ();
 sg13g2_decap_8 FILLER_73_275 ();
 sg13g2_fill_2 FILLER_73_282 ();
 sg13g2_fill_2 FILLER_73_367 ();
 sg13g2_fill_1 FILLER_73_377 ();
 sg13g2_decap_4 FILLER_73_388 ();
 sg13g2_fill_1 FILLER_73_392 ();
 sg13g2_decap_8 FILLER_73_402 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_fill_2 FILLER_74_91 ();
 sg13g2_fill_2 FILLER_74_131 ();
 sg13g2_decap_8 FILLER_74_149 ();
 sg13g2_decap_8 FILLER_74_156 ();
 sg13g2_decap_8 FILLER_74_163 ();
 sg13g2_fill_1 FILLER_74_170 ();
 sg13g2_fill_1 FILLER_74_236 ();
 sg13g2_decap_8 FILLER_74_245 ();
 sg13g2_decap_4 FILLER_74_252 ();
 sg13g2_fill_2 FILLER_74_256 ();
 sg13g2_decap_8 FILLER_74_277 ();
 sg13g2_fill_1 FILLER_74_320 ();
 sg13g2_decap_4 FILLER_74_347 ();
 sg13g2_fill_1 FILLER_74_377 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_fill_1 FILLER_75_98 ();
 sg13g2_decap_4 FILLER_75_103 ();
 sg13g2_fill_2 FILLER_75_116 ();
 sg13g2_decap_8 FILLER_75_127 ();
 sg13g2_decap_8 FILLER_75_134 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_fill_2 FILLER_75_182 ();
 sg13g2_fill_1 FILLER_75_184 ();
 sg13g2_decap_8 FILLER_75_238 ();
 sg13g2_fill_1 FILLER_75_245 ();
 sg13g2_fill_1 FILLER_75_272 ();
 sg13g2_decap_8 FILLER_75_296 ();
 sg13g2_decap_4 FILLER_75_303 ();
 sg13g2_fill_2 FILLER_75_307 ();
 sg13g2_fill_2 FILLER_75_314 ();
 sg13g2_fill_1 FILLER_75_316 ();
 sg13g2_decap_4 FILLER_75_322 ();
 sg13g2_fill_1 FILLER_75_326 ();
 sg13g2_fill_1 FILLER_75_337 ();
 sg13g2_fill_2 FILLER_75_347 ();
 sg13g2_fill_1 FILLER_75_349 ();
 sg13g2_fill_2 FILLER_75_369 ();
 sg13g2_fill_1 FILLER_75_371 ();
 sg13g2_fill_2 FILLER_75_381 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_fill_1 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_117 ();
 sg13g2_decap_8 FILLER_76_124 ();
 sg13g2_fill_2 FILLER_76_131 ();
 sg13g2_fill_2 FILLER_76_162 ();
 sg13g2_fill_1 FILLER_76_164 ();
 sg13g2_fill_1 FILLER_76_170 ();
 sg13g2_fill_2 FILLER_76_197 ();
 sg13g2_fill_1 FILLER_76_199 ();
 sg13g2_fill_1 FILLER_76_210 ();
 sg13g2_fill_1 FILLER_76_237 ();
 sg13g2_fill_2 FILLER_76_266 ();
 sg13g2_fill_1 FILLER_76_268 ();
 sg13g2_fill_2 FILLER_76_298 ();
 sg13g2_fill_2 FILLER_76_319 ();
 sg13g2_fill_1 FILLER_76_321 ();
 sg13g2_fill_1 FILLER_76_348 ();
 sg13g2_fill_1 FILLER_76_362 ();
 sg13g2_decap_4 FILLER_76_403 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_fill_2 FILLER_77_126 ();
 sg13g2_fill_1 FILLER_77_128 ();
 sg13g2_fill_2 FILLER_77_158 ();
 sg13g2_fill_2 FILLER_77_258 ();
 sg13g2_fill_1 FILLER_77_304 ();
 sg13g2_fill_1 FILLER_77_367 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_fill_1 FILLER_78_144 ();
 sg13g2_decap_4 FILLER_78_196 ();
 sg13g2_fill_1 FILLER_78_209 ();
 sg13g2_decap_8 FILLER_78_236 ();
 sg13g2_fill_1 FILLER_78_243 ();
 sg13g2_fill_1 FILLER_78_270 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_fill_2 FILLER_79_133 ();
 sg13g2_fill_1 FILLER_79_135 ();
 sg13g2_fill_2 FILLER_79_144 ();
 sg13g2_fill_2 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_173 ();
 sg13g2_fill_2 FILLER_79_180 ();
 sg13g2_fill_1 FILLER_79_182 ();
 sg13g2_fill_2 FILLER_79_209 ();
 sg13g2_fill_2 FILLER_79_267 ();
 sg13g2_fill_1 FILLER_79_269 ();
 sg13g2_fill_2 FILLER_79_340 ();
 sg13g2_fill_2 FILLER_79_355 ();
 sg13g2_fill_1 FILLER_79_357 ();
 sg13g2_fill_2 FILLER_79_367 ();
 sg13g2_decap_4 FILLER_79_403 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_fill_2 FILLER_80_148 ();
 sg13g2_fill_1 FILLER_80_159 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_fill_2 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_4 FILLER_80_215 ();
 sg13g2_fill_2 FILLER_80_246 ();
 sg13g2_fill_2 FILLER_80_261 ();
 sg13g2_fill_1 FILLER_80_268 ();
 sg13g2_fill_1 FILLER_80_304 ();
 sg13g2_fill_2 FILLER_80_315 ();
 sg13g2_fill_2 FILLER_80_352 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net25;
 assign uio_out[1] = net26;
 assign uio_out[2] = net27;
 assign uio_out[3] = net28;
 assign uio_out[4] = net29;
 assign uio_out[5] = net30;
 assign uio_out[6] = net31;
 assign uio_out[7] = net32;
endmodule

module tt_um_edwintorok (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire audio;
 wire \generated._1000[0] ;
 wire \generated._100[0] ;
 wire \generated._100[1] ;
 wire \generated._100[2] ;
 wire \generated._100[3] ;
 wire \generated._100[4] ;
 wire \generated._100[5] ;
 wire \generated._100[6] ;
 wire \generated._100[7] ;
 wire \generated._100[8] ;
 wire \generated._100[9] ;
 wire \generated._1023[3] ;
 wire \generated._1023[4] ;
 wire \generated._1023[5] ;
 wire \generated._1023[6] ;
 wire \generated._1023[7] ;
 wire \generated._1023[8] ;
 wire \generated._1023[9] ;
 wire \generated._1024[0] ;
 wire \generated._1024[1] ;
 wire \generated._1024[2] ;
 wire \generated._1024[3] ;
 wire \generated._1024[4] ;
 wire \generated._1024[5] ;
 wire \generated._1024[6] ;
 wire \generated._1024[7] ;
 wire \generated._1024[8] ;
 wire \generated._1024[9] ;
 wire \generated._1025[0] ;
 wire \generated._1073[3] ;
 wire \generated._1073[4] ;
 wire \generated._1073[5] ;
 wire \generated._1073[6] ;
 wire \generated._1073[7] ;
 wire \generated._1073[8] ;
 wire \generated._1073[9] ;
 wire \generated._1074[0] ;
 wire \generated._1074[1] ;
 wire \generated._1074[2] ;
 wire \generated._1074[3] ;
 wire \generated._1074[4] ;
 wire \generated._1074[5] ;
 wire \generated._1074[6] ;
 wire \generated._1074[7] ;
 wire \generated._1074[8] ;
 wire \generated._1074[9] ;
 wire \generated._1076[0] ;
 wire \generated._1078[0] ;
 wire \generated._1078[1] ;
 wire \generated._1078[2] ;
 wire \generated._1078[3] ;
 wire \generated._1084[0] ;
 wire \generated._1084[1] ;
 wire \generated._1084[2] ;
 wire \generated._1084[3] ;
 wire \generated._1084[4] ;
 wire \generated._1084[5] ;
 wire \generated._1084[6] ;
 wire \generated._1084[7] ;
 wire \generated._1084[8] ;
 wire \generated._1084[9] ;
 wire \generated._1087[0] ;
 wire \generated._1118[0] ;
 wire \generated._1148[0] ;
 wire \generated._115 ;
 wire \generated._123 ;
 wire \generated._165[4] ;
 wire \generated._16[0] ;
 wire \generated._16[1] ;
 wire \generated._16[2] ;
 wire \generated._16[3] ;
 wire \generated._16[4] ;
 wire \generated._21[0] ;
 wire \generated._21[1] ;
 wire \generated._21[2] ;
 wire \generated._21[3] ;
 wire \generated._21[4] ;
 wire \generated._221[0] ;
 wire \generated._221[1] ;
 wire \generated._221[2] ;
 wire \generated._221[3] ;
 wire \generated._28[0] ;
 wire \generated._28[1] ;
 wire \generated._28[2] ;
 wire \generated._28[3] ;
 wire \generated._301[0] ;
 wire \generated._328[0] ;
 wire \generated._33[0] ;
 wire \generated._33[1] ;
 wire \generated._33[2] ;
 wire \generated._33[3] ;
 wire \generated._33[4] ;
 wire \generated._33[5] ;
 wire \generated._33[6] ;
 wire \generated._346[0] ;
 wire \generated._346[1] ;
 wire \generated._346[2] ;
 wire \generated._346[3] ;
 wire \generated._346[4] ;
 wire \generated._346[5] ;
 wire \generated._353[0] ;
 wire \generated._357[0] ;
 wire \generated._357[1] ;
 wire \generated._357[2] ;
 wire \generated._357[3] ;
 wire \generated._357[4] ;
 wire \generated._371 ;
 wire \generated._373[0] ;
 wire \generated._373[1] ;
 wire \generated._373[2] ;
 wire \generated._373[3] ;
 wire \generated._373[4] ;
 wire \generated._373[5] ;
 wire \generated._373[6] ;
 wire \generated._373[7] ;
 wire \generated._373[8] ;
 wire \generated._378 ;
 wire \generated._379 ;
 wire \generated._380 ;
 wire \generated._381[0] ;
 wire \generated._381[1] ;
 wire \generated._381[2] ;
 wire \generated._381[3] ;
 wire \generated._381[4] ;
 wire \generated._381[5] ;
 wire \generated._381[6] ;
 wire \generated._381[7] ;
 wire \generated._394[0] ;
 wire \generated._394[1] ;
 wire \generated._394[2] ;
 wire \generated._394[3] ;
 wire \generated._394[4] ;
 wire \generated._394[5] ;
 wire \generated._394[6] ;
 wire \generated._394[7] ;
 wire \generated._394[8] ;
 wire \generated._394[9] ;
 wire \generated._395[0] ;
 wire \generated._406[1] ;
 wire \generated._406[2] ;
 wire \generated._406[3] ;
 wire \generated._406[4] ;
 wire \generated._406[5] ;
 wire \generated._406[6] ;
 wire \generated._406[7] ;
 wire \generated._425[1] ;
 wire \generated._434[10] ;
 wire \generated._434[11] ;
 wire \generated._434[12] ;
 wire \generated._434[13] ;
 wire \generated._434[14] ;
 wire \generated._434[15] ;
 wire \generated._434[16] ;
 wire \generated._434[17] ;
 wire \generated._434[18] ;
 wire \generated._434[19] ;
 wire \generated._481[0] ;
 wire \generated._481[1] ;
 wire \generated._481[2] ;
 wire \generated._481[3] ;
 wire \generated._481[4] ;
 wire \generated._481[5] ;
 wire \generated._481[6] ;
 wire \generated._481[7] ;
 wire \generated._481[8] ;
 wire \generated._481[9] ;
 wire \generated._485[0] ;
 wire \generated._487[0] ;
 wire \generated._487[1] ;
 wire \generated._487[2] ;
 wire \generated._487[3] ;
 wire \generated._501[0] ;
 wire \generated._503 ;
 wire \generated._505[0] ;
 wire \generated._505[1] ;
 wire \generated._505[2] ;
 wire \generated._505[3] ;
 wire \generated._505[4] ;
 wire \generated._505[5] ;
 wire \generated._505[6] ;
 wire \generated._505[7] ;
 wire \generated._505[8] ;
 wire \generated._509 ;
 wire \generated._510 ;
 wire \generated._511 ;
 wire \generated._512[0] ;
 wire \generated._512[1] ;
 wire \generated._512[2] ;
 wire \generated._512[3] ;
 wire \generated._512[4] ;
 wire \generated._512[5] ;
 wire \generated._512[6] ;
 wire \generated._512[7] ;
 wire \generated._561[0] ;
 wire \generated._561[1] ;
 wire \generated._561[2] ;
 wire \generated._561[3] ;
 wire \generated._561[4] ;
 wire \generated._561[5] ;
 wire \generated._561[6] ;
 wire \generated._561[7] ;
 wire \generated._561[8] ;
 wire \generated._561[9] ;
 wire \generated._562[0] ;
 wire \generated._562[1] ;
 wire \generated._562[2] ;
 wire \generated._562[3] ;
 wire \generated._562[4] ;
 wire \generated._562[5] ;
 wire \generated._562[6] ;
 wire \generated._562[7] ;
 wire \generated._562[8] ;
 wire \generated._562[9] ;
 wire \generated._563[0] ;
 wire \generated._614[0] ;
 wire \generated._614[1] ;
 wire \generated._614[2] ;
 wire \generated._614[3] ;
 wire \generated._614[4] ;
 wire \generated._614[5] ;
 wire \generated._63[0] ;
 wire \generated._63[1] ;
 wire \generated._63[2] ;
 wire \generated._63[3] ;
 wire \generated._64[0] ;
 wire \generated._65[2] ;
 wire \generated._65[3] ;
 wire \generated._65[4] ;
 wire \generated._65[5] ;
 wire \generated._65[6] ;
 wire \generated._66[1] ;
 wire \generated._66[2] ;
 wire \generated._66[3] ;
 wire \generated._66[4] ;
 wire \generated._66[5] ;
 wire \generated._66[6] ;
 wire \generated._66[7] ;
 wire \generated._66[8] ;
 wire \generated._66[9] ;
 wire \generated._695[0] ;
 wire \generated._695[1] ;
 wire \generated._695[2] ;
 wire \generated._695[3] ;
 wire \generated._695[4] ;
 wire \generated._695[5] ;
 wire \generated._695[6] ;
 wire \generated._695[7] ;
 wire \generated._695[8] ;
 wire \generated._695[9] ;
 wire \generated._698[0] ;
 wire \generated._69[0] ;
 wire \generated._69[1] ;
 wire \generated._69[2] ;
 wire \generated._69[3] ;
 wire \generated._69[4] ;
 wire \generated._69[5] ;
 wire \generated._69[6] ;
 wire \generated._69[7] ;
 wire \generated._69[8] ;
 wire \generated._69[9] ;
 wire \generated._71[0] ;
 wire \generated._71[1] ;
 wire \generated._71[2] ;
 wire \generated._71[3] ;
 wire \generated._77[0] ;
 wire \generated._843 ;
 wire \generated._844 ;
 wire \generated._889[3] ;
 wire \generated._889[4] ;
 wire \generated._889[5] ;
 wire \generated._889[6] ;
 wire \generated._889[7] ;
 wire \generated._889[8] ;
 wire \generated._889[9] ;
 wire \generated._891[0] ;
 wire \generated._938[3] ;
 wire \generated._938[4] ;
 wire \generated._938[5] ;
 wire \generated._938[6] ;
 wire \generated._938[7] ;
 wire \generated._938[8] ;
 wire \generated._938[9] ;
 wire \generated._941[0] ;
 wire \generated._969 ;
 wire \generated._970 ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_leaf_0_clk;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net1;
 wire net2;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net750;
 wire net751;
 wire net752;
 wire net753;

 sg13g2_inv_1 _3587_ (.Y(_2830_),
    .A(net348));
 sg13g2_inv_1 _3588_ (.Y(_2831_),
    .A(net318));
 sg13g2_inv_1 _3589_ (.Y(_2832_),
    .A(net329));
 sg13g2_inv_1 _3590_ (.Y(_2833_),
    .A(net418));
 sg13g2_inv_1 _3591_ (.Y(_2834_),
    .A(net265));
 sg13g2_inv_2 _3592_ (.Y(_2835_),
    .A(\generated._221[3] ));
 sg13g2_inv_4 _3593_ (.A(net727),
    .Y(_2836_));
 sg13g2_inv_1 _3594_ (.Y(_2837_),
    .A(net729));
 sg13g2_inv_1 _3595_ (.Y(_2838_),
    .A(net379));
 sg13g2_inv_1 _3596_ (.Y(_2839_),
    .A(_0089_));
 sg13g2_inv_2 _3597_ (.Y(_2840_),
    .A(net667));
 sg13g2_inv_1 _3598_ (.Y(_2841_),
    .A(_0093_));
 sg13g2_inv_1 _3599_ (.Y(_2842_),
    .A(_0094_));
 sg13g2_inv_1 _3600_ (.Y(_2843_),
    .A(net420));
 sg13g2_inv_1 _3601_ (.Y(_2844_),
    .A(net748));
 sg13g2_inv_1 _3602_ (.Y(_2845_),
    .A(net720));
 sg13g2_inv_1 _3603_ (.Y(_2846_),
    .A(\generated._21[0] ));
 sg13g2_inv_1 _3604_ (.Y(_2847_),
    .A(net299));
 sg13g2_inv_1 _3605_ (.Y(_2848_),
    .A(_0019_));
 sg13g2_inv_1 _3606_ (.Y(_2849_),
    .A(_0038_));
 sg13g2_inv_1 _3607_ (.Y(_2850_),
    .A(_0039_));
 sg13g2_inv_1 _3608_ (.Y(_2851_),
    .A(_0041_));
 sg13g2_inv_1 _3609_ (.Y(_2852_),
    .A(_0042_));
 sg13g2_inv_1 _3610_ (.Y(_2853_),
    .A(_0043_));
 sg13g2_inv_1 _3611_ (.Y(_2854_),
    .A(net684));
 sg13g2_inv_1 _3612_ (.Y(_2855_),
    .A(net480));
 sg13g2_inv_1 _3613_ (.Y(_2856_),
    .A(_0050_));
 sg13g2_inv_1 _3614_ (.Y(_2857_),
    .A(_0054_));
 sg13g2_inv_1 _3615_ (.Y(_2858_),
    .A(\generated._394[7] ));
 sg13g2_inv_1 _3616_ (.Y(_2859_),
    .A(\generated._512[4] ));
 sg13g2_inv_1 _3617_ (.Y(_2860_),
    .A(_0063_));
 sg13g2_inv_2 _3618_ (.Y(_2861_),
    .A(_0064_));
 sg13g2_inv_1 _3619_ (.Y(_2862_),
    .A(_0073_));
 sg13g2_inv_1 _3620_ (.Y(_2863_),
    .A(net415));
 sg13g2_inv_2 _3621_ (.Y(_2864_),
    .A(net671));
 sg13g2_inv_1 _3622_ (.Y(_2865_),
    .A(\generated._373[7] ));
 sg13g2_inv_1 _3623_ (.Y(_2866_),
    .A(\generated._1084[3] ));
 sg13g2_inv_1 _3624_ (.Y(_2867_),
    .A(\generated._1084[4] ));
 sg13g2_inv_1 _3625_ (.Y(_2868_),
    .A(\generated._65[2] ));
 sg13g2_inv_1 _3626_ (.Y(_2869_),
    .A(net744));
 sg13g2_inv_1 _3627_ (.Y(_2870_),
    .A(\generated._381[4] ));
 sg13g2_inv_1 _3628_ (.Y(_2871_),
    .A(_0085_));
 sg13g2_inv_1 _3629_ (.Y(_2872_),
    .A(_0088_));
 sg13g2_nand2_1 _3630_ (.Y(_2873_),
    .A(\generated._21[3] ),
    .B(\generated._21[4] ));
 sg13g2_nor4_2 _3631_ (.A(\generated._21[1] ),
    .B(_2846_),
    .C(\generated._21[2] ),
    .Y(_2874_),
    .D(_2873_));
 sg13g2_or4_1 _3632_ (.A(_2830_),
    .B(\generated._16[2] ),
    .C(\generated._16[1] ),
    .D(_0095_),
    .X(_2875_));
 sg13g2_o21ai_1 _3633_ (.B1(_2874_),
    .Y(_2876_),
    .A1(\generated._16[0] ),
    .A2(_2875_));
 sg13g2_nor2b_1 _3634_ (.A(net359),
    .B_N(_2876_),
    .Y(_2877_));
 sg13g2_nor2_1 _3635_ (.A(\generated._100[3] ),
    .B(net724),
    .Y(_2878_));
 sg13g2_or3_1 _3636_ (.A(\generated._100[3] ),
    .B(net723),
    .C(\generated._100[5] ),
    .X(_2879_));
 sg13g2_nor3_2 _3637_ (.A(net723),
    .B(\generated._100[5] ),
    .C(\generated._100[6] ),
    .Y(_2880_));
 sg13g2_nor4_1 _3638_ (.A(\generated._100[3] ),
    .B(net722),
    .C(net721),
    .D(net720),
    .Y(_2881_));
 sg13g2_nand2_1 _3639_ (.Y(_2882_),
    .A(_2880_),
    .B(_2881_));
 sg13g2_nor4_1 _3640_ (.A(\generated._100[1] ),
    .B(\generated._100[0] ),
    .C(\generated._100[2] ),
    .D(_2882_),
    .Y(_2883_));
 sg13g2_or4_2 _3641_ (.A(\generated._100[1] ),
    .B(\generated._100[0] ),
    .C(\generated._100[2] ),
    .D(_2882_),
    .X(_2884_));
 sg13g2_and2_1 _3642_ (.A(net359),
    .B(_2874_),
    .X(_2885_));
 sg13g2_nor3_1 _3643_ (.A(_2877_),
    .B(net623),
    .C(_2885_),
    .Y(_0227_));
 sg13g2_nor2_2 _3644_ (.A(_2874_),
    .B(net623),
    .Y(_2886_));
 sg13g2_nand2b_2 _3645_ (.Y(_2887_),
    .B(_2884_),
    .A_N(_2874_));
 sg13g2_nand2_1 _3646_ (.Y(_2888_),
    .A(net276),
    .B(_2886_));
 sg13g2_nand2b_1 _3647_ (.Y(_2889_),
    .B(_2884_),
    .A_N(_2876_));
 sg13g2_nand3_1 _3648_ (.B(net337),
    .C(net394),
    .A(net278),
    .Y(_2890_));
 sg13g2_or2_1 _3649_ (.X(_2891_),
    .B(_2890_),
    .A(_2830_));
 sg13g2_xnor2_1 _3650_ (.Y(_2892_),
    .A(_0095_),
    .B(_2891_));
 sg13g2_o21ai_1 _3651_ (.B1(_2888_),
    .Y(_0231_),
    .A1(_2889_),
    .A2(_2892_));
 sg13g2_xnor2_1 _3652_ (.Y(_2893_),
    .A(net348),
    .B(_2890_));
 sg13g2_a21oi_1 _3653_ (.A1(net277),
    .A2(_2893_),
    .Y(_0003_),
    .B1(_0227_));
 sg13g2_and2_1 _3654_ (.A(\generated._357[1] ),
    .B(net271),
    .X(_2894_));
 sg13g2_nor2_1 _3655_ (.A(\generated._357[3] ),
    .B(\generated._357[2] ),
    .Y(_2895_));
 sg13g2_nand3_1 _3656_ (.B(_2894_),
    .C(_2895_),
    .A(\generated._357[4] ),
    .Y(_2896_));
 sg13g2_inv_1 _3657_ (.Y(_2897_),
    .A(_2896_));
 sg13g2_or2_1 _3658_ (.X(_2898_),
    .B(\generated._346[0] ),
    .A(\generated._346[1] ));
 sg13g2_nand2b_1 _3659_ (.Y(_2899_),
    .B(\generated._346[5] ),
    .A_N(\generated._346[4] ));
 sg13g2_nor4_1 _3660_ (.A(\generated._346[3] ),
    .B(\generated._346[2] ),
    .C(_2898_),
    .D(_2899_),
    .Y(_2900_));
 sg13g2_nor2_1 _3661_ (.A(_2896_),
    .B(_2900_),
    .Y(_2901_));
 sg13g2_nand2_2 _3662_ (.Y(_2902_),
    .A(net313),
    .B(\generated._346[0] ));
 sg13g2_nor2_1 _3663_ (.A(_0097_),
    .B(_2902_),
    .Y(_2903_));
 sg13g2_xnor2_1 _3664_ (.Y(_2904_),
    .A(net532),
    .B(_2903_));
 sg13g2_a22oi_1 _3665_ (.Y(_2905_),
    .B1(_2901_),
    .B2(_2904_),
    .A2(_2896_),
    .A1(net316));
 sg13g2_a21oi_1 _3666_ (.A1(net472),
    .A2(_2897_),
    .Y(_2906_),
    .B1(net624));
 sg13g2_nor2_2 _3667_ (.A(net625),
    .B(_2897_),
    .Y(_2907_));
 sg13g2_nand2_1 _3668_ (.Y(_2908_),
    .A(_2884_),
    .B(_2896_));
 sg13g2_or2_1 _3669_ (.X(_2909_),
    .B(_2900_),
    .A(net624));
 sg13g2_o21ai_1 _3670_ (.B1(_2906_),
    .Y(_2910_),
    .A1(\generated._346[0] ),
    .A2(_2901_));
 sg13g2_inv_1 _3671_ (.Y(_0245_),
    .A(_2910_));
 sg13g2_nor2_1 _3672_ (.A(net317),
    .B(_2910_),
    .Y(_0004_));
 sg13g2_and4_1 _3673_ (.A(_2884_),
    .B(_2897_),
    .C(_2898_),
    .D(_2902_),
    .X(_2911_));
 sg13g2_a21oi_2 _3674_ (.B1(_2911_),
    .Y(_2912_),
    .A2(_2907_),
    .A1(_2847_));
 sg13g2_nor2_1 _3675_ (.A(net317),
    .B(_2912_),
    .Y(_0005_));
 sg13g2_xor2_1 _3676_ (.B(_2902_),
    .A(_0097_),
    .X(_2913_));
 sg13g2_a22oi_1 _3677_ (.Y(_2914_),
    .B1(_2901_),
    .B2(_2913_),
    .A2(_2896_),
    .A1(net384));
 sg13g2_nor2_1 _3678_ (.A(net624),
    .B(net317),
    .Y(_0248_));
 sg13g2_nor2_1 _3679_ (.A(net624),
    .B(net385),
    .Y(_0247_));
 sg13g2_nor3_1 _3680_ (.A(net624),
    .B(net317),
    .C(net385),
    .Y(_0006_));
 sg13g2_nand2_1 _3681_ (.Y(_2915_),
    .A(net316),
    .B(\generated._346[2] ));
 sg13g2_nor3_1 _3682_ (.A(_2896_),
    .B(_2902_),
    .C(_2915_),
    .Y(_2916_));
 sg13g2_and2_1 _3683_ (.A(net341),
    .B(_2916_),
    .X(_2917_));
 sg13g2_o21ai_1 _3684_ (.B1(_2884_),
    .Y(_2918_),
    .A1(net341),
    .A2(_2916_));
 sg13g2_nor2_2 _3685_ (.A(_2917_),
    .B(_2918_),
    .Y(_0249_));
 sg13g2_xnor2_1 _3686_ (.Y(_2919_),
    .A(_2905_),
    .B(_0249_));
 sg13g2_nor2_1 _3687_ (.A(_2910_),
    .B(_2919_),
    .Y(_0000_));
 sg13g2_nor2_1 _3688_ (.A(_2912_),
    .B(_2919_),
    .Y(_0001_));
 sg13g2_nor2b_1 _3689_ (.A(_2919_),
    .B_N(_0247_),
    .Y(_0002_));
 sg13g2_nand2_1 _3690_ (.Y(_2920_),
    .A(net738),
    .B(net737));
 sg13g2_nor2_1 _3691_ (.A(net736),
    .B(_2920_),
    .Y(_2921_));
 sg13g2_nand2_1 _3692_ (.Y(_2922_),
    .A(net736),
    .B(net737));
 sg13g2_xnor2_1 _3693_ (.Y(_2923_),
    .A(net736),
    .B(net737));
 sg13g2_a21oi_1 _3694_ (.A1(_2920_),
    .A2(_2923_),
    .Y(_2924_),
    .B1(_2921_));
 sg13g2_nand2_1 _3695_ (.Y(_2925_),
    .A(net688),
    .B(\generated._66[7] ));
 sg13g2_xor2_1 _3696_ (.B(net734),
    .A(net688),
    .X(_2926_));
 sg13g2_a21oi_1 _3697_ (.A1(_2924_),
    .A2(_2926_),
    .Y(_2927_),
    .B1(_2921_));
 sg13g2_nor2_1 _3698_ (.A(net734),
    .B(_2922_),
    .Y(_2928_));
 sg13g2_nand2_1 _3699_ (.Y(_2929_),
    .A(net734),
    .B(net735));
 sg13g2_xnor2_1 _3700_ (.Y(_2930_),
    .A(net734),
    .B(net736));
 sg13g2_a21oi_1 _3701_ (.A1(_2922_),
    .A2(_2930_),
    .Y(_2931_),
    .B1(_2928_));
 sg13g2_nand2_1 _3702_ (.Y(_2932_),
    .A(net740),
    .B(\generated._66[8] ));
 sg13g2_xor2_1 _3703_ (.B(net733),
    .A(net740),
    .X(_2933_));
 sg13g2_xnor2_1 _3704_ (.Y(_2934_),
    .A(_2931_),
    .B(_2933_));
 sg13g2_nor2_1 _3705_ (.A(_2927_),
    .B(_2934_),
    .Y(_2935_));
 sg13g2_xor2_1 _3706_ (.B(_2934_),
    .A(_2927_),
    .X(_2936_));
 sg13g2_nor2b_1 _3707_ (.A(_2925_),
    .B_N(_2936_),
    .Y(_2937_));
 sg13g2_a21oi_1 _3708_ (.A1(_2931_),
    .A2(_2933_),
    .Y(_2938_),
    .B1(_2928_));
 sg13g2_xor2_1 _3709_ (.B(net732),
    .A(net738),
    .X(_2939_));
 sg13g2_nand2_1 _3710_ (.Y(_2940_),
    .A(net733),
    .B(net735));
 sg13g2_nand2_1 _3711_ (.Y(_2941_),
    .A(net733),
    .B(net734));
 sg13g2_nor2_1 _3712_ (.A(net733),
    .B(net734),
    .Y(_2942_));
 sg13g2_nand2b_1 _3713_ (.Y(_2943_),
    .B(_2941_),
    .A_N(net735));
 sg13g2_o21ai_1 _3714_ (.B1(_2940_),
    .Y(_2944_),
    .A1(_2942_),
    .A2(_2943_));
 sg13g2_xor2_1 _3715_ (.B(_2944_),
    .A(_2939_),
    .X(_2945_));
 sg13g2_nand2b_1 _3716_ (.Y(_2946_),
    .B(_2945_),
    .A_N(_2938_));
 sg13g2_xnor2_1 _3717_ (.Y(_2947_),
    .A(_2938_),
    .B(_2945_));
 sg13g2_nand2b_1 _3718_ (.Y(_2948_),
    .B(_2947_),
    .A_N(_2932_));
 sg13g2_xnor2_1 _3719_ (.Y(_2949_),
    .A(_2932_),
    .B(_2947_));
 sg13g2_o21ai_1 _3720_ (.B1(_2949_),
    .Y(_2950_),
    .A1(_2935_),
    .A2(_2937_));
 sg13g2_or3_1 _3721_ (.A(_2935_),
    .B(_2937_),
    .C(_2949_),
    .X(_2951_));
 sg13g2_and2_1 _3722_ (.A(_2950_),
    .B(_2951_),
    .X(_2952_));
 sg13g2_nand2_1 _3723_ (.Y(_2953_),
    .A(net740),
    .B(net739));
 sg13g2_nor2_1 _3724_ (.A(\generated._66[5] ),
    .B(_2953_),
    .Y(_2954_));
 sg13g2_nand2_1 _3725_ (.Y(_2955_),
    .A(\generated._66[1] ),
    .B(net735));
 sg13g2_xor2_1 _3726_ (.B(net735),
    .A(net689),
    .X(_2956_));
 sg13g2_xnor2_1 _3727_ (.Y(_2957_),
    .A(net739),
    .B(net737));
 sg13g2_a21oi_2 _3728_ (.B1(_2954_),
    .Y(_2958_),
    .A2(_2957_),
    .A1(_2953_));
 sg13g2_a21oi_1 _3729_ (.A1(_2956_),
    .A2(_2958_),
    .Y(_2959_),
    .B1(_2954_));
 sg13g2_xnor2_1 _3730_ (.Y(_2960_),
    .A(_2924_),
    .B(_2926_));
 sg13g2_xor2_1 _3731_ (.B(_2960_),
    .A(_2959_),
    .X(_2961_));
 sg13g2_nand2b_1 _3732_ (.Y(_2962_),
    .B(_2961_),
    .A_N(_2955_));
 sg13g2_o21ai_1 _3733_ (.B1(_2962_),
    .Y(_2963_),
    .A1(_2959_),
    .A2(_2960_));
 sg13g2_xnor2_1 _3734_ (.Y(_2964_),
    .A(_2925_),
    .B(_2936_));
 sg13g2_nand2_1 _3735_ (.Y(_2965_),
    .A(\generated._425[1] ),
    .B(net737));
 sg13g2_nand2_1 _3736_ (.Y(_2966_),
    .A(net688),
    .B(\generated._66[3] ));
 sg13g2_nor2_1 _3737_ (.A(net739),
    .B(_2966_),
    .Y(_2967_));
 sg13g2_xnor2_1 _3738_ (.Y(_2968_),
    .A(\generated._425[1] ),
    .B(net737));
 sg13g2_nand2b_1 _3739_ (.Y(_2969_),
    .B(\generated._66[3] ),
    .A_N(net688));
 sg13g2_xor2_1 _3740_ (.B(_2969_),
    .A(net738),
    .X(_2970_));
 sg13g2_nor2_1 _3741_ (.A(_2968_),
    .B(_2970_),
    .Y(_2971_));
 sg13g2_nor2_1 _3742_ (.A(_2967_),
    .B(_2971_),
    .Y(_2972_));
 sg13g2_xnor2_1 _3743_ (.Y(_2973_),
    .A(_2956_),
    .B(_2958_));
 sg13g2_nor2_1 _3744_ (.A(_2972_),
    .B(_2973_),
    .Y(_2974_));
 sg13g2_xnor2_1 _3745_ (.Y(_2975_),
    .A(_2972_),
    .B(_2973_));
 sg13g2_or2_1 _3746_ (.X(_2976_),
    .B(_2975_),
    .A(_2965_));
 sg13g2_nand2_1 _3747_ (.Y(_2977_),
    .A(net689),
    .B(net688));
 sg13g2_nor2_1 _3748_ (.A(net740),
    .B(_2977_),
    .Y(_2978_));
 sg13g2_xor2_1 _3749_ (.B(net740),
    .A(net688),
    .X(_2979_));
 sg13g2_a21oi_1 _3750_ (.A1(net689),
    .A2(net688),
    .Y(_2980_),
    .B1(_2979_));
 sg13g2_nor2_1 _3751_ (.A(_2978_),
    .B(_2980_),
    .Y(_2981_));
 sg13g2_a21oi_1 _3752_ (.A1(net738),
    .A2(_2981_),
    .Y(_2982_),
    .B1(_2978_));
 sg13g2_xnor2_1 _3753_ (.Y(_2983_),
    .A(_2968_),
    .B(_2970_));
 sg13g2_nand2_1 _3754_ (.Y(_2984_),
    .A(_2982_),
    .B(_2983_));
 sg13g2_nor2b_1 _3755_ (.A(\generated._425[1] ),
    .B_N(net689),
    .Y(_2985_));
 sg13g2_nand2b_1 _3756_ (.Y(_2986_),
    .B(net689),
    .A_N(net688));
 sg13g2_a22oi_1 _3757_ (.Y(_2987_),
    .B1(_2986_),
    .B2(_2966_),
    .A2(_2985_),
    .A1(_2969_));
 sg13g2_xor2_1 _3758_ (.B(_2981_),
    .A(net738),
    .X(_2988_));
 sg13g2_nand2_1 _3759_ (.Y(_2989_),
    .A(_2987_),
    .B(_2988_));
 sg13g2_o21ai_1 _3760_ (.B1(_2989_),
    .Y(_2990_),
    .A1(_2982_),
    .A2(_2983_));
 sg13g2_nand3_1 _3761_ (.B(_2984_),
    .C(_2990_),
    .A(_2976_),
    .Y(_2991_));
 sg13g2_a21oi_1 _3762_ (.A1(_2965_),
    .A2(_2975_),
    .Y(_2992_),
    .B1(_2991_));
 sg13g2_nand2_1 _3763_ (.Y(_2993_),
    .A(\generated._425[1] ),
    .B(net689));
 sg13g2_or2_1 _3764_ (.X(_2994_),
    .B(_2988_),
    .A(_2987_));
 sg13g2_mux2_1 _3765_ (.A0(\generated._425[1] ),
    .A1(_2985_),
    .S(net740),
    .X(_2995_));
 sg13g2_nand4_1 _3766_ (.B(_2984_),
    .C(_2994_),
    .A(\generated._66[2] ),
    .Y(_2996_),
    .D(_2995_));
 sg13g2_o21ai_1 _3767_ (.B1(_2993_),
    .Y(_2997_),
    .A1(_2990_),
    .A2(_2996_));
 sg13g2_nand4_1 _3768_ (.B(net738),
    .C(_2958_),
    .A(_2839_),
    .Y(_2998_),
    .D(_2979_));
 sg13g2_nand2b_1 _3769_ (.Y(_2999_),
    .B(_2998_),
    .A_N(_2993_));
 sg13g2_nand3_1 _3770_ (.B(_2997_),
    .C(_2999_),
    .A(_2956_),
    .Y(_3000_));
 sg13g2_nor2b_1 _3771_ (.A(_2974_),
    .B_N(_2976_),
    .Y(_3001_));
 sg13g2_xor2_1 _3772_ (.B(_2961_),
    .A(_2955_),
    .X(_3002_));
 sg13g2_nand2_1 _3773_ (.Y(_3003_),
    .A(_3001_),
    .B(_3002_));
 sg13g2_nand2_1 _3774_ (.Y(_3004_),
    .A(_2963_),
    .B(_2964_));
 sg13g2_o21ai_1 _3775_ (.B1(_3000_),
    .Y(_3005_),
    .A1(_3001_),
    .A2(_3002_));
 sg13g2_nor2_1 _3776_ (.A(_2992_),
    .B(_3005_),
    .Y(_3006_));
 sg13g2_o21ai_1 _3777_ (.B1(_3003_),
    .Y(_3007_),
    .A1(_2963_),
    .A2(_2964_));
 sg13g2_o21ai_1 _3778_ (.B1(_3004_),
    .Y(_3008_),
    .A1(_3006_),
    .A2(_3007_));
 sg13g2_nand2_1 _3779_ (.Y(_3009_),
    .A(_2952_),
    .B(_3008_));
 sg13g2_nor2_1 _3780_ (.A(_2952_),
    .B(_3008_),
    .Y(_3010_));
 sg13g2_nor3_2 _3781_ (.A(\generated._1078[0] ),
    .B(\generated._1078[1] ),
    .C(\generated._1078[3] ),
    .Y(_3011_));
 sg13g2_nor2b_1 _3782_ (.A(net456),
    .B_N(_3011_),
    .Y(_3012_));
 sg13g2_nand2b_1 _3783_ (.Y(_3013_),
    .B(_3011_),
    .A_N(\generated._1078[2] ));
 sg13g2_nand2_1 _3784_ (.Y(_3014_),
    .A(_3009_),
    .B(net654));
 sg13g2_nor4_1 _3785_ (.A(\generated._1074[5] ),
    .B(\generated._1074[4] ),
    .C(\generated._1074[2] ),
    .D(\generated._1074[1] ),
    .Y(_3015_));
 sg13g2_or4_1 _3786_ (.A(\generated._1074[9] ),
    .B(\generated._1074[8] ),
    .C(\generated._1074[7] ),
    .D(\generated._1074[6] ),
    .X(_3016_));
 sg13g2_nor3_1 _3787_ (.A(\generated._1074[0] ),
    .B(\generated._1074[3] ),
    .C(_3016_),
    .Y(_3017_));
 sg13g2_a21oi_1 _3788_ (.A1(_3015_),
    .A2(_3017_),
    .Y(_3018_),
    .B1(_0107_));
 sg13g2_mux2_1 _3789_ (.A0(_0092_),
    .A1(_0103_),
    .S(net707),
    .X(_3019_));
 sg13g2_nor2_2 _3790_ (.A(net707),
    .B(net701),
    .Y(_3020_));
 sg13g2_nand2_1 _3791_ (.Y(_3021_),
    .A(_0106_),
    .B(_3020_));
 sg13g2_nor2b_2 _3792_ (.A(net701),
    .B_N(net710),
    .Y(_3022_));
 sg13g2_a22oi_1 _3793_ (.Y(_3023_),
    .B1(_3022_),
    .B2(_0091_),
    .A2(_3019_),
    .A1(net701));
 sg13g2_nand2_1 _3794_ (.Y(_3024_),
    .A(_3021_),
    .B(_3023_));
 sg13g2_nor2b_1 _3795_ (.A(net710),
    .B_N(_0091_),
    .Y(_3025_));
 sg13g2_a21oi_1 _3796_ (.A1(net710),
    .A2(_0092_),
    .Y(_3026_),
    .B1(_3025_));
 sg13g2_and2_1 _3797_ (.A(\generated._1024[1] ),
    .B(_3022_),
    .X(_3027_));
 sg13g2_a221oi_1 _3798_ (.B2(net701),
    .C1(_3027_),
    .B1(_3026_),
    .A1(\generated._1024[0] ),
    .Y(_3028_),
    .A2(_3020_));
 sg13g2_nand2_1 _3799_ (.Y(_3029_),
    .A(_3024_),
    .B(_3028_));
 sg13g2_nand2_1 _3800_ (.Y(_3030_),
    .A(net618),
    .B(_3029_));
 sg13g2_mux2_1 _3801_ (.A0(_0103_),
    .A1(_0104_),
    .S(net707),
    .X(_3031_));
 sg13g2_nand2_1 _3802_ (.Y(_3032_),
    .A(net702),
    .B(_3031_));
 sg13g2_o21ai_1 _3803_ (.B1(_3032_),
    .Y(_3033_),
    .A1(net702),
    .A2(_3026_));
 sg13g2_xor2_1 _3804_ (.B(_3033_),
    .A(_3030_),
    .X(_3034_));
 sg13g2_nor2b_1 _3805_ (.A(_3034_),
    .B_N(\generated._1074[2] ),
    .Y(_3035_));
 sg13g2_nor2b_1 _3806_ (.A(_3028_),
    .B_N(net618),
    .Y(_3036_));
 sg13g2_xnor2_1 _3807_ (.Y(_3037_),
    .A(_3024_),
    .B(_3036_));
 sg13g2_nor2_1 _3808_ (.A(_0109_),
    .B(_3037_),
    .Y(_3038_));
 sg13g2_nor2_1 _3809_ (.A(\generated._1074[0] ),
    .B(_3028_),
    .Y(_3039_));
 sg13g2_xnor2_1 _3810_ (.Y(_3040_),
    .A(net475),
    .B(_3037_));
 sg13g2_nor2_1 _3811_ (.A(_3039_),
    .B(_3040_),
    .Y(_3041_));
 sg13g2_nor2_1 _3812_ (.A(_3038_),
    .B(_3041_),
    .Y(_3042_));
 sg13g2_xor2_1 _3813_ (.B(_3034_),
    .A(net461),
    .X(_3043_));
 sg13g2_nor2b_1 _3814_ (.A(_3042_),
    .B_N(_3043_),
    .Y(_3044_));
 sg13g2_nand3_1 _3815_ (.B(_3028_),
    .C(_3033_),
    .A(_3024_),
    .Y(_3045_));
 sg13g2_nand2_1 _3816_ (.Y(_3046_),
    .A(net619),
    .B(_3045_));
 sg13g2_nor2_1 _3817_ (.A(net701),
    .B(_3019_),
    .Y(_3047_));
 sg13g2_nor2b_1 _3818_ (.A(net708),
    .B_N(_0104_),
    .Y(_3048_));
 sg13g2_a21oi_2 _3819_ (.B1(_3048_),
    .Y(_3049_),
    .A2(_0105_),
    .A1(net708));
 sg13g2_a21oi_1 _3820_ (.A1(net705),
    .A2(_3049_),
    .Y(_3050_),
    .B1(_3047_));
 sg13g2_xnor2_1 _3821_ (.Y(_3051_),
    .A(_3046_),
    .B(_3050_));
 sg13g2_nand2b_1 _3822_ (.Y(_3052_),
    .B(_3051_),
    .A_N(_0102_));
 sg13g2_xnor2_1 _3823_ (.Y(_3053_),
    .A(_0102_),
    .B(_3051_));
 sg13g2_o21ai_1 _3824_ (.B1(_3053_),
    .Y(_3054_),
    .A1(_3035_),
    .A2(_3044_));
 sg13g2_or3_1 _3825_ (.A(_3035_),
    .B(_3044_),
    .C(_3053_),
    .X(_3055_));
 sg13g2_nand3_1 _3826_ (.B(_3054_),
    .C(_3055_),
    .A(net651),
    .Y(_3056_));
 sg13g2_o21ai_1 _3827_ (.B1(_3056_),
    .Y(\generated._1073[3] ),
    .A1(_3010_),
    .A2(_3014_));
 sg13g2_and2_1 _3828_ (.A(_2946_),
    .B(_2948_),
    .X(_3057_));
 sg13g2_nor2_1 _3829_ (.A(net733),
    .B(_2929_),
    .Y(_3058_));
 sg13g2_a21o_1 _3830_ (.A2(_2944_),
    .A1(_2939_),
    .B1(_3058_),
    .X(_3059_));
 sg13g2_nand2_1 _3831_ (.Y(_3060_),
    .A(net732),
    .B(net737));
 sg13g2_xor2_1 _3832_ (.B(net737),
    .A(net732),
    .X(_3061_));
 sg13g2_xnor2_1 _3833_ (.Y(_3062_),
    .A(net733),
    .B(net732));
 sg13g2_and2_1 _3834_ (.A(_2941_),
    .B(_3062_),
    .X(_3063_));
 sg13g2_nor2_1 _3835_ (.A(net731),
    .B(_2941_),
    .Y(_3064_));
 sg13g2_nor2_1 _3836_ (.A(_3063_),
    .B(_3064_),
    .Y(_3065_));
 sg13g2_xor2_1 _3837_ (.B(_3065_),
    .A(_3061_),
    .X(_3066_));
 sg13g2_xor2_1 _3838_ (.B(_3066_),
    .A(_3059_),
    .X(_3067_));
 sg13g2_and3_1 _3839_ (.X(_3068_),
    .A(net738),
    .B(net731),
    .C(_3067_));
 sg13g2_a21oi_1 _3840_ (.A1(net738),
    .A2(net731),
    .Y(_3069_),
    .B1(_3067_));
 sg13g2_or2_1 _3841_ (.X(_3070_),
    .B(_3069_),
    .A(_3068_));
 sg13g2_nor2_1 _3842_ (.A(_3057_),
    .B(_3070_),
    .Y(_3071_));
 sg13g2_xnor2_1 _3843_ (.Y(_3072_),
    .A(_3057_),
    .B(_3070_));
 sg13g2_nand3_1 _3844_ (.B(_3009_),
    .C(_3072_),
    .A(_2950_),
    .Y(_3073_));
 sg13g2_a21oi_1 _3845_ (.A1(_2950_),
    .A2(_3009_),
    .Y(_3074_),
    .B1(_3072_));
 sg13g2_nand3b_1 _3846_ (.B(net654),
    .C(_3073_),
    .Y(_3075_),
    .A_N(_3074_));
 sg13g2_nand2b_1 _3847_ (.Y(_3076_),
    .B(_3050_),
    .A_N(_3045_));
 sg13g2_nand2_1 _3848_ (.Y(_3077_),
    .A(net620),
    .B(_3076_));
 sg13g2_nor2_1 _3849_ (.A(net705),
    .B(_3031_),
    .Y(_3078_));
 sg13g2_nor2b_1 _3850_ (.A(net708),
    .B_N(_0105_),
    .Y(_3079_));
 sg13g2_a21oi_1 _3851_ (.A1(net708),
    .A2(_0111_),
    .Y(_3080_),
    .B1(_3079_));
 sg13g2_a21oi_1 _3852_ (.A1(net705),
    .A2(_3080_),
    .Y(_3081_),
    .B1(_3078_));
 sg13g2_xnor2_1 _3853_ (.Y(_3082_),
    .A(_3077_),
    .B(_3081_));
 sg13g2_xor2_1 _3854_ (.B(_3082_),
    .A(net432),
    .X(_3083_));
 sg13g2_a21oi_1 _3855_ (.A1(_3052_),
    .A2(_3054_),
    .Y(_3084_),
    .B1(_3083_));
 sg13g2_nand3_1 _3856_ (.B(_3054_),
    .C(_3083_),
    .A(_3052_),
    .Y(_3085_));
 sg13g2_nand2_1 _3857_ (.Y(_3086_),
    .A(net651),
    .B(_3085_));
 sg13g2_o21ai_1 _3858_ (.B1(_3075_),
    .Y(\generated._1073[4] ),
    .A1(_3084_),
    .A2(_3086_));
 sg13g2_nor2_1 _3859_ (.A(_3071_),
    .B(_3074_),
    .Y(_3087_));
 sg13g2_a21oi_1 _3860_ (.A1(_3059_),
    .A2(_3066_),
    .Y(_3088_),
    .B1(_3068_));
 sg13g2_a21oi_1 _3861_ (.A1(_3061_),
    .A2(_3065_),
    .Y(_3089_),
    .B1(_3064_));
 sg13g2_o21ai_1 _3862_ (.B1(net731),
    .Y(_3090_),
    .A1(net733),
    .A2(net735));
 sg13g2_nand2b_1 _3863_ (.Y(_3091_),
    .B(_2940_),
    .A_N(_3090_));
 sg13g2_o21ai_1 _3864_ (.B1(_3091_),
    .Y(_3092_),
    .A1(net735),
    .A2(net731));
 sg13g2_nor2_1 _3865_ (.A(_3089_),
    .B(_3092_),
    .Y(_3093_));
 sg13g2_xor2_1 _3866_ (.B(_3092_),
    .A(_3089_),
    .X(_3094_));
 sg13g2_nor2b_1 _3867_ (.A(_3060_),
    .B_N(_3094_),
    .Y(_3095_));
 sg13g2_xnor2_1 _3868_ (.Y(_3096_),
    .A(_3060_),
    .B(_3094_));
 sg13g2_nor2b_1 _3869_ (.A(_3088_),
    .B_N(_3096_),
    .Y(_3097_));
 sg13g2_xor2_1 _3870_ (.B(_3096_),
    .A(_3088_),
    .X(_3098_));
 sg13g2_nor2_1 _3871_ (.A(_3087_),
    .B(_3098_),
    .Y(_3099_));
 sg13g2_a21o_1 _3872_ (.A2(_3098_),
    .A1(_3087_),
    .B1(net650),
    .X(_3100_));
 sg13g2_a21oi_1 _3873_ (.A1(\generated._1074[4] ),
    .A2(_3082_),
    .Y(_3101_),
    .B1(_3084_));
 sg13g2_nor2b_1 _3874_ (.A(_3076_),
    .B_N(_3081_),
    .Y(_3102_));
 sg13g2_nand2b_1 _3875_ (.Y(_3103_),
    .B(net620),
    .A_N(_3102_));
 sg13g2_mux2_1 _3876_ (.A0(_0111_),
    .A1(_0113_),
    .S(net708),
    .X(_3104_));
 sg13g2_nand2_1 _3877_ (.Y(_3105_),
    .A(net704),
    .B(_3104_));
 sg13g2_o21ai_1 _3878_ (.B1(_3105_),
    .Y(_3106_),
    .A1(net705),
    .A2(_3049_));
 sg13g2_xnor2_1 _3879_ (.Y(_3107_),
    .A(_3103_),
    .B(_3106_));
 sg13g2_nand2b_1 _3880_ (.Y(_3108_),
    .B(_3107_),
    .A_N(_0112_));
 sg13g2_xnor2_1 _3881_ (.Y(_3109_),
    .A(_0112_),
    .B(_3107_));
 sg13g2_nand2b_1 _3882_ (.Y(_3110_),
    .B(_3101_),
    .A_N(_3109_));
 sg13g2_nand2b_1 _3883_ (.Y(_3111_),
    .B(_3109_),
    .A_N(_3101_));
 sg13g2_nand3_1 _3884_ (.B(_3110_),
    .C(_3111_),
    .A(net650),
    .Y(_3112_));
 sg13g2_o21ai_1 _3885_ (.B1(_3112_),
    .Y(\generated._1073[5] ),
    .A1(_3099_),
    .A2(_3100_));
 sg13g2_xnor2_1 _3886_ (.Y(_3113_),
    .A(net734),
    .B(_3090_));
 sg13g2_o21ai_1 _3887_ (.B1(_3113_),
    .Y(_3114_),
    .A1(_3093_),
    .A2(_3095_));
 sg13g2_or3_1 _3888_ (.A(_3093_),
    .B(_3095_),
    .C(_3113_),
    .X(_3115_));
 sg13g2_and2_1 _3889_ (.A(_3114_),
    .B(_3115_),
    .X(_3116_));
 sg13g2_or2_1 _3890_ (.X(_3117_),
    .B(_3116_),
    .A(_3097_));
 sg13g2_and2_1 _3891_ (.A(_3097_),
    .B(_3116_),
    .X(_3118_));
 sg13g2_inv_1 _3892_ (.Y(_3119_),
    .A(_3118_));
 sg13g2_nand2_1 _3893_ (.Y(_3120_),
    .A(_3099_),
    .B(_3116_));
 sg13g2_a21oi_1 _3894_ (.A1(_3099_),
    .A2(_3117_),
    .Y(_3121_),
    .B1(_3118_));
 sg13g2_a21oi_1 _3895_ (.A1(_3117_),
    .A2(_3119_),
    .Y(_3122_),
    .B1(_3099_));
 sg13g2_nand2_1 _3896_ (.Y(_3123_),
    .A(net654),
    .B(_3120_));
 sg13g2_and2_1 _3897_ (.A(_3108_),
    .B(_3111_),
    .X(_3124_));
 sg13g2_nand2_1 _3898_ (.Y(_3125_),
    .A(_3102_),
    .B(_3106_));
 sg13g2_nand2_1 _3899_ (.Y(_3126_),
    .A(net621),
    .B(_3125_));
 sg13g2_mux2_1 _3900_ (.A0(_0113_),
    .A1(_0115_),
    .S(net708),
    .X(_3127_));
 sg13g2_nand2_1 _3901_ (.Y(_3128_),
    .A(net706),
    .B(_3127_));
 sg13g2_o21ai_1 _3902_ (.B1(_3128_),
    .Y(_3129_),
    .A1(net704),
    .A2(_3080_));
 sg13g2_xnor2_1 _3903_ (.Y(_3130_),
    .A(_3126_),
    .B(_3129_));
 sg13g2_xor2_1 _3904_ (.B(_3130_),
    .A(_0114_),
    .X(_3131_));
 sg13g2_a21oi_1 _3905_ (.A1(_3124_),
    .A2(_3131_),
    .Y(_3132_),
    .B1(net654));
 sg13g2_o21ai_1 _3906_ (.B1(_3132_),
    .Y(_3133_),
    .A1(_3124_),
    .A2(_3131_));
 sg13g2_o21ai_1 _3907_ (.B1(_3133_),
    .Y(\generated._1073[6] ),
    .A1(_3122_),
    .A2(_3123_));
 sg13g2_nand2_1 _3908_ (.Y(_3134_),
    .A(\generated._1074[6] ),
    .B(_3130_));
 sg13g2_o21ai_1 _3909_ (.B1(_3134_),
    .Y(_3135_),
    .A1(_3124_),
    .A2(_3131_));
 sg13g2_nor2b_1 _3910_ (.A(net706),
    .B_N(_3104_),
    .Y(_3136_));
 sg13g2_a21oi_2 _3911_ (.B1(_3136_),
    .Y(_3137_),
    .A2(_0115_),
    .A1(net706));
 sg13g2_nand3_1 _3912_ (.B(_3106_),
    .C(_3129_),
    .A(_3102_),
    .Y(_3138_));
 sg13g2_nand2_1 _3913_ (.Y(_3139_),
    .A(net621),
    .B(_3138_));
 sg13g2_xor2_1 _3914_ (.B(_3139_),
    .A(_3137_),
    .X(_3140_));
 sg13g2_xnor2_1 _3915_ (.Y(_3141_),
    .A(_0016_),
    .B(_3140_));
 sg13g2_nand2_1 _3916_ (.Y(_3142_),
    .A(_3135_),
    .B(_3141_));
 sg13g2_o21ai_1 _3917_ (.B1(net650),
    .Y(_3143_),
    .A1(_3135_),
    .A2(_3141_));
 sg13g2_nand2b_1 _3918_ (.Y(_3144_),
    .B(_3142_),
    .A_N(_3143_));
 sg13g2_or2_1 _3919_ (.X(_3145_),
    .B(_3063_),
    .A(_3058_));
 sg13g2_xor2_1 _3920_ (.B(_3145_),
    .A(_3114_),
    .X(_3146_));
 sg13g2_xor2_1 _3921_ (.B(_3146_),
    .A(_3121_),
    .X(_3147_));
 sg13g2_o21ai_1 _3922_ (.B1(_3144_),
    .Y(\generated._1073[7] ),
    .A1(net650),
    .A2(_3147_));
 sg13g2_nand2_1 _3923_ (.Y(_3148_),
    .A(net530),
    .B(_3140_));
 sg13g2_nor2b_1 _3924_ (.A(net706),
    .B_N(_3127_),
    .Y(_3149_));
 sg13g2_a21oi_1 _3925_ (.A1(net706),
    .A2(_0115_),
    .Y(_3150_),
    .B1(_3149_));
 sg13g2_o21ai_1 _3926_ (.B1(net620),
    .Y(_3151_),
    .A1(_3137_),
    .A2(_3138_));
 sg13g2_xor2_1 _3927_ (.B(_3151_),
    .A(_3150_),
    .X(_3152_));
 sg13g2_xor2_1 _3928_ (.B(_3152_),
    .A(_0017_),
    .X(_3153_));
 sg13g2_a21oi_1 _3929_ (.A1(_3142_),
    .A2(_3148_),
    .Y(_3154_),
    .B1(_3153_));
 sg13g2_nand3_1 _3930_ (.B(_3148_),
    .C(_3153_),
    .A(_3142_),
    .Y(_3155_));
 sg13g2_nand2b_1 _3931_ (.Y(_3156_),
    .B(_3155_),
    .A_N(_3154_));
 sg13g2_nor2b_1 _3932_ (.A(_3120_),
    .B_N(_3146_),
    .Y(_3157_));
 sg13g2_nor2_1 _3933_ (.A(_2942_),
    .B(_3090_),
    .Y(_3158_));
 sg13g2_a21oi_1 _3934_ (.A1(_3114_),
    .A2(_3119_),
    .Y(_3159_),
    .B1(_3145_));
 sg13g2_nor4_1 _3935_ (.A(net650),
    .B(_3157_),
    .C(_3158_),
    .D(_3159_),
    .Y(_3160_));
 sg13g2_a21oi_1 _3936_ (.A1(net650),
    .A2(_3156_),
    .Y(\generated._1073[8] ),
    .B1(_3160_));
 sg13g2_nor2_1 _3937_ (.A(net731),
    .B(net649),
    .Y(_3161_));
 sg13g2_a21oi_1 _3938_ (.A1(\generated._1074[8] ),
    .A2(_3152_),
    .Y(_3162_),
    .B1(_3154_));
 sg13g2_nor2_1 _3939_ (.A(_0115_),
    .B(net620),
    .Y(_3163_));
 sg13g2_nor3_1 _3940_ (.A(_3137_),
    .B(_3138_),
    .C(_3150_),
    .Y(_3164_));
 sg13g2_xnor2_1 _3941_ (.Y(_3165_),
    .A(\generated._1024[9] ),
    .B(_3164_));
 sg13g2_a21oi_1 _3942_ (.A1(net620),
    .A2(_3165_),
    .Y(_3166_),
    .B1(_3163_));
 sg13g2_xor2_1 _3943_ (.B(_3166_),
    .A(_0107_),
    .X(_3167_));
 sg13g2_xnor2_1 _3944_ (.Y(_3168_),
    .A(_3162_),
    .B(_3167_));
 sg13g2_a21oi_1 _3945_ (.A1(net650),
    .A2(_3168_),
    .Y(\generated._1073[9] ),
    .B1(_3161_));
 sg13g2_or3_1 _3946_ (.A(\generated._406[3] ),
    .B(\generated._406[2] ),
    .C(net750),
    .X(_3169_));
 sg13g2_o21ai_1 _3947_ (.B1(\generated._406[3] ),
    .Y(_3170_),
    .A1(\generated._406[2] ),
    .A2(\generated._406[1] ));
 sg13g2_a21oi_2 _3948_ (.B1(net649),
    .Y(_3171_),
    .A2(_3170_),
    .A1(net751));
 sg13g2_nor2b_1 _3949_ (.A(net707),
    .B_N(_0108_),
    .Y(_3172_));
 sg13g2_a21oi_1 _3950_ (.A1(net707),
    .A2(_0102_),
    .Y(_3173_),
    .B1(_3172_));
 sg13g2_nand2_1 _3951_ (.Y(_3174_),
    .A(net701),
    .B(_3173_));
 sg13g2_a22oi_1 _3952_ (.Y(_3175_),
    .B1(_3022_),
    .B2(\generated._1074[1] ),
    .A2(_3020_),
    .A1(\generated._1074[0] ));
 sg13g2_nand2_1 _3953_ (.Y(_3176_),
    .A(_3174_),
    .B(_3175_));
 sg13g2_and2_1 _3954_ (.A(net357),
    .B(_3176_),
    .X(_3177_));
 sg13g2_mux2_1 _3955_ (.A0(_0102_),
    .A1(_0110_),
    .S(net709),
    .X(_3178_));
 sg13g2_nand2_1 _3956_ (.Y(_3179_),
    .A(_0108_),
    .B(_3022_));
 sg13g2_a22oi_1 _3957_ (.Y(_3180_),
    .B1(_3178_),
    .B2(net702),
    .A2(_3020_),
    .A1(_0109_));
 sg13g2_nand2_1 _3958_ (.Y(_3181_),
    .A(_3179_),
    .B(_3180_));
 sg13g2_nand2_1 _3959_ (.Y(_3182_),
    .A(net618),
    .B(_3176_));
 sg13g2_xor2_1 _3960_ (.B(_3182_),
    .A(_3181_),
    .X(_3183_));
 sg13g2_xnor2_1 _3961_ (.Y(_3184_),
    .A(net410),
    .B(_3183_));
 sg13g2_and2_1 _3962_ (.A(_3177_),
    .B(_3184_),
    .X(_3185_));
 sg13g2_a21o_1 _3963_ (.A2(_3183_),
    .A1(\generated._1024[1] ),
    .B1(_3185_),
    .X(_3186_));
 sg13g2_nand3_1 _3964_ (.B(_3175_),
    .C(_3181_),
    .A(_3174_),
    .Y(_3187_));
 sg13g2_nand2_1 _3965_ (.Y(_3188_),
    .A(net618),
    .B(_3187_));
 sg13g2_mux2_1 _3966_ (.A0(_0110_),
    .A1(_0112_),
    .S(net709),
    .X(_3189_));
 sg13g2_nand2_1 _3967_ (.Y(_3190_),
    .A(net702),
    .B(_3189_));
 sg13g2_o21ai_1 _3968_ (.B1(_3190_),
    .Y(_3191_),
    .A1(net701),
    .A2(_3173_));
 sg13g2_xor2_1 _3969_ (.B(_3191_),
    .A(_3188_),
    .X(_3192_));
 sg13g2_xor2_1 _3970_ (.B(_3192_),
    .A(net429),
    .X(_3193_));
 sg13g2_nand2_1 _3971_ (.Y(_3194_),
    .A(_3186_),
    .B(_3193_));
 sg13g2_nand2b_1 _3972_ (.Y(_3195_),
    .B(_3192_),
    .A_N(_0091_));
 sg13g2_nand2b_1 _3973_ (.Y(_3196_),
    .B(_3191_),
    .A_N(_3187_));
 sg13g2_nand2_1 _3974_ (.Y(_3197_),
    .A(net618),
    .B(_3196_));
 sg13g2_nor2_1 _3975_ (.A(net701),
    .B(_3178_),
    .Y(_3198_));
 sg13g2_nor2b_1 _3976_ (.A(net709),
    .B_N(_0112_),
    .Y(_3199_));
 sg13g2_a21oi_1 _3977_ (.A1(net708),
    .A2(_0114_),
    .Y(_3200_),
    .B1(_3199_));
 sg13g2_a21oi_1 _3978_ (.A1(net705),
    .A2(_3200_),
    .Y(_3201_),
    .B1(_3198_));
 sg13g2_xor2_1 _3979_ (.B(_3201_),
    .A(_3197_),
    .X(_3202_));
 sg13g2_xnor2_1 _3980_ (.Y(_3203_),
    .A(\generated._1024[3] ),
    .B(_3202_));
 sg13g2_and3_1 _3981_ (.X(_3204_),
    .A(_3194_),
    .B(_3195_),
    .C(_3203_));
 sg13g2_a21oi_1 _3982_ (.A1(_3194_),
    .A2(_3195_),
    .Y(_3205_),
    .B1(_3203_));
 sg13g2_or2_1 _3983_ (.X(_3206_),
    .B(_3205_),
    .A(_3204_));
 sg13g2_a21oi_1 _3984_ (.A1(net648),
    .A2(_3206_),
    .Y(\generated._1023[3] ),
    .B1(_3171_));
 sg13g2_nand2b_1 _3985_ (.Y(_3207_),
    .B(_3170_),
    .A_N(\generated._406[4] ));
 sg13g2_xnor2_1 _3986_ (.Y(_3208_),
    .A(net362),
    .B(_3170_));
 sg13g2_a21oi_1 _3987_ (.A1(\generated._1024[3] ),
    .A2(_3202_),
    .Y(_3209_),
    .B1(_3205_));
 sg13g2_nand2b_1 _3988_ (.Y(_3210_),
    .B(_3201_),
    .A_N(_3196_));
 sg13g2_nand2_1 _3989_ (.Y(_3211_),
    .A(net618),
    .B(_3210_));
 sg13g2_nor2_1 _3990_ (.A(net705),
    .B(_3189_),
    .Y(_3212_));
 sg13g2_nor2b_1 _3991_ (.A(net709),
    .B_N(_0114_),
    .Y(_3213_));
 sg13g2_a21oi_1 _3992_ (.A1(net709),
    .A2(_0016_),
    .Y(_3214_),
    .B1(_3213_));
 sg13g2_a21oi_1 _3993_ (.A1(net705),
    .A2(_3214_),
    .Y(_3215_),
    .B1(_3212_));
 sg13g2_xnor2_1 _3994_ (.Y(_3216_),
    .A(_3211_),
    .B(_3215_));
 sg13g2_xnor2_1 _3995_ (.Y(_3217_),
    .A(net539),
    .B(_3216_));
 sg13g2_nor2b_1 _3996_ (.A(_3209_),
    .B_N(_3217_),
    .Y(_3218_));
 sg13g2_xnor2_1 _3997_ (.Y(_3219_),
    .A(_3209_),
    .B(_3217_));
 sg13g2_nand2_1 _3998_ (.Y(_3220_),
    .A(net648),
    .B(_3219_));
 sg13g2_o21ai_1 _3999_ (.B1(_3220_),
    .Y(\generated._1023[4] ),
    .A1(net648),
    .A2(_3208_));
 sg13g2_and2_1 _4000_ (.A(\generated._406[5] ),
    .B(_3207_),
    .X(_3221_));
 sg13g2_xor2_1 _4001_ (.B(_3207_),
    .A(net310),
    .X(_3222_));
 sg13g2_nand2_1 _4002_ (.Y(_3223_),
    .A(net654),
    .B(_3222_));
 sg13g2_nor2_1 _4003_ (.A(net511),
    .B(_3216_),
    .Y(_3224_));
 sg13g2_nor2_1 _4004_ (.A(_3218_),
    .B(_3224_),
    .Y(_3225_));
 sg13g2_nor2b_1 _4005_ (.A(_3210_),
    .B_N(_3215_),
    .Y(_3226_));
 sg13g2_nand2b_1 _4006_ (.Y(_3227_),
    .B(net620),
    .A_N(_3226_));
 sg13g2_mux2_1 _4007_ (.A0(_0016_),
    .A1(_0017_),
    .S(net709),
    .X(_3228_));
 sg13g2_nand2_1 _4008_ (.Y(_3229_),
    .A(net704),
    .B(_3228_));
 sg13g2_o21ai_1 _4009_ (.B1(_3229_),
    .Y(_3230_),
    .A1(net705),
    .A2(_3200_));
 sg13g2_xnor2_1 _4010_ (.Y(_3231_),
    .A(_3227_),
    .B(_3230_));
 sg13g2_inv_1 _4011_ (.Y(_3232_),
    .A(_3231_));
 sg13g2_xor2_1 _4012_ (.B(_3231_),
    .A(\generated._1024[5] ),
    .X(_3233_));
 sg13g2_nor2_1 _4013_ (.A(_3225_),
    .B(_3233_),
    .Y(_3234_));
 sg13g2_a21o_1 _4014_ (.A2(_3233_),
    .A1(_3225_),
    .B1(net652),
    .X(_3235_));
 sg13g2_o21ai_1 _4015_ (.B1(_3223_),
    .Y(\generated._1023[5] ),
    .A1(net512),
    .A2(_3235_));
 sg13g2_xnor2_1 _4016_ (.Y(_3236_),
    .A(net329),
    .B(_3221_));
 sg13g2_a21oi_1 _4017_ (.A1(\generated._1024[5] ),
    .A2(_3232_),
    .Y(_3237_),
    .B1(_3234_));
 sg13g2_nand2_1 _4018_ (.Y(_3238_),
    .A(_3226_),
    .B(_3230_));
 sg13g2_nand2_1 _4019_ (.Y(_3239_),
    .A(net620),
    .B(_3238_));
 sg13g2_mux2_1 _4020_ (.A0(_0017_),
    .A1(_0107_),
    .S(net708),
    .X(_0281_));
 sg13g2_nand2_1 _4021_ (.Y(_0282_),
    .A(net704),
    .B(_0281_));
 sg13g2_o21ai_1 _4022_ (.B1(_0282_),
    .Y(_0283_),
    .A1(net704),
    .A2(_3214_));
 sg13g2_xnor2_1 _4023_ (.Y(_0284_),
    .A(_3239_),
    .B(_0283_));
 sg13g2_xnor2_1 _4024_ (.Y(_0285_),
    .A(net510),
    .B(_0284_));
 sg13g2_nor2b_1 _4025_ (.A(_3237_),
    .B_N(_0285_),
    .Y(_0286_));
 sg13g2_xnor2_1 _4026_ (.Y(_0287_),
    .A(_3237_),
    .B(_0285_));
 sg13g2_nand2_1 _4027_ (.Y(_0288_),
    .A(net648),
    .B(_0287_));
 sg13g2_o21ai_1 _4028_ (.B1(_0288_),
    .Y(\generated._1023[6] ),
    .A1(net649),
    .A2(_3236_));
 sg13g2_nand3_1 _4029_ (.B(\generated._406[6] ),
    .C(_3221_),
    .A(net318),
    .Y(_0289_));
 sg13g2_a21o_1 _4030_ (.A2(_3221_),
    .A1(net329),
    .B1(net318),
    .X(_0290_));
 sg13g2_nand2_2 _4031_ (.Y(_0291_),
    .A(_0289_),
    .B(_0290_));
 sg13g2_nor2_1 _4032_ (.A(_0105_),
    .B(_0284_),
    .Y(_0292_));
 sg13g2_nor2b_1 _4033_ (.A(net706),
    .B_N(_3228_),
    .Y(_0293_));
 sg13g2_a21oi_2 _4034_ (.B1(_0293_),
    .Y(_0294_),
    .A2(_0107_),
    .A1(net704));
 sg13g2_nand3_1 _4035_ (.B(_3230_),
    .C(_0283_),
    .A(_3226_),
    .Y(_0295_));
 sg13g2_nand2_1 _4036_ (.Y(_0296_),
    .A(net621),
    .B(_0295_));
 sg13g2_xor2_1 _4037_ (.B(_0296_),
    .A(_0294_),
    .X(_0297_));
 sg13g2_xnor2_1 _4038_ (.Y(_0298_),
    .A(net478),
    .B(_0297_));
 sg13g2_o21ai_1 _4039_ (.B1(_0298_),
    .Y(_0299_),
    .A1(_0286_),
    .A2(_0292_));
 sg13g2_or3_1 _4040_ (.A(_0286_),
    .B(_0292_),
    .C(_0298_),
    .X(_0300_));
 sg13g2_nand3_1 _4041_ (.B(net479),
    .C(_0300_),
    .A(net649),
    .Y(_0301_));
 sg13g2_o21ai_1 _4042_ (.B1(_0301_),
    .Y(\generated._1023[7] ),
    .A1(net649),
    .A2(_0291_));
 sg13g2_nor2_1 _4043_ (.A(net649),
    .B(_0289_),
    .Y(_0302_));
 sg13g2_o21ai_1 _4044_ (.B1(_0299_),
    .Y(_0303_),
    .A1(net516),
    .A2(_0297_));
 sg13g2_nor2b_1 _4045_ (.A(net704),
    .B_N(_0281_),
    .Y(_0304_));
 sg13g2_a21oi_1 _4046_ (.A1(net704),
    .A2(_0107_),
    .Y(_0305_),
    .B1(_0304_));
 sg13g2_o21ai_1 _4047_ (.B1(net621),
    .Y(_0306_),
    .A1(_0294_),
    .A2(_0295_));
 sg13g2_xor2_1 _4048_ (.B(_0306_),
    .A(_0305_),
    .X(_0307_));
 sg13g2_xor2_1 _4049_ (.B(_0307_),
    .A(\generated._1024[8] ),
    .X(_0308_));
 sg13g2_inv_1 _4050_ (.Y(_0309_),
    .A(_0308_));
 sg13g2_xnor2_1 _4051_ (.Y(_0310_),
    .A(_0303_),
    .B(_0309_));
 sg13g2_a21oi_1 _4052_ (.A1(net649),
    .A2(net517),
    .Y(\generated._1023[8] ),
    .B1(_0302_));
 sg13g2_nor2_1 _4053_ (.A(net542),
    .B(_0307_),
    .Y(_0311_));
 sg13g2_a21oi_1 _4054_ (.A1(_0303_),
    .A2(_0309_),
    .Y(_0312_),
    .B1(_0311_));
 sg13g2_nor3_1 _4055_ (.A(_0294_),
    .B(_0295_),
    .C(_0305_),
    .Y(_0313_));
 sg13g2_o21ai_1 _4056_ (.B1(net620),
    .Y(_0314_),
    .A1(\generated._1074[9] ),
    .A2(_0313_));
 sg13g2_a21oi_1 _4057_ (.A1(\generated._1074[9] ),
    .A2(_0313_),
    .Y(_0315_),
    .B1(_0314_));
 sg13g2_nor2_1 _4058_ (.A(_0107_),
    .B(_0315_),
    .Y(_0316_));
 sg13g2_xor2_1 _4059_ (.B(_0316_),
    .A(\generated._1024[9] ),
    .X(_0317_));
 sg13g2_xnor2_1 _4060_ (.Y(_0318_),
    .A(_0312_),
    .B(_0317_));
 sg13g2_a21o_1 _4061_ (.A2(_0318_),
    .A1(net649),
    .B1(_0302_),
    .X(\generated._1023[9] ));
 sg13g2_a21o_2 _4062_ (.A2(_2879_),
    .A1(\generated._100[6] ),
    .B1(net722),
    .X(_0319_));
 sg13g2_nand2_1 _4063_ (.Y(_0320_),
    .A(net721),
    .B(_0319_));
 sg13g2_a21oi_1 _4064_ (.A1(net721),
    .A2(_0319_),
    .Y(_0321_),
    .B1(net720));
 sg13g2_nand2_1 _4065_ (.Y(_0322_),
    .A(_2845_),
    .B(_0320_));
 sg13g2_and4_1 _4066_ (.A(\generated._221[1] ),
    .B(\generated._221[0] ),
    .C(net728),
    .D(net729),
    .X(_0323_));
 sg13g2_and2_1 _4067_ (.A(net730),
    .B(_0323_),
    .X(_0324_));
 sg13g2_nor2_1 _4068_ (.A(\generated._221[3] ),
    .B(\generated._221[2] ),
    .Y(_0325_));
 sg13g2_a21oi_2 _4069_ (.B1(\generated._221[2] ),
    .Y(_0326_),
    .A2(_0323_),
    .A1(net730));
 sg13g2_and2_2 _4070_ (.A(_2835_),
    .B(_0326_),
    .X(_0327_));
 sg13g2_and2_1 _4071_ (.A(net617),
    .B(_0327_),
    .X(_0328_));
 sg13g2_xnor2_1 _4072_ (.Y(_0329_),
    .A(\generated._100[3] ),
    .B(net724));
 sg13g2_nand2_1 _4073_ (.Y(_0330_),
    .A(net601),
    .B(_0329_));
 sg13g2_a221oi_1 _4074_ (.B2(_2835_),
    .C1(net720),
    .B1(_0326_),
    .A1(net721),
    .Y(_0331_),
    .A2(_0319_));
 sg13g2_nand2b_2 _4075_ (.Y(_0332_),
    .B(net617),
    .A_N(_0327_));
 sg13g2_nor3_2 _4076_ (.A(\generated._71[0] ),
    .B(\generated._71[1] ),
    .C(net400),
    .Y(_0333_));
 sg13g2_nor2b_1 _4077_ (.A(net452),
    .B_N(_0333_),
    .Y(_0334_));
 sg13g2_nand2b_2 _4078_ (.Y(_0335_),
    .B(_0333_),
    .A_N(\generated._71[2] ));
 sg13g2_xor2_1 _4079_ (.B(net730),
    .A(net729),
    .X(_0336_));
 sg13g2_a221oi_1 _4080_ (.B2(net603),
    .C1(net640),
    .B1(_0336_),
    .A1(net724),
    .Y(_0337_),
    .A2(net612));
 sg13g2_nor4_1 _4081_ (.A(\generated._69[5] ),
    .B(\generated._69[4] ),
    .C(\generated._69[2] ),
    .D(\generated._69[1] ),
    .Y(_0338_));
 sg13g2_nor2_1 _4082_ (.A(\generated._69[0] ),
    .B(\generated._69[3] ),
    .Y(_0339_));
 sg13g2_nor4_1 _4083_ (.A(\generated._69[9] ),
    .B(\generated._69[8] ),
    .C(\generated._69[7] ),
    .D(\generated._69[6] ),
    .Y(_0340_));
 sg13g2_nand3_1 _4084_ (.B(_0339_),
    .C(_0340_),
    .A(_0338_),
    .Y(_0341_));
 sg13g2_nor2b_1 _4085_ (.A(_0023_),
    .B_N(_0341_),
    .Y(_0342_));
 sg13g2_nand2b_1 _4086_ (.Y(_0343_),
    .B(_0341_),
    .A_N(_0023_));
 sg13g2_nor2_1 _4087_ (.A(net698),
    .B(_0090_),
    .Y(_0344_));
 sg13g2_a21oi_1 _4088_ (.A1(net698),
    .A2(_2848_),
    .Y(_0345_),
    .B1(_0344_));
 sg13g2_nor2b_2 _4089_ (.A(net693),
    .B_N(net696),
    .Y(_0346_));
 sg13g2_nand2_1 _4090_ (.Y(_0347_),
    .A(_0089_),
    .B(_0346_));
 sg13g2_nor2_2 _4091_ (.A(net696),
    .B(net694),
    .Y(_0348_));
 sg13g2_a22oi_1 _4092_ (.Y(_0349_),
    .B1(_0348_),
    .B2(_0022_),
    .A2(_0345_),
    .A1(net692));
 sg13g2_nand2_1 _4093_ (.Y(_0350_),
    .A(_0347_),
    .B(_0349_));
 sg13g2_nor2_1 _4094_ (.A(net698),
    .B(_2839_),
    .Y(_0351_));
 sg13g2_a21oi_1 _4095_ (.A1(net698),
    .A2(_0090_),
    .Y(_0352_),
    .B1(_0351_));
 sg13g2_and2_1 _4096_ (.A(net689),
    .B(_0346_),
    .X(_0353_));
 sg13g2_a221oi_1 _4097_ (.B2(net692),
    .C1(_0353_),
    .B1(_0352_),
    .A1(\generated._425[1] ),
    .Y(_0354_),
    .A2(_0348_));
 sg13g2_a21oi_1 _4098_ (.A1(_0350_),
    .A2(_0354_),
    .Y(_0355_),
    .B1(net606));
 sg13g2_nand2_1 _4099_ (.Y(_0356_),
    .A(net697),
    .B(_0020_));
 sg13g2_o21ai_1 _4100_ (.B1(_0356_),
    .Y(_0357_),
    .A1(net697),
    .A2(_2848_));
 sg13g2_nand2_1 _4101_ (.Y(_0358_),
    .A(net692),
    .B(_0357_));
 sg13g2_o21ai_1 _4102_ (.B1(_0358_),
    .Y(_0359_),
    .A1(net692),
    .A2(_0352_));
 sg13g2_xnor2_1 _4103_ (.Y(_0360_),
    .A(_0355_),
    .B(_0359_));
 sg13g2_inv_1 _4104_ (.Y(_0361_),
    .A(_0360_));
 sg13g2_nor2_1 _4105_ (.A(net606),
    .B(_0354_),
    .Y(_0362_));
 sg13g2_xnor2_1 _4106_ (.Y(_0363_),
    .A(_0350_),
    .B(_0362_));
 sg13g2_nor2_1 _4107_ (.A(_0025_),
    .B(_0363_),
    .Y(_0364_));
 sg13g2_nor2_1 _4108_ (.A(\generated._69[0] ),
    .B(_0354_),
    .Y(_0365_));
 sg13g2_xnor2_1 _4109_ (.Y(_0366_),
    .A(net506),
    .B(_0363_));
 sg13g2_nor2_1 _4110_ (.A(_0365_),
    .B(_0366_),
    .Y(_0367_));
 sg13g2_nor2_1 _4111_ (.A(_0364_),
    .B(_0367_),
    .Y(_0368_));
 sg13g2_xor2_1 _4112_ (.B(_0360_),
    .A(net433),
    .X(_0369_));
 sg13g2_nor2b_1 _4113_ (.A(_0368_),
    .B_N(_0369_),
    .Y(_0370_));
 sg13g2_a21oi_1 _4114_ (.A1(\generated._69[2] ),
    .A2(_0361_),
    .Y(_0371_),
    .B1(_0370_));
 sg13g2_nand3_1 _4115_ (.B(_0354_),
    .C(_0359_),
    .A(_0350_),
    .Y(_0372_));
 sg13g2_nand2_1 _4116_ (.Y(_0373_),
    .A(net609),
    .B(_0372_));
 sg13g2_nor2_1 _4117_ (.A(net692),
    .B(_0345_),
    .Y(_0374_));
 sg13g2_nor2b_1 _4118_ (.A(net697),
    .B_N(_0020_),
    .Y(_0375_));
 sg13g2_a21oi_2 _4119_ (.B1(_0375_),
    .Y(_0376_),
    .A2(_0021_),
    .A1(net697));
 sg13g2_a21oi_1 _4120_ (.A1(net692),
    .A2(_0376_),
    .Y(_0377_),
    .B1(_0374_));
 sg13g2_xnor2_1 _4121_ (.Y(_0378_),
    .A(_0373_),
    .B(_0377_));
 sg13g2_nand2b_1 _4122_ (.Y(_0379_),
    .B(_0378_),
    .A_N(_0018_));
 sg13g2_xor2_1 _4123_ (.B(_0378_),
    .A(net549),
    .X(_0380_));
 sg13g2_xnor2_1 _4124_ (.Y(_0381_),
    .A(_0371_),
    .B(_0380_));
 sg13g2_a22oi_1 _4125_ (.Y(\generated._938[3] ),
    .B1(net550),
    .B2(net643),
    .A2(_0337_),
    .A1(_0330_));
 sg13g2_o21ai_1 _4126_ (.B1(_0379_),
    .Y(_0382_),
    .A1(_0371_),
    .A2(_0380_));
 sg13g2_nand2b_1 _4127_ (.Y(_0383_),
    .B(_0377_),
    .A_N(_0372_));
 sg13g2_nand2_1 _4128_ (.Y(_0384_),
    .A(net608),
    .B(_0383_));
 sg13g2_nor2_1 _4129_ (.A(net690),
    .B(_0357_),
    .Y(_0385_));
 sg13g2_nor2b_1 _4130_ (.A(net697),
    .B_N(_0021_),
    .Y(_0386_));
 sg13g2_a21oi_1 _4131_ (.A1(net697),
    .A2(_0028_),
    .Y(_0387_),
    .B1(_0386_));
 sg13g2_a21oi_1 _4132_ (.A1(net691),
    .A2(_0387_),
    .Y(_0388_),
    .B1(_0385_));
 sg13g2_xnor2_1 _4133_ (.Y(_0389_),
    .A(_0384_),
    .B(_0388_));
 sg13g2_xor2_1 _4134_ (.B(_0389_),
    .A(net519),
    .X(_0390_));
 sg13g2_nor2b_1 _4135_ (.A(_0390_),
    .B_N(_0382_),
    .Y(_0391_));
 sg13g2_xor2_1 _4136_ (.B(_0390_),
    .A(_0382_),
    .X(_0392_));
 sg13g2_xnor2_1 _4137_ (.Y(_0393_),
    .A(_0026_),
    .B(_2878_));
 sg13g2_nand3b_1 _4138_ (.B(_0026_),
    .C(\generated._100[3] ),
    .Y(_0394_),
    .A_N(net723));
 sg13g2_xnor2_1 _4139_ (.Y(_0395_),
    .A(net723),
    .B(_0026_));
 sg13g2_xor2_1 _4140_ (.B(_0026_),
    .A(net723),
    .X(_0396_));
 sg13g2_nand3_1 _4141_ (.B(net729),
    .C(\generated._614[3] ),
    .A(net728),
    .Y(_0397_));
 sg13g2_inv_1 _4142_ (.Y(_0398_),
    .A(_0397_));
 sg13g2_a21o_1 _4143_ (.A2(net730),
    .A1(net729),
    .B1(net728),
    .X(_0399_));
 sg13g2_nand2_1 _4144_ (.Y(_0400_),
    .A(_0397_),
    .B(_0399_));
 sg13g2_o21ai_1 _4145_ (.B1(net646),
    .Y(_0401_),
    .A1(net616),
    .A2(_0400_));
 sg13g2_a221oi_1 _4146_ (.B2(net612),
    .C1(_0401_),
    .B1(_0395_),
    .A1(_0328_),
    .Y(_0402_),
    .A2(_0393_));
 sg13g2_a21oi_1 _4147_ (.A1(net640),
    .A2(_0392_),
    .Y(\generated._938[4] ),
    .B1(_0402_));
 sg13g2_xor2_1 _4148_ (.B(_2879_),
    .A(\generated._100[6] ),
    .X(_0403_));
 sg13g2_or2_1 _4149_ (.X(_0404_),
    .B(_0403_),
    .A(_0394_));
 sg13g2_xor2_1 _4150_ (.B(_0403_),
    .A(_0394_),
    .X(_0405_));
 sg13g2_xnor2_1 _4151_ (.Y(_0406_),
    .A(_0394_),
    .B(_0403_));
 sg13g2_nor2_1 _4152_ (.A(net726),
    .B(_0397_),
    .Y(_0407_));
 sg13g2_xor2_1 _4153_ (.B(_0397_),
    .A(net726),
    .X(_0408_));
 sg13g2_a22oi_1 _4154_ (.Y(_0409_),
    .B1(_0408_),
    .B2(net603),
    .A2(_0403_),
    .A1(net601));
 sg13g2_o21ai_1 _4155_ (.B1(_0409_),
    .Y(_0410_),
    .A1(_0332_),
    .A2(_0406_));
 sg13g2_nand2_1 _4156_ (.Y(_0411_),
    .A(net646),
    .B(_0410_));
 sg13g2_a21o_1 _4157_ (.A2(_0389_),
    .A1(\generated._69[4] ),
    .B1(_0391_),
    .X(_0412_));
 sg13g2_nor2b_1 _4158_ (.A(_0383_),
    .B_N(_0388_),
    .Y(_0413_));
 sg13g2_nor2_1 _4159_ (.A(net607),
    .B(_0413_),
    .Y(_0414_));
 sg13g2_mux2_1 _4160_ (.A0(_0028_),
    .A1(_0030_),
    .S(net695),
    .X(_0415_));
 sg13g2_nand2_1 _4161_ (.Y(_0416_),
    .A(net690),
    .B(_0415_));
 sg13g2_o21ai_1 _4162_ (.B1(_0416_),
    .Y(_0417_),
    .A1(net691),
    .A2(_0376_));
 sg13g2_xor2_1 _4163_ (.B(_0417_),
    .A(_0414_),
    .X(_0418_));
 sg13g2_inv_1 _4164_ (.Y(_0419_),
    .A(_0418_));
 sg13g2_nand2_1 _4165_ (.Y(_0420_),
    .A(net551),
    .B(_0419_));
 sg13g2_nand2b_1 _4166_ (.Y(_0421_),
    .B(_0418_),
    .A_N(_0029_));
 sg13g2_nand2_1 _4167_ (.Y(_0422_),
    .A(_0420_),
    .B(_0421_));
 sg13g2_xor2_1 _4168_ (.B(net552),
    .A(_0412_),
    .X(_0423_));
 sg13g2_o21ai_1 _4169_ (.B1(_0411_),
    .Y(\generated._938[5] ),
    .A1(net647),
    .A2(net553));
 sg13g2_a21oi_1 _4170_ (.A1(_0413_),
    .A2(_0417_),
    .Y(_0424_),
    .B1(net607));
 sg13g2_mux2_1 _4171_ (.A0(_0030_),
    .A1(_0032_),
    .S(net695),
    .X(_0425_));
 sg13g2_nand2_1 _4172_ (.Y(_0426_),
    .A(net690),
    .B(_0425_));
 sg13g2_o21ai_1 _4173_ (.B1(_0426_),
    .Y(_0427_),
    .A1(net691),
    .A2(_0387_));
 sg13g2_xor2_1 _4174_ (.B(_0427_),
    .A(_0424_),
    .X(_0428_));
 sg13g2_xor2_1 _4175_ (.B(_0428_),
    .A(_0031_),
    .X(_0429_));
 sg13g2_nand2_1 _4176_ (.Y(_0430_),
    .A(_0412_),
    .B(_0420_));
 sg13g2_a21oi_1 _4177_ (.A1(_0421_),
    .A2(_0430_),
    .Y(_0431_),
    .B1(_0429_));
 sg13g2_nand3_1 _4178_ (.B(_0429_),
    .C(_0430_),
    .A(_0421_),
    .Y(_0432_));
 sg13g2_nand2b_1 _4179_ (.Y(_0433_),
    .B(_0432_),
    .A_N(_0431_));
 sg13g2_nand3_1 _4180_ (.B(net722),
    .C(_2879_),
    .A(\generated._100[6] ),
    .Y(_0434_));
 sg13g2_nand2_2 _4181_ (.Y(_0435_),
    .A(_0319_),
    .B(_0434_));
 sg13g2_nor2_2 _4182_ (.A(_0404_),
    .B(_0435_),
    .Y(_0436_));
 sg13g2_xor2_1 _4183_ (.B(_0435_),
    .A(_0404_),
    .X(_0437_));
 sg13g2_nand2_1 _4184_ (.Y(_0438_),
    .A(net613),
    .B(net600));
 sg13g2_nor2_1 _4185_ (.A(\generated._221[1] ),
    .B(_0398_),
    .Y(_0439_));
 sg13g2_nor2_1 _4186_ (.A(\generated._221[1] ),
    .B(\generated._221[0] ),
    .Y(_0440_));
 sg13g2_nor3_2 _4187_ (.A(_0324_),
    .B(_0439_),
    .C(_0440_),
    .Y(_0441_));
 sg13g2_a221oi_1 _4188_ (.B2(net603),
    .C1(net641),
    .B1(_0441_),
    .A1(net601),
    .Y(_0442_),
    .A2(_0435_));
 sg13g2_a22oi_1 _4189_ (.Y(\generated._938[6] ),
    .B1(_0438_),
    .B2(_0442_),
    .A2(_0433_),
    .A1(net640));
 sg13g2_a21oi_1 _4190_ (.A1(net533),
    .A2(_0428_),
    .Y(_0443_),
    .B1(_0431_));
 sg13g2_nor2b_1 _4191_ (.A(net690),
    .B_N(_0415_),
    .Y(_0444_));
 sg13g2_a21oi_2 _4192_ (.B1(_0444_),
    .Y(_0445_),
    .A2(_0032_),
    .A1(net694));
 sg13g2_nand3_1 _4193_ (.B(_0417_),
    .C(_0427_),
    .A(_0413_),
    .Y(_0446_));
 sg13g2_nand2_1 _4194_ (.Y(_0447_),
    .A(net608),
    .B(_0446_));
 sg13g2_xor2_1 _4195_ (.B(_0447_),
    .A(_0445_),
    .X(_0448_));
 sg13g2_xnor2_1 _4196_ (.Y(_0449_),
    .A(_0033_),
    .B(_0448_));
 sg13g2_nand2b_1 _4197_ (.Y(_0450_),
    .B(_0449_),
    .A_N(_0443_));
 sg13g2_xor2_1 _4198_ (.B(_0449_),
    .A(_0443_),
    .X(_0451_));
 sg13g2_xor2_1 _4199_ (.B(_0319_),
    .A(net721),
    .X(_0452_));
 sg13g2_nand2b_1 _4200_ (.Y(_0453_),
    .B(_0436_),
    .A_N(_0452_));
 sg13g2_xnor2_1 _4201_ (.Y(_0454_),
    .A(_0436_),
    .B(_0452_));
 sg13g2_xor2_1 _4202_ (.B(_0452_),
    .A(_0436_),
    .X(_0455_));
 sg13g2_and3_1 _4203_ (.X(_0456_),
    .A(\generated._221[2] ),
    .B(\generated._221[1] ),
    .C(\generated._221[0] ));
 sg13g2_nand3_1 _4204_ (.B(net342),
    .C(net360),
    .A(net486),
    .Y(_0457_));
 sg13g2_a21oi_2 _4205_ (.B1(_0326_),
    .Y(_0458_),
    .A2(_0456_),
    .A1(_0398_));
 sg13g2_inv_1 _4206_ (.Y(_0459_),
    .A(_0458_));
 sg13g2_o21ai_1 _4207_ (.B1(net646),
    .Y(_0460_),
    .A1(net616),
    .A2(_0458_));
 sg13g2_a221oi_1 _4208_ (.B2(net612),
    .C1(_0460_),
    .B1(_0454_),
    .A1(net601),
    .Y(_0461_),
    .A2(_0452_));
 sg13g2_a21oi_1 _4209_ (.A1(net642),
    .A2(net534),
    .Y(\generated._938[7] ),
    .B1(_0461_));
 sg13g2_xnor2_1 _4210_ (.Y(_0462_),
    .A(\generated._221[3] ),
    .B(_0326_));
 sg13g2_or3_1 _4211_ (.A(_0331_),
    .B(net640),
    .C(_0462_),
    .X(_0463_));
 sg13g2_nand2_1 _4212_ (.Y(_0464_),
    .A(\generated._69[7] ),
    .B(_0448_));
 sg13g2_nor2b_1 _4213_ (.A(net690),
    .B_N(_0425_),
    .Y(_0465_));
 sg13g2_a21oi_1 _4214_ (.A1(net694),
    .A2(_0032_),
    .Y(_0466_),
    .B1(_0465_));
 sg13g2_o21ai_1 _4215_ (.B1(net608),
    .Y(_0467_),
    .A1(_0445_),
    .A2(_0446_));
 sg13g2_xor2_1 _4216_ (.B(_0467_),
    .A(_0466_),
    .X(_0468_));
 sg13g2_xor2_1 _4217_ (.B(_0468_),
    .A(net424),
    .X(_0469_));
 sg13g2_nand3_1 _4218_ (.B(_0464_),
    .C(_0469_),
    .A(_0450_),
    .Y(_0470_));
 sg13g2_a21oi_1 _4219_ (.A1(_0450_),
    .A2(_0464_),
    .Y(_0471_),
    .B1(_0469_));
 sg13g2_nand2_1 _4220_ (.Y(_0472_),
    .A(net642),
    .B(_0470_));
 sg13g2_o21ai_1 _4221_ (.B1(_0463_),
    .Y(\generated._938[8] ),
    .A1(net425),
    .A2(_0472_));
 sg13g2_nor2_1 _4222_ (.A(_0327_),
    .B(net640),
    .Y(_0473_));
 sg13g2_a21oi_1 _4223_ (.A1(net483),
    .A2(_0468_),
    .Y(_0474_),
    .B1(_0471_));
 sg13g2_nor3_1 _4224_ (.A(_0445_),
    .B(_0446_),
    .C(_0466_),
    .Y(_0475_));
 sg13g2_xnor2_1 _4225_ (.Y(_0476_),
    .A(net731),
    .B(_0475_));
 sg13g2_nand2_1 _4226_ (.Y(_0477_),
    .A(_0032_),
    .B(net607));
 sg13g2_o21ai_1 _4227_ (.B1(_0477_),
    .Y(_0478_),
    .A1(net607),
    .A2(_0476_));
 sg13g2_xnor2_1 _4228_ (.Y(_0479_),
    .A(_0023_),
    .B(_0478_));
 sg13g2_xor2_1 _4229_ (.B(_0479_),
    .A(_0474_),
    .X(_0480_));
 sg13g2_a21oi_1 _4230_ (.A1(net642),
    .A2(_0480_),
    .Y(\generated._938[9] ),
    .B1(_0473_));
 sg13g2_a21o_1 _4231_ (.A2(_0329_),
    .A1(net603),
    .B1(net640),
    .X(_0481_));
 sg13g2_a221oi_1 _4232_ (.B2(_0336_),
    .C1(_0481_),
    .B1(net612),
    .A1(_2837_),
    .Y(_0482_),
    .A2(net601));
 sg13g2_nor2b_1 _4233_ (.A(net697),
    .B_N(_0024_),
    .Y(_0483_));
 sg13g2_a21oi_1 _4234_ (.A1(net697),
    .A2(_0018_),
    .Y(_0484_),
    .B1(_0483_));
 sg13g2_nand2_1 _4235_ (.Y(_0485_),
    .A(net692),
    .B(_0484_));
 sg13g2_a22oi_1 _4236_ (.Y(_0486_),
    .B1(_0348_),
    .B2(\generated._69[0] ),
    .A2(_0346_),
    .A1(\generated._69[1] ));
 sg13g2_nand2_2 _4237_ (.Y(_0487_),
    .A(_0485_),
    .B(_0486_));
 sg13g2_and2_1 _4238_ (.A(\generated._425[1] ),
    .B(_0487_),
    .X(_0488_));
 sg13g2_mux2_1 _4239_ (.A0(_0018_),
    .A1(_0027_),
    .S(net696),
    .X(_0489_));
 sg13g2_nand2_1 _4240_ (.Y(_0490_),
    .A(_0024_),
    .B(_0346_));
 sg13g2_a22oi_1 _4241_ (.Y(_0491_),
    .B1(_0489_),
    .B2(net693),
    .A2(_0348_),
    .A1(_0025_));
 sg13g2_nand2_1 _4242_ (.Y(_0492_),
    .A(_0490_),
    .B(_0491_));
 sg13g2_nand2_1 _4243_ (.Y(_0493_),
    .A(_0342_),
    .B(_0487_));
 sg13g2_xor2_1 _4244_ (.B(_0493_),
    .A(_0492_),
    .X(_0494_));
 sg13g2_xnor2_1 _4245_ (.Y(_0495_),
    .A(net444),
    .B(_0494_));
 sg13g2_nand2_1 _4246_ (.Y(_0496_),
    .A(_0488_),
    .B(_0495_));
 sg13g2_nand2_1 _4247_ (.Y(_0497_),
    .A(net689),
    .B(_0494_));
 sg13g2_nand3_1 _4248_ (.B(_0486_),
    .C(_0492_),
    .A(_0485_),
    .Y(_0498_));
 sg13g2_nand2_1 _4249_ (.Y(_0499_),
    .A(net609),
    .B(_0498_));
 sg13g2_mux2_1 _4250_ (.A0(_0027_),
    .A1(_0029_),
    .S(net696),
    .X(_0500_));
 sg13g2_nand2_1 _4251_ (.Y(_0501_),
    .A(net693),
    .B(_0500_));
 sg13g2_o21ai_1 _4252_ (.B1(_0501_),
    .Y(_0502_),
    .A1(net692),
    .A2(_0484_));
 sg13g2_xor2_1 _4253_ (.B(_0502_),
    .A(_0499_),
    .X(_0503_));
 sg13g2_xnor2_1 _4254_ (.Y(_0504_),
    .A(\generated._66[2] ),
    .B(_0503_));
 sg13g2_a21o_1 _4255_ (.A2(_0497_),
    .A1(_0496_),
    .B1(_0504_),
    .X(_0505_));
 sg13g2_nand2_1 _4256_ (.Y(_0506_),
    .A(_2839_),
    .B(_0503_));
 sg13g2_nand2b_1 _4257_ (.Y(_0507_),
    .B(_0502_),
    .A_N(_0498_));
 sg13g2_nand2_1 _4258_ (.Y(_0508_),
    .A(net608),
    .B(_0507_));
 sg13g2_nor2_1 _4259_ (.A(net693),
    .B(_0489_),
    .Y(_0509_));
 sg13g2_nor2b_1 _4260_ (.A(net695),
    .B_N(_0029_),
    .Y(_0510_));
 sg13g2_a21oi_1 _4261_ (.A1(net696),
    .A2(_0031_),
    .Y(_0511_),
    .B1(_0510_));
 sg13g2_a21oi_1 _4262_ (.A1(net693),
    .A2(_0511_),
    .Y(_0512_),
    .B1(_0509_));
 sg13g2_xor2_1 _4263_ (.B(_0512_),
    .A(_0508_),
    .X(_0513_));
 sg13g2_xnor2_1 _4264_ (.Y(_0514_),
    .A(net740),
    .B(_0513_));
 sg13g2_a21oi_1 _4265_ (.A1(_0505_),
    .A2(_0506_),
    .Y(_0515_),
    .B1(_0514_));
 sg13g2_and3_1 _4266_ (.X(_0516_),
    .A(_0505_),
    .B(_0506_),
    .C(_0514_));
 sg13g2_o21ai_1 _4267_ (.B1(net644),
    .Y(_0517_),
    .A1(_0515_),
    .A2(_0516_));
 sg13g2_nor2b_1 _4268_ (.A(_0482_),
    .B_N(_0517_),
    .Y(\generated._889[3] ));
 sg13g2_a21oi_1 _4269_ (.A1(net740),
    .A2(_0513_),
    .Y(_0518_),
    .B1(_0515_));
 sg13g2_nand2b_1 _4270_ (.Y(_0519_),
    .B(_0512_),
    .A_N(_0507_));
 sg13g2_nand2_1 _4271_ (.Y(_0520_),
    .A(net608),
    .B(_0519_));
 sg13g2_nor2_1 _4272_ (.A(net693),
    .B(_0500_),
    .Y(_0521_));
 sg13g2_nor2b_1 _4273_ (.A(net695),
    .B_N(_0031_),
    .Y(_0522_));
 sg13g2_a21oi_1 _4274_ (.A1(net696),
    .A2(_0033_),
    .Y(_0523_),
    .B1(_0522_));
 sg13g2_a21oi_1 _4275_ (.A1(net693),
    .A2(_0523_),
    .Y(_0524_),
    .B1(_0521_));
 sg13g2_xor2_1 _4276_ (.B(_0524_),
    .A(_0520_),
    .X(_0525_));
 sg13g2_xnor2_1 _4277_ (.Y(_0526_),
    .A(net739),
    .B(_0525_));
 sg13g2_nor2_1 _4278_ (.A(_0518_),
    .B(_0526_),
    .Y(_0527_));
 sg13g2_xnor2_1 _4279_ (.Y(_0528_),
    .A(_0518_),
    .B(_0526_));
 sg13g2_nand3_1 _4280_ (.B(_0397_),
    .C(_0399_),
    .A(net612),
    .Y(_0529_));
 sg13g2_a221oi_1 _4281_ (.B2(net603),
    .C1(net641),
    .B1(_0393_),
    .A1(_2836_),
    .Y(_0530_),
    .A2(net601));
 sg13g2_a22oi_1 _4282_ (.Y(\generated._889[4] ),
    .B1(_0529_),
    .B2(_0530_),
    .A2(_0528_),
    .A1(net644));
 sg13g2_nand2_1 _4283_ (.Y(_0531_),
    .A(net726),
    .B(net601));
 sg13g2_a22oi_1 _4284_ (.Y(_0532_),
    .B1(_0408_),
    .B2(net612),
    .A2(_0403_),
    .A1(net602));
 sg13g2_a21oi_1 _4285_ (.A1(_0531_),
    .A2(_0532_),
    .Y(_0533_),
    .B1(net644));
 sg13g2_a21oi_1 _4286_ (.A1(_2848_),
    .A2(_0525_),
    .Y(_0534_),
    .B1(_0527_));
 sg13g2_nor2b_1 _4287_ (.A(_0519_),
    .B_N(_0524_),
    .Y(_0535_));
 sg13g2_nor2_1 _4288_ (.A(net606),
    .B(_0535_),
    .Y(_0536_));
 sg13g2_mux2_1 _4289_ (.A0(_0033_),
    .A1(_0034_),
    .S(net695),
    .X(_0537_));
 sg13g2_nand2_1 _4290_ (.Y(_0538_),
    .A(net691),
    .B(_0537_));
 sg13g2_o21ai_1 _4291_ (.B1(_0538_),
    .Y(_0539_),
    .A1(net691),
    .A2(_0511_));
 sg13g2_xor2_1 _4292_ (.B(_0539_),
    .A(_0536_),
    .X(_0540_));
 sg13g2_inv_1 _4293_ (.Y(_0541_),
    .A(_0540_));
 sg13g2_nor2_1 _4294_ (.A(\generated._66[5] ),
    .B(_0541_),
    .Y(_0542_));
 sg13g2_nand2_1 _4295_ (.Y(_0543_),
    .A(\generated._66[5] ),
    .B(_0541_));
 sg13g2_nor2b_1 _4296_ (.A(_0542_),
    .B_N(_0543_),
    .Y(_0544_));
 sg13g2_xnor2_1 _4297_ (.Y(_0545_),
    .A(_0534_),
    .B(_0544_));
 sg13g2_a21o_1 _4298_ (.A2(_0545_),
    .A1(net643),
    .B1(_0533_),
    .X(\generated._889[5] ));
 sg13g2_o21ai_1 _4299_ (.B1(_0543_),
    .Y(_0546_),
    .A1(_0534_),
    .A2(_0542_));
 sg13g2_a21oi_1 _4300_ (.A1(_0535_),
    .A2(_0539_),
    .Y(_0547_),
    .B1(net606));
 sg13g2_mux2_1 _4301_ (.A0(_0034_),
    .A1(_0023_),
    .S(net695),
    .X(_0548_));
 sg13g2_nand2_1 _4302_ (.Y(_0549_),
    .A(net691),
    .B(_0548_));
 sg13g2_o21ai_1 _4303_ (.B1(_0549_),
    .Y(_0550_),
    .A1(net691),
    .A2(_0523_));
 sg13g2_xor2_1 _4304_ (.B(_0550_),
    .A(_0547_),
    .X(_0551_));
 sg13g2_xor2_1 _4305_ (.B(_0551_),
    .A(net735),
    .X(_0552_));
 sg13g2_nor2b_1 _4306_ (.A(_0552_),
    .B_N(_0546_),
    .Y(_0553_));
 sg13g2_xor2_1 _4307_ (.B(_0552_),
    .A(_0546_),
    .X(_0554_));
 sg13g2_nand2_1 _4308_ (.Y(_0555_),
    .A(net612),
    .B(_0441_));
 sg13g2_nor2b_2 _4309_ (.A(_0441_),
    .B_N(_0407_),
    .Y(_0556_));
 sg13g2_xnor2_1 _4310_ (.Y(_0557_),
    .A(_0407_),
    .B(_0441_));
 sg13g2_a221oi_1 _4311_ (.B2(net601),
    .C1(net640),
    .B1(_0557_),
    .A1(net602),
    .Y(_0558_),
    .A2(_0435_));
 sg13g2_a22oi_1 _4312_ (.Y(\generated._889[6] ),
    .B1(_0555_),
    .B2(_0558_),
    .A2(_0554_),
    .A1(net644));
 sg13g2_nand2_1 _4313_ (.Y(_0559_),
    .A(_0328_),
    .B(_0556_));
 sg13g2_a221oi_1 _4314_ (.B2(net612),
    .C1(net640),
    .B1(_0459_),
    .A1(net720),
    .Y(_0560_),
    .A2(_0452_));
 sg13g2_nor2_1 _4315_ (.A(_0021_),
    .B(_0551_),
    .Y(_0561_));
 sg13g2_nor2b_1 _4316_ (.A(net694),
    .B_N(_0537_),
    .Y(_0562_));
 sg13g2_a21oi_2 _4317_ (.B1(_0562_),
    .Y(_0563_),
    .A2(_0023_),
    .A1(net690));
 sg13g2_nand3_1 _4318_ (.B(_0539_),
    .C(_0550_),
    .A(_0535_),
    .Y(_0564_));
 sg13g2_nand2_1 _4319_ (.Y(_0565_),
    .A(net608),
    .B(_0564_));
 sg13g2_xor2_1 _4320_ (.B(_0565_),
    .A(_0563_),
    .X(_0566_));
 sg13g2_xnor2_1 _4321_ (.Y(_0567_),
    .A(net734),
    .B(_0566_));
 sg13g2_o21ai_1 _4322_ (.B1(_0567_),
    .Y(_0568_),
    .A1(_0553_),
    .A2(_0561_));
 sg13g2_or3_1 _4323_ (.A(_0553_),
    .B(_0561_),
    .C(_0567_),
    .X(_0569_));
 sg13g2_nand2_1 _4324_ (.Y(_0570_),
    .A(_0568_),
    .B(_0569_));
 sg13g2_a22oi_1 _4325_ (.Y(\generated._889[7] ),
    .B1(_0570_),
    .B2(net641),
    .A2(_0560_),
    .A1(_0559_));
 sg13g2_xnor2_1 _4326_ (.Y(_0571_),
    .A(_2845_),
    .B(_0320_));
 sg13g2_o21ai_1 _4327_ (.B1(_0320_),
    .Y(_0572_),
    .A1(_2835_),
    .A2(_0326_));
 sg13g2_nand3_1 _4328_ (.B(_0571_),
    .C(_0572_),
    .A(net647),
    .Y(_0573_));
 sg13g2_o21ai_1 _4329_ (.B1(_0568_),
    .Y(_0574_),
    .A1(net547),
    .A2(_0566_));
 sg13g2_nor2b_1 _4330_ (.A(net690),
    .B_N(_0548_),
    .Y(_0575_));
 sg13g2_a21oi_1 _4331_ (.A1(net690),
    .A2(_0023_),
    .Y(_0576_),
    .B1(_0575_));
 sg13g2_o21ai_1 _4332_ (.B1(net608),
    .Y(_0577_),
    .A1(_0563_),
    .A2(_0564_));
 sg13g2_xor2_1 _4333_ (.B(_0577_),
    .A(_0576_),
    .X(_0578_));
 sg13g2_xnor2_1 _4334_ (.Y(_0579_),
    .A(net733),
    .B(_0578_));
 sg13g2_and2_1 _4335_ (.A(_0574_),
    .B(_0579_),
    .X(_0580_));
 sg13g2_o21ai_1 _4336_ (.B1(net643),
    .Y(_0581_),
    .A1(_0574_),
    .A2(_0579_));
 sg13g2_o21ai_1 _4337_ (.B1(_0573_),
    .Y(\generated._889[8] ),
    .A1(_0580_),
    .A2(_0581_));
 sg13g2_nor2_1 _4338_ (.A(net409),
    .B(_0578_),
    .Y(_0582_));
 sg13g2_nor2_1 _4339_ (.A(_0580_),
    .B(_0582_),
    .Y(_0583_));
 sg13g2_nor3_1 _4340_ (.A(_0563_),
    .B(_0564_),
    .C(_0576_),
    .Y(_0584_));
 sg13g2_o21ai_1 _4341_ (.B1(net608),
    .Y(_0585_),
    .A1(\generated._69[9] ),
    .A2(_0584_));
 sg13g2_a21oi_1 _4342_ (.A1(\generated._69[9] ),
    .A2(_0584_),
    .Y(_0586_),
    .B1(_0585_));
 sg13g2_nor2_1 _4343_ (.A(_0023_),
    .B(_0586_),
    .Y(_0587_));
 sg13g2_xnor2_1 _4344_ (.Y(_0588_),
    .A(net731),
    .B(_0587_));
 sg13g2_o21ai_1 _4345_ (.B1(net643),
    .Y(_0589_),
    .A1(_0583_),
    .A2(_0588_));
 sg13g2_a21oi_1 _4346_ (.A1(_0583_),
    .A2(_0588_),
    .Y(\generated._889[9] ),
    .B1(_0589_));
 sg13g2_nor3_2 _4347_ (.A(\generated._63[1] ),
    .B(\generated._63[0] ),
    .C(\generated._63[3] ),
    .Y(_0590_));
 sg13g2_nor2b_1 _4348_ (.A(\generated._63[2] ),
    .B_N(_0590_),
    .Y(_0591_));
 sg13g2_nand2b_2 _4349_ (.Y(_0592_),
    .B(_0590_),
    .A_N(\generated._63[2] ));
 sg13g2_xnor2_1 _4350_ (.Y(_0593_),
    .A(net326),
    .B(net614));
 sg13g2_nand2_2 _4351_ (.Y(_0594_),
    .A(net679),
    .B(net673));
 sg13g2_inv_1 _4352_ (.Y(_0595_),
    .A(_0594_));
 sg13g2_xnor2_1 _4353_ (.Y(_0596_),
    .A(net374),
    .B(_0594_));
 sg13g2_nor2_1 _4354_ (.A(net635),
    .B(_0596_),
    .Y(_0597_));
 sg13g2_a21oi_1 _4355_ (.A1(net635),
    .A2(_0593_),
    .Y(\generated._695[0] ),
    .B1(_0597_));
 sg13g2_nand2_1 _4356_ (.Y(_0598_),
    .A(net679),
    .B(net656));
 sg13g2_xnor2_1 _4357_ (.Y(_0599_),
    .A(net673),
    .B(net684));
 sg13g2_nor2_1 _4358_ (.A(net679),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_a21oi_2 _4359_ (.B1(_0600_),
    .Y(_0601_),
    .A2(net656),
    .A1(net679));
 sg13g2_nor2_2 _4360_ (.A(_0595_),
    .B(_0601_),
    .Y(_0602_));
 sg13g2_nor2_1 _4361_ (.A(net509),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_xnor2_1 _4362_ (.Y(_0604_),
    .A(_0044_),
    .B(_0602_));
 sg13g2_nand3_1 _4363_ (.B(_0594_),
    .C(_0604_),
    .A(net374),
    .Y(_0605_));
 sg13g2_a21oi_1 _4364_ (.A1(net374),
    .A2(_0594_),
    .Y(_0606_),
    .B1(_0604_));
 sg13g2_nor2_1 _4365_ (.A(net634),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_nand2_1 _4366_ (.Y(_0608_),
    .A(net375),
    .B(_0607_));
 sg13g2_nor2b_2 _4367_ (.A(net616),
    .B_N(_0037_),
    .Y(_0609_));
 sg13g2_nand2_2 _4368_ (.Y(_0610_),
    .A(_0037_),
    .B(net602));
 sg13g2_xnor2_1 _4369_ (.Y(_0611_),
    .A(\generated._434[11] ),
    .B(net610));
 sg13g2_a22oi_1 _4370_ (.Y(_0612_),
    .B1(_0611_),
    .B2(\generated._434[10] ),
    .A2(_0332_),
    .A1(_2853_));
 sg13g2_xnor2_1 _4371_ (.Y(_0613_),
    .A(\generated._434[13] ),
    .B(net610));
 sg13g2_xnor2_1 _4372_ (.Y(_0614_),
    .A(\generated._434[12] ),
    .B(net610));
 sg13g2_nand2b_1 _4373_ (.Y(_0615_),
    .B(_0614_),
    .A_N(_0613_));
 sg13g2_o21ai_1 _4374_ (.B1(\generated._434[13] ),
    .Y(_0616_),
    .A1(_2852_),
    .A2(net610));
 sg13g2_o21ai_1 _4375_ (.B1(_0616_),
    .Y(_0617_),
    .A1(_0612_),
    .A2(_0615_));
 sg13g2_xor2_1 _4376_ (.B(net611),
    .A(\generated._434[17] ),
    .X(_0618_));
 sg13g2_xnor2_1 _4377_ (.Y(_0619_),
    .A(_0039_),
    .B(net611));
 sg13g2_xnor2_1 _4378_ (.Y(_0620_),
    .A(\generated._434[14] ),
    .B(net611));
 sg13g2_xor2_1 _4379_ (.B(net610),
    .A(_0040_),
    .X(_0621_));
 sg13g2_and4_1 _4380_ (.A(_0618_),
    .B(_0619_),
    .C(_0620_),
    .D(_0621_),
    .X(_0622_));
 sg13g2_o21ai_1 _4381_ (.B1(net611),
    .Y(_0623_),
    .A1(\generated._434[17] ),
    .A2(\generated._434[16] ));
 sg13g2_a21oi_1 _4382_ (.A1(_0040_),
    .A2(_0041_),
    .Y(_0624_),
    .B1(net610));
 sg13g2_nand3_1 _4383_ (.B(_0619_),
    .C(_0624_),
    .A(_0618_),
    .Y(_0625_));
 sg13g2_nand2_1 _4384_ (.Y(_0626_),
    .A(_0623_),
    .B(_0625_));
 sg13g2_a21oi_1 _4385_ (.A1(_0617_),
    .A2(_0622_),
    .Y(_0627_),
    .B1(_0626_));
 sg13g2_xor2_1 _4386_ (.B(net613),
    .A(\generated._434[18] ),
    .X(_0628_));
 sg13g2_nor2_1 _4387_ (.A(_0627_),
    .B(_0628_),
    .Y(_0629_));
 sg13g2_xnor2_1 _4388_ (.Y(_0630_),
    .A(\generated._434[19] ),
    .B(net613));
 sg13g2_a21oi_1 _4389_ (.A1(_0037_),
    .A2(_0038_),
    .Y(_0631_),
    .B1(net613));
 sg13g2_nand2b_1 _4390_ (.Y(_0632_),
    .B(_0630_),
    .A_N(_0631_));
 sg13g2_inv_1 _4391_ (.Y(_0633_),
    .A(_0632_));
 sg13g2_o21ai_1 _4392_ (.B1(_0633_),
    .Y(_0634_),
    .A1(_0627_),
    .A2(_0628_));
 sg13g2_nand3b_1 _4393_ (.B(_0332_),
    .C(\generated._434[19] ),
    .Y(_0635_),
    .A_N(_0037_));
 sg13g2_nand2_1 _4394_ (.Y(_0636_),
    .A(_0634_),
    .B(_0635_));
 sg13g2_and3_1 _4395_ (.X(_0637_),
    .A(net616),
    .B(_0634_),
    .C(_0635_));
 sg13g2_nand3_1 _4396_ (.B(_0634_),
    .C(_0635_),
    .A(net616),
    .Y(_0638_));
 sg13g2_nor2_1 _4397_ (.A(_0609_),
    .B(net573),
    .Y(_0639_));
 sg13g2_nand2_2 _4398_ (.Y(_0640_),
    .A(_0610_),
    .B(net571));
 sg13g2_nor2_1 _4399_ (.A(_0043_),
    .B(net614),
    .Y(_0641_));
 sg13g2_xor2_1 _4400_ (.B(_0611_),
    .A(\generated._434[10] ),
    .X(_0642_));
 sg13g2_a21oi_1 _4401_ (.A1(net614),
    .A2(_0642_),
    .Y(_0643_),
    .B1(_0641_));
 sg13g2_nor2_1 _4402_ (.A(_0639_),
    .B(_0643_),
    .Y(_0644_));
 sg13g2_xnor2_1 _4403_ (.Y(_0645_),
    .A(_0640_),
    .B(_0643_));
 sg13g2_and2_1 _4404_ (.A(_0593_),
    .B(_0645_),
    .X(_0646_));
 sg13g2_o21ai_1 _4405_ (.B1(net634),
    .Y(_0647_),
    .A1(_0593_),
    .A2(_0645_));
 sg13g2_o21ai_1 _4406_ (.B1(_0608_),
    .Y(\generated._695[1] ),
    .A1(_0646_),
    .A2(_0647_));
 sg13g2_nor2_1 _4407_ (.A(_0042_),
    .B(net614),
    .Y(_0648_));
 sg13g2_nand2b_1 _4408_ (.Y(_0649_),
    .B(_0614_),
    .A_N(_0612_));
 sg13g2_xnor2_1 _4409_ (.Y(_0650_),
    .A(_0612_),
    .B(_0614_));
 sg13g2_a21oi_1 _4410_ (.A1(net614),
    .A2(_0650_),
    .Y(_0651_),
    .B1(_0648_));
 sg13g2_xnor2_1 _4411_ (.Y(_0652_),
    .A(_0640_),
    .B(_0651_));
 sg13g2_o21ai_1 _4412_ (.B1(_0652_),
    .Y(_0653_),
    .A1(_0644_),
    .A2(_0646_));
 sg13g2_nor3_1 _4413_ (.A(_0644_),
    .B(_0646_),
    .C(_0652_),
    .Y(_0654_));
 sg13g2_nand3b_1 _4414_ (.B(net634),
    .C(_0653_),
    .Y(_0655_),
    .A_N(_0654_));
 sg13g2_nor2b_2 _4415_ (.A(net673),
    .B_N(net679),
    .Y(_0656_));
 sg13g2_o21ai_1 _4416_ (.B1(_0598_),
    .Y(_0657_),
    .A1(net656),
    .A2(_0656_));
 sg13g2_nand2_1 _4417_ (.Y(_0658_),
    .A(\generated._505[2] ),
    .B(_0657_));
 sg13g2_xor2_1 _4418_ (.B(_0657_),
    .A(\generated._505[2] ),
    .X(_0659_));
 sg13g2_nor3_1 _4419_ (.A(_0603_),
    .B(_0606_),
    .C(_0659_),
    .Y(_0660_));
 sg13g2_o21ai_1 _4420_ (.B1(_0659_),
    .Y(_0661_),
    .A1(_0603_),
    .A2(_0606_));
 sg13g2_nand2_1 _4421_ (.Y(_0662_),
    .A(net633),
    .B(_0661_));
 sg13g2_o21ai_1 _4422_ (.B1(_0655_),
    .Y(\generated._695[2] ),
    .A1(_0660_),
    .A2(_0662_));
 sg13g2_nor2_1 _4423_ (.A(\generated._434[19] ),
    .B(net616),
    .Y(_0663_));
 sg13g2_or2_1 _4424_ (.X(_0664_),
    .B(net616),
    .A(\generated._434[19] ));
 sg13g2_nor2_2 _4425_ (.A(net573),
    .B(net597),
    .Y(_0665_));
 sg13g2_nand2_2 _4426_ (.Y(_0666_),
    .A(net571),
    .B(net596));
 sg13g2_o21ai_1 _4427_ (.B1(_0653_),
    .Y(_0667_),
    .A1(_0651_),
    .A2(_0665_));
 sg13g2_nor2_1 _4428_ (.A(_0045_),
    .B(net615),
    .Y(_0668_));
 sg13g2_o21ai_1 _4429_ (.B1(_0649_),
    .Y(_0669_),
    .A1(_0042_),
    .A2(net610));
 sg13g2_xnor2_1 _4430_ (.Y(_0670_),
    .A(_0613_),
    .B(_0669_));
 sg13g2_a21oi_1 _4431_ (.A1(net614),
    .A2(_0670_),
    .Y(_0671_),
    .B1(_0668_));
 sg13g2_nand2b_1 _4432_ (.Y(_0672_),
    .B(net569),
    .A_N(_0671_));
 sg13g2_xnor2_1 _4433_ (.Y(_0673_),
    .A(net569),
    .B(_0671_));
 sg13g2_nand2_1 _4434_ (.Y(_0674_),
    .A(_0667_),
    .B(_0673_));
 sg13g2_o21ai_1 _4435_ (.B1(net634),
    .Y(_0675_),
    .A1(_0667_),
    .A2(_0673_));
 sg13g2_nand2b_1 _4436_ (.Y(_0676_),
    .B(_0674_),
    .A_N(_0675_));
 sg13g2_nor2_1 _4437_ (.A(net566),
    .B(_0602_),
    .Y(_0677_));
 sg13g2_xnor2_1 _4438_ (.Y(_0678_),
    .A(net449),
    .B(_0602_));
 sg13g2_nand3_1 _4439_ (.B(_0661_),
    .C(_0678_),
    .A(_0658_),
    .Y(_0679_));
 sg13g2_a21oi_1 _4440_ (.A1(_0658_),
    .A2(_0661_),
    .Y(_0680_),
    .B1(_0678_));
 sg13g2_nand2_1 _4441_ (.Y(_0681_),
    .A(net633),
    .B(_0679_));
 sg13g2_o21ai_1 _4442_ (.B1(_0676_),
    .Y(\generated._695[3] ),
    .A1(net450),
    .A2(_0681_));
 sg13g2_nor2_1 _4443_ (.A(_0041_),
    .B(net614),
    .Y(_0682_));
 sg13g2_xor2_1 _4444_ (.B(_0620_),
    .A(_0617_),
    .X(_0683_));
 sg13g2_a21oi_2 _4445_ (.B1(_0682_),
    .Y(_0684_),
    .A2(_0683_),
    .A1(net614));
 sg13g2_xnor2_1 _4446_ (.Y(_0685_),
    .A(net569),
    .B(_0684_));
 sg13g2_nand3_1 _4447_ (.B(_0674_),
    .C(_0685_),
    .A(_0672_),
    .Y(_0686_));
 sg13g2_a21o_1 _4448_ (.A2(_0674_),
    .A1(_0672_),
    .B1(_0685_),
    .X(_0687_));
 sg13g2_nand3_1 _4449_ (.B(_0686_),
    .C(_0687_),
    .A(net634),
    .Y(_0688_));
 sg13g2_nor2_1 _4450_ (.A(_0677_),
    .B(_0680_),
    .Y(_0689_));
 sg13g2_and3_1 _4451_ (.X(_0690_),
    .A(\generated._505[4] ),
    .B(_0594_),
    .C(_0601_));
 sg13g2_a21oi_1 _4452_ (.A1(_0594_),
    .A2(_0601_),
    .Y(_0691_),
    .B1(\generated._505[4] ));
 sg13g2_or2_1 _4453_ (.X(_0692_),
    .B(_0691_),
    .A(_0690_));
 sg13g2_nor2_1 _4454_ (.A(_0689_),
    .B(_0692_),
    .Y(_0693_));
 sg13g2_a21o_1 _4455_ (.A2(_0692_),
    .A1(_0689_),
    .B1(net634),
    .X(_0694_));
 sg13g2_o21ai_1 _4456_ (.B1(_0688_),
    .Y(\generated._695[4] ),
    .A1(_0693_),
    .A2(_0694_));
 sg13g2_nand2b_1 _4457_ (.Y(_0695_),
    .B(\generated._505[5] ),
    .A_N(_0599_));
 sg13g2_xnor2_1 _4458_ (.Y(_0696_),
    .A(\generated._505[5] ),
    .B(_0599_));
 sg13g2_o21ai_1 _4459_ (.B1(_0696_),
    .Y(_0697_),
    .A1(_0690_),
    .A2(_0693_));
 sg13g2_or3_1 _4460_ (.A(_0690_),
    .B(_0693_),
    .C(_0696_),
    .X(_0698_));
 sg13g2_a21oi_1 _4461_ (.A1(_0697_),
    .A2(_0698_),
    .Y(_0699_),
    .B1(net634));
 sg13g2_o21ai_1 _4462_ (.B1(_0687_),
    .Y(_0700_),
    .A1(_0665_),
    .A2(_0684_));
 sg13g2_nand2_1 _4463_ (.Y(_0701_),
    .A(_0040_),
    .B(net602));
 sg13g2_a22oi_1 _4464_ (.Y(_0702_),
    .B1(_0617_),
    .B2(_0620_),
    .A2(_0332_),
    .A1(_2851_));
 sg13g2_xnor2_1 _4465_ (.Y(_0703_),
    .A(_0621_),
    .B(_0702_));
 sg13g2_o21ai_1 _4466_ (.B1(_0701_),
    .Y(_0704_),
    .A1(net602),
    .A2(_0703_));
 sg13g2_nor2_1 _4467_ (.A(net569),
    .B(_0704_),
    .Y(_0705_));
 sg13g2_nand2_1 _4468_ (.Y(_0706_),
    .A(net569),
    .B(_0704_));
 sg13g2_nor2b_1 _4469_ (.A(_0705_),
    .B_N(_0706_),
    .Y(_0707_));
 sg13g2_xnor2_1 _4470_ (.Y(_0708_),
    .A(_0700_),
    .B(_0707_));
 sg13g2_a21oi_1 _4471_ (.A1(net634),
    .A2(_0708_),
    .Y(\generated._695[5] ),
    .B1(_0699_));
 sg13g2_a21oi_1 _4472_ (.A1(_0700_),
    .A2(_0706_),
    .Y(_0709_),
    .B1(_0705_));
 sg13g2_nor2_1 _4473_ (.A(_0039_),
    .B(net617),
    .Y(_0710_));
 sg13g2_a21oi_1 _4474_ (.A1(_0617_),
    .A2(_0620_),
    .Y(_0711_),
    .B1(_0624_));
 sg13g2_a21oi_1 _4475_ (.A1(_0040_),
    .A2(net610),
    .Y(_0712_),
    .B1(_0711_));
 sg13g2_xor2_1 _4476_ (.B(_0712_),
    .A(_0619_),
    .X(_0713_));
 sg13g2_a21oi_2 _4477_ (.B1(_0710_),
    .Y(_0714_),
    .A2(_0713_),
    .A1(net615));
 sg13g2_xnor2_1 _4478_ (.Y(_0715_),
    .A(_0666_),
    .B(_0714_));
 sg13g2_or2_1 _4479_ (.X(_0716_),
    .B(_0715_),
    .A(_0709_));
 sg13g2_a21oi_1 _4480_ (.A1(_0709_),
    .A2(_0715_),
    .Y(_0717_),
    .B1(net633));
 sg13g2_nand2_1 _4481_ (.Y(_0718_),
    .A(_0716_),
    .B(_0717_));
 sg13g2_nor2b_1 _4482_ (.A(_0601_),
    .B_N(\generated._505[6] ),
    .Y(_0719_));
 sg13g2_xor2_1 _4483_ (.B(_0601_),
    .A(net514),
    .X(_0720_));
 sg13g2_nand3_1 _4484_ (.B(_0697_),
    .C(_0720_),
    .A(_0695_),
    .Y(_0721_));
 sg13g2_a21oi_1 _4485_ (.A1(_0695_),
    .A2(_0697_),
    .Y(_0722_),
    .B1(_0720_));
 sg13g2_nand2_1 _4486_ (.Y(_0723_),
    .A(net632),
    .B(_0721_));
 sg13g2_o21ai_1 _4487_ (.B1(_0718_),
    .Y(\generated._695[6] ),
    .A1(_0722_),
    .A2(_0723_));
 sg13g2_o21ai_1 _4488_ (.B1(_0716_),
    .Y(_0724_),
    .A1(_0640_),
    .A2(_0714_));
 sg13g2_a22oi_1 _4489_ (.Y(_0725_),
    .B1(_0619_),
    .B2(_0712_),
    .A2(net611),
    .A1(\generated._434[16] ));
 sg13g2_xnor2_1 _4490_ (.Y(_0726_),
    .A(_0618_),
    .B(_0725_));
 sg13g2_nand2_1 _4491_ (.Y(_0727_),
    .A(net617),
    .B(_0726_));
 sg13g2_o21ai_1 _4492_ (.B1(_0727_),
    .Y(_0728_),
    .A1(_0047_),
    .A2(net615));
 sg13g2_xnor2_1 _4493_ (.Y(_0729_),
    .A(_0665_),
    .B(_0728_));
 sg13g2_inv_1 _4494_ (.Y(_0730_),
    .A(_0729_));
 sg13g2_xnor2_1 _4495_ (.Y(_0731_),
    .A(_0724_),
    .B(_0730_));
 sg13g2_or2_1 _4496_ (.X(_0732_),
    .B(_0722_),
    .A(_0719_));
 sg13g2_nand2b_1 _4497_ (.Y(_0733_),
    .B(net685),
    .A_N(\generated._505[7] ));
 sg13g2_nor2b_1 _4498_ (.A(net684),
    .B_N(\generated._505[7] ),
    .Y(_0734_));
 sg13g2_xor2_1 _4499_ (.B(net540),
    .A(net684),
    .X(_0735_));
 sg13g2_xnor2_1 _4500_ (.Y(_0736_),
    .A(_0732_),
    .B(_0735_));
 sg13g2_nor2_1 _4501_ (.A(net635),
    .B(_0736_),
    .Y(_0737_));
 sg13g2_a21oi_1 _4502_ (.A1(net635),
    .A2(_0731_),
    .Y(\generated._695[7] ),
    .B1(_0737_));
 sg13g2_xor2_1 _4503_ (.B(net684),
    .A(\generated._505[8] ),
    .X(_0738_));
 sg13g2_a21oi_1 _4504_ (.A1(_0732_),
    .A2(_0733_),
    .Y(_0739_),
    .B1(_0734_));
 sg13g2_o21ai_1 _4505_ (.B1(net632),
    .Y(_0740_),
    .A1(_0738_),
    .A2(_0739_));
 sg13g2_a21o_1 _4506_ (.A2(_0739_),
    .A1(_0738_),
    .B1(_0740_),
    .X(_0741_));
 sg13g2_a22oi_1 _4507_ (.Y(_0742_),
    .B1(_0730_),
    .B2(_0724_),
    .A2(_0728_),
    .A1(net569));
 sg13g2_nand2_1 _4508_ (.Y(_0743_),
    .A(_0627_),
    .B(_0628_));
 sg13g2_nor2_1 _4509_ (.A(net602),
    .B(_0629_),
    .Y(_0744_));
 sg13g2_a22oi_1 _4510_ (.Y(_0745_),
    .B1(_0743_),
    .B2(_0744_),
    .A2(net602),
    .A1(_2849_));
 sg13g2_inv_1 _4511_ (.Y(_0746_),
    .A(_0745_));
 sg13g2_xnor2_1 _4512_ (.Y(_0747_),
    .A(net569),
    .B(_0745_));
 sg13g2_nor2_1 _4513_ (.A(_0742_),
    .B(_0747_),
    .Y(_0748_));
 sg13g2_a21o_1 _4514_ (.A2(_0747_),
    .A1(_0742_),
    .B1(net633),
    .X(_0749_));
 sg13g2_o21ai_1 _4515_ (.B1(_0741_),
    .Y(\generated._695[8] ),
    .A1(_0748_),
    .A2(_0749_));
 sg13g2_a21oi_1 _4516_ (.A1(net383),
    .A2(net656),
    .Y(_0750_),
    .B1(_0740_));
 sg13g2_a21oi_1 _4517_ (.A1(_0666_),
    .A2(_0746_),
    .Y(_0751_),
    .B1(_0748_));
 sg13g2_a21oi_1 _4518_ (.A1(_2849_),
    .A2(_0332_),
    .Y(_0752_),
    .B1(_0629_));
 sg13g2_xnor2_1 _4519_ (.Y(_0753_),
    .A(_0630_),
    .B(_0752_));
 sg13g2_a21oi_1 _4520_ (.A1(_0636_),
    .A2(_0753_),
    .Y(_0754_),
    .B1(net602));
 sg13g2_o21ai_1 _4521_ (.B1(_0754_),
    .Y(_0755_),
    .A1(_0636_),
    .A2(_0753_));
 sg13g2_xnor2_1 _4522_ (.Y(_0756_),
    .A(_0751_),
    .B(_0755_));
 sg13g2_a21o_1 _4523_ (.A2(_0756_),
    .A1(net635),
    .B1(_0750_),
    .X(\generated._695[9] ));
 sg13g2_or3_1 _4524_ (.A(net658),
    .B(\generated._394[2] ),
    .C(\generated._394[1] ),
    .X(_0757_));
 sg13g2_or2_1 _4525_ (.X(_0758_),
    .B(_0757_),
    .A(\generated._394[3] ));
 sg13g2_or2_2 _4526_ (.X(_0759_),
    .B(_0758_),
    .A(\generated._394[4] ));
 sg13g2_xnor2_1 _4527_ (.Y(_0760_),
    .A(\generated._394[5] ),
    .B(_0759_));
 sg13g2_nor2b_1 _4528_ (.A(net715),
    .B_N(_0049_),
    .Y(_0761_));
 sg13g2_a21oi_2 _4529_ (.B1(_0761_),
    .Y(_0762_),
    .A2(_0760_),
    .A1(net714));
 sg13g2_nand2_1 _4530_ (.Y(_0763_),
    .A(\generated._394[0] ),
    .B(_0762_));
 sg13g2_xnor2_1 _4531_ (.Y(_0764_),
    .A(_2843_),
    .B(_0762_));
 sg13g2_nor2_1 _4532_ (.A(_0048_),
    .B(net714),
    .Y(_0765_));
 sg13g2_nand2_1 _4533_ (.Y(_0766_),
    .A(\generated._394[4] ),
    .B(_0758_));
 sg13g2_nand3_1 _4534_ (.B(_0759_),
    .C(_0766_),
    .A(net714),
    .Y(_0767_));
 sg13g2_nor2b_2 _4535_ (.A(_0765_),
    .B_N(_0767_),
    .Y(_0768_));
 sg13g2_nand2b_2 _4536_ (.Y(_0769_),
    .B(_0767_),
    .A_N(_0765_));
 sg13g2_nand2_1 _4537_ (.Y(_0770_),
    .A(\generated._394[3] ),
    .B(_0757_));
 sg13g2_nand3_1 _4538_ (.B(_0758_),
    .C(_0770_),
    .A(net714),
    .Y(_0771_));
 sg13g2_o21ai_1 _4539_ (.B1(_0771_),
    .Y(_0772_),
    .A1(net714),
    .A2(_0050_));
 sg13g2_inv_1 _4540_ (.Y(_0773_),
    .A(_0772_));
 sg13g2_o21ai_1 _4541_ (.B1(\generated._394[2] ),
    .Y(_0774_),
    .A1(net658),
    .A2(\generated._394[1] ));
 sg13g2_nand3_1 _4542_ (.B(_0757_),
    .C(_0774_),
    .A(net714),
    .Y(_0775_));
 sg13g2_o21ai_1 _4543_ (.B1(_0775_),
    .Y(_0776_),
    .A1(net714),
    .A2(_0053_));
 sg13g2_nand2b_1 _4544_ (.Y(_0777_),
    .B(_0772_),
    .A_N(_0776_));
 sg13g2_xnor2_1 _4545_ (.Y(_0778_),
    .A(_0769_),
    .B(_0777_));
 sg13g2_xor2_1 _4546_ (.B(_0778_),
    .A(_0764_),
    .X(_0779_));
 sg13g2_nor2_1 _4547_ (.A(net715),
    .B(_0052_),
    .Y(_0780_));
 sg13g2_xor2_1 _4548_ (.B(\generated._394[1] ),
    .A(net658),
    .X(_0781_));
 sg13g2_a21oi_2 _4549_ (.B1(_0780_),
    .Y(_0782_),
    .A2(_0781_),
    .A1(net714));
 sg13g2_nand2_1 _4550_ (.Y(_0783_),
    .A(_0773_),
    .B(_0776_));
 sg13g2_nor2_1 _4551_ (.A(_0782_),
    .B(_0783_),
    .Y(_0784_));
 sg13g2_nor2_1 _4552_ (.A(_0779_),
    .B(_0784_),
    .Y(_0785_));
 sg13g2_and2_1 _4553_ (.A(_0776_),
    .B(_0782_),
    .X(_0786_));
 sg13g2_xor2_1 _4554_ (.B(_0786_),
    .A(_0772_),
    .X(_0787_));
 sg13g2_a21oi_1 _4555_ (.A1(_0769_),
    .A2(_0787_),
    .Y(_0788_),
    .B1(_0784_));
 sg13g2_nor2b_2 _4556_ (.A(_0788_),
    .B_N(_0779_),
    .Y(_0789_));
 sg13g2_xnor2_1 _4557_ (.Y(_0790_),
    .A(_0769_),
    .B(_0787_));
 sg13g2_nor3_1 _4558_ (.A(_0785_),
    .B(_0789_),
    .C(_0790_),
    .Y(_0791_));
 sg13g2_and2_1 _4559_ (.A(_0772_),
    .B(_0776_),
    .X(_0792_));
 sg13g2_nor2_1 _4560_ (.A(net658),
    .B(_0782_),
    .Y(_0793_));
 sg13g2_nand2_1 _4561_ (.Y(_0794_),
    .A(_0792_),
    .B(_0793_));
 sg13g2_nand3_1 _4562_ (.B(_0773_),
    .C(_0786_),
    .A(net658),
    .Y(_0795_));
 sg13g2_nand2_1 _4563_ (.Y(_0796_),
    .A(_0794_),
    .B(_0795_));
 sg13g2_nor2_1 _4564_ (.A(net590),
    .B(_0768_),
    .Y(_0797_));
 sg13g2_and2_1 _4565_ (.A(_0784_),
    .B(_0797_),
    .X(_0798_));
 sg13g2_a22oi_1 _4566_ (.Y(_0799_),
    .B1(_0798_),
    .B2(net658),
    .A2(_0796_),
    .A1(_0791_));
 sg13g2_a21oi_1 _4567_ (.A1(_2843_),
    .A2(_0777_),
    .Y(_0800_),
    .B1(_0782_));
 sg13g2_or2_1 _4568_ (.X(_0801_),
    .B(_0800_),
    .A(_0786_));
 sg13g2_nand3_1 _4569_ (.B(_0791_),
    .C(_0801_),
    .A(_0783_),
    .Y(_0802_));
 sg13g2_a22oi_1 _4570_ (.Y(_0803_),
    .B1(_0792_),
    .B2(_0768_),
    .A2(_0778_),
    .A1(_0764_));
 sg13g2_o21ai_1 _4571_ (.B1(\generated._394[6] ),
    .Y(_0804_),
    .A1(\generated._394[5] ),
    .A2(_0759_));
 sg13g2_nor3_2 _4572_ (.A(\generated._394[5] ),
    .B(\generated._394[6] ),
    .C(_0759_),
    .Y(_0805_));
 sg13g2_nand3b_1 _4573_ (.B(net715),
    .C(_0804_),
    .Y(_0806_),
    .A_N(_0805_));
 sg13g2_o21ai_1 _4574_ (.B1(_0806_),
    .Y(_0807_),
    .A1(net715),
    .A2(_0051_));
 sg13g2_nand2b_1 _4575_ (.Y(_0808_),
    .B(net583),
    .A_N(_0782_));
 sg13g2_xor2_1 _4576_ (.B(_0807_),
    .A(_0782_),
    .X(_0809_));
 sg13g2_nor2_1 _4577_ (.A(_0768_),
    .B(_0772_),
    .Y(_0810_));
 sg13g2_xnor2_1 _4578_ (.Y(_0811_),
    .A(net590),
    .B(_0810_));
 sg13g2_nor2_1 _4579_ (.A(_0809_),
    .B(_0811_),
    .Y(_0812_));
 sg13g2_xnor2_1 _4580_ (.Y(_0813_),
    .A(_0809_),
    .B(_0811_));
 sg13g2_nor2_1 _4581_ (.A(_0803_),
    .B(_0813_),
    .Y(_0814_));
 sg13g2_xor2_1 _4582_ (.B(_0813_),
    .A(_0803_),
    .X(_0815_));
 sg13g2_nor2b_1 _4583_ (.A(_0763_),
    .B_N(_0815_),
    .Y(_0816_));
 sg13g2_xnor2_1 _4584_ (.Y(_0817_),
    .A(_0763_),
    .B(_0815_));
 sg13g2_nand2_1 _4585_ (.Y(_0818_),
    .A(_0789_),
    .B(_0817_));
 sg13g2_xor2_1 _4586_ (.B(_0817_),
    .A(_0789_),
    .X(_0819_));
 sg13g2_nor2b_1 _4587_ (.A(_0802_),
    .B_N(_0819_),
    .Y(_0820_));
 sg13g2_xnor2_1 _4588_ (.Y(_0821_),
    .A(_0802_),
    .B(_0819_));
 sg13g2_nor2b_1 _4589_ (.A(_0799_),
    .B_N(_0821_),
    .Y(_0822_));
 sg13g2_xor2_1 _4590_ (.B(_0821_),
    .A(_0799_),
    .X(_0823_));
 sg13g2_nand2_1 _4591_ (.Y(_0824_),
    .A(net682),
    .B(_0055_));
 sg13g2_o21ai_1 _4592_ (.B1(_0824_),
    .Y(_0825_),
    .A1(net680),
    .A2(_2857_));
 sg13g2_nor2b_1 _4593_ (.A(_0825_),
    .B_N(net676),
    .Y(_0826_));
 sg13g2_nor2_2 _4594_ (.A(net679),
    .B(net673),
    .Y(_0827_));
 sg13g2_a221oi_1 _4595_ (.B2(net686),
    .C1(_0826_),
    .B1(_0827_),
    .A1(\generated._512[0] ),
    .Y(_0828_),
    .A2(_0656_));
 sg13g2_or2_1 _4596_ (.X(_0829_),
    .B(_0828_),
    .A(net700));
 sg13g2_a21oi_1 _4597_ (.A1(net700),
    .A2(_0828_),
    .Y(_0830_),
    .B1(net637));
 sg13g2_a22oi_1 _4598_ (.Y(\generated._561[0] ),
    .B1(_0829_),
    .B2(_0830_),
    .A2(_0823_),
    .A1(net637));
 sg13g2_nor2_1 _4599_ (.A(_0814_),
    .B(_0816_),
    .Y(_0831_));
 sg13g2_a21oi_1 _4600_ (.A1(_0772_),
    .A2(_0797_),
    .Y(_0832_),
    .B1(_0812_));
 sg13g2_nand2_1 _4601_ (.Y(_0833_),
    .A(_2858_),
    .B(_0805_));
 sg13g2_o21ai_1 _4602_ (.B1(net713),
    .Y(_0834_),
    .A1(_2858_),
    .A2(_0805_));
 sg13g2_nand2b_1 _4603_ (.Y(_0835_),
    .B(_0833_),
    .A_N(_0834_));
 sg13g2_o21ai_1 _4604_ (.B1(_0835_),
    .Y(_0836_),
    .A1(net713),
    .A2(_0056_));
 sg13g2_inv_1 _4605_ (.Y(_0837_),
    .A(_0836_));
 sg13g2_nand2_1 _4606_ (.Y(_0838_),
    .A(_0776_),
    .B(_0836_));
 sg13g2_xnor2_1 _4607_ (.Y(_0839_),
    .A(_0776_),
    .B(_0836_));
 sg13g2_and2_1 _4608_ (.A(net590),
    .B(_0768_),
    .X(_0840_));
 sg13g2_xnor2_1 _4609_ (.Y(_0841_),
    .A(net583),
    .B(_0840_));
 sg13g2_nor2_1 _4610_ (.A(_0839_),
    .B(_0841_),
    .Y(_0842_));
 sg13g2_xnor2_1 _4611_ (.Y(_0843_),
    .A(_0839_),
    .B(_0841_));
 sg13g2_or2_1 _4612_ (.X(_0844_),
    .B(_0843_),
    .A(_0832_));
 sg13g2_xnor2_1 _4613_ (.Y(_0845_),
    .A(_0832_),
    .B(_0843_));
 sg13g2_xor2_1 _4614_ (.B(_0845_),
    .A(_0808_),
    .X(_0846_));
 sg13g2_nand2b_1 _4615_ (.Y(_0847_),
    .B(_0846_),
    .A_N(_0831_));
 sg13g2_xor2_1 _4616_ (.B(_0846_),
    .A(_0831_),
    .X(_0848_));
 sg13g2_xor2_1 _4617_ (.B(_0848_),
    .A(_0818_),
    .X(_0849_));
 sg13g2_or3_1 _4618_ (.A(_0820_),
    .B(_0822_),
    .C(_0849_),
    .X(_0850_));
 sg13g2_o21ai_1 _4619_ (.B1(_0849_),
    .Y(_0851_),
    .A1(_0820_),
    .A2(_0822_));
 sg13g2_nand3_1 _4620_ (.B(_0850_),
    .C(_0851_),
    .A(net636),
    .Y(_0852_));
 sg13g2_mux2_1 _4621_ (.A0(_0055_),
    .A1(_0059_),
    .S(net680),
    .X(_0853_));
 sg13g2_nand2_1 _4622_ (.Y(_0854_),
    .A(_0058_),
    .B(_0827_));
 sg13g2_a22oi_1 _4623_ (.Y(_0855_),
    .B1(_0853_),
    .B2(net677),
    .A2(_0656_),
    .A1(_0054_));
 sg13g2_nand2_1 _4624_ (.Y(_0856_),
    .A(_0854_),
    .B(_0855_));
 sg13g2_nor2_1 _4625_ (.A(net657),
    .B(_0828_),
    .Y(_0857_));
 sg13g2_xnor2_1 _4626_ (.Y(_0858_),
    .A(_0856_),
    .B(_0857_));
 sg13g2_nor2_1 _4627_ (.A(_0057_),
    .B(_0858_),
    .Y(_0859_));
 sg13g2_xor2_1 _4628_ (.B(_0858_),
    .A(net561),
    .X(_0860_));
 sg13g2_and2_1 _4629_ (.A(_0829_),
    .B(_0860_),
    .X(_0861_));
 sg13g2_o21ai_1 _4630_ (.B1(_0592_),
    .Y(_0862_),
    .A1(_0829_),
    .A2(_0860_));
 sg13g2_o21ai_1 _4631_ (.B1(_0852_),
    .Y(\generated._561[1] ),
    .A1(_0861_),
    .A2(_0862_));
 sg13g2_o21ai_1 _4632_ (.B1(_0851_),
    .Y(_0863_),
    .A1(_0818_),
    .A2(_0848_));
 sg13g2_o21ai_1 _4633_ (.B1(_0844_),
    .Y(_0864_),
    .A1(_0808_),
    .A2(_0845_));
 sg13g2_nand3b_1 _4634_ (.B(_0769_),
    .C(net590),
    .Y(_0865_),
    .A_N(_0807_));
 sg13g2_nor2b_1 _4635_ (.A(_0842_),
    .B_N(_0865_),
    .Y(_0866_));
 sg13g2_nor2_1 _4636_ (.A(net713),
    .B(_0060_),
    .Y(_0867_));
 sg13g2_nor2_1 _4637_ (.A(\generated._394[8] ),
    .B(_0833_),
    .Y(_0868_));
 sg13g2_xor2_1 _4638_ (.B(_0833_),
    .A(\generated._394[8] ),
    .X(_0869_));
 sg13g2_a21oi_1 _4639_ (.A1(net713),
    .A2(_0869_),
    .Y(_0870_),
    .B1(_0867_));
 sg13g2_inv_1 _4640_ (.Y(_0871_),
    .A(_0870_));
 sg13g2_xnor2_1 _4641_ (.Y(_0872_),
    .A(_0772_),
    .B(net579));
 sg13g2_nand2b_1 _4642_ (.Y(_0873_),
    .B(net583),
    .A_N(net590));
 sg13g2_xnor2_1 _4643_ (.Y(_0874_),
    .A(_0836_),
    .B(_0873_));
 sg13g2_nand2_1 _4644_ (.Y(_0875_),
    .A(_0872_),
    .B(_0874_));
 sg13g2_xor2_1 _4645_ (.B(_0874_),
    .A(_0872_),
    .X(_0876_));
 sg13g2_inv_1 _4646_ (.Y(_0877_),
    .A(_0876_));
 sg13g2_xnor2_1 _4647_ (.Y(_0878_),
    .A(_0866_),
    .B(_0876_));
 sg13g2_nand2b_1 _4648_ (.Y(_0879_),
    .B(_0878_),
    .A_N(_0838_));
 sg13g2_xnor2_1 _4649_ (.Y(_0880_),
    .A(_0838_),
    .B(_0878_));
 sg13g2_nand2_1 _4650_ (.Y(_0881_),
    .A(_0864_),
    .B(_0880_));
 sg13g2_xnor2_1 _4651_ (.Y(_0882_),
    .A(_0864_),
    .B(_0880_));
 sg13g2_nor2_1 _4652_ (.A(_0847_),
    .B(_0882_),
    .Y(_0883_));
 sg13g2_xor2_1 _4653_ (.B(_0882_),
    .A(_0847_),
    .X(_0884_));
 sg13g2_and2_1 _4654_ (.A(_0863_),
    .B(_0884_),
    .X(_0885_));
 sg13g2_o21ai_1 _4655_ (.B1(net636),
    .Y(_0886_),
    .A1(_0863_),
    .A2(_0884_));
 sg13g2_nor2_1 _4656_ (.A(_0859_),
    .B(_0861_),
    .Y(_0887_));
 sg13g2_a21oi_1 _4657_ (.A1(_0828_),
    .A2(_0856_),
    .Y(_0888_),
    .B1(net657));
 sg13g2_mux2_1 _4658_ (.A0(_0059_),
    .A1(_0062_),
    .S(net682),
    .X(_0889_));
 sg13g2_mux2_1 _4659_ (.A0(_0825_),
    .A1(_0889_),
    .S(net676),
    .X(_0890_));
 sg13g2_xnor2_1 _4660_ (.Y(_0891_),
    .A(_0888_),
    .B(_0890_));
 sg13g2_xnor2_1 _4661_ (.Y(_0892_),
    .A(_0061_),
    .B(_0891_));
 sg13g2_nor2_1 _4662_ (.A(_0887_),
    .B(_0892_),
    .Y(_0893_));
 sg13g2_a21oi_1 _4663_ (.A1(_0887_),
    .A2(_0892_),
    .Y(_0894_),
    .B1(net637));
 sg13g2_nand2b_2 _4664_ (.Y(_0895_),
    .B(_0894_),
    .A_N(_0893_));
 sg13g2_o21ai_1 _4665_ (.B1(_0895_),
    .Y(\generated._561[2] ),
    .A1(_0885_),
    .A2(_0886_));
 sg13g2_o21ai_1 _4666_ (.B1(_0879_),
    .Y(_0896_),
    .A1(_0866_),
    .A2(_0877_));
 sg13g2_nand2_1 _4667_ (.Y(_0897_),
    .A(net590),
    .B(net583));
 sg13g2_o21ai_1 _4668_ (.B1(_0875_),
    .Y(_0898_),
    .A1(_0836_),
    .A2(_0897_));
 sg13g2_xnor2_1 _4669_ (.Y(_0899_),
    .A(\generated._394[9] ),
    .B(_0868_));
 sg13g2_mux2_2 _4670_ (.A0(_2860_),
    .A1(_0899_),
    .S(net713),
    .X(_0900_));
 sg13g2_nand2_1 _4671_ (.Y(_0901_),
    .A(_0769_),
    .B(net577));
 sg13g2_xnor2_1 _4672_ (.Y(_0902_),
    .A(_0768_),
    .B(net577));
 sg13g2_nor2_1 _4673_ (.A(net583),
    .B(_0837_),
    .Y(_0903_));
 sg13g2_xnor2_1 _4674_ (.Y(_0904_),
    .A(net579),
    .B(_0903_));
 sg13g2_nand2_1 _4675_ (.Y(_0905_),
    .A(_0902_),
    .B(_0904_));
 sg13g2_xor2_1 _4676_ (.B(_0904_),
    .A(_0902_),
    .X(_0906_));
 sg13g2_xnor2_1 _4677_ (.Y(_0907_),
    .A(_0898_),
    .B(_0906_));
 sg13g2_nor3_1 _4678_ (.A(_0773_),
    .B(net579),
    .C(_0907_),
    .Y(_0908_));
 sg13g2_o21ai_1 _4679_ (.B1(_0907_),
    .Y(_0909_),
    .A1(_0773_),
    .A2(net579));
 sg13g2_nor2b_1 _4680_ (.A(_0908_),
    .B_N(_0909_),
    .Y(_0910_));
 sg13g2_nand2_1 _4681_ (.Y(_0911_),
    .A(_0896_),
    .B(_0910_));
 sg13g2_xnor2_1 _4682_ (.Y(_0912_),
    .A(_0896_),
    .B(_0910_));
 sg13g2_nor2_1 _4683_ (.A(_0881_),
    .B(_0912_),
    .Y(_0913_));
 sg13g2_xor2_1 _4684_ (.B(_0912_),
    .A(_0881_),
    .X(_0914_));
 sg13g2_nor3_1 _4685_ (.A(_0883_),
    .B(_0885_),
    .C(_0914_),
    .Y(_0915_));
 sg13g2_o21ai_1 _4686_ (.B1(_0914_),
    .Y(_0916_),
    .A1(_0883_),
    .A2(_0885_));
 sg13g2_nor2b_2 _4687_ (.A(_0915_),
    .B_N(_0916_),
    .Y(_0917_));
 sg13g2_nor2b_1 _4688_ (.A(_0891_),
    .B_N(\generated._562[2] ),
    .Y(_0918_));
 sg13g2_or2_1 _4689_ (.X(_0919_),
    .B(_0918_),
    .A(_0893_));
 sg13g2_nand3_1 _4690_ (.B(_0856_),
    .C(_0890_),
    .A(_0828_),
    .Y(_0920_));
 sg13g2_nand2_1 _4691_ (.Y(_0921_),
    .A(net685),
    .B(_0920_));
 sg13g2_nor2_1 _4692_ (.A(net676),
    .B(_0853_),
    .Y(_0922_));
 sg13g2_nor2b_1 _4693_ (.A(net680),
    .B_N(_0062_),
    .Y(_0923_));
 sg13g2_a21oi_1 _4694_ (.A1(net682),
    .A2(_0065_),
    .Y(_0924_),
    .B1(_0923_));
 sg13g2_a21oi_1 _4695_ (.A1(net676),
    .A2(_0924_),
    .Y(_0925_),
    .B1(_0922_));
 sg13g2_xnor2_1 _4696_ (.Y(_0926_),
    .A(_0921_),
    .B(_0925_));
 sg13g2_xnor2_1 _4697_ (.Y(_0927_),
    .A(_2861_),
    .B(_0926_));
 sg13g2_nor2b_1 _4698_ (.A(_0927_),
    .B_N(_0919_),
    .Y(_0928_));
 sg13g2_nor2b_1 _4699_ (.A(_0919_),
    .B_N(_0927_),
    .Y(_0929_));
 sg13g2_nor3_1 _4700_ (.A(net637),
    .B(_0928_),
    .C(_0929_),
    .Y(_0930_));
 sg13g2_a21o_1 _4701_ (.A2(_0917_),
    .A1(net637),
    .B1(_0930_),
    .X(\generated._561[3] ));
 sg13g2_nor2b_1 _4702_ (.A(_0913_),
    .B_N(_0916_),
    .Y(_0931_));
 sg13g2_a21oi_2 _4703_ (.B1(_0908_),
    .Y(_0932_),
    .A2(_0906_),
    .A1(_0898_));
 sg13g2_nand2_1 _4704_ (.Y(_0933_),
    .A(net583),
    .B(_0836_));
 sg13g2_o21ai_1 _4705_ (.B1(_0905_),
    .Y(_0934_),
    .A1(_0871_),
    .A2(_0933_));
 sg13g2_nand2_1 _4706_ (.Y(_0935_),
    .A(net590),
    .B(net577));
 sg13g2_xor2_1 _4707_ (.B(net577),
    .A(net590),
    .X(_0936_));
 sg13g2_nor3_1 _4708_ (.A(_0837_),
    .B(net579),
    .C(net577),
    .Y(_0937_));
 sg13g2_nand2_1 _4709_ (.Y(_0938_),
    .A(net579),
    .B(net577));
 sg13g2_and2_1 _4710_ (.A(_0837_),
    .B(net577),
    .X(_0939_));
 sg13g2_o21ai_1 _4711_ (.B1(_0938_),
    .Y(_0940_),
    .A1(net579),
    .A2(_0939_));
 sg13g2_nor2b_1 _4712_ (.A(_0937_),
    .B_N(_0940_),
    .Y(_0941_));
 sg13g2_xor2_1 _4713_ (.B(_0941_),
    .A(_0936_),
    .X(_0942_));
 sg13g2_nand2_1 _4714_ (.Y(_0943_),
    .A(_0934_),
    .B(_0942_));
 sg13g2_xnor2_1 _4715_ (.Y(_0944_),
    .A(_0934_),
    .B(_0942_));
 sg13g2_xor2_1 _4716_ (.B(_0944_),
    .A(_0901_),
    .X(_0945_));
 sg13g2_nand2b_1 _4717_ (.Y(_0946_),
    .B(_0945_),
    .A_N(_0932_));
 sg13g2_xnor2_1 _4718_ (.Y(_0947_),
    .A(_0932_),
    .B(_0945_));
 sg13g2_nor2b_1 _4719_ (.A(_0911_),
    .B_N(_0947_),
    .Y(_0948_));
 sg13g2_xnor2_1 _4720_ (.Y(_0949_),
    .A(_0911_),
    .B(_0947_));
 sg13g2_nor2b_1 _4721_ (.A(_0931_),
    .B_N(_0949_),
    .Y(_0950_));
 sg13g2_xnor2_1 _4722_ (.Y(_0951_),
    .A(_0931_),
    .B(_0949_));
 sg13g2_a21oi_1 _4723_ (.A1(_2861_),
    .A2(_0926_),
    .Y(_0952_),
    .B1(_0928_));
 sg13g2_nand2b_1 _4724_ (.Y(_0953_),
    .B(_0925_),
    .A_N(_0920_));
 sg13g2_nand2_1 _4725_ (.Y(_0954_),
    .A(net685),
    .B(_0953_));
 sg13g2_nor2_1 _4726_ (.A(net676),
    .B(_0889_),
    .Y(_0955_));
 sg13g2_nor2b_1 _4727_ (.A(net681),
    .B_N(_0065_),
    .Y(_0956_));
 sg13g2_a21oi_1 _4728_ (.A1(net681),
    .A2(_0067_),
    .Y(_0957_),
    .B1(_0956_));
 sg13g2_a21oi_1 _4729_ (.A1(net675),
    .A2(_0957_),
    .Y(_0958_),
    .B1(_0955_));
 sg13g2_xnor2_1 _4730_ (.Y(_0959_),
    .A(_0954_),
    .B(_0958_));
 sg13g2_xor2_1 _4731_ (.B(_0959_),
    .A(_0066_),
    .X(_0960_));
 sg13g2_or2_1 _4732_ (.X(_0961_),
    .B(_0960_),
    .A(_0952_));
 sg13g2_a21oi_1 _4733_ (.A1(_0952_),
    .A2(_0960_),
    .Y(_0962_),
    .B1(net636));
 sg13g2_a22oi_1 _4734_ (.Y(_0963_),
    .B1(_0961_),
    .B2(_0962_),
    .A2(_0951_),
    .A1(net636));
 sg13g2_inv_1 _4735_ (.Y(\generated._561[4] ),
    .A(_0963_));
 sg13g2_nor2_1 _4736_ (.A(_0948_),
    .B(_0950_),
    .Y(_0964_));
 sg13g2_o21ai_1 _4737_ (.B1(_0943_),
    .Y(_0965_),
    .A1(_0901_),
    .A2(_0944_));
 sg13g2_a21oi_1 _4738_ (.A1(_0936_),
    .A2(_0940_),
    .Y(_0966_),
    .B1(_0937_));
 sg13g2_xor2_1 _4739_ (.B(_0938_),
    .A(net583),
    .X(_0967_));
 sg13g2_xor2_1 _4740_ (.B(_0967_),
    .A(_0966_),
    .X(_0968_));
 sg13g2_nand2b_1 _4741_ (.Y(_0969_),
    .B(_0968_),
    .A_N(_0935_));
 sg13g2_xnor2_1 _4742_ (.Y(_0970_),
    .A(_0935_),
    .B(_0968_));
 sg13g2_nand2_1 _4743_ (.Y(_0971_),
    .A(_0965_),
    .B(_0970_));
 sg13g2_xnor2_1 _4744_ (.Y(_0972_),
    .A(_0965_),
    .B(_0970_));
 sg13g2_nor2_1 _4745_ (.A(_0946_),
    .B(_0972_),
    .Y(_0973_));
 sg13g2_xor2_1 _4746_ (.B(_0972_),
    .A(_0946_),
    .X(_0974_));
 sg13g2_nor3_1 _4747_ (.A(_0948_),
    .B(_0950_),
    .C(_0974_),
    .Y(_0975_));
 sg13g2_nor2b_1 _4748_ (.A(_0964_),
    .B_N(_0974_),
    .Y(_0976_));
 sg13g2_nor3_1 _4749_ (.A(net632),
    .B(_0975_),
    .C(_0976_),
    .Y(_0977_));
 sg13g2_nand2_1 _4750_ (.Y(_0978_),
    .A(\generated._562[4] ),
    .B(_0959_));
 sg13g2_nor2b_1 _4751_ (.A(_0953_),
    .B_N(_0958_),
    .Y(_0979_));
 sg13g2_nor2_1 _4752_ (.A(net656),
    .B(_0979_),
    .Y(_0980_));
 sg13g2_mux2_1 _4753_ (.A0(_0067_),
    .A1(_0069_),
    .S(net681),
    .X(_0981_));
 sg13g2_nand2_1 _4754_ (.Y(_0982_),
    .A(net675),
    .B(_0981_));
 sg13g2_o21ai_1 _4755_ (.B1(_0982_),
    .Y(_0983_),
    .A1(net675),
    .A2(_0924_));
 sg13g2_xor2_1 _4756_ (.B(_0983_),
    .A(_0980_),
    .X(_0984_));
 sg13g2_nand2b_1 _4757_ (.Y(_0985_),
    .B(_0984_),
    .A_N(_0068_));
 sg13g2_xor2_1 _4758_ (.B(_0984_),
    .A(_0068_),
    .X(_0986_));
 sg13g2_a21o_1 _4759_ (.A2(_0978_),
    .A1(_0961_),
    .B1(_0986_),
    .X(_0987_));
 sg13g2_nand3_1 _4760_ (.B(_0978_),
    .C(_0986_),
    .A(_0961_),
    .Y(_0988_));
 sg13g2_nand3_1 _4761_ (.B(_0987_),
    .C(_0988_),
    .A(net632),
    .Y(_0989_));
 sg13g2_nand2b_1 _4762_ (.Y(\generated._561[5] ),
    .B(_0989_),
    .A_N(_0977_));
 sg13g2_o21ai_1 _4763_ (.B1(_0969_),
    .Y(_0990_),
    .A1(_0966_),
    .A2(_0967_));
 sg13g2_o21ai_1 _4764_ (.B1(net577),
    .Y(_0991_),
    .A1(net583),
    .A2(_0871_));
 sg13g2_xnor2_1 _4765_ (.Y(_0992_),
    .A(_0836_),
    .B(_0991_));
 sg13g2_nand2_1 _4766_ (.Y(_0993_),
    .A(_0990_),
    .B(_0992_));
 sg13g2_xor2_1 _4767_ (.B(_0992_),
    .A(_0990_),
    .X(_0994_));
 sg13g2_inv_1 _4768_ (.Y(_0995_),
    .A(_0994_));
 sg13g2_xnor2_1 _4769_ (.Y(_0996_),
    .A(_0971_),
    .B(_0994_));
 sg13g2_o21ai_1 _4770_ (.B1(_0996_),
    .Y(_0997_),
    .A1(_0973_),
    .A2(_0976_));
 sg13g2_or3_1 _4771_ (.A(_0973_),
    .B(_0976_),
    .C(_0996_),
    .X(_0998_));
 sg13g2_nand3_1 _4772_ (.B(_0997_),
    .C(_0998_),
    .A(net636),
    .Y(_0999_));
 sg13g2_a21oi_1 _4773_ (.A1(_0979_),
    .A2(_0983_),
    .Y(_1000_),
    .B1(net656));
 sg13g2_mux2_1 _4774_ (.A0(_0069_),
    .A1(_0071_),
    .S(net681),
    .X(_1001_));
 sg13g2_nand2_1 _4775_ (.Y(_1002_),
    .A(net678),
    .B(_1001_));
 sg13g2_o21ai_1 _4776_ (.B1(_1002_),
    .Y(_1003_),
    .A1(net675),
    .A2(_0957_));
 sg13g2_xor2_1 _4777_ (.B(_1003_),
    .A(_1000_),
    .X(_1004_));
 sg13g2_xor2_1 _4778_ (.B(_1004_),
    .A(_0070_),
    .X(_1005_));
 sg13g2_nand3_1 _4779_ (.B(_0987_),
    .C(_1005_),
    .A(_0985_),
    .Y(_1006_));
 sg13g2_a21oi_1 _4780_ (.A1(_0985_),
    .A2(_0987_),
    .Y(_1007_),
    .B1(_1005_));
 sg13g2_nand2_1 _4781_ (.Y(_1008_),
    .A(net632),
    .B(_1006_));
 sg13g2_o21ai_1 _4782_ (.B1(_0999_),
    .Y(\generated._561[6] ),
    .A1(_1007_),
    .A2(_1008_));
 sg13g2_o21ai_1 _4783_ (.B1(_0997_),
    .Y(_1009_),
    .A1(_0971_),
    .A2(_0995_));
 sg13g2_o21ai_1 _4784_ (.B1(_0940_),
    .Y(_1010_),
    .A1(_0871_),
    .A2(_0933_));
 sg13g2_nor2_1 _4785_ (.A(_0993_),
    .B(_1010_),
    .Y(_1011_));
 sg13g2_xor2_1 _4786_ (.B(_1010_),
    .A(_0993_),
    .X(_1012_));
 sg13g2_a21oi_1 _4787_ (.A1(_1009_),
    .A2(_1012_),
    .Y(_1013_),
    .B1(net632));
 sg13g2_o21ai_1 _4788_ (.B1(_1013_),
    .Y(_1014_),
    .A1(_1009_),
    .A2(_1012_));
 sg13g2_a21oi_1 _4789_ (.A1(\generated._562[6] ),
    .A2(_1004_),
    .Y(_1015_),
    .B1(_1007_));
 sg13g2_nor2b_1 _4790_ (.A(net673),
    .B_N(_0981_),
    .Y(_1016_));
 sg13g2_a21oi_2 _4791_ (.B1(_1016_),
    .Y(_1017_),
    .A2(_0071_),
    .A1(net674));
 sg13g2_nand3_1 _4792_ (.B(_0983_),
    .C(_1003_),
    .A(_0979_),
    .Y(_1018_));
 sg13g2_nand2_1 _4793_ (.Y(_1019_),
    .A(net684),
    .B(_1018_));
 sg13g2_xor2_1 _4794_ (.B(_1019_),
    .A(_1017_),
    .X(_1020_));
 sg13g2_xnor2_1 _4795_ (.Y(_1021_),
    .A(_0072_),
    .B(_1020_));
 sg13g2_nor2b_1 _4796_ (.A(_1015_),
    .B_N(_1021_),
    .Y(_1022_));
 sg13g2_xor2_1 _4797_ (.B(_1021_),
    .A(_1015_),
    .X(_1023_));
 sg13g2_o21ai_1 _4798_ (.B1(_1014_),
    .Y(\generated._561[7] ),
    .A1(net636),
    .A2(_1023_));
 sg13g2_a21oi_1 _4799_ (.A1(\generated._562[7] ),
    .A2(_1020_),
    .Y(_1024_),
    .B1(_1022_));
 sg13g2_nor2b_1 _4800_ (.A(net674),
    .B_N(_1001_),
    .Y(_1025_));
 sg13g2_a21oi_1 _4801_ (.A1(net674),
    .A2(_0071_),
    .Y(_1026_),
    .B1(_1025_));
 sg13g2_o21ai_1 _4802_ (.B1(net684),
    .Y(_1027_),
    .A1(_1017_),
    .A2(_1018_));
 sg13g2_xor2_1 _4803_ (.B(_1027_),
    .A(_1026_),
    .X(_1028_));
 sg13g2_xnor2_1 _4804_ (.Y(_1029_),
    .A(_2862_),
    .B(_1028_));
 sg13g2_nor2_1 _4805_ (.A(_1024_),
    .B(_1029_),
    .Y(_1030_));
 sg13g2_xnor2_1 _4806_ (.Y(_1031_),
    .A(_1024_),
    .B(_1029_));
 sg13g2_nand2_1 _4807_ (.Y(_1032_),
    .A(net579),
    .B(_0933_));
 sg13g2_a21oi_2 _4808_ (.B1(_1011_),
    .Y(_1033_),
    .A2(_1032_),
    .A1(_0900_));
 sg13g2_a22oi_1 _4809_ (.Y(\generated._561[8] ),
    .B1(_1033_),
    .B2(_1013_),
    .A2(_1031_),
    .A1(net632));
 sg13g2_a21oi_1 _4810_ (.A1(net562),
    .A2(_1028_),
    .Y(_1034_),
    .B1(_1030_));
 sg13g2_nor3_1 _4811_ (.A(_1017_),
    .B(_1018_),
    .C(_1026_),
    .Y(_1035_));
 sg13g2_xnor2_1 _4812_ (.Y(_1036_),
    .A(\generated._511 ),
    .B(_1035_));
 sg13g2_nor2_1 _4813_ (.A(net656),
    .B(_1036_),
    .Y(_1037_));
 sg13g2_a21oi_1 _4814_ (.A1(net656),
    .A2(_0071_),
    .Y(_1038_),
    .B1(_1037_));
 sg13g2_xnor2_1 _4815_ (.Y(_1039_),
    .A(_0074_),
    .B(_1038_));
 sg13g2_o21ai_1 _4816_ (.B1(net632),
    .Y(_1040_),
    .A1(_1034_),
    .A2(_1039_));
 sg13g2_a21oi_1 _4817_ (.A1(_1034_),
    .A2(_1039_),
    .Y(_1041_),
    .B1(_1040_));
 sg13g2_a21o_1 _4818_ (.A2(_0900_),
    .A1(net636),
    .B1(_1041_),
    .X(\generated._561[9] ));
 sg13g2_nor3_2 _4819_ (.A(\generated._487[1] ),
    .B(\generated._487[0] ),
    .C(\generated._487[3] ),
    .Y(_1042_));
 sg13g2_nor2b_1 _4820_ (.A(\generated._487[2] ),
    .B_N(_1042_),
    .Y(_1043_));
 sg13g2_nand2b_2 _4821_ (.Y(_1044_),
    .B(_1042_),
    .A_N(\generated._487[2] ));
 sg13g2_nor2_1 _4822_ (.A(net296),
    .B(_1044_),
    .Y(_1045_));
 sg13g2_nand2_2 _4823_ (.Y(_1046_),
    .A(net667),
    .B(net664));
 sg13g2_inv_1 _4824_ (.Y(_1047_),
    .A(_1046_));
 sg13g2_xor2_1 _4825_ (.B(_1046_),
    .A(_0076_),
    .X(_1048_));
 sg13g2_a21oi_1 _4826_ (.A1(_1044_),
    .A2(_1048_),
    .Y(\generated._481[0] ),
    .B1(net297));
 sg13g2_nor2b_1 _4827_ (.A(net717),
    .B_N(\generated._1084[1] ),
    .Y(_1049_));
 sg13g2_nand2b_1 _4828_ (.Y(_1050_),
    .B(net717),
    .A_N(\generated._1084[1] ));
 sg13g2_nand2b_1 _4829_ (.Y(_1051_),
    .B(_1050_),
    .A_N(_1049_));
 sg13g2_o21ai_1 _4830_ (.B1(net629),
    .Y(_1052_),
    .A1(net296),
    .A2(_1051_));
 sg13g2_a21o_1 _4831_ (.A2(_1051_),
    .A1(net296),
    .B1(_1052_),
    .X(_1053_));
 sg13g2_nor2_1 _4832_ (.A(_2840_),
    .B(net671),
    .Y(_1054_));
 sg13g2_xor2_1 _4833_ (.B(net671),
    .A(net664),
    .X(_1055_));
 sg13g2_a21oi_2 _4834_ (.B1(_1054_),
    .Y(_1056_),
    .A2(_1055_),
    .A1(_2840_));
 sg13g2_nor2_2 _4835_ (.A(_1047_),
    .B(_1056_),
    .Y(_1057_));
 sg13g2_nor2_1 _4836_ (.A(_0077_),
    .B(_1057_),
    .Y(_1058_));
 sg13g2_xnor2_1 _4837_ (.Y(_1059_),
    .A(_0077_),
    .B(_1057_));
 sg13g2_a21oi_1 _4838_ (.A1(net398),
    .A2(_1046_),
    .Y(_1060_),
    .B1(_1059_));
 sg13g2_nand3_1 _4839_ (.B(_1046_),
    .C(_1059_),
    .A(net398),
    .Y(_1061_));
 sg13g2_nand2_1 _4840_ (.Y(_1062_),
    .A(_1044_),
    .B(_1061_));
 sg13g2_o21ai_1 _4841_ (.B1(_1053_),
    .Y(\generated._481[1] ),
    .A1(_1060_),
    .A2(_1062_));
 sg13g2_nand2b_1 _4842_ (.Y(_1063_),
    .B(net422),
    .A_N(net717));
 sg13g2_xor2_1 _4843_ (.B(\generated._1084[2] ),
    .A(net717),
    .X(_1064_));
 sg13g2_o21ai_1 _4844_ (.B1(_1050_),
    .Y(_1065_),
    .A1(net335),
    .A2(_1049_));
 sg13g2_or2_1 _4845_ (.X(_1066_),
    .B(_1065_),
    .A(_1064_));
 sg13g2_xnor2_1 _4846_ (.Y(_1067_),
    .A(_1064_),
    .B(_1065_));
 sg13g2_nor2_2 _4847_ (.A(_2840_),
    .B(net664),
    .Y(_1068_));
 sg13g2_nor2_1 _4848_ (.A(_2864_),
    .B(_1068_),
    .Y(_1069_));
 sg13g2_or2_1 _4849_ (.X(_1070_),
    .B(_1069_),
    .A(_1054_));
 sg13g2_nand2_1 _4850_ (.Y(_1071_),
    .A(\generated._373[2] ),
    .B(_1070_));
 sg13g2_xor2_1 _4851_ (.B(_1070_),
    .A(\generated._373[2] ),
    .X(_1072_));
 sg13g2_o21ai_1 _4852_ (.B1(_1072_),
    .Y(_1073_),
    .A1(_1058_),
    .A2(_1060_));
 sg13g2_or3_1 _4853_ (.A(_1058_),
    .B(_1060_),
    .C(_1072_),
    .X(_1074_));
 sg13g2_nand3_1 _4854_ (.B(_1073_),
    .C(_1074_),
    .A(net627),
    .Y(_1075_));
 sg13g2_o21ai_1 _4855_ (.B1(_1075_),
    .Y(\generated._481[2] ),
    .A1(net627),
    .A2(_1067_));
 sg13g2_xnor2_1 _4856_ (.Y(_1076_),
    .A(net717),
    .B(\generated._1084[3] ));
 sg13g2_nand3_1 _4857_ (.B(_1066_),
    .C(_1076_),
    .A(_1063_),
    .Y(_1077_));
 sg13g2_a21oi_1 _4858_ (.A1(_1063_),
    .A2(_1066_),
    .Y(_1078_),
    .B1(_1076_));
 sg13g2_nand2_1 _4859_ (.Y(_1079_),
    .A(net629),
    .B(_1077_));
 sg13g2_and2_1 _4860_ (.A(_1071_),
    .B(_1073_),
    .X(_1080_));
 sg13g2_nor2_1 _4861_ (.A(net468),
    .B(_1057_),
    .Y(_1081_));
 sg13g2_xnor2_1 _4862_ (.Y(_1082_),
    .A(net468),
    .B(_1057_));
 sg13g2_nor2_1 _4863_ (.A(_1080_),
    .B(_1082_),
    .Y(_1083_));
 sg13g2_a21oi_1 _4864_ (.A1(_1080_),
    .A2(_1082_),
    .Y(_1084_),
    .B1(net629));
 sg13g2_nand2b_1 _4865_ (.Y(_1085_),
    .B(_1084_),
    .A_N(_1083_));
 sg13g2_o21ai_1 _4866_ (.B1(_1085_),
    .Y(\generated._481[3] ),
    .A1(_1078_),
    .A2(_1079_));
 sg13g2_a21oi_1 _4867_ (.A1(net717),
    .A2(\generated._1084[3] ),
    .Y(_1086_),
    .B1(_1078_));
 sg13g2_xor2_1 _4868_ (.B(net544),
    .A(net717),
    .X(_1087_));
 sg13g2_or2_1 _4869_ (.X(_1088_),
    .B(_1087_),
    .A(_1086_));
 sg13g2_a21oi_1 _4870_ (.A1(_1086_),
    .A2(_1087_),
    .Y(_1089_),
    .B1(net627));
 sg13g2_nor2_1 _4871_ (.A(_1081_),
    .B(_1083_),
    .Y(_1090_));
 sg13g2_nand3_1 _4872_ (.B(_1046_),
    .C(_1056_),
    .A(net560),
    .Y(_1091_));
 sg13g2_a21o_1 _4873_ (.A2(_1056_),
    .A1(_1046_),
    .B1(net753),
    .X(_1092_));
 sg13g2_nand2_1 _4874_ (.Y(_1093_),
    .A(_1091_),
    .B(_1092_));
 sg13g2_or2_1 _4875_ (.X(_1094_),
    .B(_1093_),
    .A(_1090_));
 sg13g2_a21oi_1 _4876_ (.A1(_1090_),
    .A2(_1093_),
    .Y(_1095_),
    .B1(net629));
 sg13g2_a22oi_1 _4877_ (.Y(_1096_),
    .B1(_1094_),
    .B2(_1095_),
    .A2(_1089_),
    .A1(_1088_));
 sg13g2_inv_1 _4878_ (.Y(\generated._481[4] ),
    .A(_1096_));
 sg13g2_nand2_1 _4879_ (.Y(_1097_),
    .A(_1091_),
    .B(_1094_));
 sg13g2_nor2_1 _4880_ (.A(\generated._373[5] ),
    .B(_1055_),
    .Y(_1098_));
 sg13g2_and2_1 _4881_ (.A(\generated._373[5] ),
    .B(_1055_),
    .X(_1099_));
 sg13g2_nor2_1 _4882_ (.A(_1098_),
    .B(_1099_),
    .Y(_1100_));
 sg13g2_o21ai_1 _4883_ (.B1(_1088_),
    .Y(_1101_),
    .A1(net717),
    .A2(_2867_));
 sg13g2_nor2b_1 _4884_ (.A(net718),
    .B_N(\generated._1084[5] ),
    .Y(_1102_));
 sg13g2_nand2b_1 _4885_ (.Y(_1103_),
    .B(net718),
    .A_N(\generated._1084[5] ));
 sg13g2_nand2b_1 _4886_ (.Y(_1104_),
    .B(_1103_),
    .A_N(_1102_));
 sg13g2_xnor2_1 _4887_ (.Y(_1105_),
    .A(_1101_),
    .B(_1104_));
 sg13g2_nand2_1 _4888_ (.Y(_1106_),
    .A(net629),
    .B(_1105_));
 sg13g2_xnor2_1 _4889_ (.Y(_1107_),
    .A(_1097_),
    .B(_1100_));
 sg13g2_o21ai_1 _4890_ (.B1(_1106_),
    .Y(\generated._481[5] ),
    .A1(net629),
    .A2(_1107_));
 sg13g2_xor2_1 _4891_ (.B(\generated._1084[6] ),
    .A(net718),
    .X(_1108_));
 sg13g2_o21ai_1 _4892_ (.B1(_1103_),
    .Y(_1109_),
    .A1(_1101_),
    .A2(_1102_));
 sg13g2_inv_1 _4893_ (.Y(_1110_),
    .A(_1109_));
 sg13g2_nor2b_1 _4894_ (.A(_1109_),
    .B_N(_1108_),
    .Y(_1111_));
 sg13g2_o21ai_1 _4895_ (.B1(net629),
    .Y(_1112_),
    .A1(_1108_),
    .A2(_1110_));
 sg13g2_nand2b_1 _4896_ (.Y(_1113_),
    .B(\generated._373[6] ),
    .A_N(_1056_));
 sg13g2_xnor2_1 _4897_ (.Y(_1114_),
    .A(\generated._373[6] ),
    .B(_1056_));
 sg13g2_a21oi_1 _4898_ (.A1(_1091_),
    .A2(_1094_),
    .Y(_1115_),
    .B1(_1098_));
 sg13g2_o21ai_1 _4899_ (.B1(_1114_),
    .Y(_1116_),
    .A1(_1099_),
    .A2(_1115_));
 sg13g2_or3_1 _4900_ (.A(_1099_),
    .B(_1114_),
    .C(_1115_),
    .X(_1117_));
 sg13g2_nand3_1 _4901_ (.B(_1116_),
    .C(_1117_),
    .A(net627),
    .Y(_1118_));
 sg13g2_o21ai_1 _4902_ (.B1(_1118_),
    .Y(\generated._481[6] ),
    .A1(_1111_),
    .A2(_1112_));
 sg13g2_xnor2_1 _4903_ (.Y(_1119_),
    .A(net718),
    .B(\generated._1084[7] ));
 sg13g2_a21oi_1 _4904_ (.A1(net718),
    .A2(\generated._1084[6] ),
    .Y(_1120_),
    .B1(_1111_));
 sg13g2_xnor2_1 _4905_ (.Y(_1121_),
    .A(net671),
    .B(net496));
 sg13g2_nand3_1 _4906_ (.B(_1116_),
    .C(_1121_),
    .A(_1113_),
    .Y(_1122_));
 sg13g2_a21oi_1 _4907_ (.A1(_1113_),
    .A2(_1116_),
    .Y(_1123_),
    .B1(_1121_));
 sg13g2_nor2_1 _4908_ (.A(net630),
    .B(_1123_),
    .Y(_1124_));
 sg13g2_xnor2_1 _4909_ (.Y(_1125_),
    .A(_1119_),
    .B(_1120_));
 sg13g2_a22oi_1 _4910_ (.Y(\generated._481[7] ),
    .B1(_1125_),
    .B2(net629),
    .A2(_1124_),
    .A1(net497));
 sg13g2_xnor2_1 _4911_ (.Y(_1126_),
    .A(net415),
    .B(net671));
 sg13g2_a22oi_1 _4912_ (.Y(_1127_),
    .B1(_1113_),
    .B2(_1116_),
    .A2(_2865_),
    .A1(net671));
 sg13g2_a21o_1 _4913_ (.A2(net529),
    .A1(_2864_),
    .B1(_1127_),
    .X(_1128_));
 sg13g2_a21oi_1 _4914_ (.A1(_1126_),
    .A2(_1128_),
    .Y(_1129_),
    .B1(net630));
 sg13g2_o21ai_1 _4915_ (.B1(_1129_),
    .Y(_1130_),
    .A1(_1126_),
    .A2(_1128_));
 sg13g2_o21ai_1 _4916_ (.B1(net718),
    .Y(_1131_),
    .A1(\generated._1084[6] ),
    .A2(\generated._1084[7] ));
 sg13g2_o21ai_1 _4917_ (.B1(_1111_),
    .Y(_1132_),
    .A1(net718),
    .A2(\generated._1084[7] ));
 sg13g2_and2_1 _4918_ (.A(_1131_),
    .B(_1132_),
    .X(_1133_));
 sg13g2_nor2b_1 _4919_ (.A(net719),
    .B_N(\generated._1084[8] ),
    .Y(_1134_));
 sg13g2_xor2_1 _4920_ (.B(\generated._1084[8] ),
    .A(net719),
    .X(_1135_));
 sg13g2_and2_1 _4921_ (.A(_1133_),
    .B(_1135_),
    .X(_1136_));
 sg13g2_o21ai_1 _4922_ (.B1(net630),
    .Y(_1137_),
    .A1(_1133_),
    .A2(_1135_));
 sg13g2_o21ai_1 _4923_ (.B1(_1130_),
    .Y(\generated._481[8] ),
    .A1(_1136_),
    .A2(_1137_));
 sg13g2_o21ai_1 _4924_ (.B1(_1129_),
    .Y(_1138_),
    .A1(_2863_),
    .A2(net671));
 sg13g2_o21ai_1 _4925_ (.B1(net416),
    .Y(\generated._481[9] ),
    .A1(_1134_),
    .A2(_1137_));
 sg13g2_nor2b_1 _4926_ (.A(_2910_),
    .B_N(_0249_),
    .Y(_0116_));
 sg13g2_nor2b_1 _4927_ (.A(_2912_),
    .B_N(_0249_),
    .Y(_0117_));
 sg13g2_nor3_1 _4928_ (.A(net385),
    .B(_2917_),
    .C(_2918_),
    .Y(_0118_));
 sg13g2_nand2_1 _4929_ (.Y(_1139_),
    .A(net722),
    .B(net720));
 sg13g2_nor2_1 _4930_ (.A(net721),
    .B(_1139_),
    .Y(_1140_));
 sg13g2_and3_1 _4931_ (.X(_1141_),
    .A(net723),
    .B(\generated._100[5] ),
    .C(\generated._100[6] ));
 sg13g2_nor4_2 _4932_ (.A(net721),
    .B(_2880_),
    .C(_1139_),
    .Y(_1142_),
    .D(_1141_));
 sg13g2_nor2_1 _4933_ (.A(net742),
    .B(_1142_),
    .Y(_0279_));
 sg13g2_nand2_1 _4934_ (.Y(_1143_),
    .A(net728),
    .B(_0456_));
 sg13g2_nand4_1 _4935_ (.B(net727),
    .C(net730),
    .A(_2835_),
    .Y(_1144_),
    .D(net379));
 sg13g2_nor4_1 _4936_ (.A(net729),
    .B(net350),
    .C(_0457_),
    .D(_1144_),
    .Y(_1145_));
 sg13g2_nor2_1 _4937_ (.A(net741),
    .B(_1145_),
    .Y(_0280_));
 sg13g2_a21oi_1 _4938_ (.A1(_1142_),
    .A2(_1145_),
    .Y(_0119_),
    .B1(net741));
 sg13g2_o21ai_1 _4939_ (.B1(net720),
    .Y(_1146_),
    .A1(net722),
    .A2(net721));
 sg13g2_nand4_1 _4940_ (.B(net748),
    .C(_1143_),
    .A(_2835_),
    .Y(_1147_),
    .D(_1146_));
 sg13g2_nor4_1 _4941_ (.A(\generated._221[1] ),
    .B(\generated._221[0] ),
    .C(net727),
    .D(net729),
    .Y(_1148_));
 sg13g2_nand3b_1 _4942_ (.B(_0325_),
    .C(_1148_),
    .Y(_1149_),
    .A_N(net730));
 sg13g2_a21oi_1 _4943_ (.A1(_0399_),
    .A2(_0456_),
    .Y(_1150_),
    .B1(\generated._221[3] ));
 sg13g2_nand2_2 _4944_ (.Y(_1151_),
    .A(_1149_),
    .B(_1150_));
 sg13g2_nand3_1 _4945_ (.B(net720),
    .C(_1141_),
    .A(\generated._100[3] ),
    .Y(_1152_));
 sg13g2_nand3_1 _4946_ (.B(_1146_),
    .C(_1152_),
    .A(_2882_),
    .Y(_1153_));
 sg13g2_nor2_1 _4947_ (.A(_1151_),
    .B(_1153_),
    .Y(_1154_));
 sg13g2_mux2_1 _4948_ (.A0(net726),
    .A1(\generated._1148[0] ),
    .S(_1151_),
    .X(_1155_));
 sg13g2_nand2b_1 _4949_ (.Y(_1156_),
    .B(_1155_),
    .A_N(_1154_));
 sg13g2_and2_1 _4950_ (.A(net744),
    .B(_1156_),
    .X(_1157_));
 sg13g2_nand2b_2 _4951_ (.Y(_1158_),
    .B(_0325_),
    .A_N(_0323_));
 sg13g2_nor2_1 _4952_ (.A(\generated._28[3] ),
    .B(\generated._28[1] ),
    .Y(_1159_));
 sg13g2_o21ai_1 _4953_ (.B1(_1154_),
    .Y(_1160_),
    .A1(_1158_),
    .A2(_1159_));
 sg13g2_nand2b_2 _4954_ (.Y(_1161_),
    .B(_1158_),
    .A_N(\generated._346[5] ));
 sg13g2_nor2_1 _4955_ (.A(net557),
    .B(_1161_),
    .Y(_1162_));
 sg13g2_o21ai_1 _4956_ (.B1(_1157_),
    .Y(_1163_),
    .A1(_1160_),
    .A2(_1162_));
 sg13g2_nand2_2 _4957_ (.Y(_1164_),
    .A(net687),
    .B(\generated._1087[0] ));
 sg13g2_or2_1 _4958_ (.X(_1165_),
    .B(\generated._1087[0] ),
    .A(net687));
 sg13g2_nand3_1 _4959_ (.B(_1164_),
    .C(_1165_),
    .A(\generated._65[4] ),
    .Y(_1166_));
 sg13g2_a21o_1 _4960_ (.A2(_1165_),
    .A1(_1164_),
    .B1(\generated._65[4] ),
    .X(_1167_));
 sg13g2_nand2_2 _4961_ (.Y(_1168_),
    .A(_1166_),
    .B(_1167_));
 sg13g2_nand2_1 _4962_ (.Y(_1169_),
    .A(\generated._65[3] ),
    .B(\generated._65[2] ));
 sg13g2_nor2_1 _4963_ (.A(\generated._1087[0] ),
    .B(\generated._165[4] ),
    .Y(_1170_));
 sg13g2_xor2_1 _4964_ (.B(\generated._165[4] ),
    .A(\generated._1087[0] ),
    .X(_1171_));
 sg13g2_xnor2_1 _4965_ (.Y(_1172_),
    .A(\generated._65[4] ),
    .B(_1171_));
 sg13g2_nor2_1 _4966_ (.A(_1164_),
    .B(_1172_),
    .Y(_1173_));
 sg13g2_xor2_1 _4967_ (.B(_1172_),
    .A(_1164_),
    .X(_1174_));
 sg13g2_xnor2_1 _4968_ (.Y(_1175_),
    .A(\generated._65[5] ),
    .B(_1174_));
 sg13g2_nor2_1 _4969_ (.A(_1166_),
    .B(_1175_),
    .Y(_1176_));
 sg13g2_xnor2_1 _4970_ (.Y(_1177_),
    .A(_1166_),
    .B(_1175_));
 sg13g2_nor3_1 _4971_ (.A(_1168_),
    .B(_1169_),
    .C(_1177_),
    .Y(_1178_));
 sg13g2_o21ai_1 _4972_ (.B1(_1177_),
    .Y(_1179_),
    .A1(_1168_),
    .A2(_1169_));
 sg13g2_nor2b_1 _4973_ (.A(_1178_),
    .B_N(_1179_),
    .Y(_1180_));
 sg13g2_inv_1 _4974_ (.Y(_1181_),
    .A(_1180_));
 sg13g2_nand2_1 _4975_ (.Y(_1182_),
    .A(\generated._65[2] ),
    .B(\generated._165[4] ));
 sg13g2_nor3_1 _4976_ (.A(net687),
    .B(_1168_),
    .C(_1182_),
    .Y(_1183_));
 sg13g2_nand2_1 _4977_ (.Y(_1184_),
    .A(\generated._1087[0] ),
    .B(\generated._65[2] ));
 sg13g2_nor2_1 _4978_ (.A(_1165_),
    .B(_1182_),
    .Y(_1185_));
 sg13g2_nor2_1 _4979_ (.A(net687),
    .B(\generated._165[4] ),
    .Y(_1186_));
 sg13g2_or2_1 _4980_ (.X(_1187_),
    .B(\generated._165[4] ),
    .A(net687));
 sg13g2_nor2_1 _4981_ (.A(\generated._65[2] ),
    .B(_1187_),
    .Y(_1188_));
 sg13g2_nor2_1 _4982_ (.A(_1185_),
    .B(_1188_),
    .Y(_1189_));
 sg13g2_nor2_1 _4983_ (.A(_2868_),
    .B(_1186_),
    .Y(_1190_));
 sg13g2_xor2_1 _4984_ (.B(_1190_),
    .A(_1168_),
    .X(_1191_));
 sg13g2_nor3_1 _4985_ (.A(_1185_),
    .B(_1188_),
    .C(_1191_),
    .Y(_1192_));
 sg13g2_nor2_1 _4986_ (.A(_1183_),
    .B(_1192_),
    .Y(_1193_));
 sg13g2_xnor2_1 _4987_ (.Y(_1194_),
    .A(_1180_),
    .B(_1193_));
 sg13g2_o21ai_1 _4988_ (.B1(_1163_),
    .Y(_1195_),
    .A1(net1),
    .A2(_1194_));
 sg13g2_nor2_1 _4989_ (.A(_0007_),
    .B(_1161_),
    .Y(_1196_));
 sg13g2_o21ai_1 _4990_ (.B1(_1157_),
    .Y(_1197_),
    .A1(_1160_),
    .A2(_1196_));
 sg13g2_xnor2_1 _4991_ (.Y(_1198_),
    .A(_1189_),
    .B(_1191_));
 sg13g2_o21ai_1 _4992_ (.B1(_1197_),
    .Y(_1199_),
    .A1(net1),
    .A2(_1198_));
 sg13g2_nor2_1 _4993_ (.A(_0009_),
    .B(_1161_),
    .Y(_1200_));
 sg13g2_o21ai_1 _4994_ (.B1(_1157_),
    .Y(_1201_),
    .A1(_1160_),
    .A2(_1200_));
 sg13g2_nand4_1 _4995_ (.B(\generated._1087[0] ),
    .C(_2868_),
    .A(net687),
    .Y(_1202_),
    .D(\generated._165[4] ));
 sg13g2_nor3_1 _4996_ (.A(_1181_),
    .B(_1191_),
    .C(_1202_),
    .Y(_1203_));
 sg13g2_nor4_1 _4997_ (.A(net687),
    .B(_1168_),
    .C(_1177_),
    .D(_1182_),
    .Y(_1204_));
 sg13g2_nor3_1 _4998_ (.A(_1178_),
    .B(_1203_),
    .C(_1204_),
    .Y(_1205_));
 sg13g2_nand3_1 _4999_ (.B(_1192_),
    .C(_1202_),
    .A(_1180_),
    .Y(_1206_));
 sg13g2_a21oi_1 _5000_ (.A1(\generated._65[5] ),
    .A2(_1174_),
    .Y(_1207_),
    .B1(_1173_));
 sg13g2_a21oi_1 _5001_ (.A1(\generated._65[4] ),
    .A2(_1171_),
    .Y(_1208_),
    .B1(_1170_));
 sg13g2_xnor2_1 _5002_ (.Y(_1209_),
    .A(\generated._65[5] ),
    .B(\generated._65[6] ));
 sg13g2_xnor2_1 _5003_ (.Y(_1210_),
    .A(\generated._65[2] ),
    .B(_1209_));
 sg13g2_xnor2_1 _5004_ (.Y(_1211_),
    .A(_1208_),
    .B(_1210_));
 sg13g2_xnor2_1 _5005_ (.Y(_1212_),
    .A(_1207_),
    .B(_1211_));
 sg13g2_xnor2_1 _5006_ (.Y(_1213_),
    .A(_1176_),
    .B(_1212_));
 sg13g2_xnor2_1 _5007_ (.Y(_1214_),
    .A(_1206_),
    .B(_1213_));
 sg13g2_xnor2_1 _5008_ (.Y(_1215_),
    .A(_1205_),
    .B(_1214_));
 sg13g2_o21ai_1 _5009_ (.B1(_1201_),
    .Y(_1216_),
    .A1(net744),
    .A2(_1215_));
 sg13g2_mux2_1 _5010_ (.A0(_1216_),
    .A1(_1199_),
    .S(_1195_),
    .X(_1217_));
 sg13g2_nor2_1 _5011_ (.A(_1147_),
    .B(_1217_),
    .Y(_0120_));
 sg13g2_a21oi_1 _5012_ (.A1(_1195_),
    .A2(_1216_),
    .Y(_0121_),
    .B1(_1147_));
 sg13g2_nor4_1 _5013_ (.A(_2835_),
    .B(\generated._221[2] ),
    .C(\generated._614[1] ),
    .D(\generated._614[0] ),
    .Y(_1218_));
 sg13g2_nand4_1 _5014_ (.B(\generated._614[2] ),
    .C(_1148_),
    .A(\generated._614[3] ),
    .Y(_1219_),
    .D(_1218_));
 sg13g2_and3_1 _5015_ (.X(_1220_),
    .A(\generated._100[1] ),
    .B(net354),
    .C(net285));
 sg13g2_and2_2 _5016_ (.A(\generated._100[3] ),
    .B(_1220_),
    .X(_1221_));
 sg13g2_nand3_1 _5017_ (.B(_1140_),
    .C(_1221_),
    .A(_2880_),
    .Y(_1222_));
 sg13g2_nor2b_2 _5018_ (.A(_1222_),
    .B_N(_1219_),
    .Y(_1223_));
 sg13g2_nand4_1 _5019_ (.B(_2880_),
    .C(_1140_),
    .A(\generated._614[0] ),
    .Y(_1224_),
    .D(_1221_));
 sg13g2_o21ai_1 _5020_ (.B1(_1224_),
    .Y(_1225_),
    .A1(net427),
    .A2(_1223_));
 sg13g2_nor2_1 _5021_ (.A(net742),
    .B(_1225_),
    .Y(_0122_));
 sg13g2_o21ai_1 _5022_ (.B1(net748),
    .Y(_1226_),
    .A1(_2838_),
    .A2(_1224_));
 sg13g2_a21oi_1 _5023_ (.A1(_2838_),
    .A2(_1224_),
    .Y(_0123_),
    .B1(_1226_));
 sg13g2_and3_1 _5024_ (.X(_1227_),
    .A(\generated._614[2] ),
    .B(\generated._614[1] ),
    .C(\generated._614[0] ));
 sg13g2_nand3_1 _5025_ (.B(\generated._614[1] ),
    .C(\generated._614[0] ),
    .A(\generated._614[2] ),
    .Y(_1228_));
 sg13g2_a22oi_1 _5026_ (.Y(_1229_),
    .B1(_1223_),
    .B2(_1228_),
    .A2(net605),
    .A1(net350));
 sg13g2_a21oi_1 _5027_ (.A1(\generated._614[1] ),
    .A2(\generated._614[0] ),
    .Y(_1230_),
    .B1(net350));
 sg13g2_nor3_1 _5028_ (.A(net742),
    .B(_1229_),
    .C(net351),
    .Y(_0124_));
 sg13g2_o21ai_1 _5029_ (.B1(net748),
    .Y(_1231_),
    .A1(net730),
    .A2(_1227_));
 sg13g2_nand2_1 _5030_ (.Y(_1232_),
    .A(net413),
    .B(_1227_));
 sg13g2_a22oi_1 _5031_ (.Y(_1233_),
    .B1(_1223_),
    .B2(_1232_),
    .A2(net605),
    .A1(net730));
 sg13g2_nor2_1 _5032_ (.A(_1231_),
    .B(_1233_),
    .Y(_0125_));
 sg13g2_nor2_1 _5033_ (.A(net605),
    .B(_1232_),
    .Y(_1234_));
 sg13g2_o21ai_1 _5034_ (.B1(net748),
    .Y(_1235_),
    .A1(net267),
    .A2(_1234_));
 sg13g2_a21oi_1 _5035_ (.A1(net267),
    .A2(_1234_),
    .Y(_0126_),
    .B1(_1235_));
 sg13g2_a21oi_1 _5036_ (.A1(net729),
    .A2(_1234_),
    .Y(_1236_),
    .B1(net727));
 sg13g2_nor2_1 _5037_ (.A(_0397_),
    .B(_1228_),
    .Y(_1237_));
 sg13g2_nor2b_1 _5038_ (.A(net605),
    .B_N(_1237_),
    .Y(_1238_));
 sg13g2_nor3_1 _5039_ (.A(net741),
    .B(net412),
    .C(_1238_),
    .Y(_0127_));
 sg13g2_xnor2_1 _5040_ (.Y(_1239_),
    .A(net726),
    .B(_1237_));
 sg13g2_a22oi_1 _5041_ (.Y(_1240_),
    .B1(_1223_),
    .B2(_1239_),
    .A2(net605),
    .A1(net360));
 sg13g2_nor2_1 _5042_ (.A(net741),
    .B(net361),
    .Y(_0128_));
 sg13g2_nand2_1 _5043_ (.Y(_1241_),
    .A(_0324_),
    .B(_1227_));
 sg13g2_nor2_1 _5044_ (.A(net605),
    .B(_1241_),
    .Y(_1242_));
 sg13g2_a21oi_1 _5045_ (.A1(\generated._221[0] ),
    .A2(_1238_),
    .Y(_1243_),
    .B1(net342));
 sg13g2_nor3_1 _5046_ (.A(net741),
    .B(_1242_),
    .C(net343),
    .Y(_0129_));
 sg13g2_nor2_1 _5047_ (.A(net294),
    .B(_1241_),
    .Y(_1244_));
 sg13g2_nand2b_1 _5048_ (.Y(_1245_),
    .B(_1223_),
    .A_N(_1244_));
 sg13g2_a21oi_1 _5049_ (.A1(net294),
    .A2(_1241_),
    .Y(_1246_),
    .B1(_1245_));
 sg13g2_a21oi_1 _5050_ (.A1(\generated._221[2] ),
    .A2(net605),
    .Y(_1247_),
    .B1(_1246_));
 sg13g2_nor2_1 _5051_ (.A(net741),
    .B(net295),
    .Y(_0130_));
 sg13g2_xnor2_1 _5052_ (.Y(_1248_),
    .A(net314),
    .B(_1244_));
 sg13g2_a22oi_1 _5053_ (.Y(_1249_),
    .B1(_1223_),
    .B2(_1248_),
    .A2(net605),
    .A1(\generated._221[3] ));
 sg13g2_nor2_1 _5054_ (.A(net741),
    .B(net315),
    .Y(_0131_));
 sg13g2_o21ai_1 _5055_ (.B1(net648),
    .Y(_1250_),
    .A1(net357),
    .A2(_3176_));
 sg13g2_nor2_1 _5056_ (.A(_3177_),
    .B(_1250_),
    .Y(_0132_));
 sg13g2_o21ai_1 _5057_ (.B1(net651),
    .Y(_1251_),
    .A1(_3177_),
    .A2(_3184_));
 sg13g2_nor2_1 _5058_ (.A(_3185_),
    .B(_1251_),
    .Y(_0133_));
 sg13g2_o21ai_1 _5059_ (.B1(net651),
    .Y(_1252_),
    .A1(_3186_),
    .A2(_3193_));
 sg13g2_nor2b_1 _5060_ (.A(net430),
    .B_N(_3194_),
    .Y(_0134_));
 sg13g2_nand2_2 _5061_ (.Y(_1253_),
    .A(net695),
    .B(net694));
 sg13g2_inv_1 _5062_ (.Y(_1254_),
    .A(_1253_));
 sg13g2_xor2_1 _5063_ (.B(_1253_),
    .A(net326),
    .X(_1255_));
 sg13g2_nor2_1 _5064_ (.A(net645),
    .B(_1255_),
    .Y(_0135_));
 sg13g2_xnor2_1 _5065_ (.Y(_1256_),
    .A(net606),
    .B(_0348_));
 sg13g2_nor2_2 _5066_ (.A(_1254_),
    .B(_1256_),
    .Y(_1257_));
 sg13g2_xnor2_1 _5067_ (.Y(_1258_),
    .A(_0043_),
    .B(_1257_));
 sg13g2_a21oi_1 _5068_ (.A1(net369),
    .A2(_1253_),
    .Y(_1259_),
    .B1(_1258_));
 sg13g2_and3_1 _5069_ (.X(_1260_),
    .A(net369),
    .B(_1253_),
    .C(_1258_));
 sg13g2_nor3_1 _5070_ (.A(net645),
    .B(net370),
    .C(_1260_),
    .Y(_0136_));
 sg13g2_a21oi_1 _5071_ (.A1(\generated._434[11] ),
    .A2(_1257_),
    .Y(_1261_),
    .B1(_1260_));
 sg13g2_nand2_1 _5072_ (.Y(_1262_),
    .A(net695),
    .B(net606));
 sg13g2_o21ai_1 _5073_ (.B1(_1262_),
    .Y(_1263_),
    .A1(net606),
    .A2(_0346_));
 sg13g2_xor2_1 _5074_ (.B(_1263_),
    .A(net498),
    .X(_1264_));
 sg13g2_nor2_1 _5075_ (.A(_1261_),
    .B(_1264_),
    .Y(_1265_));
 sg13g2_a21oi_1 _5076_ (.A1(_1261_),
    .A2(_1264_),
    .Y(_1266_),
    .B1(net645));
 sg13g2_nor2b_1 _5077_ (.A(net499),
    .B_N(_1266_),
    .Y(_0137_));
 sg13g2_nand2_1 _5078_ (.Y(_1267_),
    .A(net565),
    .B(_1257_));
 sg13g2_xnor2_1 _5079_ (.Y(_1268_),
    .A(net487),
    .B(_1257_));
 sg13g2_nor2_1 _5080_ (.A(_0042_),
    .B(_1263_),
    .Y(_1269_));
 sg13g2_nor2_1 _5081_ (.A(_1265_),
    .B(_1269_),
    .Y(_1270_));
 sg13g2_o21ai_1 _5082_ (.B1(net642),
    .Y(_1271_),
    .A1(_1268_),
    .A2(_1270_));
 sg13g2_a21oi_1 _5083_ (.A1(_1268_),
    .A2(_1270_),
    .Y(_0138_),
    .B1(_1271_));
 sg13g2_o21ai_1 _5084_ (.B1(_1267_),
    .Y(_1272_),
    .A1(_1268_),
    .A2(_1270_));
 sg13g2_nand2_1 _5085_ (.Y(_1273_),
    .A(_1253_),
    .B(_1256_));
 sg13g2_xor2_1 _5086_ (.B(_1273_),
    .A(net446),
    .X(_1274_));
 sg13g2_nor2_1 _5087_ (.A(_1272_),
    .B(_1274_),
    .Y(_1275_));
 sg13g2_nand2_1 _5088_ (.Y(_1276_),
    .A(_1272_),
    .B(_1274_));
 sg13g2_inv_1 _5089_ (.Y(_1277_),
    .A(_1276_));
 sg13g2_nor3_1 _5090_ (.A(net645),
    .B(_1275_),
    .C(_1277_),
    .Y(_0139_));
 sg13g2_a21oi_1 _5091_ (.A1(_2851_),
    .A2(_1273_),
    .Y(_1278_),
    .B1(_1277_));
 sg13g2_xnor2_1 _5092_ (.Y(_1279_),
    .A(net694),
    .B(net609));
 sg13g2_nand2_1 _5093_ (.Y(_1280_),
    .A(net752),
    .B(_1279_));
 sg13g2_nor2_1 _5094_ (.A(\generated._434[15] ),
    .B(_1279_),
    .Y(_1281_));
 sg13g2_xnor2_1 _5095_ (.Y(_1282_),
    .A(net470),
    .B(_1279_));
 sg13g2_xnor2_1 _5096_ (.Y(_1283_),
    .A(_1278_),
    .B(_1282_));
 sg13g2_nor2_1 _5097_ (.A(net645),
    .B(net471),
    .Y(_0140_));
 sg13g2_o21ai_1 _5098_ (.B1(_1280_),
    .Y(_1284_),
    .A1(_1278_),
    .A2(_1281_));
 sg13g2_xor2_1 _5099_ (.B(_1256_),
    .A(net463),
    .X(_1285_));
 sg13g2_nor2_1 _5100_ (.A(_1284_),
    .B(_1285_),
    .Y(_1286_));
 sg13g2_and2_1 _5101_ (.A(_1284_),
    .B(_1285_),
    .X(_1287_));
 sg13g2_nor3_1 _5102_ (.A(net645),
    .B(net464),
    .C(_1287_),
    .Y(_0141_));
 sg13g2_a21oi_1 _5103_ (.A1(_2850_),
    .A2(_1256_),
    .Y(_1288_),
    .B1(_1287_));
 sg13g2_xnor2_1 _5104_ (.Y(_1289_),
    .A(net554),
    .B(net609));
 sg13g2_nor2_1 _5105_ (.A(_1288_),
    .B(_1289_),
    .Y(_1290_));
 sg13g2_a21oi_1 _5106_ (.A1(_1288_),
    .A2(_1289_),
    .Y(_1291_),
    .B1(net645));
 sg13g2_nor2b_1 _5107_ (.A(_1290_),
    .B_N(net555),
    .Y(_0142_));
 sg13g2_a21oi_1 _5108_ (.A1(_2855_),
    .A2(net609),
    .Y(_1292_),
    .B1(_1290_));
 sg13g2_xnor2_1 _5109_ (.Y(_1293_),
    .A(\generated._434[18] ),
    .B(net609));
 sg13g2_nor2_1 _5110_ (.A(_1292_),
    .B(_1293_),
    .Y(_1294_));
 sg13g2_a21oi_1 _5111_ (.A1(_1292_),
    .A2(_1293_),
    .Y(_1295_),
    .B1(net646));
 sg13g2_nor2b_1 _5112_ (.A(net481),
    .B_N(_1295_),
    .Y(_0143_));
 sg13g2_nand3_1 _5113_ (.B(net606),
    .C(_1290_),
    .A(\generated._434[18] ),
    .Y(_1296_));
 sg13g2_nand2_1 _5114_ (.Y(_1297_),
    .A(_0038_),
    .B(net609));
 sg13g2_o21ai_1 _5115_ (.B1(_1296_),
    .Y(_1298_),
    .A1(_1294_),
    .A2(_1297_));
 sg13g2_o21ai_1 _5116_ (.B1(net641),
    .Y(_1299_),
    .A1(net331),
    .A2(_1298_));
 sg13g2_a21oi_1 _5117_ (.A1(net331),
    .A2(_1298_),
    .Y(_0144_),
    .B1(_1299_));
 sg13g2_and2_1 _5118_ (.A(net723),
    .B(_1221_),
    .X(_1300_));
 sg13g2_nor3_1 _5119_ (.A(\generated._100[5] ),
    .B(\generated._100[6] ),
    .C(net722),
    .Y(_1301_));
 sg13g2_nand4_1 _5120_ (.B(net564),
    .C(_1300_),
    .A(net280),
    .Y(_1302_),
    .D(_1301_));
 sg13g2_nand2_2 _5121_ (.Y(_1303_),
    .A(net748),
    .B(_1302_));
 sg13g2_and3_1 _5122_ (.X(_0145_),
    .A(net748),
    .B(net254),
    .C(_1302_));
 sg13g2_xnor2_1 _5123_ (.Y(_1304_),
    .A(\generated._100[1] ),
    .B(net354));
 sg13g2_nor2_1 _5124_ (.A(_1303_),
    .B(net355),
    .Y(_0146_));
 sg13g2_a21oi_1 _5125_ (.A1(\generated._100[1] ),
    .A2(\generated._100[0] ),
    .Y(_1305_),
    .B1(net285));
 sg13g2_nor3_1 _5126_ (.A(net743),
    .B(_1220_),
    .C(net286),
    .Y(_0147_));
 sg13g2_o21ai_1 _5127_ (.B1(net748),
    .Y(_1306_),
    .A1(net442),
    .A2(_1220_));
 sg13g2_nor2_1 _5128_ (.A(_1221_),
    .B(net443),
    .Y(_0148_));
 sg13g2_nor2_1 _5129_ (.A(net723),
    .B(_1221_),
    .Y(_1307_));
 sg13g2_nor3_1 _5130_ (.A(net743),
    .B(_1300_),
    .C(_1307_),
    .Y(_0149_));
 sg13g2_xnor2_1 _5131_ (.Y(_1308_),
    .A(net388),
    .B(_1300_));
 sg13g2_nor2_1 _5132_ (.A(_1303_),
    .B(_1308_),
    .Y(_0150_));
 sg13g2_a21oi_1 _5133_ (.A1(\generated._100[5] ),
    .A2(_1300_),
    .Y(_1309_),
    .B1(net381));
 sg13g2_and2_1 _5134_ (.A(_1141_),
    .B(_1221_),
    .X(_1310_));
 sg13g2_nor3_1 _5135_ (.A(_1303_),
    .B(net382),
    .C(_1310_),
    .Y(_0151_));
 sg13g2_xnor2_1 _5136_ (.Y(_1311_),
    .A(net302),
    .B(_1310_));
 sg13g2_nor2_1 _5137_ (.A(_1303_),
    .B(_1311_),
    .Y(_0152_));
 sg13g2_and3_1 _5138_ (.X(_1312_),
    .A(net722),
    .B(net280),
    .C(_1310_));
 sg13g2_a21oi_1 _5139_ (.A1(net722),
    .A2(_1310_),
    .Y(_1313_),
    .B1(net280));
 sg13g2_nor3_1 _5140_ (.A(_1303_),
    .B(_1312_),
    .C(net281),
    .Y(_0153_));
 sg13g2_a21oi_1 _5141_ (.A1(net366),
    .A2(_1312_),
    .Y(_1314_),
    .B1(_1303_));
 sg13g2_o21ai_1 _5142_ (.B1(_1314_),
    .Y(_1315_),
    .A1(net366),
    .A2(_1312_));
 sg13g2_inv_1 _5143_ (.Y(_0154_),
    .A(_1315_));
 sg13g2_and2_1 _5144_ (.A(net707),
    .B(net703),
    .X(_1316_));
 sg13g2_nand2_1 _5145_ (.Y(_1317_),
    .A(net707),
    .B(net703));
 sg13g2_xnor2_1 _5146_ (.Y(_1318_),
    .A(net296),
    .B(_1316_));
 sg13g2_nor2_1 _5147_ (.A(net652),
    .B(_1318_),
    .Y(_0155_));
 sg13g2_xnor2_1 _5148_ (.Y(_1319_),
    .A(net619),
    .B(_3020_));
 sg13g2_inv_1 _5149_ (.Y(_1320_),
    .A(_1319_));
 sg13g2_nand2_1 _5150_ (.Y(_1321_),
    .A(_1317_),
    .B(_1319_));
 sg13g2_and3_1 _5151_ (.X(_1322_),
    .A(\generated._1084[1] ),
    .B(_1317_),
    .C(_1319_));
 sg13g2_xnor2_1 _5152_ (.Y(_1323_),
    .A(\generated._1084[1] ),
    .B(_1321_));
 sg13g2_a21oi_1 _5153_ (.A1(net335),
    .A2(_1317_),
    .Y(_1324_),
    .B1(_1323_));
 sg13g2_and3_1 _5154_ (.X(_1325_),
    .A(net335),
    .B(_1317_),
    .C(_1323_));
 sg13g2_nor3_1 _5155_ (.A(net652),
    .B(net336),
    .C(_1325_),
    .Y(_0156_));
 sg13g2_or2_1 _5156_ (.X(_1326_),
    .B(_1325_),
    .A(_1322_));
 sg13g2_nand2_1 _5157_ (.Y(_1327_),
    .A(net618),
    .B(_3022_));
 sg13g2_o21ai_1 _5158_ (.B1(_1327_),
    .Y(_1328_),
    .A1(net707),
    .A2(net618));
 sg13g2_xor2_1 _5159_ (.B(_1328_),
    .A(net422),
    .X(_1329_));
 sg13g2_nor2_1 _5160_ (.A(_1326_),
    .B(_1329_),
    .Y(_1330_));
 sg13g2_and2_1 _5161_ (.A(_1326_),
    .B(_1329_),
    .X(_1331_));
 sg13g2_nor3_1 _5162_ (.A(net652),
    .B(_1330_),
    .C(_1331_),
    .Y(_0157_));
 sg13g2_a21oi_1 _5163_ (.A1(net422),
    .A2(_1328_),
    .Y(_1332_),
    .B1(_1331_));
 sg13g2_xnor2_1 _5164_ (.Y(_1333_),
    .A(_2866_),
    .B(_1321_));
 sg13g2_or2_1 _5165_ (.X(_1334_),
    .B(_1333_),
    .A(_1332_));
 sg13g2_nand2_1 _5166_ (.Y(_1335_),
    .A(net648),
    .B(_1334_));
 sg13g2_a21oi_1 _5167_ (.A1(_1332_),
    .A2(_1333_),
    .Y(_0158_),
    .B1(_1335_));
 sg13g2_o21ai_1 _5168_ (.B1(_1334_),
    .Y(_1336_),
    .A1(_2866_),
    .A2(_1321_));
 sg13g2_nor2_1 _5169_ (.A(_1316_),
    .B(_1319_),
    .Y(_1337_));
 sg13g2_nor2_1 _5170_ (.A(_2867_),
    .B(_1337_),
    .Y(_1338_));
 sg13g2_xnor2_1 _5171_ (.Y(_1339_),
    .A(net505),
    .B(_1337_));
 sg13g2_nor2_1 _5172_ (.A(_1336_),
    .B(_1339_),
    .Y(_1340_));
 sg13g2_nand2_1 _5173_ (.Y(_1341_),
    .A(_1336_),
    .B(_1339_));
 sg13g2_inv_1 _5174_ (.Y(_1342_),
    .A(_1341_));
 sg13g2_nor3_1 _5175_ (.A(net652),
    .B(_1340_),
    .C(_1342_),
    .Y(_0159_));
 sg13g2_nor2_1 _5176_ (.A(_1338_),
    .B(_1342_),
    .Y(_1343_));
 sg13g2_xnor2_1 _5177_ (.Y(_1344_),
    .A(net703),
    .B(net619));
 sg13g2_xor2_1 _5178_ (.B(_1344_),
    .A(net465),
    .X(_1345_));
 sg13g2_nor2b_1 _5179_ (.A(_1345_),
    .B_N(_1343_),
    .Y(_1346_));
 sg13g2_nor2b_1 _5180_ (.A(_1343_),
    .B_N(_1345_),
    .Y(_1347_));
 sg13g2_nor3_1 _5181_ (.A(net652),
    .B(_1346_),
    .C(_1347_),
    .Y(_0160_));
 sg13g2_a21oi_1 _5182_ (.A1(net465),
    .A2(_1344_),
    .Y(_1348_),
    .B1(_1347_));
 sg13g2_xor2_1 _5183_ (.B(_1319_),
    .A(\generated._1084[6] ),
    .X(_1349_));
 sg13g2_and2_1 _5184_ (.A(_1348_),
    .B(_1349_),
    .X(_1350_));
 sg13g2_nor2_1 _5185_ (.A(_1348_),
    .B(_1349_),
    .Y(_1351_));
 sg13g2_nor3_1 _5186_ (.A(net653),
    .B(_1350_),
    .C(_1351_),
    .Y(_0161_));
 sg13g2_a21o_1 _5187_ (.A2(_1320_),
    .A1(\generated._1084[6] ),
    .B1(_1351_),
    .X(_1352_));
 sg13g2_nand2_1 _5188_ (.Y(_1353_),
    .A(net527),
    .B(net619));
 sg13g2_xor2_1 _5189_ (.B(net619),
    .A(net527),
    .X(_1354_));
 sg13g2_o21ai_1 _5190_ (.B1(net648),
    .Y(_1355_),
    .A1(_1352_),
    .A2(_1354_));
 sg13g2_a21oi_1 _5191_ (.A1(_1352_),
    .A2(_1354_),
    .Y(_0162_),
    .B1(_1355_));
 sg13g2_xnor2_1 _5192_ (.Y(_1356_),
    .A(net428),
    .B(net622));
 sg13g2_o21ai_1 _5193_ (.B1(_1352_),
    .Y(_1357_),
    .A1(\generated._1084[7] ),
    .A2(net619));
 sg13g2_and3_1 _5194_ (.X(_1358_),
    .A(_1353_),
    .B(_1356_),
    .C(_1357_));
 sg13g2_a21oi_1 _5195_ (.A1(_1353_),
    .A2(_1357_),
    .Y(_1359_),
    .B1(_1356_));
 sg13g2_nor3_1 _5196_ (.A(net652),
    .B(_1358_),
    .C(_1359_),
    .Y(_0163_));
 sg13g2_a21oi_1 _5197_ (.A1(net428),
    .A2(net622),
    .Y(_1360_),
    .B1(_1359_));
 sg13g2_xnor2_1 _5198_ (.Y(_1361_),
    .A(net719),
    .B(net622));
 sg13g2_o21ai_1 _5199_ (.B1(net648),
    .Y(_1362_),
    .A1(_1360_),
    .A2(_1361_));
 sg13g2_a21oi_1 _5200_ (.A1(_1360_),
    .A2(_1361_),
    .Y(_0164_),
    .B1(_1362_));
 sg13g2_nand2_1 _5201_ (.Y(_1363_),
    .A(net456),
    .B(_3011_));
 sg13g2_and3_1 _5202_ (.X(_0165_),
    .A(net747),
    .B(net262),
    .C(_1363_));
 sg13g2_o21ai_1 _5203_ (.B1(net747),
    .Y(_1364_),
    .A1(net333),
    .A2(\generated._1078[1] ));
 sg13g2_a21oi_1 _5204_ (.A1(net333),
    .A2(\generated._1078[1] ),
    .Y(_0166_),
    .B1(_1364_));
 sg13g2_nand3_1 _5205_ (.B(\generated._1078[1] ),
    .C(\generated._1078[2] ),
    .A(net333),
    .Y(_1365_));
 sg13g2_a21o_1 _5206_ (.A2(\generated._1078[1] ),
    .A1(net333),
    .B1(net456),
    .X(_1366_));
 sg13g2_and4_1 _5207_ (.A(net747),
    .B(_1363_),
    .C(_1365_),
    .D(net457),
    .X(_0167_));
 sg13g2_xnor2_1 _5208_ (.Y(_1367_),
    .A(net391),
    .B(_1365_));
 sg13g2_and3_1 _5209_ (.X(_0168_),
    .A(net747),
    .B(_1363_),
    .C(net392));
 sg13g2_xor2_1 _5210_ (.B(_3028_),
    .A(net390),
    .X(_1368_));
 sg13g2_nor2_1 _5211_ (.A(net653),
    .B(_1368_),
    .Y(_0169_));
 sg13g2_a21oi_1 _5212_ (.A1(_3039_),
    .A2(_3040_),
    .Y(_1369_),
    .B1(net653));
 sg13g2_nor2b_1 _5213_ (.A(_3041_),
    .B_N(net476),
    .Y(_0170_));
 sg13g2_nor3_1 _5214_ (.A(_3038_),
    .B(_3041_),
    .C(_3043_),
    .Y(_1370_));
 sg13g2_nor3_1 _5215_ (.A(net653),
    .B(_3044_),
    .C(net462),
    .Y(_0171_));
 sg13g2_and2_1 _5216_ (.A(net251),
    .B(net651),
    .X(_0172_));
 sg13g2_nor3_1 _5217_ (.A(net652),
    .B(_3020_),
    .C(_1316_),
    .Y(_0173_));
 sg13g2_nor4_1 _5218_ (.A(\generated._614[2] ),
    .B(\generated._614[1] ),
    .C(\generated._614[0] ),
    .D(_1149_),
    .Y(_1371_));
 sg13g2_and2_2 _5219_ (.A(net623),
    .B(_1371_),
    .X(_1372_));
 sg13g2_o21ai_1 _5220_ (.B1(net747),
    .Y(_1373_),
    .A1(\generated._1000[0] ),
    .A2(_1372_));
 sg13g2_a21oi_1 _5221_ (.A1(_2834_),
    .A2(_1372_),
    .Y(_0174_),
    .B1(_1373_));
 sg13g2_a21oi_1 _5222_ (.A1(\generated._1000[0] ),
    .A2(_1372_),
    .Y(_1374_),
    .B1(net303));
 sg13g2_nand3_1 _5223_ (.B(\generated._1000[0] ),
    .C(_1372_),
    .A(net303),
    .Y(_1375_));
 sg13g2_nand2_1 _5224_ (.Y(_1376_),
    .A(net747),
    .B(_1375_));
 sg13g2_nor2_1 _5225_ (.A(net304),
    .B(_1376_),
    .Y(_0175_));
 sg13g2_and2_1 _5226_ (.A(_2833_),
    .B(_1375_),
    .X(_1377_));
 sg13g2_nor2_1 _5227_ (.A(_2833_),
    .B(_1375_),
    .Y(_1378_));
 sg13g2_nor3_1 _5228_ (.A(net743),
    .B(net419),
    .C(_1378_),
    .Y(_0176_));
 sg13g2_and2_1 _5229_ (.A(net371),
    .B(_1378_),
    .X(_1379_));
 sg13g2_o21ai_1 _5230_ (.B1(net745),
    .Y(_1380_),
    .A1(net371),
    .A2(_1378_));
 sg13g2_nor2_1 _5231_ (.A(_1379_),
    .B(net372),
    .Y(_0177_));
 sg13g2_xnor2_1 _5232_ (.Y(_1381_),
    .A(net362),
    .B(_1379_));
 sg13g2_nor2_1 _5233_ (.A(net743),
    .B(net363),
    .Y(_0178_));
 sg13g2_a21oi_1 _5234_ (.A1(\generated._406[4] ),
    .A2(_1379_),
    .Y(_1382_),
    .B1(net310));
 sg13g2_nand3_1 _5235_ (.B(\generated._406[4] ),
    .C(_1379_),
    .A(net310),
    .Y(_1383_));
 sg13g2_nand2_1 _5236_ (.Y(_1384_),
    .A(net745),
    .B(_1383_));
 sg13g2_nor2_1 _5237_ (.A(net311),
    .B(_1384_),
    .Y(_0179_));
 sg13g2_or2_1 _5238_ (.X(_1385_),
    .B(_1383_),
    .A(_2832_));
 sg13g2_nand2_1 _5239_ (.Y(_1386_),
    .A(net745),
    .B(_1385_));
 sg13g2_a21oi_1 _5240_ (.A1(_2832_),
    .A2(_1383_),
    .Y(_0180_),
    .B1(_1386_));
 sg13g2_o21ai_1 _5241_ (.B1(net745),
    .Y(_1387_),
    .A1(_2831_),
    .A2(_1385_));
 sg13g2_a21oi_1 _5242_ (.A1(_2831_),
    .A2(_1385_),
    .Y(_0181_),
    .B1(_1387_));
 sg13g2_nand2_1 _5243_ (.Y(_1388_),
    .A(net452),
    .B(_0333_));
 sg13g2_and3_1 _5244_ (.X(_0182_),
    .A(net746),
    .B(net256),
    .C(_1388_));
 sg13g2_o21ai_1 _5245_ (.B1(net746),
    .Y(_1389_),
    .A1(net306),
    .A2(\generated._71[1] ));
 sg13g2_a21oi_1 _5246_ (.A1(net306),
    .A2(\generated._71[1] ),
    .Y(_0183_),
    .B1(_1389_));
 sg13g2_nand3_1 _5247_ (.B(\generated._71[1] ),
    .C(\generated._71[2] ),
    .A(net306),
    .Y(_1390_));
 sg13g2_a21o_1 _5248_ (.A2(\generated._71[1] ),
    .A1(net306),
    .B1(net452),
    .X(_1391_));
 sg13g2_and4_1 _5249_ (.A(net746),
    .B(_1388_),
    .C(_1390_),
    .D(net453),
    .X(_0184_));
 sg13g2_xnor2_1 _5250_ (.Y(_1392_),
    .A(net400),
    .B(_1390_));
 sg13g2_and3_1 _5251_ (.X(_0185_),
    .A(net746),
    .B(_1388_),
    .C(net401));
 sg13g2_nand2_1 _5252_ (.Y(_1393_),
    .A(net376),
    .B(_0590_));
 sg13g2_and3_1 _5253_ (.X(_0186_),
    .A(net746),
    .B(net258),
    .C(_1393_));
 sg13g2_o21ai_1 _5254_ (.B1(net746),
    .Y(_1394_),
    .A1(net300),
    .A2(\generated._63[0] ));
 sg13g2_a21oi_1 _5255_ (.A1(net300),
    .A2(\generated._63[0] ),
    .Y(_0187_),
    .B1(_1394_));
 sg13g2_nand3_1 _5256_ (.B(\generated._63[0] ),
    .C(net376),
    .A(net300),
    .Y(_1395_));
 sg13g2_a21o_1 _5257_ (.A2(net445),
    .A1(net300),
    .B1(net376),
    .X(_1396_));
 sg13g2_and4_1 _5258_ (.A(net746),
    .B(_1393_),
    .C(_1395_),
    .D(_1396_),
    .X(_0188_));
 sg13g2_xnor2_1 _5259_ (.Y(_1397_),
    .A(net403),
    .B(_1395_));
 sg13g2_and3_1 _5260_ (.X(_0189_),
    .A(net746),
    .B(_1393_),
    .C(net404));
 sg13g2_xor2_1 _5261_ (.B(_0354_),
    .A(net364),
    .X(_1398_));
 sg13g2_nor2_1 _5262_ (.A(net647),
    .B(_1398_),
    .Y(_0190_));
 sg13g2_a21oi_1 _5263_ (.A1(_0365_),
    .A2(_0366_),
    .Y(_1399_),
    .B1(net647));
 sg13g2_nor2b_1 _5264_ (.A(_0367_),
    .B_N(net507),
    .Y(_0191_));
 sg13g2_nor3_1 _5265_ (.A(_0364_),
    .B(_0367_),
    .C(_0369_),
    .Y(_1400_));
 sg13g2_nor3_1 _5266_ (.A(net647),
    .B(_0370_),
    .C(net434),
    .Y(_0192_));
 sg13g2_and2_1 _5267_ (.A(net252),
    .B(net643),
    .X(_0193_));
 sg13g2_nor3_1 _5268_ (.A(net645),
    .B(_0348_),
    .C(_1254_),
    .Y(_0194_));
 sg13g2_o21ai_1 _5269_ (.B1(net643),
    .Y(_1401_),
    .A1(net431),
    .A2(_0487_));
 sg13g2_nor2_1 _5270_ (.A(_0488_),
    .B(_1401_),
    .Y(_0195_));
 sg13g2_o21ai_1 _5271_ (.B1(net643),
    .Y(_1402_),
    .A1(_0488_),
    .A2(_0495_));
 sg13g2_nor2b_1 _5272_ (.A(_1402_),
    .B_N(_0496_),
    .Y(_0196_));
 sg13g2_nand3_1 _5273_ (.B(_0497_),
    .C(_0504_),
    .A(_0496_),
    .Y(_1403_));
 sg13g2_and3_1 _5274_ (.X(_0197_),
    .A(net643),
    .B(_0505_),
    .C(_1403_));
 sg13g2_nor3_2 _5275_ (.A(net686),
    .B(\generated._512[0] ),
    .C(\generated._512[1] ),
    .Y(_1404_));
 sg13g2_nand2b_2 _5276_ (.Y(_1405_),
    .B(_1404_),
    .A_N(\generated._512[2] ));
 sg13g2_xnor2_1 _5277_ (.Y(_1406_),
    .A(\generated._512[3] ),
    .B(_1405_));
 sg13g2_nand3_1 _5278_ (.B(net571),
    .C(_0664_),
    .A(_0059_),
    .Y(_1407_));
 sg13g2_o21ai_1 _5279_ (.B1(_1406_),
    .Y(_1408_),
    .A1(net573),
    .A2(_0663_));
 sg13g2_and2_2 _5280_ (.A(_1407_),
    .B(_1408_),
    .X(_1409_));
 sg13g2_nand3_1 _5281_ (.B(_1407_),
    .C(_1408_),
    .A(net594),
    .Y(_1410_));
 sg13g2_xor2_1 _5282_ (.B(_1404_),
    .A(\generated._512[2] ),
    .X(_1411_));
 sg13g2_nor3_2 _5283_ (.A(_0055_),
    .B(net573),
    .C(net597),
    .Y(_1412_));
 sg13g2_a21oi_2 _5284_ (.B1(_1411_),
    .Y(_1413_),
    .A2(net596),
    .A1(net571));
 sg13g2_or2_1 _5285_ (.X(_1414_),
    .B(_1413_),
    .A(_1412_));
 sg13g2_nor2_2 _5286_ (.A(_1412_),
    .B(_1413_),
    .Y(_1415_));
 sg13g2_o21ai_1 _5287_ (.B1(net598),
    .Y(_1416_),
    .A1(_1412_),
    .A2(_1413_));
 sg13g2_nand3_1 _5288_ (.B(_1407_),
    .C(_1408_),
    .A(net598),
    .Y(_1417_));
 sg13g2_o21ai_1 _5289_ (.B1(net594),
    .Y(_1418_),
    .A1(_1412_),
    .A2(_1413_));
 sg13g2_or2_1 _5290_ (.X(_1419_),
    .B(_1416_),
    .A(_1410_));
 sg13g2_nor3_2 _5291_ (.A(\generated._512[3] ),
    .B(\generated._512[4] ),
    .C(_1405_),
    .Y(_1420_));
 sg13g2_o21ai_1 _5292_ (.B1(\generated._512[4] ),
    .Y(_1421_),
    .A1(\generated._512[3] ),
    .A2(_1405_));
 sg13g2_nand2b_1 _5293_ (.Y(_1422_),
    .B(_1421_),
    .A_N(_1420_));
 sg13g2_nor3_1 _5294_ (.A(_0062_),
    .B(net573),
    .C(net597),
    .Y(_1423_));
 sg13g2_a21oi_1 _5295_ (.A1(_0638_),
    .A2(net596),
    .Y(_1424_),
    .B1(_1422_));
 sg13g2_or2_2 _5296_ (.X(_1425_),
    .B(_1424_),
    .A(_1423_));
 sg13g2_nand2_1 _5297_ (.Y(_1426_),
    .A(_0405_),
    .B(_1425_));
 sg13g2_and2_1 _5298_ (.A(_1417_),
    .B(_1418_),
    .X(_1427_));
 sg13g2_xor2_1 _5299_ (.B(_1418_),
    .A(_1417_),
    .X(_1428_));
 sg13g2_o21ai_1 _5300_ (.B1(_1419_),
    .Y(_1429_),
    .A1(_1426_),
    .A2(_1427_));
 sg13g2_nor2b_1 _5301_ (.A(\generated._512[5] ),
    .B_N(_1420_),
    .Y(_1430_));
 sg13g2_xor2_1 _5302_ (.B(_1420_),
    .A(\generated._512[5] ),
    .X(_1431_));
 sg13g2_nor3_1 _5303_ (.A(_0065_),
    .B(net573),
    .C(net597),
    .Y(_1432_));
 sg13g2_a21oi_1 _5304_ (.A1(_0638_),
    .A2(net596),
    .Y(_1433_),
    .B1(_1431_));
 sg13g2_or2_2 _5305_ (.X(_1434_),
    .B(_1433_),
    .A(_1432_));
 sg13g2_nand2_1 _5306_ (.Y(_1435_),
    .A(_0405_),
    .B(_1434_));
 sg13g2_o21ai_1 _5307_ (.B1(net594),
    .Y(_1436_),
    .A1(_1423_),
    .A2(_1424_));
 sg13g2_o21ai_1 _5308_ (.B1(net598),
    .Y(_1437_),
    .A1(_1423_),
    .A2(_1424_));
 sg13g2_or2_1 _5309_ (.X(_1438_),
    .B(_1436_),
    .A(_1417_));
 sg13g2_and2_1 _5310_ (.A(_1410_),
    .B(_1437_),
    .X(_1439_));
 sg13g2_xor2_1 _5311_ (.B(_1437_),
    .A(_1410_),
    .X(_1440_));
 sg13g2_xnor2_1 _5312_ (.Y(_1441_),
    .A(_1435_),
    .B(_1440_));
 sg13g2_and2_1 _5313_ (.A(_1429_),
    .B(_1441_),
    .X(_1442_));
 sg13g2_or2_1 _5314_ (.X(_1443_),
    .B(_1441_),
    .A(_1429_));
 sg13g2_xnor2_1 _5315_ (.Y(_1444_),
    .A(_1429_),
    .B(_1441_));
 sg13g2_a21oi_1 _5316_ (.A1(_2845_),
    .A2(_0436_),
    .Y(_1445_),
    .B1(net616));
 sg13g2_inv_2 _5317_ (.Y(_1446_),
    .A(net588));
 sg13g2_o21ai_1 _5318_ (.B1(\generated._512[1] ),
    .Y(_1447_),
    .A1(net686),
    .A2(\generated._512[0] ));
 sg13g2_nand2b_1 _5319_ (.Y(_1448_),
    .B(_1447_),
    .A_N(_1404_));
 sg13g2_nor3_2 _5320_ (.A(_0054_),
    .B(net573),
    .C(net597),
    .Y(_1449_));
 sg13g2_a21oi_2 _5321_ (.B1(_1448_),
    .Y(_1450_),
    .A2(net596),
    .A1(net571));
 sg13g2_or2_2 _5322_ (.X(_1451_),
    .B(_1450_),
    .A(_1449_));
 sg13g2_nor2_1 _5323_ (.A(_1449_),
    .B(_1450_),
    .Y(_1452_));
 sg13g2_nor2_1 _5324_ (.A(_1446_),
    .B(_1452_),
    .Y(_1453_));
 sg13g2_nand2b_1 _5325_ (.Y(_1454_),
    .B(_1430_),
    .A_N(\generated._512[6] ));
 sg13g2_xor2_1 _5326_ (.B(_1430_),
    .A(\generated._512[6] ),
    .X(_1455_));
 sg13g2_nand3_1 _5327_ (.B(net571),
    .C(net596),
    .A(_0067_),
    .Y(_1456_));
 sg13g2_o21ai_1 _5328_ (.B1(_1455_),
    .Y(_1457_),
    .A1(_0637_),
    .A2(net597));
 sg13g2_nand2_2 _5329_ (.Y(_1458_),
    .A(_1456_),
    .B(_1457_));
 sg13g2_xor2_1 _5330_ (.B(_0571_),
    .A(_0453_),
    .X(_1459_));
 sg13g2_nor2b_2 _5331_ (.A(_1458_),
    .B_N(net581),
    .Y(_1460_));
 sg13g2_nor2_1 _5332_ (.A(_0396_),
    .B(_1415_),
    .Y(_1461_));
 sg13g2_nor2_1 _5333_ (.A(_0396_),
    .B(_1458_),
    .Y(_1462_));
 sg13g2_nand2_1 _5334_ (.Y(_1463_),
    .A(_1414_),
    .B(net582));
 sg13g2_xnor2_1 _5335_ (.Y(_1464_),
    .A(_1462_),
    .B(_1463_));
 sg13g2_xor2_1 _5336_ (.B(_1464_),
    .A(_1453_),
    .X(_1465_));
 sg13g2_a21oi_1 _5337_ (.A1(_1443_),
    .A2(_1465_),
    .Y(_1466_),
    .B1(_1442_));
 sg13g2_o21ai_1 _5338_ (.B1(_1438_),
    .Y(_1467_),
    .A1(_1435_),
    .A2(_1439_));
 sg13g2_nor2_1 _5339_ (.A(_0406_),
    .B(_1458_),
    .Y(_1468_));
 sg13g2_nand2_1 _5340_ (.Y(_1469_),
    .A(net594),
    .B(_1434_));
 sg13g2_o21ai_1 _5341_ (.B1(net598),
    .Y(_1470_),
    .A1(_1432_),
    .A2(_1433_));
 sg13g2_nor2_1 _5342_ (.A(_1436_),
    .B(_1470_),
    .Y(_1471_));
 sg13g2_xor2_1 _5343_ (.B(_1470_),
    .A(_1436_),
    .X(_1472_));
 sg13g2_xor2_1 _5344_ (.B(_1472_),
    .A(_1468_),
    .X(_1473_));
 sg13g2_and2_1 _5345_ (.A(_1467_),
    .B(_1473_),
    .X(_1474_));
 sg13g2_or2_1 _5346_ (.X(_1475_),
    .B(_1473_),
    .A(_1467_));
 sg13g2_xnor2_1 _5347_ (.Y(_1476_),
    .A(_1467_),
    .B(_1473_));
 sg13g2_nand2_1 _5348_ (.Y(_1477_),
    .A(_1414_),
    .B(net589));
 sg13g2_nand2_1 _5349_ (.Y(_1478_),
    .A(net655),
    .B(_1409_));
 sg13g2_nor2_1 _5350_ (.A(\generated._512[7] ),
    .B(_1454_),
    .Y(_1479_));
 sg13g2_xnor2_1 _5351_ (.Y(_1480_),
    .A(\generated._512[7] ),
    .B(_1454_));
 sg13g2_nor3_1 _5352_ (.A(_0069_),
    .B(_0637_),
    .C(net597),
    .Y(_1481_));
 sg13g2_a21oi_1 _5353_ (.A1(_0638_),
    .A2(_0664_),
    .Y(_1482_),
    .B1(_1480_));
 sg13g2_or2_2 _5354_ (.X(_1483_),
    .B(_1482_),
    .A(_1481_));
 sg13g2_nand2_1 _5355_ (.Y(_1484_),
    .A(net581),
    .B(_1483_));
 sg13g2_nand2_1 _5356_ (.Y(_1485_),
    .A(_1409_),
    .B(net581));
 sg13g2_nand2_1 _5357_ (.Y(_1486_),
    .A(net655),
    .B(_1483_));
 sg13g2_xor2_1 _5358_ (.B(_1486_),
    .A(_1485_),
    .X(_1487_));
 sg13g2_nand2b_1 _5359_ (.Y(_1488_),
    .B(_1487_),
    .A_N(_1477_));
 sg13g2_xnor2_1 _5360_ (.Y(_1489_),
    .A(_1477_),
    .B(_1487_));
 sg13g2_xnor2_1 _5361_ (.Y(_1490_),
    .A(_1476_),
    .B(_1489_));
 sg13g2_nand2b_1 _5362_ (.Y(_1491_),
    .B(_1490_),
    .A_N(_1466_));
 sg13g2_nor2_1 _5363_ (.A(net589),
    .B(_1452_),
    .Y(_1492_));
 sg13g2_a221oi_1 _5364_ (.B2(_1453_),
    .C1(_1492_),
    .B1(_1464_),
    .A1(_1460_),
    .Y(_1493_),
    .A2(_1461_));
 sg13g2_nor2b_1 _5365_ (.A(_1490_),
    .B_N(_1466_),
    .Y(_1494_));
 sg13g2_xnor2_1 _5366_ (.Y(_1495_),
    .A(_1466_),
    .B(_1490_));
 sg13g2_o21ai_1 _5367_ (.B1(_1491_),
    .Y(_1496_),
    .A1(_1493_),
    .A2(_1494_));
 sg13g2_o21ai_1 _5368_ (.B1(_1488_),
    .Y(_1497_),
    .A1(_1485_),
    .A2(_1486_));
 sg13g2_nand2_1 _5369_ (.Y(_1498_),
    .A(_1415_),
    .B(_1446_));
 sg13g2_o21ai_1 _5370_ (.B1(_1498_),
    .Y(_1499_),
    .A1(_1409_),
    .A2(_1446_));
 sg13g2_nor2b_1 _5371_ (.A(_1499_),
    .B_N(_1497_),
    .Y(_1500_));
 sg13g2_xnor2_1 _5372_ (.Y(_1501_),
    .A(_1497_),
    .B(_1499_));
 sg13g2_a21oi_1 _5373_ (.A1(_1475_),
    .A2(_1489_),
    .Y(_1502_),
    .B1(_1474_));
 sg13g2_a21o_1 _5374_ (.A2(_1472_),
    .A1(_1468_),
    .B1(_1471_),
    .X(_1503_));
 sg13g2_nand3_1 _5375_ (.B(_1456_),
    .C(_1457_),
    .A(net594),
    .Y(_1504_));
 sg13g2_nor2b_1 _5376_ (.A(_1458_),
    .B_N(net599),
    .Y(_1505_));
 sg13g2_nor2_2 _5377_ (.A(_1470_),
    .B(_1504_),
    .Y(_1506_));
 sg13g2_xnor2_1 _5378_ (.Y(_1507_),
    .A(_1469_),
    .B(_1505_));
 sg13g2_and2_1 _5379_ (.A(_1503_),
    .B(_1507_),
    .X(_1508_));
 sg13g2_or2_1 _5380_ (.X(_1509_),
    .B(_1507_),
    .A(_1503_));
 sg13g2_xnor2_1 _5381_ (.Y(_1510_),
    .A(_1503_),
    .B(_1507_));
 sg13g2_nand2_1 _5382_ (.Y(_1511_),
    .A(_1425_),
    .B(net581));
 sg13g2_xor2_1 _5383_ (.B(_1479_),
    .A(\generated._511 ),
    .X(_1512_));
 sg13g2_a21o_1 _5384_ (.A2(net596),
    .A1(net571),
    .B1(_1512_),
    .X(_1513_));
 sg13g2_mux2_2 _5385_ (.A0(_0071_),
    .A1(_1512_),
    .S(_0666_),
    .X(_1514_));
 sg13g2_o21ai_1 _5386_ (.B1(_1513_),
    .Y(_1515_),
    .A1(_0071_),
    .A2(_0666_));
 sg13g2_nor2_1 _5387_ (.A(_0406_),
    .B(_1514_),
    .Y(_1516_));
 sg13g2_nand2_2 _5388_ (.Y(_1517_),
    .A(_0405_),
    .B(net568));
 sg13g2_nand2_1 _5389_ (.Y(_1518_),
    .A(_0405_),
    .B(_1483_));
 sg13g2_nor2_2 _5390_ (.A(_0396_),
    .B(_1514_),
    .Y(_1519_));
 sg13g2_nand2_2 _5391_ (.Y(_1520_),
    .A(net655),
    .B(net568));
 sg13g2_xnor2_1 _5392_ (.Y(_1521_),
    .A(_1518_),
    .B(_1519_));
 sg13g2_nand2b_1 _5393_ (.Y(_1522_),
    .B(_1521_),
    .A_N(_1511_));
 sg13g2_xnor2_1 _5394_ (.Y(_1523_),
    .A(_1511_),
    .B(_1521_));
 sg13g2_xnor2_1 _5395_ (.Y(_1524_),
    .A(_1510_),
    .B(_1523_));
 sg13g2_nor2b_1 _5396_ (.A(_1502_),
    .B_N(_1524_),
    .Y(_1525_));
 sg13g2_xnor2_1 _5397_ (.Y(_1526_),
    .A(_1502_),
    .B(_1524_));
 sg13g2_xor2_1 _5398_ (.B(_1526_),
    .A(_1501_),
    .X(_1527_));
 sg13g2_nand2_1 _5399_ (.Y(_1528_),
    .A(_1496_),
    .B(_1527_));
 sg13g2_a21oi_1 _5400_ (.A1(_1501_),
    .A2(_1526_),
    .Y(_1529_),
    .B1(_1525_));
 sg13g2_nand2_1 _5401_ (.Y(_1530_),
    .A(_1409_),
    .B(_1446_));
 sg13g2_o21ai_1 _5402_ (.B1(_1522_),
    .Y(_1531_),
    .A1(_1486_),
    .A2(_1517_));
 sg13g2_nand2b_1 _5403_ (.Y(_1532_),
    .B(_1531_),
    .A_N(_1530_));
 sg13g2_xor2_1 _5404_ (.B(_1531_),
    .A(_1530_),
    .X(_1533_));
 sg13g2_a21oi_2 _5405_ (.B1(_1508_),
    .Y(_1534_),
    .A2(_1523_),
    .A1(_1509_));
 sg13g2_o21ai_1 _5406_ (.B1(net598),
    .Y(_1535_),
    .A1(_1481_),
    .A2(_1482_));
 sg13g2_nor2_1 _5407_ (.A(_1504_),
    .B(_1535_),
    .Y(_1536_));
 sg13g2_xor2_1 _5408_ (.B(_1535_),
    .A(_1504_),
    .X(_1537_));
 sg13g2_xnor2_1 _5409_ (.Y(_1538_),
    .A(_1517_),
    .B(_1537_));
 sg13g2_and2_1 _5410_ (.A(_1506_),
    .B(_1538_),
    .X(_1539_));
 sg13g2_or2_1 _5411_ (.X(_1540_),
    .B(_1538_),
    .A(_1506_));
 sg13g2_xnor2_1 _5412_ (.Y(_1541_),
    .A(_1506_),
    .B(_1538_));
 sg13g2_nand2_1 _5413_ (.Y(_1542_),
    .A(_1425_),
    .B(net588));
 sg13g2_and2_1 _5414_ (.A(net581),
    .B(_1519_),
    .X(_1543_));
 sg13g2_nand2_1 _5415_ (.Y(_1544_),
    .A(_1434_),
    .B(net581));
 sg13g2_xnor2_1 _5416_ (.Y(_1545_),
    .A(_1519_),
    .B(_1544_));
 sg13g2_xnor2_1 _5417_ (.Y(_1546_),
    .A(_1542_),
    .B(_1545_));
 sg13g2_xnor2_1 _5418_ (.Y(_1547_),
    .A(_1541_),
    .B(_1546_));
 sg13g2_nand2b_1 _5419_ (.Y(_1548_),
    .B(_1547_),
    .A_N(_1534_));
 sg13g2_xnor2_1 _5420_ (.Y(_1549_),
    .A(_1534_),
    .B(_1547_));
 sg13g2_nand2b_1 _5421_ (.Y(_1550_),
    .B(_1549_),
    .A_N(_1533_));
 sg13g2_xnor2_1 _5422_ (.Y(_1551_),
    .A(_1533_),
    .B(_1549_));
 sg13g2_nor2b_1 _5423_ (.A(_1529_),
    .B_N(_1551_),
    .Y(_1552_));
 sg13g2_xnor2_1 _5424_ (.Y(_1553_),
    .A(_1529_),
    .B(_1551_));
 sg13g2_xnor2_1 _5425_ (.Y(_1554_),
    .A(_1500_),
    .B(_1553_));
 sg13g2_nor2_1 _5426_ (.A(_1528_),
    .B(_1554_),
    .Y(_1555_));
 sg13g2_xor2_1 _5427_ (.B(_1554_),
    .A(_1528_),
    .X(_1556_));
 sg13g2_xor2_1 _5428_ (.B(_1527_),
    .A(_1496_),
    .X(_1557_));
 sg13g2_inv_1 _5429_ (.Y(_1558_),
    .A(_1557_));
 sg13g2_o21ai_1 _5430_ (.B1(net598),
    .Y(_1559_),
    .A1(_1449_),
    .A2(_1450_));
 sg13g2_o21ai_1 _5431_ (.B1(net594),
    .Y(_1560_),
    .A1(_1449_),
    .A2(_1450_));
 sg13g2_or2_1 _5432_ (.X(_1561_),
    .B(_1559_),
    .A(_1418_));
 sg13g2_nand2_1 _5433_ (.Y(_1562_),
    .A(_0405_),
    .B(_1409_));
 sg13g2_and2_1 _5434_ (.A(_1416_),
    .B(_1560_),
    .X(_1563_));
 sg13g2_xor2_1 _5435_ (.B(_1560_),
    .A(_1416_),
    .X(_1564_));
 sg13g2_o21ai_1 _5436_ (.B1(_1561_),
    .Y(_1565_),
    .A1(_1562_),
    .A2(_1563_));
 sg13g2_xnor2_1 _5437_ (.Y(_1566_),
    .A(_1426_),
    .B(_1428_));
 sg13g2_and2_1 _5438_ (.A(_1565_),
    .B(_1566_),
    .X(_1567_));
 sg13g2_or2_1 _5439_ (.X(_1568_),
    .B(_1566_),
    .A(_1565_));
 sg13g2_xnor2_1 _5440_ (.Y(_1569_),
    .A(_1565_),
    .B(_1566_));
 sg13g2_xnor2_1 _5441_ (.Y(_1570_),
    .A(net686),
    .B(\generated._512[0] ));
 sg13g2_o21ai_1 _5442_ (.B1(_1570_),
    .Y(_1571_),
    .A1(net573),
    .A2(net597));
 sg13g2_nand3_1 _5443_ (.B(net571),
    .C(net596),
    .A(_0058_),
    .Y(_1572_));
 sg13g2_and2_2 _5444_ (.A(_1571_),
    .B(_1572_),
    .X(_1573_));
 sg13g2_nand2_1 _5445_ (.Y(_1574_),
    .A(net589),
    .B(_1573_));
 sg13g2_and4_1 _5446_ (.A(net655),
    .B(_1434_),
    .C(_1451_),
    .D(net582),
    .X(_1575_));
 sg13g2_a22oi_1 _5447_ (.Y(_1576_),
    .B1(_1451_),
    .B2(net581),
    .A2(_1434_),
    .A1(net655));
 sg13g2_nor2_1 _5448_ (.A(_1575_),
    .B(_1576_),
    .Y(_1577_));
 sg13g2_xnor2_1 _5449_ (.Y(_1578_),
    .A(_1574_),
    .B(_1577_));
 sg13g2_a21oi_2 _5450_ (.B1(_1567_),
    .Y(_1579_),
    .A2(_1578_),
    .A1(_1568_));
 sg13g2_xnor2_1 _5451_ (.Y(_1580_),
    .A(_1444_),
    .B(_1465_));
 sg13g2_nor2b_1 _5452_ (.A(_1579_),
    .B_N(_1580_),
    .Y(_1581_));
 sg13g2_nand2_1 _5453_ (.Y(_1582_),
    .A(net589),
    .B(_1576_));
 sg13g2_a21oi_1 _5454_ (.A1(_1573_),
    .A2(_1582_),
    .Y(_1583_),
    .B1(_1575_));
 sg13g2_inv_1 _5455_ (.Y(_1584_),
    .A(_1583_));
 sg13g2_xnor2_1 _5456_ (.Y(_1585_),
    .A(_1579_),
    .B(_1580_));
 sg13g2_a21oi_2 _5457_ (.B1(_1581_),
    .Y(_1586_),
    .A2(_1585_),
    .A1(_1584_));
 sg13g2_xnor2_1 _5458_ (.Y(_1587_),
    .A(_1493_),
    .B(_1495_));
 sg13g2_nand2b_1 _5459_ (.Y(_1588_),
    .B(_1587_),
    .A_N(_1586_));
 sg13g2_nand3_1 _5460_ (.B(_1571_),
    .C(_1572_),
    .A(net598),
    .Y(_1589_));
 sg13g2_nor2_1 _5461_ (.A(_0080_),
    .B(_0455_),
    .Y(_1590_));
 sg13g2_nand2b_1 _5462_ (.Y(_1591_),
    .B(_1590_),
    .A_N(_1589_));
 sg13g2_nand2_1 _5463_ (.Y(_1592_),
    .A(_0405_),
    .B(_1451_));
 sg13g2_a21oi_1 _5464_ (.A1(net600),
    .A2(_1573_),
    .Y(_1593_),
    .B1(_1590_));
 sg13g2_xnor2_1 _5465_ (.Y(_1594_),
    .A(_1589_),
    .B(_1590_));
 sg13g2_o21ai_1 _5466_ (.B1(_1591_),
    .Y(_1595_),
    .A1(_1592_),
    .A2(_1593_));
 sg13g2_nor2_1 _5467_ (.A(_0406_),
    .B(_1415_),
    .Y(_1596_));
 sg13g2_nand3_1 _5468_ (.B(_1571_),
    .C(_1572_),
    .A(net594),
    .Y(_1597_));
 sg13g2_nor2_1 _5469_ (.A(_1560_),
    .B(_1589_),
    .Y(_1598_));
 sg13g2_xor2_1 _5470_ (.B(_1597_),
    .A(_1559_),
    .X(_1599_));
 sg13g2_xor2_1 _5471_ (.B(_1599_),
    .A(_1596_),
    .X(_1600_));
 sg13g2_nand2_1 _5472_ (.Y(_1601_),
    .A(_1595_),
    .B(_1600_));
 sg13g2_xnor2_1 _5473_ (.Y(_1602_),
    .A(_1595_),
    .B(_1600_));
 sg13g2_nand2_1 _5474_ (.Y(_1603_),
    .A(\generated._64[0] ),
    .B(net582));
 sg13g2_or2_1 _5475_ (.X(_1604_),
    .B(_1603_),
    .A(_1478_));
 sg13g2_xnor2_1 _5476_ (.Y(_1605_),
    .A(_1478_),
    .B(_1603_));
 sg13g2_nor2_1 _5477_ (.A(_1602_),
    .B(_1605_),
    .Y(_1606_));
 sg13g2_o21ai_1 _5478_ (.B1(_1601_),
    .Y(_1607_),
    .A1(_1602_),
    .A2(_1605_));
 sg13g2_a21o_1 _5479_ (.A2(_1599_),
    .A1(_1596_),
    .B1(_1598_),
    .X(_1608_));
 sg13g2_xnor2_1 _5480_ (.Y(_1609_),
    .A(_1562_),
    .B(_1564_));
 sg13g2_nand2_1 _5481_ (.Y(_1610_),
    .A(_1608_),
    .B(_1609_));
 sg13g2_xnor2_1 _5482_ (.Y(_1611_),
    .A(_1608_),
    .B(_1609_));
 sg13g2_nand2_1 _5483_ (.Y(_1612_),
    .A(\generated._64[0] ),
    .B(net589));
 sg13g2_and4_1 _5484_ (.A(_0395_),
    .B(_1425_),
    .C(net582),
    .D(_1573_),
    .X(_1613_));
 sg13g2_a22oi_1 _5485_ (.Y(_1614_),
    .B1(net582),
    .B2(_1573_),
    .A2(_1425_),
    .A1(net655));
 sg13g2_nor2_1 _5486_ (.A(_1613_),
    .B(_1614_),
    .Y(_1615_));
 sg13g2_xor2_1 _5487_ (.B(_1615_),
    .A(_1612_),
    .X(_1616_));
 sg13g2_xnor2_1 _5488_ (.Y(_1617_),
    .A(_1611_),
    .B(_1616_));
 sg13g2_nand2b_1 _5489_ (.Y(_1618_),
    .B(_1607_),
    .A_N(_1617_));
 sg13g2_nand2_1 _5490_ (.Y(_1619_),
    .A(net589),
    .B(_1614_));
 sg13g2_a21oi_1 _5491_ (.A1(\generated._64[0] ),
    .A2(_1619_),
    .Y(_1620_),
    .B1(_1613_));
 sg13g2_o21ai_1 _5492_ (.B1(_1610_),
    .Y(_1621_),
    .A1(_1611_),
    .A2(_1616_));
 sg13g2_xnor2_1 _5493_ (.Y(_1622_),
    .A(_1569_),
    .B(_1578_));
 sg13g2_nand2_1 _5494_ (.Y(_1623_),
    .A(_1621_),
    .B(_1622_));
 sg13g2_xnor2_1 _5495_ (.Y(_1624_),
    .A(_1621_),
    .B(_1622_));
 sg13g2_xnor2_1 _5496_ (.Y(_1625_),
    .A(_1620_),
    .B(_1624_));
 sg13g2_xor2_1 _5497_ (.B(_1617_),
    .A(_1607_),
    .X(_1626_));
 sg13g2_and2_1 _5498_ (.A(_1602_),
    .B(_1605_),
    .X(_1627_));
 sg13g2_and4_1 _5499_ (.A(net686),
    .B(_0405_),
    .C(net600),
    .D(_1573_),
    .X(_1628_));
 sg13g2_xnor2_1 _5500_ (.Y(_1629_),
    .A(_1592_),
    .B(_1594_));
 sg13g2_or2_1 _5501_ (.X(_1630_),
    .B(_1629_),
    .A(_1628_));
 sg13g2_a22oi_1 _5502_ (.Y(_1631_),
    .B1(_1573_),
    .B2(_0405_),
    .A2(net600),
    .A1(net686));
 sg13g2_a21oi_1 _5503_ (.A1(net686),
    .A2(net599),
    .Y(_1632_),
    .B1(_0080_));
 sg13g2_o21ai_1 _5504_ (.B1(net655),
    .Y(_1633_),
    .A1(_1451_),
    .A2(_1632_));
 sg13g2_nor2_1 _5505_ (.A(_1631_),
    .B(_1633_),
    .Y(_1634_));
 sg13g2_nand2_1 _5506_ (.Y(_1635_),
    .A(_0080_),
    .B(_1628_));
 sg13g2_a21o_1 _5507_ (.A2(_1635_),
    .A1(_1634_),
    .B1(_1461_),
    .X(_1636_));
 sg13g2_and2_1 _5508_ (.A(_1628_),
    .B(_1629_),
    .X(_1637_));
 sg13g2_a221oi_1 _5509_ (.B2(_1630_),
    .C1(_1637_),
    .B1(_1636_),
    .A1(_1414_),
    .Y(_1638_),
    .A2(_1634_));
 sg13g2_or3_1 _5510_ (.A(_1606_),
    .B(_1627_),
    .C(_1638_),
    .X(_1639_));
 sg13g2_nand4_1 _5511_ (.B(_1634_),
    .C(_1635_),
    .A(_1461_),
    .Y(_1640_),
    .D(_1637_));
 sg13g2_a22oi_1 _5512_ (.Y(_1641_),
    .B1(_1639_),
    .B2(_1640_),
    .A2(_1626_),
    .A1(_1604_));
 sg13g2_o21ai_1 _5513_ (.B1(_1623_),
    .Y(_1642_),
    .A1(_1620_),
    .A2(_1624_));
 sg13g2_xnor2_1 _5514_ (.Y(_1643_),
    .A(_1583_),
    .B(_1585_));
 sg13g2_and2_1 _5515_ (.A(_1642_),
    .B(_1643_),
    .X(_1644_));
 sg13g2_or2_1 _5516_ (.X(_1645_),
    .B(_1626_),
    .A(_1604_));
 sg13g2_or2_1 _5517_ (.X(_1646_),
    .B(_1643_),
    .A(_1642_));
 sg13g2_nand2b_1 _5518_ (.Y(_1647_),
    .B(_1586_),
    .A_N(_1587_));
 sg13g2_nor2_1 _5519_ (.A(_1558_),
    .B(_1588_),
    .Y(_1648_));
 sg13g2_xnor2_1 _5520_ (.Y(_1649_),
    .A(_1586_),
    .B(_1587_));
 sg13g2_nand4_1 _5521_ (.B(_1588_),
    .C(_1646_),
    .A(_1557_),
    .Y(_1650_),
    .D(_1647_));
 sg13g2_a21oi_1 _5522_ (.A1(_1618_),
    .A2(_1645_),
    .Y(_1651_),
    .B1(_1625_));
 sg13g2_nand2_1 _5523_ (.Y(_1652_),
    .A(_1618_),
    .B(_1625_));
 sg13g2_and2_1 _5524_ (.A(_1641_),
    .B(_1645_),
    .X(_1653_));
 sg13g2_a221oi_1 _5525_ (.B2(_1653_),
    .C1(_1651_),
    .B1(_1652_),
    .A1(_1644_),
    .Y(_1654_),
    .A2(_1649_));
 sg13g2_nor2_1 _5526_ (.A(_1650_),
    .B(_1654_),
    .Y(_1655_));
 sg13g2_o21ai_1 _5527_ (.B1(_1556_),
    .Y(_1656_),
    .A1(_1648_),
    .A2(_1655_));
 sg13g2_or3_1 _5528_ (.A(_1556_),
    .B(_1648_),
    .C(_1655_),
    .X(_1657_));
 sg13g2_and2_1 _5529_ (.A(_1656_),
    .B(_1657_),
    .X(_1658_));
 sg13g2_and2_1 _5530_ (.A(_0458_),
    .B(_0556_),
    .X(_1659_));
 sg13g2_nor2_1 _5531_ (.A(_0462_),
    .B(_1659_),
    .Y(_1660_));
 sg13g2_a21oi_2 _5532_ (.B1(_1660_),
    .Y(_1661_),
    .A2(_1659_),
    .A1(_2835_));
 sg13g2_inv_1 _5533_ (.Y(_1662_),
    .A(net576));
 sg13g2_nor3_2 _5534_ (.A(net700),
    .B(\generated._562[1] ),
    .C(\generated._562[2] ),
    .Y(_1663_));
 sg13g2_nand2b_2 _5535_ (.Y(_1664_),
    .B(_1663_),
    .A_N(\generated._562[3] ));
 sg13g2_xor2_1 _5536_ (.B(_1663_),
    .A(\generated._562[3] ),
    .X(_1665_));
 sg13g2_o21ai_1 _5537_ (.B1(_0064_),
    .Y(_1666_),
    .A1(_0609_),
    .A2(net574));
 sg13g2_nand3_1 _5538_ (.B(net572),
    .C(_1665_),
    .A(_0610_),
    .Y(_1667_));
 sg13g2_and2_1 _5539_ (.A(_1666_),
    .B(_1667_),
    .X(_1668_));
 sg13g2_a21o_2 _5540_ (.A2(_1659_),
    .A1(_2835_),
    .B1(_0327_),
    .X(_1669_));
 sg13g2_inv_1 _5541_ (.Y(_1670_),
    .A(net578));
 sg13g2_o21ai_1 _5542_ (.B1(\generated._562[2] ),
    .Y(_1671_),
    .A1(net700),
    .A2(\generated._562[1] ));
 sg13g2_nand2b_1 _5543_ (.Y(_1672_),
    .B(_1671_),
    .A_N(_1663_));
 sg13g2_o21ai_1 _5544_ (.B1(_0061_),
    .Y(_1673_),
    .A1(_0609_),
    .A2(net574));
 sg13g2_nand3_1 _5545_ (.B(net572),
    .C(_1672_),
    .A(_0610_),
    .Y(_1674_));
 sg13g2_and2_1 _5546_ (.A(_1673_),
    .B(_1674_),
    .X(_1675_));
 sg13g2_a22oi_1 _5547_ (.Y(_1676_),
    .B1(net578),
    .B2(_1675_),
    .A2(_1668_),
    .A1(net576));
 sg13g2_xnor2_1 _5548_ (.Y(_1677_),
    .A(\generated._562[4] ),
    .B(_1664_));
 sg13g2_o21ai_1 _5549_ (.B1(_0066_),
    .Y(_1678_),
    .A1(_0609_),
    .A2(net574));
 sg13g2_nand3_1 _5550_ (.B(net572),
    .C(_1677_),
    .A(_0610_),
    .Y(_1679_));
 sg13g2_nand2_1 _5551_ (.Y(_1680_),
    .A(_1678_),
    .B(_1679_));
 sg13g2_and2_1 _5552_ (.A(_1678_),
    .B(_1679_),
    .X(_1681_));
 sg13g2_xnor2_1 _5553_ (.Y(_1682_),
    .A(_0459_),
    .B(_0556_));
 sg13g2_nand3_1 _5554_ (.B(_1679_),
    .C(net580),
    .A(_1678_),
    .Y(_1683_));
 sg13g2_nand3_1 _5555_ (.B(_1666_),
    .C(_1667_),
    .A(net591),
    .Y(_1684_));
 sg13g2_nand3_1 _5556_ (.B(_1678_),
    .C(_1679_),
    .A(net591),
    .Y(_1685_));
 sg13g2_nand3_1 _5557_ (.B(_1667_),
    .C(net580),
    .A(_1666_),
    .Y(_1686_));
 sg13g2_or2_1 _5558_ (.X(_1687_),
    .B(_1684_),
    .A(_1683_));
 sg13g2_nor3_2 _5559_ (.A(\generated._562[4] ),
    .B(\generated._562[5] ),
    .C(_1664_),
    .Y(_1688_));
 sg13g2_o21ai_1 _5560_ (.B1(\generated._562[5] ),
    .Y(_1689_),
    .A1(\generated._562[4] ),
    .A2(_1664_));
 sg13g2_nand2b_1 _5561_ (.Y(_1690_),
    .B(_1689_),
    .A_N(_1688_));
 sg13g2_o21ai_1 _5562_ (.B1(_0068_),
    .Y(_1691_),
    .A1(_0609_),
    .A2(net574));
 sg13g2_nand3_1 _5563_ (.B(net572),
    .C(_1690_),
    .A(_0610_),
    .Y(_1692_));
 sg13g2_nand2_2 _5564_ (.Y(_1693_),
    .A(_1691_),
    .B(_1692_));
 sg13g2_nand3_1 _5565_ (.B(_1691_),
    .C(_1692_),
    .A(net725),
    .Y(_1694_));
 sg13g2_xnor2_1 _5566_ (.Y(_1695_),
    .A(_1685_),
    .B(_1686_));
 sg13g2_o21ai_1 _5567_ (.B1(_1687_),
    .Y(_1696_),
    .A1(_1694_),
    .A2(_1695_));
 sg13g2_nor2b_1 _5568_ (.A(\generated._562[6] ),
    .B_N(_1688_),
    .Y(_1697_));
 sg13g2_xor2_1 _5569_ (.B(_1688_),
    .A(\generated._562[6] ),
    .X(_1698_));
 sg13g2_o21ai_1 _5570_ (.B1(_0070_),
    .Y(_1699_),
    .A1(_0609_),
    .A2(net574));
 sg13g2_nand3_1 _5571_ (.B(net572),
    .C(_1698_),
    .A(_0610_),
    .Y(_1700_));
 sg13g2_and2_1 _5572_ (.A(_1699_),
    .B(_1700_),
    .X(_1701_));
 sg13g2_nand2_1 _5573_ (.Y(_1702_),
    .A(net725),
    .B(_1701_));
 sg13g2_nand3_1 _5574_ (.B(_1691_),
    .C(_1692_),
    .A(net580),
    .Y(_1703_));
 sg13g2_nand3_1 _5575_ (.B(_1691_),
    .C(_1692_),
    .A(net591),
    .Y(_1704_));
 sg13g2_or2_1 _5576_ (.X(_1705_),
    .B(_1703_),
    .A(_1685_));
 sg13g2_and2_1 _5577_ (.A(_1683_),
    .B(_1704_),
    .X(_1706_));
 sg13g2_xor2_1 _5578_ (.B(_1704_),
    .A(_1683_),
    .X(_1707_));
 sg13g2_xnor2_1 _5579_ (.Y(_1708_),
    .A(_1702_),
    .B(_1707_));
 sg13g2_nand2_1 _5580_ (.Y(_1709_),
    .A(_1696_),
    .B(_1708_));
 sg13g2_xnor2_1 _5581_ (.Y(_1710_),
    .A(_1696_),
    .B(_1708_));
 sg13g2_or2_1 _5582_ (.X(_1711_),
    .B(_1710_),
    .A(_1676_));
 sg13g2_a22oi_1 _5583_ (.Y(_1712_),
    .B1(_1681_),
    .B2(net576),
    .A2(net578),
    .A1(_1668_));
 sg13g2_o21ai_1 _5584_ (.B1(_1705_),
    .Y(_1713_),
    .A1(_1702_),
    .A2(_1706_));
 sg13g2_nand2b_1 _5585_ (.Y(_1714_),
    .B(_1697_),
    .A_N(\generated._562[7] ));
 sg13g2_xor2_1 _5586_ (.B(_1697_),
    .A(\generated._562[7] ),
    .X(_1715_));
 sg13g2_nand3_1 _5587_ (.B(net572),
    .C(_1715_),
    .A(_0610_),
    .Y(_1716_));
 sg13g2_o21ai_1 _5588_ (.B1(_0072_),
    .Y(_1717_),
    .A1(_0609_),
    .A2(net574));
 sg13g2_nand2_2 _5589_ (.Y(_1718_),
    .A(_1716_),
    .B(_1717_));
 sg13g2_inv_1 _5590_ (.Y(_1719_),
    .A(_1718_));
 sg13g2_nand3_1 _5591_ (.B(_1716_),
    .C(_1717_),
    .A(net725),
    .Y(_1720_));
 sg13g2_nand3_1 _5592_ (.B(_1699_),
    .C(_1700_),
    .A(net580),
    .Y(_1721_));
 sg13g2_nand3_1 _5593_ (.B(_1699_),
    .C(_1700_),
    .A(net592),
    .Y(_1722_));
 sg13g2_or2_1 _5594_ (.X(_1723_),
    .B(_1721_),
    .A(_1704_));
 sg13g2_and2_1 _5595_ (.A(_1703_),
    .B(_1722_),
    .X(_1724_));
 sg13g2_xor2_1 _5596_ (.B(_1722_),
    .A(_1703_),
    .X(_1725_));
 sg13g2_xnor2_1 _5597_ (.Y(_1726_),
    .A(_1720_),
    .B(_1725_));
 sg13g2_nand2_1 _5598_ (.Y(_1727_),
    .A(_1713_),
    .B(_1726_));
 sg13g2_xnor2_1 _5599_ (.Y(_1728_),
    .A(_1713_),
    .B(_1726_));
 sg13g2_or2_1 _5600_ (.X(_1729_),
    .B(_1728_),
    .A(_1712_));
 sg13g2_xnor2_1 _5601_ (.Y(_1730_),
    .A(_1712_),
    .B(_1728_));
 sg13g2_nor2_1 _5602_ (.A(_1711_),
    .B(_1730_),
    .Y(_1731_));
 sg13g2_nor2_1 _5603_ (.A(\generated._562[8] ),
    .B(_1714_),
    .Y(_1732_));
 sg13g2_xor2_1 _5604_ (.B(_1714_),
    .A(\generated._562[8] ),
    .X(_1733_));
 sg13g2_mux2_2 _5605_ (.A0(_2862_),
    .A1(_1733_),
    .S(net569),
    .X(_1734_));
 sg13g2_and2_1 _5606_ (.A(_2836_),
    .B(_1734_),
    .X(_1735_));
 sg13g2_nand3_1 _5607_ (.B(_1708_),
    .C(_1735_),
    .A(_1696_),
    .Y(_1736_));
 sg13g2_xnor2_1 _5608_ (.Y(_1737_),
    .A(_1709_),
    .B(_1735_));
 sg13g2_xor2_1 _5609_ (.B(_1730_),
    .A(_1711_),
    .X(_1738_));
 sg13g2_a21oi_1 _5610_ (.A1(_1737_),
    .A2(_1738_),
    .Y(_1739_),
    .B1(_1731_));
 sg13g2_xnor2_1 _5611_ (.Y(_1740_),
    .A(\generated._562[9] ),
    .B(_1732_));
 sg13g2_nor2_1 _5612_ (.A(_0640_),
    .B(_1740_),
    .Y(_1741_));
 sg13g2_a21oi_2 _5613_ (.B1(_1741_),
    .Y(_1742_),
    .A2(_0640_),
    .A1(_0074_));
 sg13g2_and2_2 _5614_ (.A(_2836_),
    .B(net567),
    .X(_1743_));
 sg13g2_nand2_2 _5615_ (.Y(_1744_),
    .A(_2836_),
    .B(net567));
 sg13g2_nand3_1 _5616_ (.B(_1726_),
    .C(_1743_),
    .A(_1713_),
    .Y(_1745_));
 sg13g2_xnor2_1 _5617_ (.Y(_1746_),
    .A(_1727_),
    .B(_1743_));
 sg13g2_nand2_1 _5618_ (.Y(_1747_),
    .A(net578),
    .B(_1681_));
 sg13g2_o21ai_1 _5619_ (.B1(_1747_),
    .Y(_1748_),
    .A1(_1662_),
    .A2(_1693_));
 sg13g2_o21ai_1 _5620_ (.B1(_1723_),
    .Y(_1749_),
    .A1(_1720_),
    .A2(_1724_));
 sg13g2_and2_1 _5621_ (.A(net726),
    .B(_1734_),
    .X(_1750_));
 sg13g2_nor2b_1 _5622_ (.A(_1718_),
    .B_N(_1682_),
    .Y(_1751_));
 sg13g2_nand3_1 _5623_ (.B(_1716_),
    .C(_1717_),
    .A(net592),
    .Y(_1752_));
 sg13g2_nor2_1 _5624_ (.A(_1721_),
    .B(_1752_),
    .Y(_1753_));
 sg13g2_xor2_1 _5625_ (.B(_1752_),
    .A(_1721_),
    .X(_1754_));
 sg13g2_xor2_1 _5626_ (.B(_1754_),
    .A(_1750_),
    .X(_1755_));
 sg13g2_nand2_1 _5627_ (.Y(_1756_),
    .A(_1749_),
    .B(_1755_));
 sg13g2_xnor2_1 _5628_ (.Y(_1757_),
    .A(_1749_),
    .B(_1755_));
 sg13g2_nand2b_1 _5629_ (.Y(_1758_),
    .B(_1748_),
    .A_N(_1757_));
 sg13g2_xor2_1 _5630_ (.B(_1757_),
    .A(_1748_),
    .X(_1759_));
 sg13g2_nor2_1 _5631_ (.A(_1729_),
    .B(_1759_),
    .Y(_1760_));
 sg13g2_xor2_1 _5632_ (.B(_1759_),
    .A(_1729_),
    .X(_1761_));
 sg13g2_xnor2_1 _5633_ (.Y(_1762_),
    .A(_1746_),
    .B(_1761_));
 sg13g2_xor2_1 _5634_ (.B(_1762_),
    .A(_1739_),
    .X(_1763_));
 sg13g2_nand2b_1 _5635_ (.Y(_1764_),
    .B(_1763_),
    .A_N(_1736_));
 sg13g2_o21ai_1 _5636_ (.B1(_1764_),
    .Y(_1765_),
    .A1(_1739_),
    .A2(_1762_));
 sg13g2_a21oi_1 _5637_ (.A1(_1746_),
    .A2(_1761_),
    .Y(_1766_),
    .B1(_1760_));
 sg13g2_nand3_1 _5638_ (.B(_1749_),
    .C(_1755_),
    .A(_1743_),
    .Y(_1767_));
 sg13g2_xnor2_1 _5639_ (.Y(_1768_),
    .A(_1744_),
    .B(_1756_));
 sg13g2_inv_1 _5640_ (.Y(_1769_),
    .A(_1768_));
 sg13g2_nand2_1 _5641_ (.Y(_1770_),
    .A(net576),
    .B(_1701_));
 sg13g2_o21ai_1 _5642_ (.B1(_1770_),
    .Y(_1771_),
    .A1(_1670_),
    .A2(_1693_));
 sg13g2_a21oi_1 _5643_ (.A1(_1750_),
    .A2(_1754_),
    .Y(_1772_),
    .B1(_1753_));
 sg13g2_nand2_2 _5644_ (.Y(_1773_),
    .A(net726),
    .B(net567));
 sg13g2_inv_1 _5645_ (.Y(_1774_),
    .A(_1773_));
 sg13g2_nand2_1 _5646_ (.Y(_1775_),
    .A(_1682_),
    .B(_1734_));
 sg13g2_nand2_1 _5647_ (.Y(_1776_),
    .A(net592),
    .B(_1734_));
 sg13g2_nor2_1 _5648_ (.A(_1752_),
    .B(_1775_),
    .Y(_1777_));
 sg13g2_xnor2_1 _5649_ (.Y(_1778_),
    .A(_1751_),
    .B(_1776_));
 sg13g2_xnor2_1 _5650_ (.Y(_1779_),
    .A(_1773_),
    .B(_1778_));
 sg13g2_nand2b_2 _5651_ (.Y(_1780_),
    .B(_1779_),
    .A_N(_1772_));
 sg13g2_xor2_1 _5652_ (.B(_1779_),
    .A(_1772_),
    .X(_1781_));
 sg13g2_nand2b_1 _5653_ (.Y(_1782_),
    .B(_1771_),
    .A_N(_1781_));
 sg13g2_xor2_1 _5654_ (.B(_1781_),
    .A(_1771_),
    .X(_1783_));
 sg13g2_nor2_1 _5655_ (.A(_1758_),
    .B(_1783_),
    .Y(_1784_));
 sg13g2_xor2_1 _5656_ (.B(_1783_),
    .A(_1758_),
    .X(_1785_));
 sg13g2_xnor2_1 _5657_ (.Y(_1786_),
    .A(_1768_),
    .B(_1785_));
 sg13g2_inv_1 _5658_ (.Y(_1787_),
    .A(_1786_));
 sg13g2_xnor2_1 _5659_ (.Y(_1788_),
    .A(_1766_),
    .B(_1786_));
 sg13g2_nand2b_1 _5660_ (.Y(_1789_),
    .B(_1788_),
    .A_N(_1745_));
 sg13g2_xor2_1 _5661_ (.B(_1788_),
    .A(_1745_),
    .X(_1790_));
 sg13g2_nor2b_1 _5662_ (.A(_1790_),
    .B_N(_1765_),
    .Y(_1791_));
 sg13g2_xor2_1 _5663_ (.B(_1790_),
    .A(_1765_),
    .X(_1792_));
 sg13g2_xnor2_1 _5664_ (.Y(_1793_),
    .A(net700),
    .B(\generated._562[1] ));
 sg13g2_o21ai_1 _5665_ (.B1(_0057_),
    .Y(_1794_),
    .A1(_0609_),
    .A2(net574));
 sg13g2_nand3_1 _5666_ (.B(net572),
    .C(_1793_),
    .A(_0610_),
    .Y(_1795_));
 sg13g2_and2_2 _5667_ (.A(_1794_),
    .B(_1795_),
    .X(_1796_));
 sg13g2_a22oi_1 _5668_ (.Y(_1797_),
    .B1(_1796_),
    .B2(net576),
    .A2(net578),
    .A1(net700));
 sg13g2_nand3_1 _5669_ (.B(_1674_),
    .C(net580),
    .A(_1673_),
    .Y(_1798_));
 sg13g2_nand3_1 _5670_ (.B(_1673_),
    .C(_1674_),
    .A(net591),
    .Y(_1799_));
 sg13g2_nand3_1 _5671_ (.B(_1794_),
    .C(_1795_),
    .A(net580),
    .Y(_1800_));
 sg13g2_or2_1 _5672_ (.X(_1801_),
    .B(_1800_),
    .A(_1799_));
 sg13g2_nand2_1 _5673_ (.Y(_1802_),
    .A(net725),
    .B(_1668_));
 sg13g2_and2_1 _5674_ (.A(_1799_),
    .B(_1800_),
    .X(_1803_));
 sg13g2_xor2_1 _5675_ (.B(_1800_),
    .A(_1799_),
    .X(_1804_));
 sg13g2_o21ai_1 _5676_ (.B1(_1801_),
    .Y(_1805_),
    .A1(_1802_),
    .A2(_1803_));
 sg13g2_and2_1 _5677_ (.A(net725),
    .B(_1681_),
    .X(_1806_));
 sg13g2_nor2_1 _5678_ (.A(_1686_),
    .B(_1799_),
    .Y(_1807_));
 sg13g2_xor2_1 _5679_ (.B(_1798_),
    .A(_1684_),
    .X(_1808_));
 sg13g2_xor2_1 _5680_ (.B(_1808_),
    .A(_1806_),
    .X(_1809_));
 sg13g2_xnor2_1 _5681_ (.Y(_1810_),
    .A(_1805_),
    .B(_1809_));
 sg13g2_or2_1 _5682_ (.X(_1811_),
    .B(_1810_),
    .A(_1797_));
 sg13g2_xnor2_1 _5683_ (.Y(_1812_),
    .A(_1797_),
    .B(_1810_));
 sg13g2_nand2_1 _5684_ (.Y(_1813_),
    .A(\generated._562[0] ),
    .B(net576));
 sg13g2_nor2b_1 _5685_ (.A(_0079_),
    .B_N(net580),
    .Y(_1814_));
 sg13g2_and3_1 _5686_ (.X(_1815_),
    .A(net591),
    .B(_1796_),
    .C(_1814_));
 sg13g2_nand3_1 _5687_ (.B(_1796_),
    .C(_1814_),
    .A(net592),
    .Y(_1816_));
 sg13g2_nand2_1 _5688_ (.Y(_1817_),
    .A(net725),
    .B(_1675_));
 sg13g2_a21oi_1 _5689_ (.A1(net591),
    .A2(_1796_),
    .Y(_1818_),
    .B1(_1814_));
 sg13g2_nor2_1 _5690_ (.A(_1815_),
    .B(_1818_),
    .Y(_1819_));
 sg13g2_o21ai_1 _5691_ (.B1(_1816_),
    .Y(_1820_),
    .A1(_1817_),
    .A2(_1818_));
 sg13g2_xnor2_1 _5692_ (.Y(_1821_),
    .A(_1802_),
    .B(_1804_));
 sg13g2_xnor2_1 _5693_ (.Y(_1822_),
    .A(_1820_),
    .B(_1821_));
 sg13g2_nor2_1 _5694_ (.A(_1813_),
    .B(_1822_),
    .Y(_1823_));
 sg13g2_nor2b_1 _5695_ (.A(_1812_),
    .B_N(_1823_),
    .Y(_1824_));
 sg13g2_nor2_1 _5696_ (.A(net727),
    .B(_1693_),
    .Y(_1825_));
 sg13g2_nand3_1 _5697_ (.B(_1821_),
    .C(_1825_),
    .A(_1820_),
    .Y(_1826_));
 sg13g2_inv_1 _5698_ (.Y(_1827_),
    .A(_1826_));
 sg13g2_a21oi_1 _5699_ (.A1(_1820_),
    .A2(_1821_),
    .Y(_1828_),
    .B1(_1825_));
 sg13g2_nor2_1 _5700_ (.A(_1827_),
    .B(_1828_),
    .Y(_1829_));
 sg13g2_xnor2_1 _5701_ (.Y(_1830_),
    .A(_1812_),
    .B(_1823_));
 sg13g2_a21oi_1 _5702_ (.A1(_1829_),
    .A2(_1830_),
    .Y(_1831_),
    .B1(_1824_));
 sg13g2_and2_1 _5703_ (.A(_2836_),
    .B(_1701_),
    .X(_1832_));
 sg13g2_nand3_1 _5704_ (.B(_1809_),
    .C(_1832_),
    .A(_1805_),
    .Y(_1833_));
 sg13g2_inv_1 _5705_ (.Y(_1834_),
    .A(_1833_));
 sg13g2_a21oi_1 _5706_ (.A1(_1805_),
    .A2(_1809_),
    .Y(_1835_),
    .B1(_1832_));
 sg13g2_nor2_1 _5707_ (.A(_1834_),
    .B(_1835_),
    .Y(_1836_));
 sg13g2_a22oi_1 _5708_ (.Y(_1837_),
    .B1(_1796_),
    .B2(net578),
    .A2(_1675_),
    .A1(net576));
 sg13g2_a21o_1 _5709_ (.A2(_1808_),
    .A1(_1806_),
    .B1(_1807_),
    .X(_1838_));
 sg13g2_xor2_1 _5710_ (.B(_1695_),
    .A(_1694_),
    .X(_1839_));
 sg13g2_nand2_1 _5711_ (.Y(_1840_),
    .A(_1838_),
    .B(_1839_));
 sg13g2_xnor2_1 _5712_ (.Y(_1841_),
    .A(_1838_),
    .B(_1839_));
 sg13g2_or2_1 _5713_ (.X(_1842_),
    .B(_1841_),
    .A(_1837_));
 sg13g2_xnor2_1 _5714_ (.Y(_1843_),
    .A(_1837_),
    .B(_1841_));
 sg13g2_nor2_1 _5715_ (.A(_1811_),
    .B(_1843_),
    .Y(_1844_));
 sg13g2_xor2_1 _5716_ (.B(_1843_),
    .A(_1811_),
    .X(_1845_));
 sg13g2_xnor2_1 _5717_ (.Y(_1846_),
    .A(_1836_),
    .B(_1845_));
 sg13g2_nor2_1 _5718_ (.A(_1831_),
    .B(_1846_),
    .Y(_1847_));
 sg13g2_xor2_1 _5719_ (.B(_1846_),
    .A(_1831_),
    .X(_1848_));
 sg13g2_a21oi_1 _5720_ (.A1(_1827_),
    .A2(_1848_),
    .Y(_1849_),
    .B1(_1847_));
 sg13g2_a21oi_1 _5721_ (.A1(_1836_),
    .A2(_1845_),
    .Y(_1850_),
    .B1(_1844_));
 sg13g2_nor2_1 _5722_ (.A(net727),
    .B(_1718_),
    .Y(_1851_));
 sg13g2_nand3_1 _5723_ (.B(_1839_),
    .C(_1851_),
    .A(_1838_),
    .Y(_1852_));
 sg13g2_xnor2_1 _5724_ (.Y(_1853_),
    .A(_1840_),
    .B(_1851_));
 sg13g2_xnor2_1 _5725_ (.Y(_1854_),
    .A(_1676_),
    .B(_1710_));
 sg13g2_nor2_1 _5726_ (.A(_1842_),
    .B(_1854_),
    .Y(_1855_));
 sg13g2_xor2_1 _5727_ (.B(_1854_),
    .A(_1842_),
    .X(_1856_));
 sg13g2_xnor2_1 _5728_ (.Y(_1857_),
    .A(_1853_),
    .B(_1856_));
 sg13g2_nor2_1 _5729_ (.A(_1850_),
    .B(_1857_),
    .Y(_1858_));
 sg13g2_xor2_1 _5730_ (.B(_1857_),
    .A(_1850_),
    .X(_1859_));
 sg13g2_xnor2_1 _5731_ (.Y(_1860_),
    .A(_1834_),
    .B(_1859_));
 sg13g2_nor2_1 _5732_ (.A(_1849_),
    .B(_1860_),
    .Y(_1861_));
 sg13g2_nor2_1 _5733_ (.A(net727),
    .B(_1680_),
    .Y(_1862_));
 sg13g2_and4_1 _5734_ (.A(net725),
    .B(\generated._562[0] ),
    .C(net592),
    .D(_1796_),
    .X(_1863_));
 sg13g2_xnor2_1 _5735_ (.Y(_1864_),
    .A(_1817_),
    .B(_1819_));
 sg13g2_nand2_1 _5736_ (.Y(_1865_),
    .A(_1863_),
    .B(_1864_));
 sg13g2_nor3_1 _5737_ (.A(net727),
    .B(_1680_),
    .C(_1865_),
    .Y(_1866_));
 sg13g2_xor2_1 _5738_ (.B(_1830_),
    .A(_1829_),
    .X(_1867_));
 sg13g2_xnor2_1 _5739_ (.Y(_1868_),
    .A(_1862_),
    .B(_1865_));
 sg13g2_xor2_1 _5740_ (.B(_1822_),
    .A(_1813_),
    .X(_1869_));
 sg13g2_nor2_1 _5741_ (.A(_1868_),
    .B(_1869_),
    .Y(_1870_));
 sg13g2_a22oi_1 _5742_ (.Y(_1871_),
    .B1(_1796_),
    .B2(net725),
    .A2(net591),
    .A1(net700));
 sg13g2_a21oi_1 _5743_ (.A1(\generated._562[0] ),
    .A2(net591),
    .Y(_1872_),
    .B1(_0079_));
 sg13g2_o21ai_1 _5744_ (.B1(_2836_),
    .Y(_1873_),
    .A1(_1675_),
    .A2(_1872_));
 sg13g2_or2_1 _5745_ (.X(_1874_),
    .B(_1873_),
    .A(_1871_));
 sg13g2_a21o_1 _5746_ (.A2(_1863_),
    .A1(_0079_),
    .B1(_1874_),
    .X(_1875_));
 sg13g2_nand2_1 _5747_ (.Y(_1876_),
    .A(_2836_),
    .B(_1668_));
 sg13g2_nor2_1 _5748_ (.A(_1875_),
    .B(_1876_),
    .Y(_1877_));
 sg13g2_nor2_1 _5749_ (.A(_1863_),
    .B(_1864_),
    .Y(_1878_));
 sg13g2_a21oi_1 _5750_ (.A1(_1875_),
    .A2(_1876_),
    .Y(_1879_),
    .B1(_1878_));
 sg13g2_a221oi_1 _5751_ (.B2(_1865_),
    .C1(_1877_),
    .B1(_1879_),
    .A1(_1868_),
    .Y(_1880_),
    .A2(_1869_));
 sg13g2_nor2_1 _5752_ (.A(_1870_),
    .B(_1880_),
    .Y(_1881_));
 sg13g2_o21ai_1 _5753_ (.B1(_1866_),
    .Y(_1882_),
    .A1(_1867_),
    .A2(_1881_));
 sg13g2_nand2_1 _5754_ (.Y(_1883_),
    .A(_1867_),
    .B(_1881_));
 sg13g2_xnor2_1 _5755_ (.Y(_1884_),
    .A(_1827_),
    .B(_1848_));
 sg13g2_a21oi_1 _5756_ (.A1(_1882_),
    .A2(_1883_),
    .Y(_1885_),
    .B1(_1884_));
 sg13g2_a21oi_1 _5757_ (.A1(_1834_),
    .A2(_1859_),
    .Y(_1886_),
    .B1(_1858_));
 sg13g2_a21oi_1 _5758_ (.A1(_1853_),
    .A2(_1856_),
    .Y(_1887_),
    .B1(_1855_));
 sg13g2_xnor2_1 _5759_ (.Y(_1888_),
    .A(_1737_),
    .B(_1738_));
 sg13g2_nor2_1 _5760_ (.A(_1887_),
    .B(_1888_),
    .Y(_1889_));
 sg13g2_xor2_1 _5761_ (.B(_1888_),
    .A(_1887_),
    .X(_1890_));
 sg13g2_nor2b_1 _5762_ (.A(_1852_),
    .B_N(_1890_),
    .Y(_1891_));
 sg13g2_xor2_1 _5763_ (.B(_1890_),
    .A(_1852_),
    .X(_1892_));
 sg13g2_a22oi_1 _5764_ (.Y(_1893_),
    .B1(_1886_),
    .B2(_1892_),
    .A2(_1860_),
    .A1(_1849_));
 sg13g2_o21ai_1 _5765_ (.B1(_1893_),
    .Y(_1894_),
    .A1(_1861_),
    .A2(_1885_));
 sg13g2_nor2_1 _5766_ (.A(_1889_),
    .B(_1891_),
    .Y(_1895_));
 sg13g2_or2_1 _5767_ (.X(_1896_),
    .B(_1891_),
    .A(_1889_));
 sg13g2_xor2_1 _5768_ (.B(_1763_),
    .A(_1736_),
    .X(_1897_));
 sg13g2_inv_1 _5769_ (.Y(_1898_),
    .A(_1897_));
 sg13g2_nor2_1 _5770_ (.A(_1886_),
    .B(_1892_),
    .Y(_1899_));
 sg13g2_a21oi_1 _5771_ (.A1(_1896_),
    .A2(_1898_),
    .Y(_1900_),
    .B1(_1899_));
 sg13g2_a22oi_1 _5772_ (.Y(_1901_),
    .B1(_1900_),
    .B2(_1894_),
    .A2(_1897_),
    .A1(_1895_));
 sg13g2_a221oi_1 _5773_ (.B2(_1894_),
    .C1(_1792_),
    .B1(_1900_),
    .A1(_1895_),
    .Y(_1902_),
    .A2(_1897_));
 sg13g2_xnor2_1 _5774_ (.Y(_1903_),
    .A(_1792_),
    .B(_1901_));
 sg13g2_and2_1 _5775_ (.A(_1658_),
    .B(_1903_),
    .X(_1904_));
 sg13g2_o21ai_1 _5776_ (.B1(_1789_),
    .Y(_1905_),
    .A1(_1766_),
    .A2(_1787_));
 sg13g2_a21oi_1 _5777_ (.A1(_1769_),
    .A2(_1785_),
    .Y(_1906_),
    .B1(_1784_));
 sg13g2_or2_1 _5778_ (.X(_1907_),
    .B(_1780_),
    .A(_1744_));
 sg13g2_xnor2_1 _5779_ (.Y(_1908_),
    .A(_1744_),
    .B(_1780_));
 sg13g2_inv_1 _5780_ (.Y(_1909_),
    .A(_1908_));
 sg13g2_nand2_1 _5781_ (.Y(_1910_),
    .A(net578),
    .B(_1701_));
 sg13g2_o21ai_1 _5782_ (.B1(_1910_),
    .Y(_1911_),
    .A1(_1662_),
    .A2(_1718_));
 sg13g2_a21oi_1 _5783_ (.A1(_1774_),
    .A2(_1778_),
    .Y(_1912_),
    .B1(_1777_));
 sg13g2_nand2_1 _5784_ (.Y(_1913_),
    .A(net593),
    .B(net567));
 sg13g2_xor2_1 _5785_ (.B(_1913_),
    .A(_1775_),
    .X(_1914_));
 sg13g2_nand2_1 _5786_ (.Y(_1915_),
    .A(_1774_),
    .B(_1914_));
 sg13g2_xnor2_1 _5787_ (.Y(_1916_),
    .A(_1773_),
    .B(_1914_));
 sg13g2_nand2b_2 _5788_ (.Y(_1917_),
    .B(_1916_),
    .A_N(_1912_));
 sg13g2_xnor2_1 _5789_ (.Y(_1918_),
    .A(_1912_),
    .B(_1916_));
 sg13g2_nand2_1 _5790_ (.Y(_1919_),
    .A(_1911_),
    .B(_1918_));
 sg13g2_xnor2_1 _5791_ (.Y(_1920_),
    .A(_1911_),
    .B(_1918_));
 sg13g2_nor2_1 _5792_ (.A(_1782_),
    .B(_1920_),
    .Y(_1921_));
 sg13g2_xor2_1 _5793_ (.B(_1920_),
    .A(_1782_),
    .X(_1922_));
 sg13g2_xnor2_1 _5794_ (.Y(_1923_),
    .A(_1908_),
    .B(_1922_));
 sg13g2_nor2b_1 _5795_ (.A(_1906_),
    .B_N(_1923_),
    .Y(_1924_));
 sg13g2_xnor2_1 _5796_ (.Y(_1925_),
    .A(_1906_),
    .B(_1923_));
 sg13g2_nor2b_1 _5797_ (.A(_1767_),
    .B_N(_1925_),
    .Y(_1926_));
 sg13g2_xnor2_1 _5798_ (.Y(_1927_),
    .A(_1767_),
    .B(_1925_));
 sg13g2_nand2_1 _5799_ (.Y(_1928_),
    .A(_1905_),
    .B(_1927_));
 sg13g2_xor2_1 _5800_ (.B(_1927_),
    .A(_1905_),
    .X(_1929_));
 sg13g2_o21ai_1 _5801_ (.B1(_1929_),
    .Y(_1930_),
    .A1(_1791_),
    .A2(_1902_));
 sg13g2_or3_1 _5802_ (.A(_1791_),
    .B(_1902_),
    .C(_1929_),
    .X(_1931_));
 sg13g2_a21oi_2 _5803_ (.B1(_1552_),
    .Y(_1932_),
    .A2(_1553_),
    .A1(_1500_));
 sg13g2_nand2_1 _5804_ (.Y(_1933_),
    .A(_1548_),
    .B(_1550_));
 sg13g2_nand3_1 _5805_ (.B(_1520_),
    .C(_1544_),
    .A(net588),
    .Y(_1934_));
 sg13g2_a22oi_1 _5806_ (.Y(_1935_),
    .B1(_1934_),
    .B2(_1425_),
    .A2(_1543_),
    .A1(_1434_));
 sg13g2_a21oi_1 _5807_ (.A1(_1540_),
    .A2(_1546_),
    .Y(_1936_),
    .B1(_1539_));
 sg13g2_a21oi_1 _5808_ (.A1(_1516_),
    .A2(_1537_),
    .Y(_1937_),
    .B1(_1536_));
 sg13g2_nand2_1 _5809_ (.Y(_1938_),
    .A(net599),
    .B(net568));
 sg13g2_nor3_1 _5810_ (.A(_0455_),
    .B(_1514_),
    .C(_1535_),
    .Y(_1939_));
 sg13g2_a22oi_1 _5811_ (.Y(_1940_),
    .B1(net568),
    .B2(net599),
    .A2(_1483_),
    .A1(_0454_));
 sg13g2_nor2_1 _5812_ (.A(_1939_),
    .B(_1940_),
    .Y(_1941_));
 sg13g2_xnor2_1 _5813_ (.Y(_1942_),
    .A(_1517_),
    .B(_1941_));
 sg13g2_nor2b_1 _5814_ (.A(_1937_),
    .B_N(_1942_),
    .Y(_1943_));
 sg13g2_xnor2_1 _5815_ (.Y(_1944_),
    .A(_1937_),
    .B(_1942_));
 sg13g2_nand2_1 _5816_ (.Y(_1945_),
    .A(_1434_),
    .B(net588));
 sg13g2_xnor2_1 _5817_ (.Y(_1946_),
    .A(_1460_),
    .B(_1520_));
 sg13g2_xnor2_1 _5818_ (.Y(_1947_),
    .A(_1945_),
    .B(_1946_));
 sg13g2_xnor2_1 _5819_ (.Y(_1948_),
    .A(_1944_),
    .B(_1947_));
 sg13g2_xor2_1 _5820_ (.B(_1948_),
    .A(_1936_),
    .X(_1949_));
 sg13g2_nand2b_1 _5821_ (.Y(_1950_),
    .B(_1949_),
    .A_N(_1935_));
 sg13g2_xnor2_1 _5822_ (.Y(_1951_),
    .A(_1935_),
    .B(_1949_));
 sg13g2_nand2_1 _5823_ (.Y(_1952_),
    .A(_1933_),
    .B(_1951_));
 sg13g2_xnor2_1 _5824_ (.Y(_1953_),
    .A(_1933_),
    .B(_1951_));
 sg13g2_xnor2_1 _5825_ (.Y(_1954_),
    .A(_1532_),
    .B(_1953_));
 sg13g2_nor2_1 _5826_ (.A(_1932_),
    .B(_1954_),
    .Y(_1955_));
 sg13g2_xor2_1 _5827_ (.B(_1954_),
    .A(_1932_),
    .X(_1956_));
 sg13g2_inv_1 _5828_ (.Y(_1957_),
    .A(_1956_));
 sg13g2_nor2b_1 _5829_ (.A(_1555_),
    .B_N(_1656_),
    .Y(_1958_));
 sg13g2_xnor2_1 _5830_ (.Y(_1959_),
    .A(_1956_),
    .B(_1958_));
 sg13g2_and3_1 _5831_ (.X(_1960_),
    .A(_1930_),
    .B(_1931_),
    .C(_1959_));
 sg13g2_a21o_1 _5832_ (.A2(_1931_),
    .A1(_1930_),
    .B1(_1959_),
    .X(_1961_));
 sg13g2_nor2b_1 _5833_ (.A(_1960_),
    .B_N(_1961_),
    .Y(_1962_));
 sg13g2_nand2_1 _5834_ (.Y(_1963_),
    .A(\generated._406[3] ),
    .B(\generated._406[1] ));
 sg13g2_nor3_2 _5835_ (.A(\generated._406[2] ),
    .B(\generated._1000[0] ),
    .C(_1963_),
    .Y(_1964_));
 sg13g2_nand2_1 _5836_ (.Y(_1965_),
    .A(_3208_),
    .B(_1964_));
 sg13g2_xnor2_1 _5837_ (.Y(_1966_),
    .A(_3208_),
    .B(_1964_));
 sg13g2_or3_1 _5838_ (.A(net672),
    .B(\generated._381[0] ),
    .C(\generated._381[1] ),
    .X(_1967_));
 sg13g2_nor2_1 _5839_ (.A(\generated._381[2] ),
    .B(_1967_),
    .Y(_1968_));
 sg13g2_nand2b_2 _5840_ (.Y(_1969_),
    .B(_1968_),
    .A_N(\generated._381[3] ));
 sg13g2_nand2_1 _5841_ (.Y(_1970_),
    .A(\generated._381[4] ),
    .B(_1969_));
 sg13g2_nor2_1 _5842_ (.A(\generated._381[4] ),
    .B(_1969_),
    .Y(_1971_));
 sg13g2_nor2_1 _5843_ (.A(net711),
    .B(_1971_),
    .Y(_1972_));
 sg13g2_a22oi_1 _5844_ (.Y(_1973_),
    .B1(_1970_),
    .B2(_1972_),
    .A2(_2871_),
    .A1(net711));
 sg13g2_nor2_1 _5845_ (.A(net604),
    .B(_1973_),
    .Y(_1974_));
 sg13g2_xnor2_1 _5846_ (.Y(_1975_),
    .A(net672),
    .B(\generated._381[0] ));
 sg13g2_mux2_2 _5847_ (.A0(_1975_),
    .A1(_0087_),
    .S(net716),
    .X(_1976_));
 sg13g2_nor2_2 _5848_ (.A(_3222_),
    .B(_1965_),
    .Y(_1977_));
 sg13g2_nor2_2 _5849_ (.A(_0289_),
    .B(_1977_),
    .Y(_1978_));
 sg13g2_or2_1 _5850_ (.X(_1979_),
    .B(_1977_),
    .A(_0289_));
 sg13g2_nand2_1 _5851_ (.Y(_1980_),
    .A(net672),
    .B(net586));
 sg13g2_o21ai_1 _5852_ (.B1(_1980_),
    .Y(_1981_),
    .A1(_1976_),
    .A2(net586));
 sg13g2_nand2_1 _5853_ (.Y(_1982_),
    .A(_1974_),
    .B(_1981_));
 sg13g2_inv_1 _5854_ (.Y(_1983_),
    .A(_1982_));
 sg13g2_nand2_1 _5855_ (.Y(_1984_),
    .A(_3236_),
    .B(_1977_));
 sg13g2_xor2_1 _5856_ (.B(_1977_),
    .A(_3236_),
    .X(_1985_));
 sg13g2_nand2b_2 _5857_ (.Y(_1986_),
    .B(net584),
    .A_N(_1976_));
 sg13g2_xnor2_1 _5858_ (.Y(_1987_),
    .A(_0291_),
    .B(_1984_));
 sg13g2_xor2_1 _5859_ (.B(_1984_),
    .A(_0291_),
    .X(_1988_));
 sg13g2_o21ai_1 _5860_ (.B1(\generated._381[1] ),
    .Y(_1989_),
    .A1(net672),
    .A2(\generated._381[0] ));
 sg13g2_a21oi_1 _5861_ (.A1(_1967_),
    .A2(_1989_),
    .Y(_1990_),
    .B1(net712));
 sg13g2_a21oi_2 _5862_ (.B1(_1990_),
    .Y(_1991_),
    .A2(net716),
    .A1(_0093_));
 sg13g2_nand2_1 _5863_ (.Y(_1992_),
    .A(_1987_),
    .B(_1991_));
 sg13g2_nand2_1 _5864_ (.Y(_1993_),
    .A(net584),
    .B(_1991_));
 sg13g2_nor2_1 _5865_ (.A(_1986_),
    .B(_1992_),
    .Y(_1994_));
 sg13g2_xor2_1 _5866_ (.B(_1965_),
    .A(_3222_),
    .X(_1995_));
 sg13g2_nand2_1 _5867_ (.Y(_1996_),
    .A(\generated._381[2] ),
    .B(_1967_));
 sg13g2_nor2_1 _5868_ (.A(net712),
    .B(_1968_),
    .Y(_1997_));
 sg13g2_a22oi_1 _5869_ (.Y(_1998_),
    .B1(_1996_),
    .B2(_1997_),
    .A2(net712),
    .A1(_2842_));
 sg13g2_nand2b_1 _5870_ (.Y(_1999_),
    .B(net595),
    .A_N(_1998_));
 sg13g2_o21ai_1 _5871_ (.B1(_1993_),
    .Y(_2000_),
    .A1(_1976_),
    .A2(_1988_));
 sg13g2_o21ai_1 _5872_ (.B1(_2000_),
    .Y(_2001_),
    .A1(_1986_),
    .A2(_1992_));
 sg13g2_nor2_1 _5873_ (.A(_1999_),
    .B(_2001_),
    .Y(_2002_));
 sg13g2_nor2_2 _5874_ (.A(_1994_),
    .B(_2002_),
    .Y(_2003_));
 sg13g2_inv_1 _5875_ (.Y(_2004_),
    .A(_2003_));
 sg13g2_o21ai_1 _5876_ (.B1(\generated._381[3] ),
    .Y(_2005_),
    .A1(\generated._381[2] ),
    .A2(_1967_));
 sg13g2_a21oi_1 _5877_ (.A1(_1969_),
    .A2(_2005_),
    .Y(_2006_),
    .B1(net711));
 sg13g2_a21oi_2 _5878_ (.B1(_2006_),
    .Y(_2007_),
    .A2(_0086_),
    .A1(net712));
 sg13g2_nand2_1 _5879_ (.Y(_2008_),
    .A(net595),
    .B(_2007_));
 sg13g2_inv_1 _5880_ (.Y(_2009_),
    .A(_2008_));
 sg13g2_nand2b_1 _5881_ (.Y(_2010_),
    .B(_1987_),
    .A_N(_1998_));
 sg13g2_nor2b_1 _5882_ (.A(_1998_),
    .B_N(net584),
    .Y(_2011_));
 sg13g2_nor2_1 _5883_ (.A(_1993_),
    .B(_2010_),
    .Y(_2012_));
 sg13g2_xnor2_1 _5884_ (.Y(_2013_),
    .A(_1992_),
    .B(_2011_));
 sg13g2_xnor2_1 _5885_ (.Y(_2014_),
    .A(_2008_),
    .B(_2013_));
 sg13g2_xor2_1 _5886_ (.B(_2014_),
    .A(_2003_),
    .X(_2015_));
 sg13g2_xnor2_1 _5887_ (.Y(_2016_),
    .A(_1974_),
    .B(_1981_));
 sg13g2_nor2_1 _5888_ (.A(_2015_),
    .B(_2016_),
    .Y(_2017_));
 sg13g2_a21oi_1 _5889_ (.A1(_2004_),
    .A2(_2014_),
    .Y(_2018_),
    .B1(_2017_));
 sg13g2_a21oi_1 _5890_ (.A1(_2009_),
    .A2(_2013_),
    .Y(_2019_),
    .B1(_2012_));
 sg13g2_nor2b_1 _5891_ (.A(_1973_),
    .B_N(net595),
    .Y(_2020_));
 sg13g2_nand2_1 _5892_ (.Y(_2021_),
    .A(net584),
    .B(_2007_));
 sg13g2_nor2_1 _5893_ (.A(_2010_),
    .B(_2021_),
    .Y(_2022_));
 sg13g2_xor2_1 _5894_ (.B(_2021_),
    .A(_2010_),
    .X(_2023_));
 sg13g2_xnor2_1 _5895_ (.Y(_2024_),
    .A(_2020_),
    .B(_2023_));
 sg13g2_nor2_1 _5896_ (.A(_2019_),
    .B(_2024_),
    .Y(_2025_));
 sg13g2_xor2_1 _5897_ (.B(_2024_),
    .A(_2019_),
    .X(_2026_));
 sg13g2_nor3_1 _5898_ (.A(\generated._381[5] ),
    .B(\generated._381[4] ),
    .C(_1969_),
    .Y(_2027_));
 sg13g2_xnor2_1 _5899_ (.Y(_2028_),
    .A(\generated._381[5] ),
    .B(_1971_));
 sg13g2_nor2_1 _5900_ (.A(net711),
    .B(_2028_),
    .Y(_2029_));
 sg13g2_a21oi_2 _5901_ (.B1(_2029_),
    .Y(_2030_),
    .A2(_0084_),
    .A1(net712));
 sg13g2_nand2b_1 _5902_ (.Y(_2031_),
    .B(_2030_),
    .A_N(net604));
 sg13g2_nor2_1 _5903_ (.A(_1976_),
    .B(net587),
    .Y(_2032_));
 sg13g2_a21oi_1 _5904_ (.A1(net587),
    .A2(_1991_),
    .Y(_2033_),
    .B1(_2032_));
 sg13g2_nor2_1 _5905_ (.A(_2031_),
    .B(_2033_),
    .Y(_2034_));
 sg13g2_xor2_1 _5906_ (.B(_2033_),
    .A(_2031_),
    .X(_2035_));
 sg13g2_xnor2_1 _5907_ (.Y(_2036_),
    .A(_2026_),
    .B(_2035_));
 sg13g2_nor2_1 _5908_ (.A(_2018_),
    .B(_2036_),
    .Y(_2037_));
 sg13g2_xor2_1 _5909_ (.B(_2036_),
    .A(_2018_),
    .X(_2038_));
 sg13g2_xnor2_1 _5910_ (.Y(_2039_),
    .A(_1982_),
    .B(_2038_));
 sg13g2_nor2b_1 _5911_ (.A(net604),
    .B_N(_2007_),
    .Y(_2040_));
 sg13g2_and3_1 _5912_ (.X(_2041_),
    .A(\generated._501[0] ),
    .B(net587),
    .C(_2040_));
 sg13g2_nor3_1 _5913_ (.A(_0088_),
    .B(_1986_),
    .C(_1988_),
    .Y(_2042_));
 sg13g2_nand2_1 _5914_ (.Y(_2043_),
    .A(_1991_),
    .B(net595));
 sg13g2_o21ai_1 _5915_ (.B1(_1986_),
    .Y(_2044_),
    .A1(_0088_),
    .A2(_1988_));
 sg13g2_nand2b_1 _5916_ (.Y(_2045_),
    .B(_2044_),
    .A_N(_2042_));
 sg13g2_nor2_1 _5917_ (.A(_2043_),
    .B(_2045_),
    .Y(_2046_));
 sg13g2_nor2_1 _5918_ (.A(_2042_),
    .B(_2046_),
    .Y(_2047_));
 sg13g2_xor2_1 _5919_ (.B(_2001_),
    .A(_1999_),
    .X(_2048_));
 sg13g2_o21ai_1 _5920_ (.B1(_2048_),
    .Y(_2049_),
    .A1(_2042_),
    .A2(_2046_));
 sg13g2_a21oi_1 _5921_ (.A1(net672),
    .A2(net587),
    .Y(_2050_),
    .B1(_2040_));
 sg13g2_or2_1 _5922_ (.X(_2051_),
    .B(_2050_),
    .A(_2041_));
 sg13g2_xnor2_1 _5923_ (.Y(_2052_),
    .A(_2047_),
    .B(_2048_));
 sg13g2_nand2b_1 _5924_ (.Y(_2053_),
    .B(_2052_),
    .A_N(_2051_));
 sg13g2_and2_1 _5925_ (.A(_2049_),
    .B(_2053_),
    .X(_2054_));
 sg13g2_xnor2_1 _5926_ (.Y(_2055_),
    .A(_2015_),
    .B(_2016_));
 sg13g2_nor2_1 _5927_ (.A(_2054_),
    .B(_2055_),
    .Y(_2056_));
 sg13g2_xor2_1 _5928_ (.B(_2055_),
    .A(_2054_),
    .X(_2057_));
 sg13g2_nor2_1 _5929_ (.A(_2041_),
    .B(_2057_),
    .Y(_2058_));
 sg13g2_xnor2_1 _5930_ (.Y(_2059_),
    .A(_2051_),
    .B(_2052_));
 sg13g2_nor2b_1 _5931_ (.A(_1976_),
    .B_N(net595),
    .Y(_2060_));
 sg13g2_a21oi_1 _5932_ (.A1(net672),
    .A2(net584),
    .Y(_2061_),
    .B1(_2060_));
 sg13g2_nand3_1 _5933_ (.B(net584),
    .C(_2060_),
    .A(net672),
    .Y(_2062_));
 sg13g2_a22oi_1 _5934_ (.Y(_2063_),
    .B1(_2062_),
    .B2(_1991_),
    .A2(_2060_),
    .A1(_2872_));
 sg13g2_nor2_1 _5935_ (.A(_1991_),
    .B(_2062_),
    .Y(_2064_));
 sg13g2_or4_1 _5936_ (.A(net604),
    .B(_2061_),
    .C(_2063_),
    .D(_2064_),
    .X(_2065_));
 sg13g2_nor2_1 _5937_ (.A(_1998_),
    .B(_2065_),
    .Y(_2066_));
 sg13g2_xnor2_1 _5938_ (.Y(_2067_),
    .A(_2043_),
    .B(_2045_));
 sg13g2_nor2_1 _5939_ (.A(_2062_),
    .B(_2067_),
    .Y(_2068_));
 sg13g2_a21oi_1 _5940_ (.A1(_2066_),
    .A2(_2068_),
    .Y(_2069_),
    .B1(_2059_));
 sg13g2_nand2_1 _5941_ (.Y(_2070_),
    .A(_2062_),
    .B(_2067_));
 sg13g2_nor2_1 _5942_ (.A(_2066_),
    .B(_2070_),
    .Y(_2071_));
 sg13g2_o21ai_1 _5943_ (.B1(_2065_),
    .Y(_2072_),
    .A1(net604),
    .A2(_1998_));
 sg13g2_nor2_1 _5944_ (.A(_2068_),
    .B(_2072_),
    .Y(_2073_));
 sg13g2_nor4_1 _5945_ (.A(_2058_),
    .B(_2069_),
    .C(_2071_),
    .D(_2073_),
    .Y(_2074_));
 sg13g2_a21o_1 _5946_ (.A2(_2057_),
    .A1(_2041_),
    .B1(_2074_),
    .X(_2075_));
 sg13g2_o21ai_1 _5947_ (.B1(_2056_),
    .Y(_2076_),
    .A1(_2039_),
    .A2(_2074_));
 sg13g2_a21oi_1 _5948_ (.A1(_1983_),
    .A2(_2038_),
    .Y(_2077_),
    .B1(_2037_));
 sg13g2_a21oi_1 _5949_ (.A1(_2026_),
    .A2(_2035_),
    .Y(_2078_),
    .B1(_2025_));
 sg13g2_a21oi_1 _5950_ (.A1(_2020_),
    .A2(_2023_),
    .Y(_2079_),
    .B1(_2022_));
 sg13g2_nand2_1 _5951_ (.Y(_2080_),
    .A(net595),
    .B(_2030_));
 sg13g2_inv_1 _5952_ (.Y(_2081_),
    .A(_2080_));
 sg13g2_nand2b_1 _5953_ (.Y(_2082_),
    .B(_1987_),
    .A_N(_1973_));
 sg13g2_nor2b_1 _5954_ (.A(_1973_),
    .B_N(net584),
    .Y(_2083_));
 sg13g2_nor2_1 _5955_ (.A(_2021_),
    .B(_2082_),
    .Y(_2084_));
 sg13g2_a21oi_1 _5956_ (.A1(_1987_),
    .A2(_2007_),
    .Y(_2085_),
    .B1(_2083_));
 sg13g2_nor2_1 _5957_ (.A(_2084_),
    .B(_2085_),
    .Y(_2086_));
 sg13g2_xnor2_1 _5958_ (.Y(_2087_),
    .A(_2080_),
    .B(_2086_));
 sg13g2_nand2b_1 _5959_ (.Y(_2088_),
    .B(_2087_),
    .A_N(_2079_));
 sg13g2_xnor2_1 _5960_ (.Y(_2089_),
    .A(_2079_),
    .B(_2087_));
 sg13g2_nand2b_1 _5961_ (.Y(_2090_),
    .B(\generated._381[6] ),
    .A_N(_2027_));
 sg13g2_nand2b_1 _5962_ (.Y(_2091_),
    .B(_2027_),
    .A_N(\generated._381[6] ));
 sg13g2_a21oi_1 _5963_ (.A1(_2090_),
    .A2(_2091_),
    .Y(_2092_),
    .B1(net711));
 sg13g2_a21oi_2 _5964_ (.B1(_2092_),
    .Y(_2093_),
    .A2(_0083_),
    .A1(net711));
 sg13g2_nand2b_1 _5965_ (.Y(_2094_),
    .B(_2093_),
    .A_N(net604));
 sg13g2_nor2_1 _5966_ (.A(net586),
    .B(_1998_),
    .Y(_2095_));
 sg13g2_a21oi_1 _5967_ (.A1(net586),
    .A2(_1991_),
    .Y(_2096_),
    .B1(_2095_));
 sg13g2_or2_1 _5968_ (.X(_2097_),
    .B(_2096_),
    .A(_2094_));
 sg13g2_xor2_1 _5969_ (.B(_2096_),
    .A(_2094_),
    .X(_2098_));
 sg13g2_nand2_1 _5970_ (.Y(_2099_),
    .A(_2089_),
    .B(_2098_));
 sg13g2_xnor2_1 _5971_ (.Y(_2100_),
    .A(_2089_),
    .B(_2098_));
 sg13g2_or2_1 _5972_ (.X(_2101_),
    .B(_2100_),
    .A(_2078_));
 sg13g2_xor2_1 _5973_ (.B(_2100_),
    .A(_2078_),
    .X(_2102_));
 sg13g2_nand2_1 _5974_ (.Y(_2103_),
    .A(_2034_),
    .B(_2102_));
 sg13g2_xnor2_1 _5975_ (.Y(_2104_),
    .A(_2034_),
    .B(_2102_));
 sg13g2_o21ai_1 _5976_ (.B1(_2076_),
    .Y(_2105_),
    .A1(_2077_),
    .A2(_2104_));
 sg13g2_a21oi_1 _5977_ (.A1(_2039_),
    .A2(_2075_),
    .Y(_2106_),
    .B1(_2105_));
 sg13g2_and2_1 _5978_ (.A(_2088_),
    .B(_2099_),
    .X(_2107_));
 sg13g2_a21oi_1 _5979_ (.A1(_2081_),
    .A2(_2086_),
    .Y(_2108_),
    .B1(_2084_));
 sg13g2_nand2_1 _5980_ (.Y(_2109_),
    .A(_1995_),
    .B(_2093_));
 sg13g2_inv_1 _5981_ (.Y(_2110_),
    .A(_2109_));
 sg13g2_nand2_1 _5982_ (.Y(_2111_),
    .A(net585),
    .B(_2030_));
 sg13g2_nor2_1 _5983_ (.A(_2082_),
    .B(_2111_),
    .Y(_2112_));
 sg13g2_xor2_1 _5984_ (.B(_2111_),
    .A(_2082_),
    .X(_2113_));
 sg13g2_xnor2_1 _5985_ (.Y(_2114_),
    .A(_2109_),
    .B(_2113_));
 sg13g2_nand2b_1 _5986_ (.Y(_2115_),
    .B(_2114_),
    .A_N(_2108_));
 sg13g2_xnor2_1 _5987_ (.Y(_2116_),
    .A(_2108_),
    .B(_2114_));
 sg13g2_nor2_1 _5988_ (.A(\generated._381[7] ),
    .B(_2091_),
    .Y(_2117_));
 sg13g2_xor2_1 _5989_ (.B(_2091_),
    .A(\generated._381[7] ),
    .X(_2118_));
 sg13g2_nand2_1 _5990_ (.Y(_2119_),
    .A(net711),
    .B(_0082_));
 sg13g2_o21ai_1 _5991_ (.B1(_2119_),
    .Y(_2120_),
    .A1(net711),
    .A2(_2118_));
 sg13g2_nor2_1 _5992_ (.A(net604),
    .B(_2120_),
    .Y(_2121_));
 sg13g2_nand2_1 _5993_ (.Y(_2122_),
    .A(net587),
    .B(_2007_));
 sg13g2_o21ai_1 _5994_ (.B1(_2122_),
    .Y(_2123_),
    .A1(net587),
    .A2(_1998_));
 sg13g2_nor2_1 _5995_ (.A(_1979_),
    .B(_2120_),
    .Y(_2124_));
 sg13g2_and2_1 _5996_ (.A(_2121_),
    .B(_2123_),
    .X(_2125_));
 sg13g2_xor2_1 _5997_ (.B(_2123_),
    .A(_2121_),
    .X(_2126_));
 sg13g2_nand2_1 _5998_ (.Y(_2127_),
    .A(_2116_),
    .B(_2126_));
 sg13g2_xnor2_1 _5999_ (.Y(_2128_),
    .A(_2116_),
    .B(_2126_));
 sg13g2_or2_1 _6000_ (.X(_2129_),
    .B(_2128_),
    .A(_2107_));
 sg13g2_xor2_1 _6001_ (.B(_2128_),
    .A(_2107_),
    .X(_2130_));
 sg13g2_nand2b_1 _6002_ (.Y(_2131_),
    .B(_2130_),
    .A_N(_2097_));
 sg13g2_nand3_1 _6003_ (.B(_2007_),
    .C(_2125_),
    .A(net586),
    .Y(_2132_));
 sg13g2_inv_1 _6004_ (.Y(_2133_),
    .A(_2132_));
 sg13g2_a21oi_1 _6005_ (.A1(net586),
    .A2(_2007_),
    .Y(_2134_),
    .B1(_2125_));
 sg13g2_or2_1 _6006_ (.X(_2135_),
    .B(_2134_),
    .A(_2133_));
 sg13g2_inv_1 _6007_ (.Y(_2136_),
    .A(_2135_));
 sg13g2_and2_1 _6008_ (.A(_2115_),
    .B(_2127_),
    .X(_2137_));
 sg13g2_a21oi_1 _6009_ (.A1(_2110_),
    .A2(_2113_),
    .Y(_2138_),
    .B1(_2112_));
 sg13g2_nand2_1 _6010_ (.Y(_2139_),
    .A(_1987_),
    .B(_2093_));
 sg13g2_and2_1 _6011_ (.A(net585),
    .B(_2093_),
    .X(_2140_));
 sg13g2_nor2_1 _6012_ (.A(_2111_),
    .B(_2139_),
    .Y(_2141_));
 sg13g2_a21oi_1 _6013_ (.A1(_1987_),
    .A2(_2030_),
    .Y(_2142_),
    .B1(_2140_));
 sg13g2_nor2_1 _6014_ (.A(_2141_),
    .B(_2142_),
    .Y(_2143_));
 sg13g2_nor2b_1 _6015_ (.A(_2138_),
    .B_N(_2143_),
    .Y(_2144_));
 sg13g2_xnor2_1 _6016_ (.Y(_2145_),
    .A(_2138_),
    .B(_2143_));
 sg13g2_xor2_1 _6017_ (.B(_2117_),
    .A(\generated._380 ),
    .X(_2146_));
 sg13g2_nand2b_1 _6018_ (.Y(_2147_),
    .B(net713),
    .A_N(_0081_));
 sg13g2_o21ai_1 _6019_ (.B1(_2147_),
    .Y(_2148_),
    .A1(net713),
    .A2(_2146_));
 sg13g2_inv_1 _6020_ (.Y(_2149_),
    .A(_2148_));
 sg13g2_and2_1 _6021_ (.A(net595),
    .B(net575),
    .X(_2150_));
 sg13g2_nand2_2 _6022_ (.Y(_2151_),
    .A(net595),
    .B(net575));
 sg13g2_nand2b_1 _6023_ (.Y(_2152_),
    .B(_1995_),
    .A_N(_2120_));
 sg13g2_nand2b_1 _6024_ (.Y(_2153_),
    .B(net575),
    .A_N(_1966_));
 sg13g2_xnor2_1 _6025_ (.Y(_2154_),
    .A(_2152_),
    .B(net570));
 sg13g2_nor3_1 _6026_ (.A(_1973_),
    .B(net586),
    .C(_2154_),
    .Y(_2155_));
 sg13g2_o21ai_1 _6027_ (.B1(_2154_),
    .Y(_2156_),
    .A1(_1973_),
    .A2(net586));
 sg13g2_nand2b_1 _6028_ (.Y(_2157_),
    .B(_2156_),
    .A_N(_2155_));
 sg13g2_inv_1 _6029_ (.Y(_2158_),
    .A(_2157_));
 sg13g2_xor2_1 _6030_ (.B(_2157_),
    .A(_2145_),
    .X(_2159_));
 sg13g2_nor2_1 _6031_ (.A(_2137_),
    .B(_2159_),
    .Y(_2160_));
 sg13g2_xor2_1 _6032_ (.B(_2159_),
    .A(_2137_),
    .X(_2161_));
 sg13g2_xnor2_1 _6033_ (.Y(_2162_),
    .A(_2136_),
    .B(_2161_));
 sg13g2_a21oi_1 _6034_ (.A1(_2129_),
    .A2(_2131_),
    .Y(_2163_),
    .B1(_2162_));
 sg13g2_xor2_1 _6035_ (.B(_2130_),
    .A(_2097_),
    .X(_2164_));
 sg13g2_a21oi_1 _6036_ (.A1(_2101_),
    .A2(_2103_),
    .Y(_2165_),
    .B1(_2164_));
 sg13g2_or2_1 _6037_ (.X(_2166_),
    .B(_2165_),
    .A(_2163_));
 sg13g2_nand3_1 _6038_ (.B(_2131_),
    .C(_2162_),
    .A(_2129_),
    .Y(_2167_));
 sg13g2_nand2_1 _6039_ (.Y(_2168_),
    .A(_2077_),
    .B(_2104_));
 sg13g2_nand3_1 _6040_ (.B(_2103_),
    .C(_2164_),
    .A(_2101_),
    .Y(_2169_));
 sg13g2_nand3_1 _6041_ (.B(_2168_),
    .C(_2169_),
    .A(_2167_),
    .Y(_2170_));
 sg13g2_nor3_1 _6042_ (.A(_2106_),
    .B(_2166_),
    .C(_2170_),
    .Y(_2171_));
 sg13g2_a21oi_1 _6043_ (.A1(_2136_),
    .A2(_2161_),
    .Y(_2172_),
    .B1(_2160_));
 sg13g2_a21oi_1 _6044_ (.A1(_2121_),
    .A2(_2150_),
    .Y(_2173_),
    .B1(_2155_));
 sg13g2_a21oi_1 _6045_ (.A1(_2145_),
    .A2(_2158_),
    .Y(_2174_),
    .B1(_2144_));
 sg13g2_nor2_1 _6046_ (.A(_1988_),
    .B(_2120_),
    .Y(_2175_));
 sg13g2_nor2b_1 _6047_ (.A(_2120_),
    .B_N(net585),
    .Y(_2176_));
 sg13g2_xnor2_1 _6048_ (.Y(_2177_),
    .A(_2139_),
    .B(_2176_));
 sg13g2_xnor2_1 _6049_ (.Y(_2178_),
    .A(_2151_),
    .B(_2177_));
 sg13g2_xnor2_1 _6050_ (.Y(_2179_),
    .A(_2141_),
    .B(_2178_));
 sg13g2_nor2_1 _6051_ (.A(_1973_),
    .B(net587),
    .Y(_2180_));
 sg13g2_a21oi_1 _6052_ (.A1(_1978_),
    .A2(_2030_),
    .Y(_2181_),
    .B1(_2180_));
 sg13g2_or2_1 _6053_ (.X(_2182_),
    .B(_2181_),
    .A(_2153_));
 sg13g2_xor2_1 _6054_ (.B(_2181_),
    .A(net570),
    .X(_2183_));
 sg13g2_nor2b_1 _6055_ (.A(_2179_),
    .B_N(_2183_),
    .Y(_2184_));
 sg13g2_xnor2_1 _6056_ (.Y(_2185_),
    .A(_2179_),
    .B(_2183_));
 sg13g2_nand2b_1 _6057_ (.Y(_2186_),
    .B(_2185_),
    .A_N(_2174_));
 sg13g2_xnor2_1 _6058_ (.Y(_2187_),
    .A(_2174_),
    .B(_2185_));
 sg13g2_inv_1 _6059_ (.Y(_2188_),
    .A(_2187_));
 sg13g2_xnor2_1 _6060_ (.Y(_2189_),
    .A(_2173_),
    .B(_2187_));
 sg13g2_nor2b_1 _6061_ (.A(_2172_),
    .B_N(_2189_),
    .Y(_2190_));
 sg13g2_xnor2_1 _6062_ (.Y(_2191_),
    .A(_2172_),
    .B(_2189_));
 sg13g2_xnor2_1 _6063_ (.Y(_2192_),
    .A(_2132_),
    .B(_2191_));
 sg13g2_nand2_1 _6064_ (.Y(_2193_),
    .A(_2165_),
    .B(_2167_));
 sg13g2_nand2_1 _6065_ (.Y(_2194_),
    .A(_2166_),
    .B(_2167_));
 sg13g2_xnor2_1 _6066_ (.Y(_2195_),
    .A(_2192_),
    .B(_2194_));
 sg13g2_xnor2_1 _6067_ (.Y(_2196_),
    .A(_2171_),
    .B(_2195_));
 sg13g2_nand2b_1 _6068_ (.Y(_2197_),
    .B(_2196_),
    .A_N(_1904_));
 sg13g2_o21ai_1 _6069_ (.B1(_2197_),
    .Y(_2198_),
    .A1(_1658_),
    .A2(_1903_));
 sg13g2_nand2_1 _6070_ (.Y(_2199_),
    .A(_2163_),
    .B(_2192_));
 sg13g2_a21oi_1 _6071_ (.A1(_2133_),
    .A2(_2191_),
    .Y(_2200_),
    .B1(_2190_));
 sg13g2_o21ai_1 _6072_ (.B1(_2186_),
    .Y(_2201_),
    .A1(_2173_),
    .A2(_2188_));
 sg13g2_a21o_1 _6073_ (.A2(_2178_),
    .A1(_2141_),
    .B1(_2184_),
    .X(_2202_));
 sg13g2_a22oi_1 _6074_ (.Y(_2203_),
    .B1(_2177_),
    .B2(_2150_),
    .A2(_2175_),
    .A1(_2140_));
 sg13g2_and2_1 _6075_ (.A(net585),
    .B(net575),
    .X(_2204_));
 sg13g2_and2_1 _6076_ (.A(_2175_),
    .B(_2204_),
    .X(_2205_));
 sg13g2_xnor2_1 _6077_ (.Y(_2206_),
    .A(_2175_),
    .B(_2204_));
 sg13g2_nor2_1 _6078_ (.A(_2151_),
    .B(_2206_),
    .Y(_2207_));
 sg13g2_xnor2_1 _6079_ (.Y(_2208_),
    .A(_2151_),
    .B(_2206_));
 sg13g2_xor2_1 _6080_ (.B(_2208_),
    .A(_2203_),
    .X(_2209_));
 sg13g2_mux2_1 _6081_ (.A0(_2030_),
    .A1(_2093_),
    .S(_1978_),
    .X(_2210_));
 sg13g2_nor2b_1 _6082_ (.A(net570),
    .B_N(_2210_),
    .Y(_2211_));
 sg13g2_xnor2_1 _6083_ (.Y(_2212_),
    .A(net570),
    .B(_2210_));
 sg13g2_nand2_1 _6084_ (.Y(_2213_),
    .A(_2209_),
    .B(_2212_));
 sg13g2_xnor2_1 _6085_ (.Y(_2214_),
    .A(_2209_),
    .B(_2212_));
 sg13g2_nand2b_1 _6086_ (.Y(_2215_),
    .B(_2202_),
    .A_N(_2214_));
 sg13g2_xor2_1 _6087_ (.B(_2214_),
    .A(_2202_),
    .X(_2216_));
 sg13g2_xor2_1 _6088_ (.B(_2216_),
    .A(_2182_),
    .X(_2217_));
 sg13g2_nand2_1 _6089_ (.Y(_2218_),
    .A(_2201_),
    .B(_2217_));
 sg13g2_xnor2_1 _6090_ (.Y(_2219_),
    .A(_2201_),
    .B(_2217_));
 sg13g2_nor2_1 _6091_ (.A(_2200_),
    .B(_2219_),
    .Y(_2220_));
 sg13g2_xor2_1 _6092_ (.B(_2219_),
    .A(_2200_),
    .X(_2221_));
 sg13g2_nand2b_1 _6093_ (.Y(_2222_),
    .B(_2221_),
    .A_N(_2199_));
 sg13g2_xnor2_1 _6094_ (.Y(_2223_),
    .A(_2199_),
    .B(_2221_));
 sg13g2_nor2_1 _6095_ (.A(_2163_),
    .B(_2193_),
    .Y(_2224_));
 sg13g2_a22oi_1 _6096_ (.Y(_2225_),
    .B1(_2224_),
    .B2(_2192_),
    .A2(_2195_),
    .A1(_2171_));
 sg13g2_nand2b_1 _6097_ (.Y(_2226_),
    .B(_2223_),
    .A_N(_2225_));
 sg13g2_xnor2_1 _6098_ (.Y(_2227_),
    .A(_2223_),
    .B(_2225_));
 sg13g2_nand2_1 _6099_ (.Y(_2228_),
    .A(_1962_),
    .B(_2227_));
 sg13g2_nor2_1 _6100_ (.A(_1962_),
    .B(_2227_),
    .Y(_2229_));
 sg13g2_a221oi_1 _6101_ (.B2(_2228_),
    .C1(_2229_),
    .B1(_2198_),
    .A1(_1904_),
    .Y(_2230_),
    .A2(_1962_));
 sg13g2_o21ai_1 _6102_ (.B1(_2215_),
    .Y(_2231_),
    .A1(_2182_),
    .A2(_2216_));
 sg13g2_o21ai_1 _6103_ (.B1(_2213_),
    .Y(_2232_),
    .A1(_2203_),
    .A2(_2208_));
 sg13g2_o21ai_1 _6104_ (.B1(net575),
    .Y(_2233_),
    .A1(net584),
    .A2(_1987_));
 sg13g2_a21oi_1 _6105_ (.A1(_1987_),
    .A2(_2204_),
    .Y(_2234_),
    .B1(_2233_));
 sg13g2_xnor2_1 _6106_ (.Y(_2235_),
    .A(_2151_),
    .B(_2234_));
 sg13g2_o21ai_1 _6107_ (.B1(_2235_),
    .Y(_2236_),
    .A1(_2205_),
    .A2(_2207_));
 sg13g2_or3_1 _6108_ (.A(_2205_),
    .B(_2207_),
    .C(_2235_),
    .X(_2237_));
 sg13g2_nand2_1 _6109_ (.Y(_2238_),
    .A(_2236_),
    .B(_2237_));
 sg13g2_a21oi_1 _6110_ (.A1(_1979_),
    .A2(_2093_),
    .Y(_2239_),
    .B1(_2124_));
 sg13g2_or2_1 _6111_ (.X(_2240_),
    .B(_2239_),
    .A(net570));
 sg13g2_xor2_1 _6112_ (.B(_2239_),
    .A(net570),
    .X(_2241_));
 sg13g2_inv_1 _6113_ (.Y(_2242_),
    .A(_2241_));
 sg13g2_xnor2_1 _6114_ (.Y(_2243_),
    .A(_2238_),
    .B(_2241_));
 sg13g2_xor2_1 _6115_ (.B(_2243_),
    .A(_2232_),
    .X(_2244_));
 sg13g2_and2_1 _6116_ (.A(_2211_),
    .B(_2244_),
    .X(_2245_));
 sg13g2_xnor2_1 _6117_ (.Y(_2246_),
    .A(_2211_),
    .B(_2244_));
 sg13g2_nand2b_1 _6118_ (.Y(_2247_),
    .B(_2231_),
    .A_N(_2246_));
 sg13g2_xor2_1 _6119_ (.B(_2246_),
    .A(_2231_),
    .X(_2248_));
 sg13g2_nor2_1 _6120_ (.A(_2218_),
    .B(_2248_),
    .Y(_2249_));
 sg13g2_xor2_1 _6121_ (.B(_2248_),
    .A(_2218_),
    .X(_2250_));
 sg13g2_xnor2_1 _6122_ (.Y(_2251_),
    .A(_2220_),
    .B(_2250_));
 sg13g2_a21oi_1 _6123_ (.A1(_2222_),
    .A2(_2226_),
    .Y(_2252_),
    .B1(_2251_));
 sg13g2_nand3_1 _6124_ (.B(_2226_),
    .C(_2251_),
    .A(_2222_),
    .Y(_2253_));
 sg13g2_nand2b_2 _6125_ (.Y(_2254_),
    .B(_2253_),
    .A_N(_2252_));
 sg13g2_a21o_1 _6126_ (.A2(_1961_),
    .A1(_1904_),
    .B1(_1960_),
    .X(_2255_));
 sg13g2_o21ai_1 _6127_ (.B1(_1952_),
    .Y(_2256_),
    .A1(_1532_),
    .A2(_1953_));
 sg13g2_o21ai_1 _6128_ (.B1(_1950_),
    .Y(_2257_),
    .A1(_1936_),
    .A2(_1948_));
 sg13g2_or3_1 _6129_ (.A(_1446_),
    .B(_1460_),
    .C(_1519_),
    .X(_2258_));
 sg13g2_a22oi_1 _6130_ (.Y(_2259_),
    .B1(_2258_),
    .B2(_1434_),
    .A2(_1519_),
    .A1(_1460_));
 sg13g2_a21oi_2 _6131_ (.B1(_1943_),
    .Y(_2260_),
    .A2(_1947_),
    .A1(_1944_));
 sg13g2_a21oi_2 _6132_ (.B1(_1939_),
    .Y(_2261_),
    .A2(_1941_),
    .A1(_1516_));
 sg13g2_o21ai_1 _6133_ (.B1(net568),
    .Y(_2262_),
    .A1(net598),
    .A2(net594));
 sg13g2_nor2_1 _6134_ (.A(_0455_),
    .B(_1938_),
    .Y(_2263_));
 sg13g2_nor2_1 _6135_ (.A(_2262_),
    .B(_2263_),
    .Y(_2264_));
 sg13g2_xnor2_1 _6136_ (.Y(_2265_),
    .A(_1517_),
    .B(_2264_));
 sg13g2_nor2b_2 _6137_ (.A(_2261_),
    .B_N(_2265_),
    .Y(_2266_));
 sg13g2_xnor2_1 _6138_ (.Y(_2267_),
    .A(_2261_),
    .B(_2265_));
 sg13g2_nor2_1 _6139_ (.A(_1446_),
    .B(_1458_),
    .Y(_2268_));
 sg13g2_nor2_1 _6140_ (.A(_1484_),
    .B(_1520_),
    .Y(_2269_));
 sg13g2_and2_1 _6141_ (.A(_1484_),
    .B(_1520_),
    .X(_2270_));
 sg13g2_nor2_1 _6142_ (.A(_2269_),
    .B(_2270_),
    .Y(_2271_));
 sg13g2_xor2_1 _6143_ (.B(_2271_),
    .A(_2268_),
    .X(_2272_));
 sg13g2_xnor2_1 _6144_ (.Y(_2273_),
    .A(_2267_),
    .B(_2272_));
 sg13g2_xor2_1 _6145_ (.B(_2273_),
    .A(_2260_),
    .X(_2274_));
 sg13g2_nand2b_1 _6146_ (.Y(_2275_),
    .B(_2274_),
    .A_N(_2259_));
 sg13g2_xnor2_1 _6147_ (.Y(_2276_),
    .A(_2259_),
    .B(_2274_));
 sg13g2_nand2_1 _6148_ (.Y(_2277_),
    .A(_2257_),
    .B(_2276_));
 sg13g2_xnor2_1 _6149_ (.Y(_2278_),
    .A(_2257_),
    .B(_2276_));
 sg13g2_nand2b_1 _6150_ (.Y(_2279_),
    .B(_2256_),
    .A_N(_2278_));
 sg13g2_xor2_1 _6151_ (.B(_2278_),
    .A(_2256_),
    .X(_2280_));
 sg13g2_nor3_1 _6152_ (.A(_1932_),
    .B(_1954_),
    .C(_2280_),
    .Y(_2281_));
 sg13g2_xor2_1 _6153_ (.B(_2280_),
    .A(_1955_),
    .X(_2282_));
 sg13g2_nor3_1 _6154_ (.A(_1957_),
    .B(_1958_),
    .C(_2282_),
    .Y(_2283_));
 sg13g2_o21ai_1 _6155_ (.B1(_2282_),
    .Y(_2284_),
    .A1(_1957_),
    .A2(_1958_));
 sg13g2_nor2b_1 _6156_ (.A(_2283_),
    .B_N(_2284_),
    .Y(_2285_));
 sg13g2_nor2_1 _6157_ (.A(_1924_),
    .B(_1926_),
    .Y(_2286_));
 sg13g2_a21oi_1 _6158_ (.A1(_1909_),
    .A2(_1922_),
    .Y(_2287_),
    .B1(_1921_));
 sg13g2_or2_1 _6159_ (.X(_2288_),
    .B(_1917_),
    .A(_1744_));
 sg13g2_xnor2_1 _6160_ (.Y(_2289_),
    .A(_1744_),
    .B(_1917_));
 sg13g2_inv_1 _6161_ (.Y(_2290_),
    .A(_2289_));
 sg13g2_o21ai_1 _6162_ (.B1(_1915_),
    .Y(_2291_),
    .A1(_1775_),
    .A2(_1913_));
 sg13g2_o21ai_1 _6163_ (.B1(net567),
    .Y(_2292_),
    .A1(net593),
    .A2(net580));
 sg13g2_a21oi_1 _6164_ (.A1(_0458_),
    .A2(net593),
    .Y(_2293_),
    .B1(_2292_));
 sg13g2_xnor2_1 _6165_ (.Y(_2294_),
    .A(_1773_),
    .B(_2293_));
 sg13g2_and2_1 _6166_ (.A(_2291_),
    .B(_2294_),
    .X(_2295_));
 sg13g2_xnor2_1 _6167_ (.Y(_2296_),
    .A(_2291_),
    .B(_2294_));
 sg13g2_a22oi_1 _6168_ (.Y(_2297_),
    .B1(_1734_),
    .B2(_1661_),
    .A2(_1719_),
    .A1(_1669_));
 sg13g2_or2_1 _6169_ (.X(_2298_),
    .B(_2297_),
    .A(_2296_));
 sg13g2_xnor2_1 _6170_ (.Y(_2299_),
    .A(_2296_),
    .B(_2297_));
 sg13g2_nor2_1 _6171_ (.A(_1919_),
    .B(_2299_),
    .Y(_2300_));
 sg13g2_xor2_1 _6172_ (.B(_2299_),
    .A(_1919_),
    .X(_2301_));
 sg13g2_xnor2_1 _6173_ (.Y(_2302_),
    .A(_2289_),
    .B(_2301_));
 sg13g2_inv_1 _6174_ (.Y(_2303_),
    .A(_2302_));
 sg13g2_xnor2_1 _6175_ (.Y(_2304_),
    .A(_2287_),
    .B(_2302_));
 sg13g2_nand2b_1 _6176_ (.Y(_2305_),
    .B(_2304_),
    .A_N(_1907_));
 sg13g2_xnor2_1 _6177_ (.Y(_2306_),
    .A(_1907_),
    .B(_2304_));
 sg13g2_nand2b_1 _6178_ (.Y(_2307_),
    .B(_2306_),
    .A_N(_2286_));
 sg13g2_xor2_1 _6179_ (.B(_2306_),
    .A(_2286_),
    .X(_2308_));
 sg13g2_a21o_1 _6180_ (.A2(_1930_),
    .A1(_1928_),
    .B1(_2308_),
    .X(_2309_));
 sg13g2_nand3_1 _6181_ (.B(_1930_),
    .C(_2308_),
    .A(_1928_),
    .Y(_2310_));
 sg13g2_and3_1 _6182_ (.X(_2311_),
    .A(_2285_),
    .B(_2309_),
    .C(_2310_));
 sg13g2_nand3_1 _6183_ (.B(_2309_),
    .C(_2310_),
    .A(_2285_),
    .Y(_2312_));
 sg13g2_a21o_1 _6184_ (.A2(_2310_),
    .A1(_2309_),
    .B1(_2285_),
    .X(_2313_));
 sg13g2_and3_1 _6185_ (.X(_2314_),
    .A(_2255_),
    .B(_2312_),
    .C(_2313_));
 sg13g2_a21oi_1 _6186_ (.A1(_2312_),
    .A2(_2313_),
    .Y(_2315_),
    .B1(_2255_));
 sg13g2_nor3_1 _6187_ (.A(_2254_),
    .B(_2314_),
    .C(_2315_),
    .Y(_2316_));
 sg13g2_o21ai_1 _6188_ (.B1(_2254_),
    .Y(_2317_),
    .A1(_2314_),
    .A2(_2315_));
 sg13g2_nor2b_1 _6189_ (.A(_2316_),
    .B_N(_2317_),
    .Y(_2318_));
 sg13g2_nor2_1 _6190_ (.A(_2230_),
    .B(_2318_),
    .Y(_2319_));
 sg13g2_a21oi_1 _6191_ (.A1(_2230_),
    .A2(_2318_),
    .Y(_2320_),
    .B1(net741));
 sg13g2_nor2b_1 _6192_ (.A(_2319_),
    .B_N(_2320_),
    .Y(_0198_));
 sg13g2_a21oi_1 _6193_ (.A1(_2230_),
    .A2(_2317_),
    .Y(_2321_),
    .B1(_2316_));
 sg13g2_a21oi_1 _6194_ (.A1(_2220_),
    .A2(_2250_),
    .Y(_2322_),
    .B1(_2252_));
 sg13g2_a21oi_1 _6195_ (.A1(_2232_),
    .A2(_2243_),
    .Y(_2323_),
    .B1(_2245_));
 sg13g2_o21ai_1 _6196_ (.B1(_2236_),
    .Y(_2324_),
    .A1(_2238_),
    .A2(_2242_));
 sg13g2_nor2_1 _6197_ (.A(_1978_),
    .B(_2120_),
    .Y(_2325_));
 sg13g2_a21oi_1 _6198_ (.A1(net587),
    .A2(net575),
    .Y(_2326_),
    .B1(_2325_));
 sg13g2_nor2_1 _6199_ (.A(net570),
    .B(_2326_),
    .Y(_2327_));
 sg13g2_xnor2_1 _6200_ (.Y(_2328_),
    .A(net570),
    .B(_2326_));
 sg13g2_nand2_1 _6201_ (.Y(_2329_),
    .A(_2151_),
    .B(_2233_));
 sg13g2_nand2_2 _6202_ (.Y(_2330_),
    .A(_2236_),
    .B(_2329_));
 sg13g2_xor2_1 _6203_ (.B(_2330_),
    .A(_2328_),
    .X(_2331_));
 sg13g2_xnor2_1 _6204_ (.Y(_2332_),
    .A(_2324_),
    .B(_2331_));
 sg13g2_nor2_1 _6205_ (.A(_2240_),
    .B(_2332_),
    .Y(_2333_));
 sg13g2_xnor2_1 _6206_ (.Y(_2334_),
    .A(_2240_),
    .B(_2332_));
 sg13g2_xor2_1 _6207_ (.B(_2334_),
    .A(_2323_),
    .X(_2335_));
 sg13g2_nor2b_1 _6208_ (.A(_2247_),
    .B_N(_2335_),
    .Y(_2336_));
 sg13g2_xnor2_1 _6209_ (.Y(_2337_),
    .A(_2247_),
    .B(_2335_));
 sg13g2_and2_1 _6210_ (.A(_2249_),
    .B(_2337_),
    .X(_2338_));
 sg13g2_xnor2_1 _6211_ (.Y(_2339_),
    .A(_2249_),
    .B(_2337_));
 sg13g2_xor2_1 _6212_ (.B(_2339_),
    .A(_2322_),
    .X(_2340_));
 sg13g2_a21oi_1 _6213_ (.A1(_2255_),
    .A2(_2313_),
    .Y(_2341_),
    .B1(_2311_));
 sg13g2_o21ai_1 _6214_ (.B1(_2275_),
    .Y(_2342_),
    .A1(_2260_),
    .A2(_2273_));
 sg13g2_a21oi_1 _6215_ (.A1(net588),
    .A2(_2270_),
    .Y(_2343_),
    .B1(_1458_));
 sg13g2_nor2_1 _6216_ (.A(_2269_),
    .B(_2343_),
    .Y(_2344_));
 sg13g2_a21oi_2 _6217_ (.B1(_2266_),
    .Y(_2345_),
    .A2(_2272_),
    .A1(_2267_));
 sg13g2_a21oi_2 _6218_ (.B1(_2266_),
    .Y(_2346_),
    .A2(_2262_),
    .A1(_1517_));
 sg13g2_nand2_1 _6219_ (.Y(_2347_),
    .A(net588),
    .B(_1483_));
 sg13g2_o21ai_1 _6220_ (.B1(net568),
    .Y(_2348_),
    .A1(net655),
    .A2(net581));
 sg13g2_nor2_1 _6221_ (.A(_1543_),
    .B(_2348_),
    .Y(_2349_));
 sg13g2_xnor2_1 _6222_ (.Y(_2350_),
    .A(_2347_),
    .B(_2349_));
 sg13g2_xnor2_1 _6223_ (.Y(_2351_),
    .A(_2346_),
    .B(_2350_));
 sg13g2_xor2_1 _6224_ (.B(_2351_),
    .A(_2345_),
    .X(_2352_));
 sg13g2_nand2b_1 _6225_ (.Y(_2353_),
    .B(_2352_),
    .A_N(_2344_));
 sg13g2_xnor2_1 _6226_ (.Y(_2354_),
    .A(_2344_),
    .B(_2352_));
 sg13g2_nand2_1 _6227_ (.Y(_2355_),
    .A(_2342_),
    .B(_2354_));
 sg13g2_xnor2_1 _6228_ (.Y(_2356_),
    .A(_2342_),
    .B(_2354_));
 sg13g2_nor2_1 _6229_ (.A(_2277_),
    .B(_2356_),
    .Y(_2357_));
 sg13g2_xor2_1 _6230_ (.B(_2356_),
    .A(_2277_),
    .X(_2358_));
 sg13g2_nand2b_1 _6231_ (.Y(_2359_),
    .B(_2358_),
    .A_N(_2279_));
 sg13g2_xnor2_1 _6232_ (.Y(_2360_),
    .A(_2279_),
    .B(_2358_));
 sg13g2_o21ai_1 _6233_ (.B1(_2360_),
    .Y(_2361_),
    .A1(_2281_),
    .A2(_2283_));
 sg13g2_or3_1 _6234_ (.A(_2281_),
    .B(_2283_),
    .C(_2360_),
    .X(_2362_));
 sg13g2_and2_1 _6235_ (.A(_2361_),
    .B(_2362_),
    .X(_2363_));
 sg13g2_o21ai_1 _6236_ (.B1(_2305_),
    .Y(_2364_),
    .A1(_2287_),
    .A2(_2303_));
 sg13g2_a21oi_1 _6237_ (.A1(_2290_),
    .A2(_2301_),
    .Y(_2365_),
    .B1(_2300_));
 sg13g2_nor2_1 _6238_ (.A(_1743_),
    .B(_2295_),
    .Y(_2366_));
 sg13g2_xnor2_1 _6239_ (.Y(_2367_),
    .A(_1743_),
    .B(_2295_));
 sg13g2_inv_1 _6240_ (.Y(_2368_),
    .A(_2367_));
 sg13g2_a21oi_2 _6241_ (.B1(_2295_),
    .Y(_2369_),
    .A2(_2292_),
    .A1(_1773_));
 sg13g2_and2_1 _6242_ (.A(_1669_),
    .B(_1734_),
    .X(_2370_));
 sg13g2_a21o_1 _6243_ (.A2(net567),
    .A1(_1661_),
    .B1(_2370_),
    .X(_2371_));
 sg13g2_xor2_1 _6244_ (.B(_2371_),
    .A(_2369_),
    .X(_2372_));
 sg13g2_nor2b_1 _6245_ (.A(_2298_),
    .B_N(_2372_),
    .Y(_2373_));
 sg13g2_xnor2_1 _6246_ (.Y(_2374_),
    .A(_2298_),
    .B(_2372_));
 sg13g2_xnor2_1 _6247_ (.Y(_2375_),
    .A(_2367_),
    .B(_2374_));
 sg13g2_nand2b_1 _6248_ (.Y(_2376_),
    .B(_2375_),
    .A_N(_2365_));
 sg13g2_xnor2_1 _6249_ (.Y(_2377_),
    .A(_2365_),
    .B(_2375_));
 sg13g2_nand2b_1 _6250_ (.Y(_2378_),
    .B(_2377_),
    .A_N(_2288_));
 sg13g2_xnor2_1 _6251_ (.Y(_2379_),
    .A(_2288_),
    .B(_2377_));
 sg13g2_xnor2_1 _6252_ (.Y(_2380_),
    .A(_2364_),
    .B(_2379_));
 sg13g2_a21o_1 _6253_ (.A2(_2309_),
    .A1(_2307_),
    .B1(_2380_),
    .X(_2381_));
 sg13g2_nand3_1 _6254_ (.B(_2309_),
    .C(_2380_),
    .A(_2307_),
    .Y(_2382_));
 sg13g2_nand3_1 _6255_ (.B(_2381_),
    .C(_2382_),
    .A(_2363_),
    .Y(_2383_));
 sg13g2_a21oi_1 _6256_ (.A1(_2381_),
    .A2(_2382_),
    .Y(_2384_),
    .B1(_2363_));
 sg13g2_a21o_1 _6257_ (.A2(_2382_),
    .A1(_2381_),
    .B1(_2363_),
    .X(_2385_));
 sg13g2_a21oi_1 _6258_ (.A1(_2383_),
    .A2(_2385_),
    .Y(_2386_),
    .B1(_2341_));
 sg13g2_and3_1 _6259_ (.X(_2387_),
    .A(_2341_),
    .B(_2383_),
    .C(_2385_));
 sg13g2_nor3_1 _6260_ (.A(_2340_),
    .B(_2386_),
    .C(_2387_),
    .Y(_2388_));
 sg13g2_o21ai_1 _6261_ (.B1(_2340_),
    .Y(_2389_),
    .A1(_2386_),
    .A2(_2387_));
 sg13g2_nand2b_1 _6262_ (.Y(_2390_),
    .B(_2389_),
    .A_N(_2388_));
 sg13g2_o21ai_1 _6263_ (.B1(net749),
    .Y(_2391_),
    .A1(_2321_),
    .A2(_2390_));
 sg13g2_a21oi_1 _6264_ (.A1(_2321_),
    .A2(_2390_),
    .Y(_0199_),
    .B1(_2391_));
 sg13g2_o21ai_1 _6265_ (.B1(_2389_),
    .Y(_2392_),
    .A1(_2321_),
    .A2(_2388_));
 sg13g2_inv_1 _6266_ (.Y(_2393_),
    .A(_2392_));
 sg13g2_a21oi_1 _6267_ (.A1(_2324_),
    .A2(_2331_),
    .Y(_2394_),
    .B1(_2333_));
 sg13g2_o21ai_1 _6268_ (.B1(_2236_),
    .Y(_2395_),
    .A1(_2328_),
    .A2(_2330_));
 sg13g2_nand2_1 _6269_ (.Y(_2396_),
    .A(net604),
    .B(net575));
 sg13g2_xor2_1 _6270_ (.B(_2396_),
    .A(_2330_),
    .X(_2397_));
 sg13g2_xnor2_1 _6271_ (.Y(_2398_),
    .A(_2395_),
    .B(_2397_));
 sg13g2_xnor2_1 _6272_ (.Y(_2399_),
    .A(_2327_),
    .B(_2398_));
 sg13g2_o21ai_1 _6273_ (.B1(_2394_),
    .Y(_2400_),
    .A1(_2323_),
    .A2(_2334_));
 sg13g2_nor4_1 _6274_ (.A(_2336_),
    .B(_2338_),
    .C(_2399_),
    .D(_2400_),
    .Y(_2401_));
 sg13g2_o21ai_1 _6275_ (.B1(_2401_),
    .Y(_2402_),
    .A1(_2322_),
    .A2(_2339_));
 sg13g2_o21ai_1 _6276_ (.B1(_2353_),
    .Y(_2403_),
    .A1(_2345_),
    .A2(_2351_));
 sg13g2_nand2_1 _6277_ (.Y(_2404_),
    .A(net589),
    .B(_2348_));
 sg13g2_a21oi_2 _6278_ (.B1(_1543_),
    .Y(_2405_),
    .A2(_2404_),
    .A1(_1483_));
 sg13g2_a21oi_1 _6279_ (.A1(_2346_),
    .A2(_2350_),
    .Y(_2406_),
    .B1(_2266_));
 sg13g2_nand2_1 _6280_ (.Y(_2407_),
    .A(net588),
    .B(_1515_));
 sg13g2_xnor2_1 _6281_ (.Y(_2408_),
    .A(_2349_),
    .B(_2407_));
 sg13g2_xor2_1 _6282_ (.B(_2408_),
    .A(_2346_),
    .X(_2409_));
 sg13g2_nand2b_1 _6283_ (.Y(_2410_),
    .B(_2409_),
    .A_N(_2406_));
 sg13g2_xnor2_1 _6284_ (.Y(_2411_),
    .A(_2406_),
    .B(_2409_));
 sg13g2_nand2b_1 _6285_ (.Y(_2412_),
    .B(_2411_),
    .A_N(_2405_));
 sg13g2_xnor2_1 _6286_ (.Y(_2413_),
    .A(_2405_),
    .B(_2411_));
 sg13g2_xor2_1 _6287_ (.B(_2413_),
    .A(_2403_),
    .X(_2414_));
 sg13g2_nor2b_1 _6288_ (.A(_2355_),
    .B_N(_2414_),
    .Y(_2415_));
 sg13g2_xor2_1 _6289_ (.B(_2414_),
    .A(_2355_),
    .X(_2416_));
 sg13g2_nor3_1 _6290_ (.A(_2277_),
    .B(_2356_),
    .C(_2416_),
    .Y(_2417_));
 sg13g2_xor2_1 _6291_ (.B(_2416_),
    .A(_2357_),
    .X(_2418_));
 sg13g2_a21oi_1 _6292_ (.A1(_2359_),
    .A2(_2361_),
    .Y(_2419_),
    .B1(_2418_));
 sg13g2_nand3_1 _6293_ (.B(_2361_),
    .C(_2418_),
    .A(_2359_),
    .Y(_2420_));
 sg13g2_nand2b_1 _6294_ (.Y(_2421_),
    .B(_2420_),
    .A_N(_2419_));
 sg13g2_a21oi_1 _6295_ (.A1(_2368_),
    .A2(_2374_),
    .Y(_2422_),
    .B1(_2373_));
 sg13g2_o21ai_1 _6296_ (.B1(net567),
    .Y(_2423_),
    .A1(net576),
    .A2(net578));
 sg13g2_xnor2_1 _6297_ (.Y(_2424_),
    .A(_2369_),
    .B(_2423_));
 sg13g2_a21oi_1 _6298_ (.A1(_2369_),
    .A2(_2371_),
    .Y(_2425_),
    .B1(_2424_));
 sg13g2_xnor2_1 _6299_ (.Y(_2426_),
    .A(_2422_),
    .B(_2425_));
 sg13g2_xnor2_1 _6300_ (.Y(_2427_),
    .A(_2366_),
    .B(_2426_));
 sg13g2_nand3_1 _6301_ (.B(_2378_),
    .C(_2427_),
    .A(_2376_),
    .Y(_2428_));
 sg13g2_a21oi_1 _6302_ (.A1(_2364_),
    .A2(_2379_),
    .Y(_2429_),
    .B1(_2428_));
 sg13g2_and2_1 _6303_ (.A(_2381_),
    .B(_2429_),
    .X(_2430_));
 sg13g2_nor2_1 _6304_ (.A(_2421_),
    .B(_2430_),
    .Y(_2431_));
 sg13g2_xor2_1 _6305_ (.B(_2430_),
    .A(_2421_),
    .X(_2432_));
 sg13g2_o21ai_1 _6306_ (.B1(_2383_),
    .Y(_2433_),
    .A1(_2341_),
    .A2(_2384_));
 sg13g2_xnor2_1 _6307_ (.Y(_2434_),
    .A(_2432_),
    .B(_2433_));
 sg13g2_nor2b_1 _6308_ (.A(_2434_),
    .B_N(_2402_),
    .Y(_2435_));
 sg13g2_xnor2_1 _6309_ (.Y(_2436_),
    .A(_2402_),
    .B(_2434_));
 sg13g2_inv_1 _6310_ (.Y(_2437_),
    .A(_2436_));
 sg13g2_o21ai_1 _6311_ (.B1(net749),
    .Y(_2438_),
    .A1(_2393_),
    .A2(_2437_));
 sg13g2_a21oi_1 _6312_ (.A1(_2393_),
    .A2(_2437_),
    .Y(_0200_),
    .B1(_2438_));
 sg13g2_a21oi_1 _6313_ (.A1(_2392_),
    .A2(_2436_),
    .Y(_2439_),
    .B1(_2435_));
 sg13g2_a21oi_1 _6314_ (.A1(_2432_),
    .A2(_2433_),
    .Y(_2440_),
    .B1(_2431_));
 sg13g2_nand2_1 _6315_ (.Y(_2441_),
    .A(_2410_),
    .B(_2412_));
 sg13g2_o21ai_1 _6316_ (.B1(_2348_),
    .Y(_2442_),
    .A1(net588),
    .A2(_1514_));
 sg13g2_nor3_1 _6317_ (.A(_2266_),
    .B(_2346_),
    .C(_2408_),
    .Y(_2443_));
 sg13g2_a21o_1 _6318_ (.A2(_2408_),
    .A1(_2266_),
    .B1(_2443_),
    .X(_2444_));
 sg13g2_xor2_1 _6319_ (.B(_2444_),
    .A(_2442_),
    .X(_2445_));
 sg13g2_xnor2_1 _6320_ (.Y(_2446_),
    .A(_2441_),
    .B(_2445_));
 sg13g2_a21o_1 _6321_ (.A2(_2413_),
    .A1(_2403_),
    .B1(_2417_),
    .X(_2447_));
 sg13g2_nor4_2 _6322_ (.A(_2415_),
    .B(_2419_),
    .C(_2446_),
    .Y(_2448_),
    .D(_2447_));
 sg13g2_xor2_1 _6323_ (.B(_2448_),
    .A(net567),
    .X(_2449_));
 sg13g2_xnor2_1 _6324_ (.Y(_2450_),
    .A(_2440_),
    .B(_2449_));
 sg13g2_or2_1 _6325_ (.X(_2451_),
    .B(_2450_),
    .A(_2149_));
 sg13g2_xnor2_1 _6326_ (.Y(_2452_),
    .A(_2149_),
    .B(_2450_));
 sg13g2_o21ai_1 _6327_ (.B1(net749),
    .Y(_2453_),
    .A1(_2439_),
    .A2(_2452_));
 sg13g2_a21oi_1 _6328_ (.A1(_2439_),
    .A2(_2452_),
    .Y(_0201_),
    .B1(_2453_));
 sg13g2_o21ai_1 _6329_ (.B1(_2451_),
    .Y(_2454_),
    .A1(_2439_),
    .A2(_2452_));
 sg13g2_a21oi_1 _6330_ (.A1(_1742_),
    .A2(_2448_),
    .Y(_2455_),
    .B1(net568));
 sg13g2_o21ai_1 _6331_ (.B1(net568),
    .Y(_2456_),
    .A1(_1742_),
    .A2(_2448_));
 sg13g2_nand2b_1 _6332_ (.Y(_2457_),
    .B(_2456_),
    .A_N(_2440_));
 sg13g2_nor2b_1 _6333_ (.A(_2455_),
    .B_N(_2457_),
    .Y(_2458_));
 sg13g2_nor2_1 _6334_ (.A(net575),
    .B(_2458_),
    .Y(_2459_));
 sg13g2_xnor2_1 _6335_ (.Y(_2460_),
    .A(_2149_),
    .B(_2458_));
 sg13g2_a21oi_1 _6336_ (.A1(_2454_),
    .A2(_2460_),
    .Y(_2461_),
    .B1(net742));
 sg13g2_nor2_1 _6337_ (.A(_2454_),
    .B(_2460_),
    .Y(_2462_));
 sg13g2_nor2b_1 _6338_ (.A(_2462_),
    .B_N(_2461_),
    .Y(_0202_));
 sg13g2_nor2b_1 _6339_ (.A(_2459_),
    .B_N(_2461_),
    .Y(_0203_));
 sg13g2_nor2_1 _6340_ (.A(net680),
    .B(_0061_),
    .Y(_2463_));
 sg13g2_a21oi_1 _6341_ (.A1(net680),
    .A2(_2861_),
    .Y(_2464_),
    .B1(_2463_));
 sg13g2_nor2b_1 _6342_ (.A(_2464_),
    .B_N(net677),
    .Y(_2465_));
 sg13g2_a221oi_1 _6343_ (.B2(net700),
    .C1(_2465_),
    .B1(_0827_),
    .A1(\generated._562[1] ),
    .Y(_2466_),
    .A2(_0656_));
 sg13g2_xor2_1 _6344_ (.B(_2466_),
    .A(net686),
    .X(_2467_));
 sg13g2_nor2_1 _6345_ (.A(net638),
    .B(_2467_),
    .Y(_0205_));
 sg13g2_nor2_1 _6346_ (.A(net436),
    .B(_2466_),
    .Y(_2468_));
 sg13g2_nand2_1 _6347_ (.Y(_2469_),
    .A(net680),
    .B(_0066_));
 sg13g2_o21ai_1 _6348_ (.B1(_2469_),
    .Y(_2470_),
    .A1(net680),
    .A2(_2861_));
 sg13g2_nand2_1 _6349_ (.Y(_2471_),
    .A(_0057_),
    .B(_0827_));
 sg13g2_a22oi_1 _6350_ (.Y(_2472_),
    .B1(_2470_),
    .B2(net677),
    .A2(_0656_),
    .A1(_0061_));
 sg13g2_nand2_1 _6351_ (.Y(_2473_),
    .A(_2471_),
    .B(_2472_));
 sg13g2_nor2_1 _6352_ (.A(net657),
    .B(_2466_),
    .Y(_2474_));
 sg13g2_xnor2_1 _6353_ (.Y(_2475_),
    .A(_2473_),
    .B(_2474_));
 sg13g2_xnor2_1 _6354_ (.Y(_2476_),
    .A(_0058_),
    .B(_2475_));
 sg13g2_and2_1 _6355_ (.A(_2468_),
    .B(_2476_),
    .X(_2477_));
 sg13g2_o21ai_1 _6356_ (.B1(net633),
    .Y(_2478_),
    .A1(_2468_),
    .A2(_2476_));
 sg13g2_nor2_1 _6357_ (.A(_2477_),
    .B(net437),
    .Y(_0206_));
 sg13g2_a21oi_1 _6358_ (.A1(\generated._512[0] ),
    .A2(_2475_),
    .Y(_2479_),
    .B1(_2477_));
 sg13g2_a21oi_1 _6359_ (.A1(_2466_),
    .A2(_2473_),
    .Y(_2480_),
    .B1(net657));
 sg13g2_mux2_1 _6360_ (.A0(_0066_),
    .A1(_0068_),
    .S(net680),
    .X(_2481_));
 sg13g2_mux2_1 _6361_ (.A0(_2464_),
    .A1(_2481_),
    .S(net677),
    .X(_2482_));
 sg13g2_xnor2_1 _6362_ (.Y(_2483_),
    .A(_2480_),
    .B(_2482_));
 sg13g2_xnor2_1 _6363_ (.Y(_2484_),
    .A(net531),
    .B(_2483_));
 sg13g2_nor2_1 _6364_ (.A(_2479_),
    .B(_2484_),
    .Y(_2485_));
 sg13g2_a21oi_1 _6365_ (.A1(_2479_),
    .A2(_2484_),
    .Y(_2486_),
    .B1(net637));
 sg13g2_nor2b_1 _6366_ (.A(_2485_),
    .B_N(_2486_),
    .Y(_0207_));
 sg13g2_a21oi_1 _6367_ (.A1(_2857_),
    .A2(_2483_),
    .Y(_2487_),
    .B1(_2485_));
 sg13g2_nand3_1 _6368_ (.B(_2473_),
    .C(_2482_),
    .A(_2466_),
    .Y(_2488_));
 sg13g2_nand2_1 _6369_ (.Y(_2489_),
    .A(net685),
    .B(_2488_));
 sg13g2_nor2_1 _6370_ (.A(net676),
    .B(_2470_),
    .Y(_2490_));
 sg13g2_nor2b_1 _6371_ (.A(net681),
    .B_N(_0068_),
    .Y(_2491_));
 sg13g2_a21oi_1 _6372_ (.A1(net681),
    .A2(_0070_),
    .Y(_2492_),
    .B1(_2491_));
 sg13g2_a21oi_1 _6373_ (.A1(net676),
    .A2(_2492_),
    .Y(_2493_),
    .B1(_2490_));
 sg13g2_xnor2_1 _6374_ (.Y(_2494_),
    .A(_2489_),
    .B(_2493_));
 sg13g2_nor2b_1 _6375_ (.A(_2494_),
    .B_N(\generated._512[2] ),
    .Y(_2495_));
 sg13g2_xnor2_1 _6376_ (.Y(_2496_),
    .A(net493),
    .B(_2494_));
 sg13g2_nor2b_1 _6377_ (.A(_2496_),
    .B_N(_2487_),
    .Y(_2497_));
 sg13g2_nor2b_1 _6378_ (.A(_2487_),
    .B_N(_2496_),
    .Y(_2498_));
 sg13g2_nor3_1 _6379_ (.A(net637),
    .B(_2497_),
    .C(_2498_),
    .Y(_0208_));
 sg13g2_or2_1 _6380_ (.X(_2499_),
    .B(_2498_),
    .A(_2495_));
 sg13g2_nand2b_1 _6381_ (.Y(_2500_),
    .B(_2493_),
    .A_N(_2488_));
 sg13g2_nand2_1 _6382_ (.Y(_2501_),
    .A(net685),
    .B(_2500_));
 sg13g2_nor2_1 _6383_ (.A(net676),
    .B(_2481_),
    .Y(_2502_));
 sg13g2_nor2b_1 _6384_ (.A(net681),
    .B_N(_0070_),
    .Y(_2503_));
 sg13g2_a21oi_1 _6385_ (.A1(net681),
    .A2(_0072_),
    .Y(_2504_),
    .B1(_2503_));
 sg13g2_a21oi_1 _6386_ (.A1(net675),
    .A2(_2504_),
    .Y(_2505_),
    .B1(_2502_));
 sg13g2_xnor2_1 _6387_ (.Y(_2506_),
    .A(_2501_),
    .B(_2505_));
 sg13g2_xnor2_1 _6388_ (.Y(_2507_),
    .A(net541),
    .B(_2506_));
 sg13g2_nor2_1 _6389_ (.A(_2499_),
    .B(_2507_),
    .Y(_2508_));
 sg13g2_and2_1 _6390_ (.A(_2499_),
    .B(_2507_),
    .X(_2509_));
 sg13g2_nor3_1 _6391_ (.A(net637),
    .B(_2508_),
    .C(_2509_),
    .Y(_0209_));
 sg13g2_nor2_1 _6392_ (.A(net558),
    .B(_2506_),
    .Y(_2510_));
 sg13g2_nor2b_1 _6393_ (.A(_2500_),
    .B_N(_2505_),
    .Y(_2511_));
 sg13g2_nor2_1 _6394_ (.A(net657),
    .B(_2511_),
    .Y(_2512_));
 sg13g2_nor2_1 _6395_ (.A(net683),
    .B(_0072_),
    .Y(_2513_));
 sg13g2_a21oi_1 _6396_ (.A1(net683),
    .A2(_2862_),
    .Y(_2514_),
    .B1(_2513_));
 sg13g2_nand2_1 _6397_ (.Y(_2515_),
    .A(net675),
    .B(_2514_));
 sg13g2_o21ai_1 _6398_ (.B1(_2515_),
    .Y(_2516_),
    .A1(net675),
    .A2(_2492_));
 sg13g2_xor2_1 _6399_ (.B(_2516_),
    .A(_2512_),
    .X(_2517_));
 sg13g2_xnor2_1 _6400_ (.Y(_2518_),
    .A(\generated._512[4] ),
    .B(_2517_));
 sg13g2_or3_1 _6401_ (.A(_2509_),
    .B(_2510_),
    .C(_2518_),
    .X(_2519_));
 sg13g2_o21ai_1 _6402_ (.B1(_2518_),
    .Y(_2520_),
    .A1(_2509_),
    .A2(_2510_));
 sg13g2_and3_1 _6403_ (.X(_0210_),
    .A(net633),
    .B(_2519_),
    .C(_2520_));
 sg13g2_o21ai_1 _6404_ (.B1(_2520_),
    .Y(_2521_),
    .A1(_2859_),
    .A2(_2517_));
 sg13g2_a21oi_1 _6405_ (.A1(_2511_),
    .A2(_2516_),
    .Y(_2522_),
    .B1(net657));
 sg13g2_nand2_1 _6406_ (.Y(_2523_),
    .A(net679),
    .B(_0074_));
 sg13g2_o21ai_1 _6407_ (.B1(_2523_),
    .Y(_2524_),
    .A1(net679),
    .A2(_2862_));
 sg13g2_nand2_1 _6408_ (.Y(_2525_),
    .A(net678),
    .B(_2524_));
 sg13g2_o21ai_1 _6409_ (.B1(_2525_),
    .Y(_2526_),
    .A1(net675),
    .A2(_2504_));
 sg13g2_xor2_1 _6410_ (.B(_2526_),
    .A(_2522_),
    .X(_2527_));
 sg13g2_xnor2_1 _6411_ (.Y(_2528_),
    .A(net473),
    .B(_2527_));
 sg13g2_nor2_1 _6412_ (.A(_2521_),
    .B(_2528_),
    .Y(_2529_));
 sg13g2_and2_1 _6413_ (.A(_2521_),
    .B(_2528_),
    .X(_2530_));
 sg13g2_nor3_1 _6414_ (.A(net638),
    .B(net474),
    .C(_2530_),
    .Y(_0211_));
 sg13g2_nor2_1 _6415_ (.A(net503),
    .B(_2527_),
    .Y(_2531_));
 sg13g2_nor2_1 _6416_ (.A(_2530_),
    .B(_2531_),
    .Y(_2532_));
 sg13g2_nor2b_1 _6417_ (.A(net674),
    .B_N(_2514_),
    .Y(_2533_));
 sg13g2_a21oi_2 _6418_ (.B1(_2533_),
    .Y(_2534_),
    .A2(_0074_),
    .A1(net673));
 sg13g2_nand3_1 _6419_ (.B(_2516_),
    .C(_2526_),
    .A(_2511_),
    .Y(_2535_));
 sg13g2_nand2_1 _6420_ (.Y(_2536_),
    .A(net685),
    .B(_2535_));
 sg13g2_xor2_1 _6421_ (.B(_2536_),
    .A(_2534_),
    .X(_2537_));
 sg13g2_xnor2_1 _6422_ (.Y(_2538_),
    .A(\generated._512[6] ),
    .B(_2537_));
 sg13g2_nor3_1 _6423_ (.A(_2530_),
    .B(_2531_),
    .C(_2538_),
    .Y(_2539_));
 sg13g2_nor2b_1 _6424_ (.A(_2532_),
    .B_N(_2538_),
    .Y(_2540_));
 sg13g2_nor3_1 _6425_ (.A(net638),
    .B(net504),
    .C(_2540_),
    .Y(_0212_));
 sg13g2_nor2_1 _6426_ (.A(net466),
    .B(_2537_),
    .Y(_2541_));
 sg13g2_nor2_1 _6427_ (.A(_2540_),
    .B(_2541_),
    .Y(_2542_));
 sg13g2_nor2b_1 _6428_ (.A(net673),
    .B_N(_2524_),
    .Y(_2543_));
 sg13g2_a21oi_1 _6429_ (.A1(net673),
    .A2(_0074_),
    .Y(_2544_),
    .B1(_2543_));
 sg13g2_o21ai_1 _6430_ (.B1(\generated._503 ),
    .Y(_2545_),
    .A1(_2534_),
    .A2(_2535_));
 sg13g2_xor2_1 _6431_ (.B(_2545_),
    .A(_2544_),
    .X(_2546_));
 sg13g2_xnor2_1 _6432_ (.Y(_2547_),
    .A(\generated._512[7] ),
    .B(_2546_));
 sg13g2_nor3_1 _6433_ (.A(_2540_),
    .B(_2541_),
    .C(_2547_),
    .Y(_2548_));
 sg13g2_nor2b_1 _6434_ (.A(_2542_),
    .B_N(_2547_),
    .Y(_2549_));
 sg13g2_nor3_1 _6435_ (.A(net638),
    .B(net467),
    .C(_2549_),
    .Y(_0213_));
 sg13g2_nor2_1 _6436_ (.A(net489),
    .B(_2546_),
    .Y(_2550_));
 sg13g2_nor2_1 _6437_ (.A(_2549_),
    .B(_2550_),
    .Y(_2551_));
 sg13g2_nor3_1 _6438_ (.A(_2534_),
    .B(_2535_),
    .C(_2544_),
    .Y(_2552_));
 sg13g2_nor2_1 _6439_ (.A(net685),
    .B(_0074_),
    .Y(_2553_));
 sg13g2_xnor2_1 _6440_ (.Y(_2554_),
    .A(\generated._562[9] ),
    .B(_2552_));
 sg13g2_a21oi_1 _6441_ (.A1(net684),
    .A2(_2554_),
    .Y(_2555_),
    .B1(_2553_));
 sg13g2_xor2_1 _6442_ (.B(_2555_),
    .A(\generated._511 ),
    .X(_2556_));
 sg13g2_o21ai_1 _6443_ (.B1(net633),
    .Y(_2557_),
    .A1(_2551_),
    .A2(_2556_));
 sg13g2_a21oi_1 _6444_ (.A1(_2551_),
    .A2(_2556_),
    .Y(_0214_),
    .B1(_2557_));
 sg13g2_and2_1 _6445_ (.A(net249),
    .B(_0592_),
    .X(_0215_));
 sg13g2_nor3_1 _6446_ (.A(net636),
    .B(_0595_),
    .C(_0827_),
    .Y(_0216_));
 sg13g2_nor2_1 _6447_ (.A(net666),
    .B(_0053_),
    .Y(_2558_));
 sg13g2_a21oi_1 _6448_ (.A1(net665),
    .A2(_2856_),
    .Y(_2559_),
    .B1(_2558_));
 sg13g2_nor2b_1 _6449_ (.A(_2559_),
    .B_N(net662),
    .Y(_2560_));
 sg13g2_nor2_2 _6450_ (.A(net667),
    .B(net664),
    .Y(_2561_));
 sg13g2_a221oi_1 _6451_ (.B2(net658),
    .C1(_2560_),
    .B1(_2561_),
    .A1(\generated._394[1] ),
    .Y(_2562_),
    .A2(_1068_));
 sg13g2_xor2_1 _6452_ (.B(_2562_),
    .A(net339),
    .X(_2563_));
 sg13g2_nor2_1 _6453_ (.A(net631),
    .B(_2563_),
    .Y(_0217_));
 sg13g2_nor2_1 _6454_ (.A(net406),
    .B(_2562_),
    .Y(_2564_));
 sg13g2_nand2_1 _6455_ (.Y(_2565_),
    .A(net666),
    .B(_0048_));
 sg13g2_o21ai_1 _6456_ (.B1(_2565_),
    .Y(_2566_),
    .A1(net666),
    .A2(_2856_));
 sg13g2_nand2_1 _6457_ (.Y(_2567_),
    .A(_0053_),
    .B(_1068_));
 sg13g2_a22oi_1 _6458_ (.Y(_2568_),
    .B1(_2566_),
    .B2(net662),
    .A2(_2561_),
    .A1(_0052_));
 sg13g2_nand2_1 _6459_ (.Y(_2569_),
    .A(_2567_),
    .B(_2568_));
 sg13g2_nor2_1 _6460_ (.A(_2864_),
    .B(_2562_),
    .Y(_2570_));
 sg13g2_xnor2_1 _6461_ (.Y(_2571_),
    .A(_2569_),
    .B(_2570_));
 sg13g2_xnor2_1 _6462_ (.Y(_2572_),
    .A(_0087_),
    .B(_2571_));
 sg13g2_and2_1 _6463_ (.A(_2564_),
    .B(_2572_),
    .X(_2573_));
 sg13g2_o21ai_1 _6464_ (.B1(net627),
    .Y(_2574_),
    .A1(_2564_),
    .A2(_2572_));
 sg13g2_nor2_1 _6465_ (.A(_2573_),
    .B(net407),
    .Y(_0218_));
 sg13g2_a21oi_1 _6466_ (.A1(\generated._381[0] ),
    .A2(_2571_),
    .Y(_2575_),
    .B1(_2573_));
 sg13g2_a21oi_1 _6467_ (.A1(_2562_),
    .A2(_2569_),
    .Y(_2576_),
    .B1(_2864_));
 sg13g2_mux2_1 _6468_ (.A0(_0048_),
    .A1(_0049_),
    .S(net666),
    .X(_2577_));
 sg13g2_mux2_1 _6469_ (.A0(_2559_),
    .A1(_2577_),
    .S(net662),
    .X(_2578_));
 sg13g2_xnor2_1 _6470_ (.Y(_2579_),
    .A(_2576_),
    .B(_2578_));
 sg13g2_xnor2_1 _6471_ (.Y(_2580_),
    .A(net491),
    .B(_2579_));
 sg13g2_and2_1 _6472_ (.A(_2575_),
    .B(_2580_),
    .X(_2581_));
 sg13g2_nor2_1 _6473_ (.A(_2575_),
    .B(_2580_),
    .Y(_2582_));
 sg13g2_nor3_1 _6474_ (.A(net628),
    .B(net492),
    .C(_2582_),
    .Y(_0219_));
 sg13g2_a21oi_1 _6475_ (.A1(_2841_),
    .A2(_2579_),
    .Y(_2583_),
    .B1(_2582_));
 sg13g2_nand3_1 _6476_ (.B(_2569_),
    .C(_2578_),
    .A(_2562_),
    .Y(_2584_));
 sg13g2_nand2_1 _6477_ (.Y(_2585_),
    .A(net670),
    .B(_2584_));
 sg13g2_nor2_1 _6478_ (.A(net662),
    .B(_2566_),
    .Y(_2586_));
 sg13g2_and2_1 _6479_ (.A(net666),
    .B(_0051_),
    .X(_2587_));
 sg13g2_a21oi_1 _6480_ (.A1(_2840_),
    .A2(_0049_),
    .Y(_2588_),
    .B1(_2587_));
 sg13g2_a21oi_1 _6481_ (.A1(net662),
    .A2(_2588_),
    .Y(_2589_),
    .B1(_2586_));
 sg13g2_xnor2_1 _6482_ (.Y(_2590_),
    .A(_2585_),
    .B(_2589_));
 sg13g2_nor2b_1 _6483_ (.A(_2590_),
    .B_N(\generated._381[2] ),
    .Y(_2591_));
 sg13g2_xnor2_1 _6484_ (.Y(_2592_),
    .A(net520),
    .B(_2590_));
 sg13g2_nor2b_1 _6485_ (.A(_2592_),
    .B_N(_2583_),
    .Y(_2593_));
 sg13g2_nor2b_1 _6486_ (.A(_2583_),
    .B_N(_2592_),
    .Y(_2594_));
 sg13g2_nor3_1 _6487_ (.A(net628),
    .B(_2593_),
    .C(_2594_),
    .Y(_0220_));
 sg13g2_or2_1 _6488_ (.X(_2595_),
    .B(_2594_),
    .A(_2591_));
 sg13g2_nand2b_1 _6489_ (.Y(_2596_),
    .B(_2589_),
    .A_N(_2584_));
 sg13g2_nand2_1 _6490_ (.Y(_2597_),
    .A(net670),
    .B(_2596_));
 sg13g2_nor2_1 _6491_ (.A(net662),
    .B(_2577_),
    .Y(_2598_));
 sg13g2_and2_1 _6492_ (.A(net665),
    .B(_0056_),
    .X(_2599_));
 sg13g2_a21oi_1 _6493_ (.A1(_2840_),
    .A2(_0051_),
    .Y(_2600_),
    .B1(_2599_));
 sg13g2_a21oi_1 _6494_ (.A1(net660),
    .A2(_2600_),
    .Y(_2601_),
    .B1(_2598_));
 sg13g2_xnor2_1 _6495_ (.Y(_2602_),
    .A(_2597_),
    .B(_2601_));
 sg13g2_xnor2_1 _6496_ (.Y(_2603_),
    .A(net455),
    .B(_2602_));
 sg13g2_nor2_1 _6497_ (.A(_2595_),
    .B(_2603_),
    .Y(_2604_));
 sg13g2_and2_1 _6498_ (.A(_2595_),
    .B(_2603_),
    .X(_2605_));
 sg13g2_nor3_1 _6499_ (.A(net628),
    .B(_2604_),
    .C(_2605_),
    .Y(_0221_));
 sg13g2_nor2_1 _6500_ (.A(net522),
    .B(_2602_),
    .Y(_2606_));
 sg13g2_nor2b_1 _6501_ (.A(_2596_),
    .B_N(_2601_),
    .Y(_2607_));
 sg13g2_nor2_1 _6502_ (.A(_2864_),
    .B(_2607_),
    .Y(_2608_));
 sg13g2_mux2_1 _6503_ (.A0(_0056_),
    .A1(_0060_),
    .S(net665),
    .X(_2609_));
 sg13g2_nand2_1 _6504_ (.Y(_2610_),
    .A(net660),
    .B(_2609_));
 sg13g2_o21ai_1 _6505_ (.B1(_2610_),
    .Y(_2611_),
    .A1(net660),
    .A2(_2588_));
 sg13g2_xor2_1 _6506_ (.B(_2611_),
    .A(_2608_),
    .X(_2612_));
 sg13g2_xnor2_1 _6507_ (.Y(_2613_),
    .A(\generated._381[4] ),
    .B(_2612_));
 sg13g2_or3_1 _6508_ (.A(_2605_),
    .B(_2606_),
    .C(_2613_),
    .X(_2614_));
 sg13g2_o21ai_1 _6509_ (.B1(_2613_),
    .Y(_2615_),
    .A1(_2605_),
    .A2(_2606_));
 sg13g2_and3_1 _6510_ (.X(_0222_),
    .A(net626),
    .B(_2614_),
    .C(_2615_));
 sg13g2_o21ai_1 _6511_ (.B1(_2615_),
    .Y(_2616_),
    .A1(_2870_),
    .A2(_2612_));
 sg13g2_inv_1 _6512_ (.Y(_2617_),
    .A(_2616_));
 sg13g2_a21oi_1 _6513_ (.A1(_2607_),
    .A2(_2611_),
    .Y(_2618_),
    .B1(_2864_));
 sg13g2_nor2_1 _6514_ (.A(net665),
    .B(_0060_),
    .Y(_2619_));
 sg13g2_a21oi_1 _6515_ (.A1(net665),
    .A2(_2860_),
    .Y(_2620_),
    .B1(_2619_));
 sg13g2_nand2_1 _6516_ (.Y(_2621_),
    .A(net660),
    .B(_2620_));
 sg13g2_o21ai_1 _6517_ (.B1(_2621_),
    .Y(_2622_),
    .A1(net661),
    .A2(_2600_));
 sg13g2_xor2_1 _6518_ (.B(_2622_),
    .A(_2618_),
    .X(_2623_));
 sg13g2_xor2_1 _6519_ (.B(_2623_),
    .A(net559),
    .X(_2624_));
 sg13g2_nor2_1 _6520_ (.A(_2617_),
    .B(_2624_),
    .Y(_2625_));
 sg13g2_a21oi_1 _6521_ (.A1(_2617_),
    .A2(_2624_),
    .Y(_2626_),
    .B1(net628));
 sg13g2_nor2b_1 _6522_ (.A(_2625_),
    .B_N(_2626_),
    .Y(_0223_));
 sg13g2_nor2_1 _6523_ (.A(net525),
    .B(_2623_),
    .Y(_2627_));
 sg13g2_nor2_1 _6524_ (.A(_2625_),
    .B(_2627_),
    .Y(_2628_));
 sg13g2_nor2b_1 _6525_ (.A(net660),
    .B_N(_2609_),
    .Y(_2629_));
 sg13g2_a21oi_2 _6526_ (.B1(_2629_),
    .Y(_2630_),
    .A2(_0063_),
    .A1(net659));
 sg13g2_nand3_1 _6527_ (.B(_2611_),
    .C(_2622_),
    .A(_2607_),
    .Y(_2631_));
 sg13g2_nand2_1 _6528_ (.Y(_2632_),
    .A(net669),
    .B(_2631_));
 sg13g2_xor2_1 _6529_ (.B(_2632_),
    .A(_2630_),
    .X(_2633_));
 sg13g2_xnor2_1 _6530_ (.Y(_2634_),
    .A(\generated._381[6] ),
    .B(_2633_));
 sg13g2_nor3_1 _6531_ (.A(_2625_),
    .B(_2627_),
    .C(_2634_),
    .Y(_2635_));
 sg13g2_nor2b_1 _6532_ (.A(_2628_),
    .B_N(_2634_),
    .Y(_2636_));
 sg13g2_nor3_1 _6533_ (.A(net628),
    .B(net526),
    .C(_2636_),
    .Y(_0224_));
 sg13g2_nor2_1 _6534_ (.A(net523),
    .B(_2633_),
    .Y(_2637_));
 sg13g2_nor2b_1 _6535_ (.A(net659),
    .B_N(_2620_),
    .Y(_2638_));
 sg13g2_a21oi_1 _6536_ (.A1(net659),
    .A2(_0063_),
    .Y(_2639_),
    .B1(_2638_));
 sg13g2_o21ai_1 _6537_ (.B1(net669),
    .Y(_2640_),
    .A1(_2630_),
    .A2(_2631_));
 sg13g2_xor2_1 _6538_ (.B(_2640_),
    .A(_2639_),
    .X(_2641_));
 sg13g2_xnor2_1 _6539_ (.Y(_2642_),
    .A(\generated._381[7] ),
    .B(_2641_));
 sg13g2_nor3_1 _6540_ (.A(_2636_),
    .B(_2637_),
    .C(_2642_),
    .Y(_2643_));
 sg13g2_o21ai_1 _6541_ (.B1(_2642_),
    .Y(_2644_),
    .A1(_2636_),
    .A2(_2637_));
 sg13g2_nand2_1 _6542_ (.Y(_2645_),
    .A(net626),
    .B(_2644_));
 sg13g2_nor2_1 _6543_ (.A(net524),
    .B(_2645_),
    .Y(_0225_));
 sg13g2_o21ai_1 _6544_ (.B1(_2644_),
    .Y(_2646_),
    .A1(net447),
    .A2(_2641_));
 sg13g2_nor3_1 _6545_ (.A(_2630_),
    .B(_2631_),
    .C(_2639_),
    .Y(_2647_));
 sg13g2_xnor2_1 _6546_ (.Y(_2648_),
    .A(\generated._394[9] ),
    .B(_2647_));
 sg13g2_mux2_1 _6547_ (.A0(_2860_),
    .A1(_2648_),
    .S(net669),
    .X(_2649_));
 sg13g2_xor2_1 _6548_ (.B(_2649_),
    .A(\generated._380 ),
    .X(_2650_));
 sg13g2_o21ai_1 _6549_ (.B1(net626),
    .Y(_2651_),
    .A1(_2646_),
    .A2(_2650_));
 sg13g2_a21oi_1 _6550_ (.A1(_2646_),
    .A2(_2650_),
    .Y(_0226_),
    .B1(_2651_));
 sg13g2_nor2_1 _6551_ (.A(net337),
    .B(_2885_),
    .Y(_2652_));
 sg13g2_and2_1 _6552_ (.A(net337),
    .B(_2885_),
    .X(_2653_));
 sg13g2_nor3_1 _6553_ (.A(net623),
    .B(net338),
    .C(_2653_),
    .Y(_0228_));
 sg13g2_o21ai_1 _6554_ (.B1(_2884_),
    .Y(_2654_),
    .A1(net278),
    .A2(_2653_));
 sg13g2_a21oi_1 _6555_ (.A1(net278),
    .A2(_2653_),
    .Y(_0229_),
    .B1(_2654_));
 sg13g2_nand2b_1 _6556_ (.Y(_2655_),
    .B(_2893_),
    .A_N(_2889_));
 sg13g2_o21ai_1 _6557_ (.B1(_2655_),
    .Y(_0230_),
    .A1(_2830_),
    .A2(_2887_));
 sg13g2_and2_1 _6558_ (.A(\generated._33[1] ),
    .B(net288),
    .X(_2656_));
 sg13g2_and2_1 _6559_ (.A(net282),
    .B(_2656_),
    .X(_2657_));
 sg13g2_and2_1 _6560_ (.A(net274),
    .B(_2657_),
    .X(_2658_));
 sg13g2_nor2_1 _6561_ (.A(\generated._33[5] ),
    .B(\generated._33[4] ),
    .Y(_2659_));
 sg13g2_and3_2 _6562_ (.X(_2660_),
    .A(net269),
    .B(_2658_),
    .C(_2659_));
 sg13g2_nor2_2 _6563_ (.A(net623),
    .B(_2660_),
    .Y(_2661_));
 sg13g2_and2_1 _6564_ (.A(net248),
    .B(_2661_),
    .X(_0232_));
 sg13g2_nor2_1 _6565_ (.A(\generated._33[1] ),
    .B(net288),
    .Y(_2662_));
 sg13g2_nor3_1 _6566_ (.A(net625),
    .B(_2656_),
    .C(net289),
    .Y(_0233_));
 sg13g2_nor2_1 _6567_ (.A(net282),
    .B(_2656_),
    .Y(_2663_));
 sg13g2_nor3_1 _6568_ (.A(net623),
    .B(_2657_),
    .C(net283),
    .Y(_0234_));
 sg13g2_nor2_1 _6569_ (.A(net274),
    .B(_2657_),
    .Y(_2664_));
 sg13g2_nor3_1 _6570_ (.A(net623),
    .B(_2658_),
    .C(net275),
    .Y(_0235_));
 sg13g2_and2_1 _6571_ (.A(net356),
    .B(_2658_),
    .X(_2665_));
 sg13g2_o21ai_1 _6572_ (.B1(_2661_),
    .Y(_2666_),
    .A1(net356),
    .A2(_2658_));
 sg13g2_nor2_1 _6573_ (.A(_2665_),
    .B(_2666_),
    .Y(_0236_));
 sg13g2_nor2_1 _6574_ (.A(net308),
    .B(_2665_),
    .Y(_2667_));
 sg13g2_and2_1 _6575_ (.A(net308),
    .B(_2665_),
    .X(_2668_));
 sg13g2_nor4_1 _6576_ (.A(net623),
    .B(_2660_),
    .C(net309),
    .D(_2668_),
    .Y(_0237_));
 sg13g2_o21ai_1 _6577_ (.B1(_2661_),
    .Y(_2669_),
    .A1(net269),
    .A2(_2668_));
 sg13g2_a21oi_1 _6578_ (.A1(net269),
    .A2(_2668_),
    .Y(_0238_),
    .B1(_2669_));
 sg13g2_nand2_1 _6579_ (.Y(_2670_),
    .A(net439),
    .B(_1042_));
 sg13g2_and3_1 _6580_ (.X(_0239_),
    .A(net745),
    .B(net260),
    .C(_2670_));
 sg13g2_o21ai_1 _6581_ (.B1(net745),
    .Y(_2671_),
    .A1(net324),
    .A2(\generated._487[0] ));
 sg13g2_a21oi_1 _6582_ (.A1(net324),
    .A2(\generated._487[0] ),
    .Y(_0240_),
    .B1(_2671_));
 sg13g2_nand3_1 _6583_ (.B(\generated._487[0] ),
    .C(\generated._487[2] ),
    .A(net324),
    .Y(_2672_));
 sg13g2_a21o_1 _6584_ (.A2(\generated._487[0] ),
    .A1(net324),
    .B1(net439),
    .X(_2673_));
 sg13g2_and4_1 _6585_ (.A(net745),
    .B(_2670_),
    .C(_2672_),
    .D(net440),
    .X(_0241_));
 sg13g2_xnor2_1 _6586_ (.Y(_2674_),
    .A(net395),
    .B(_2672_));
 sg13g2_and3_1 _6587_ (.X(_0242_),
    .A(net745),
    .B(_2670_),
    .C(net396));
 sg13g2_and2_1 _6588_ (.A(net253),
    .B(net626),
    .X(_0243_));
 sg13g2_nor3_1 _6589_ (.A(net630),
    .B(_1047_),
    .C(_2561_),
    .Y(_0244_));
 sg13g2_a21o_1 _6590_ (.A2(_2907_),
    .A1(net313),
    .B1(_2911_),
    .X(_0246_));
 sg13g2_xnor2_1 _6591_ (.Y(_2675_),
    .A(net386),
    .B(_2917_));
 sg13g2_a21oi_1 _6592_ (.A1(_2908_),
    .A2(_2909_),
    .Y(_0250_),
    .B1(_2675_));
 sg13g2_nor2_1 _6593_ (.A(net667),
    .B(_0093_),
    .Y(_2676_));
 sg13g2_a21oi_1 _6594_ (.A1(net668),
    .A2(_2842_),
    .Y(_2677_),
    .B1(_2676_));
 sg13g2_nor2b_1 _6595_ (.A(_2677_),
    .B_N(net662),
    .Y(_2678_));
 sg13g2_a221oi_1 _6596_ (.B2(net672),
    .C1(_2678_),
    .B1(_2561_),
    .A1(\generated._381[0] ),
    .Y(_2679_),
    .A2(_1068_));
 sg13g2_nor2_1 _6597_ (.A(net658),
    .B(_2679_),
    .Y(_2680_));
 sg13g2_xnor2_1 _6598_ (.Y(_2681_),
    .A(_2843_),
    .B(_2679_));
 sg13g2_nor2_1 _6599_ (.A(net631),
    .B(_2681_),
    .Y(_0251_));
 sg13g2_nand2_1 _6600_ (.Y(_2682_),
    .A(net667),
    .B(_0086_));
 sg13g2_o21ai_1 _6601_ (.B1(_2682_),
    .Y(_2683_),
    .A1(net667),
    .A2(_2842_));
 sg13g2_nand2_1 _6602_ (.Y(_2684_),
    .A(_0087_),
    .B(_2561_));
 sg13g2_a22oi_1 _6603_ (.Y(_2685_),
    .B1(_2683_),
    .B2(net664),
    .A2(_1068_),
    .A1(_0093_));
 sg13g2_nand2_1 _6604_ (.Y(_2686_),
    .A(_2684_),
    .B(_2685_));
 sg13g2_nor2_1 _6605_ (.A(_2864_),
    .B(_2679_),
    .Y(_2687_));
 sg13g2_xnor2_1 _6606_ (.Y(_2688_),
    .A(_2686_),
    .B(_2687_));
 sg13g2_nor2_1 _6607_ (.A(net538),
    .B(_2688_),
    .Y(_2689_));
 sg13g2_xnor2_1 _6608_ (.Y(_2690_),
    .A(net538),
    .B(_2688_));
 sg13g2_nor2_1 _6609_ (.A(_2680_),
    .B(_2690_),
    .Y(_2691_));
 sg13g2_a21oi_1 _6610_ (.A1(_2680_),
    .A2(_2690_),
    .Y(_2692_),
    .B1(net628));
 sg13g2_nor2b_1 _6611_ (.A(_2691_),
    .B_N(_2692_),
    .Y(_0252_));
 sg13g2_nor2_1 _6612_ (.A(_2689_),
    .B(_2691_),
    .Y(_2693_));
 sg13g2_a21oi_1 _6613_ (.A1(_2679_),
    .A2(_2686_),
    .Y(_2694_),
    .B1(_2864_));
 sg13g2_mux2_1 _6614_ (.A0(_0086_),
    .A1(_0085_),
    .S(net667),
    .X(_2695_));
 sg13g2_mux2_1 _6615_ (.A0(_2677_),
    .A1(_2695_),
    .S(net662),
    .X(_2696_));
 sg13g2_xor2_1 _6616_ (.B(_2696_),
    .A(_2694_),
    .X(_2697_));
 sg13g2_xnor2_1 _6617_ (.Y(_2698_),
    .A(net556),
    .B(_2697_));
 sg13g2_nor2b_1 _6618_ (.A(_2693_),
    .B_N(_2698_),
    .Y(_2699_));
 sg13g2_nor3_1 _6619_ (.A(_2689_),
    .B(_2691_),
    .C(_2698_),
    .Y(_2700_));
 sg13g2_o21ai_1 _6620_ (.B1(net627),
    .Y(_0253_),
    .A1(_2699_),
    .A2(_2700_));
 sg13g2_a21o_1 _6621_ (.A2(_2697_),
    .A1(net513),
    .B1(_2699_),
    .X(_2701_));
 sg13g2_nand3_1 _6622_ (.B(_2686_),
    .C(_2696_),
    .A(_2679_),
    .Y(_2702_));
 sg13g2_nand2_1 _6623_ (.Y(_2703_),
    .A(net670),
    .B(_2702_));
 sg13g2_nor2_1 _6624_ (.A(net663),
    .B(_2683_),
    .Y(_2704_));
 sg13g2_and2_1 _6625_ (.A(net667),
    .B(_0084_),
    .X(_2705_));
 sg13g2_a21oi_1 _6626_ (.A1(_2840_),
    .A2(_0085_),
    .Y(_2706_),
    .B1(_2705_));
 sg13g2_a21oi_1 _6627_ (.A1(net663),
    .A2(_2706_),
    .Y(_2707_),
    .B1(_2704_));
 sg13g2_xnor2_1 _6628_ (.Y(_2708_),
    .A(_2703_),
    .B(_2707_));
 sg13g2_xnor2_1 _6629_ (.Y(_2709_),
    .A(_2856_),
    .B(_2708_));
 sg13g2_nor2b_1 _6630_ (.A(_2709_),
    .B_N(_2701_),
    .Y(_2710_));
 sg13g2_nor2b_1 _6631_ (.A(_2701_),
    .B_N(_2709_),
    .Y(_2711_));
 sg13g2_o21ai_1 _6632_ (.B1(net627),
    .Y(_0254_),
    .A1(_2710_),
    .A2(_2711_));
 sg13g2_a21oi_1 _6633_ (.A1(_2856_),
    .A2(_2708_),
    .Y(_2712_),
    .B1(_2710_));
 sg13g2_nand2b_1 _6634_ (.Y(_2713_),
    .B(_2707_),
    .A_N(_2702_));
 sg13g2_nand2_1 _6635_ (.Y(_2714_),
    .A(net670),
    .B(_2713_));
 sg13g2_nor2_1 _6636_ (.A(net663),
    .B(_2695_),
    .Y(_2715_));
 sg13g2_and2_1 _6637_ (.A(net665),
    .B(_0083_),
    .X(_2716_));
 sg13g2_a21oi_1 _6638_ (.A1(_2840_),
    .A2(_0084_),
    .Y(_2717_),
    .B1(_2716_));
 sg13g2_a21oi_2 _6639_ (.B1(_2715_),
    .Y(_2718_),
    .A2(_2717_),
    .A1(net660));
 sg13g2_inv_1 _6640_ (.Y(_2719_),
    .A(_2718_));
 sg13g2_xnor2_1 _6641_ (.Y(_2720_),
    .A(_2714_),
    .B(_2718_));
 sg13g2_xnor2_1 _6642_ (.Y(_2721_),
    .A(net536),
    .B(_2720_));
 sg13g2_nor2b_1 _6643_ (.A(_2712_),
    .B_N(_2721_),
    .Y(_2722_));
 sg13g2_nor2b_1 _6644_ (.A(_2721_),
    .B_N(_2712_),
    .Y(_2723_));
 sg13g2_o21ai_1 _6645_ (.B1(net626),
    .Y(_0255_),
    .A1(_2722_),
    .A2(_2723_));
 sg13g2_a21o_1 _6646_ (.A2(_2720_),
    .A1(net501),
    .B1(_2722_),
    .X(_2724_));
 sg13g2_o21ai_1 _6647_ (.B1(net670),
    .Y(_2725_),
    .A1(_2713_),
    .A2(_2719_));
 sg13g2_mux2_1 _6648_ (.A0(_0083_),
    .A1(_0082_),
    .S(net665),
    .X(_2726_));
 sg13g2_nand2_1 _6649_ (.Y(_2727_),
    .A(net661),
    .B(_2726_));
 sg13g2_o21ai_1 _6650_ (.B1(_2727_),
    .Y(_2728_),
    .A1(net660),
    .A2(_2706_));
 sg13g2_xor2_1 _6651_ (.B(_2728_),
    .A(_2725_),
    .X(_2729_));
 sg13g2_nor2_1 _6652_ (.A(_0049_),
    .B(_2729_),
    .Y(_2730_));
 sg13g2_xnor2_1 _6653_ (.Y(_2731_),
    .A(_0049_),
    .B(_2729_));
 sg13g2_nor2b_1 _6654_ (.A(_2724_),
    .B_N(_2731_),
    .Y(_2732_));
 sg13g2_nor2b_1 _6655_ (.A(_2731_),
    .B_N(_2724_),
    .Y(_2733_));
 sg13g2_nor3_1 _6656_ (.A(net628),
    .B(_2732_),
    .C(_2733_),
    .Y(_0256_));
 sg13g2_nor2_1 _6657_ (.A(_2730_),
    .B(_2733_),
    .Y(_2734_));
 sg13g2_nand3b_1 _6658_ (.B(_2718_),
    .C(_2728_),
    .Y(_2735_),
    .A_N(_2713_));
 sg13g2_nand2_1 _6659_ (.Y(_2736_),
    .A(net669),
    .B(_2735_));
 sg13g2_mux2_1 _6660_ (.A0(_0082_),
    .A1(_0081_),
    .S(net665),
    .X(_2737_));
 sg13g2_nand2_1 _6661_ (.Y(_2738_),
    .A(net659),
    .B(_2737_));
 sg13g2_o21ai_1 _6662_ (.B1(_2738_),
    .Y(_2739_),
    .A1(net661),
    .A2(_2717_));
 sg13g2_xnor2_1 _6663_ (.Y(_2740_),
    .A(_2736_),
    .B(_2739_));
 sg13g2_xor2_1 _6664_ (.B(_2740_),
    .A(net545),
    .X(_2741_));
 sg13g2_o21ai_1 _6665_ (.B1(net626),
    .Y(_2742_),
    .A1(_2734_),
    .A2(_2741_));
 sg13g2_a21oi_1 _6666_ (.A1(_2734_),
    .A2(_2741_),
    .Y(_0257_),
    .B1(_2742_));
 sg13g2_nand2_1 _6667_ (.Y(_2743_),
    .A(\generated._394[6] ),
    .B(_2740_));
 sg13g2_o21ai_1 _6668_ (.B1(_2743_),
    .Y(_2744_),
    .A1(_2734_),
    .A2(_2741_));
 sg13g2_nor2b_1 _6669_ (.A(net659),
    .B_N(_2726_),
    .Y(_2745_));
 sg13g2_a21oi_2 _6670_ (.B1(_2745_),
    .Y(_2746_),
    .A2(_0081_),
    .A1(net659));
 sg13g2_nand2b_1 _6671_ (.Y(_2747_),
    .B(_2739_),
    .A_N(_2735_));
 sg13g2_nand2_1 _6672_ (.Y(_2748_),
    .A(net669),
    .B(_2747_));
 sg13g2_xor2_1 _6673_ (.B(_2748_),
    .A(_2746_),
    .X(_2749_));
 sg13g2_xnor2_1 _6674_ (.Y(_2750_),
    .A(_0056_),
    .B(_2749_));
 sg13g2_xnor2_1 _6675_ (.Y(_2751_),
    .A(_2744_),
    .B(_2750_));
 sg13g2_nand2_1 _6676_ (.Y(_0258_),
    .A(net626),
    .B(_2751_));
 sg13g2_a22oi_1 _6677_ (.Y(_2752_),
    .B1(_2750_),
    .B2(_2744_),
    .A2(_2749_),
    .A1(net485));
 sg13g2_nor2b_1 _6678_ (.A(net659),
    .B_N(_2737_),
    .Y(_2753_));
 sg13g2_a21oi_1 _6679_ (.A1(net659),
    .A2(_0081_),
    .Y(_2754_),
    .B1(_2753_));
 sg13g2_o21ai_1 _6680_ (.B1(net669),
    .Y(_2755_),
    .A1(_2746_),
    .A2(_2747_));
 sg13g2_xor2_1 _6681_ (.B(_2755_),
    .A(_2754_),
    .X(_2756_));
 sg13g2_xnor2_1 _6682_ (.Y(_2757_),
    .A(_0060_),
    .B(_2756_));
 sg13g2_nand2b_1 _6683_ (.Y(_2758_),
    .B(_2752_),
    .A_N(_2757_));
 sg13g2_nand2b_1 _6684_ (.Y(_2759_),
    .B(_2757_),
    .A_N(_2752_));
 sg13g2_and3_1 _6685_ (.X(_0259_),
    .A(net626),
    .B(_2758_),
    .C(_2759_));
 sg13g2_nand2_1 _6686_ (.Y(_2760_),
    .A(net495),
    .B(_2756_));
 sg13g2_nor3_1 _6687_ (.A(_2746_),
    .B(_2747_),
    .C(_2754_),
    .Y(_2761_));
 sg13g2_xnor2_1 _6688_ (.Y(_2762_),
    .A(\generated._380 ),
    .B(_2761_));
 sg13g2_nor2_1 _6689_ (.A(net669),
    .B(_0081_),
    .Y(_2763_));
 sg13g2_a21oi_1 _6690_ (.A1(net669),
    .A2(_2762_),
    .Y(_2764_),
    .B1(_2763_));
 sg13g2_xnor2_1 _6691_ (.Y(_2765_),
    .A(_2860_),
    .B(_2764_));
 sg13g2_and3_1 _6692_ (.X(_2766_),
    .A(_2759_),
    .B(_2760_),
    .C(_2765_));
 sg13g2_a21oi_1 _6693_ (.A1(_2759_),
    .A2(_2760_),
    .Y(_2767_),
    .B1(_2765_));
 sg13g2_nor3_1 _6694_ (.A(net628),
    .B(_2766_),
    .C(_2767_),
    .Y(_0260_));
 sg13g2_nor2_1 _6695_ (.A(\generated._28[2] ),
    .B(\generated._28[1] ),
    .Y(_2768_));
 sg13g2_nand2_1 _6696_ (.Y(_2769_),
    .A(\generated._28[3] ),
    .B(_2768_));
 sg13g2_o21ai_1 _6697_ (.B1(_2660_),
    .Y(_2770_),
    .A1(\generated._28[0] ),
    .A2(_2769_));
 sg13g2_a21oi_1 _6698_ (.A1(_2660_),
    .A2(_2769_),
    .Y(_2771_),
    .B1(net322));
 sg13g2_and2_1 _6699_ (.A(net322),
    .B(_2660_),
    .X(_2772_));
 sg13g2_nor3_1 _6700_ (.A(net624),
    .B(net323),
    .C(_2772_),
    .Y(_0261_));
 sg13g2_and2_1 _6701_ (.A(net373),
    .B(_2772_),
    .X(_2773_));
 sg13g2_o21ai_1 _6702_ (.B1(_2884_),
    .Y(_2774_),
    .A1(net373),
    .A2(_2772_));
 sg13g2_nor2_1 _6703_ (.A(_2773_),
    .B(_2774_),
    .Y(_0262_));
 sg13g2_nand3_1 _6704_ (.B(\generated._28[1] ),
    .C(\generated._28[0] ),
    .A(\generated._28[2] ),
    .Y(_2775_));
 sg13g2_a21oi_1 _6705_ (.A1(net367),
    .A2(_2773_),
    .Y(_2776_),
    .B1(net624));
 sg13g2_o21ai_1 _6706_ (.B1(_2776_),
    .Y(_2777_),
    .A1(net367),
    .A2(_2773_));
 sg13g2_inv_1 _6707_ (.Y(_0263_),
    .A(net368));
 sg13g2_xor2_1 _6708_ (.B(_2775_),
    .A(\generated._28[3] ),
    .X(_2778_));
 sg13g2_nor3_1 _6709_ (.A(net624),
    .B(_2770_),
    .C(_2778_),
    .Y(_2779_));
 sg13g2_a21o_1 _6710_ (.A2(_2661_),
    .A1(net377),
    .B1(_2779_),
    .X(_0264_));
 sg13g2_and2_1 _6711_ (.A(net264),
    .B(_2907_),
    .X(_0265_));
 sg13g2_nor2_1 _6712_ (.A(\generated._357[1] ),
    .B(net271),
    .Y(_2780_));
 sg13g2_nor3_1 _6713_ (.A(net625),
    .B(_2894_),
    .C(net272),
    .Y(_0266_));
 sg13g2_nor2_1 _6714_ (.A(net327),
    .B(_2894_),
    .Y(_2781_));
 sg13g2_and2_1 _6715_ (.A(net327),
    .B(_2894_),
    .X(_2782_));
 sg13g2_nor3_1 _6716_ (.A(_2908_),
    .B(net328),
    .C(_2782_),
    .Y(_0267_));
 sg13g2_nand2_1 _6717_ (.Y(_2783_),
    .A(net358),
    .B(_2782_));
 sg13g2_o21ai_1 _6718_ (.B1(_2907_),
    .Y(_2784_),
    .A1(net358),
    .A2(_2782_));
 sg13g2_nor2b_1 _6719_ (.A(_2784_),
    .B_N(_2783_),
    .Y(_0268_));
 sg13g2_xor2_1 _6720_ (.B(_2783_),
    .A(net320),
    .X(_2785_));
 sg13g2_nor2_1 _6721_ (.A(_2908_),
    .B(net321),
    .Y(_0269_));
 sg13g2_and2_1 _6722_ (.A(net247),
    .B(_2886_),
    .X(_0270_));
 sg13g2_xnor2_1 _6723_ (.Y(_2786_),
    .A(\generated._21[1] ),
    .B(net344));
 sg13g2_nor2_1 _6724_ (.A(_2887_),
    .B(net345),
    .Y(_0271_));
 sg13g2_and3_1 _6725_ (.X(_2787_),
    .A(\generated._21[1] ),
    .B(net344),
    .C(net291));
 sg13g2_a21oi_1 _6726_ (.A1(\generated._21[1] ),
    .A2(\generated._21[0] ),
    .Y(_2788_),
    .B1(net291));
 sg13g2_nor3_1 _6727_ (.A(_2887_),
    .B(_2787_),
    .C(net292),
    .Y(_0272_));
 sg13g2_nand2_1 _6728_ (.Y(_2789_),
    .A(net346),
    .B(_2787_));
 sg13g2_o21ai_1 _6729_ (.B1(_2886_),
    .Y(_2790_),
    .A1(net346),
    .A2(_2787_));
 sg13g2_nor2b_1 _6730_ (.A(net347),
    .B_N(_2789_),
    .Y(_0273_));
 sg13g2_xor2_1 _6731_ (.B(_2789_),
    .A(net349),
    .X(_2791_));
 sg13g2_nor2_1 _6732_ (.A(_2887_),
    .B(_2791_),
    .Y(_0274_));
 sg13g2_nand2b_1 _6733_ (.Y(_2792_),
    .B(_1182_),
    .A_N(\generated._1087[0] ));
 sg13g2_nand2_1 _6734_ (.Y(_2793_),
    .A(net687),
    .B(\generated._165[4] ));
 sg13g2_a21oi_1 _6735_ (.A1(_1187_),
    .A2(_2793_),
    .Y(_2794_),
    .B1(_2792_));
 sg13g2_and3_1 _6736_ (.X(_2795_),
    .A(_1187_),
    .B(_2792_),
    .C(_2793_));
 sg13g2_nor3_1 _6737_ (.A(net744),
    .B(_2794_),
    .C(_2795_),
    .Y(_2796_));
 sg13g2_nor2_1 _6738_ (.A(\generated._28[3] ),
    .B(\generated._28[2] ),
    .Y(_2797_));
 sg13g2_o21ai_1 _6739_ (.B1(_1154_),
    .Y(_2798_),
    .A1(_1158_),
    .A2(_2797_));
 sg13g2_nor2_1 _6740_ (.A(_0011_),
    .B(_1161_),
    .Y(_2799_));
 sg13g2_o21ai_1 _6741_ (.B1(_1156_),
    .Y(_2800_),
    .A1(_2798_),
    .A2(_2799_));
 sg13g2_a21oi_1 _6742_ (.A1(net744),
    .A2(_2800_),
    .Y(_2801_),
    .B1(_2796_));
 sg13g2_nor2_1 _6743_ (.A(_0010_),
    .B(_1161_),
    .Y(_2802_));
 sg13g2_o21ai_1 _6744_ (.B1(_1157_),
    .Y(_2803_),
    .A1(_2798_),
    .A2(_2802_));
 sg13g2_a22oi_1 _6745_ (.Y(_2804_),
    .B1(_1184_),
    .B2(_2792_),
    .A2(_1170_),
    .A1(_2868_));
 sg13g2_o21ai_1 _6746_ (.B1(_2803_),
    .Y(_2805_),
    .A1(net744),
    .A2(_2804_));
 sg13g2_xnor2_1 _6747_ (.Y(_2806_),
    .A(\generated._65[4] ),
    .B(\generated._65[2] ));
 sg13g2_o21ai_1 _6748_ (.B1(_2793_),
    .Y(_2807_),
    .A1(_1184_),
    .A2(_1186_));
 sg13g2_xnor2_1 _6749_ (.Y(_2808_),
    .A(_2806_),
    .B(_2807_));
 sg13g2_a21oi_1 _6750_ (.A1(_1184_),
    .A2(_2795_),
    .Y(_2809_),
    .B1(_2808_));
 sg13g2_and3_1 _6751_ (.X(_2810_),
    .A(_1184_),
    .B(_2795_),
    .C(_2808_));
 sg13g2_nor3_1 _6752_ (.A(net744),
    .B(_2809_),
    .C(_2810_),
    .Y(_2811_));
 sg13g2_nor2_1 _6753_ (.A(_0012_),
    .B(_1161_),
    .Y(_2812_));
 sg13g2_o21ai_1 _6754_ (.B1(_1156_),
    .Y(_2813_),
    .A1(_2798_),
    .A2(_2812_));
 sg13g2_a21oi_1 _6755_ (.A1(net744),
    .A2(_2813_),
    .Y(_2814_),
    .B1(_2811_));
 sg13g2_mux2_1 _6756_ (.A0(_2814_),
    .A1(_2805_),
    .S(_2801_),
    .X(_2815_));
 sg13g2_nor2_1 _6757_ (.A(_1147_),
    .B(_2815_),
    .Y(_0275_));
 sg13g2_a21oi_1 _6758_ (.A1(_2801_),
    .A2(_2814_),
    .Y(_0276_),
    .B1(_1147_));
 sg13g2_nor3_1 _6759_ (.A(\generated._28[3] ),
    .B(\generated._28[0] ),
    .C(_1158_),
    .Y(_2816_));
 sg13g2_nor3_2 _6760_ (.A(_1151_),
    .B(_1153_),
    .C(_2816_),
    .Y(_2817_));
 sg13g2_o21ai_1 _6761_ (.B1(_1158_),
    .Y(_2818_),
    .A1(\generated._346[5] ),
    .A2(_0014_));
 sg13g2_nand2_1 _6762_ (.Y(_2819_),
    .A(_2817_),
    .B(_2818_));
 sg13g2_nor2_1 _6763_ (.A(_1154_),
    .B(_1155_),
    .Y(_2820_));
 sg13g2_nor2_1 _6764_ (.A(_2869_),
    .B(_2820_),
    .Y(_2821_));
 sg13g2_a21oi_1 _6765_ (.A1(_2819_),
    .A2(_2821_),
    .Y(_2822_),
    .B1(_2796_));
 sg13g2_o21ai_1 _6766_ (.B1(_1158_),
    .Y(_2823_),
    .A1(\generated._346[5] ),
    .A2(_0015_));
 sg13g2_nand2_1 _6767_ (.Y(_2824_),
    .A(_2817_),
    .B(_2823_));
 sg13g2_a21oi_1 _6768_ (.A1(_2821_),
    .A2(_2824_),
    .Y(_2825_),
    .B1(_2811_));
 sg13g2_o21ai_1 _6769_ (.B1(_1158_),
    .Y(_2826_),
    .A1(\generated._346[5] ),
    .A2(_0013_));
 sg13g2_nand2_1 _6770_ (.Y(_2827_),
    .A(_2817_),
    .B(_2826_));
 sg13g2_a22oi_1 _6771_ (.Y(_2828_),
    .B1(_2821_),
    .B2(_2827_),
    .A2(_2804_),
    .A1(_2869_));
 sg13g2_mux2_1 _6772_ (.A0(_2825_),
    .A1(_2828_),
    .S(_2822_),
    .X(_2829_));
 sg13g2_nor2_1 _6773_ (.A(_1147_),
    .B(_2829_),
    .Y(_0277_));
 sg13g2_a21oi_1 _6774_ (.A1(_2822_),
    .A2(_2825_),
    .Y(_0278_),
    .B1(_1147_));
 sg13g2_nor2b_1 _6775_ (.A(_2459_),
    .B_N(_2461_),
    .Y(_0204_));
 sg13g2_dfrbp_1 _6776_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net244),
    .D(\generated._889[3] ),
    .Q_N(_0090_),
    .Q(\generated._66[3] ));
 sg13g2_dfrbp_1 _6777_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net245),
    .D(\generated._889[4] ),
    .Q_N(_0019_),
    .Q(\generated._66[4] ));
 sg13g2_dfrbp_1 _6778_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net16),
    .D(\generated._889[5] ),
    .Q_N(_0020_),
    .Q(\generated._66[5] ));
 sg13g2_dfrbp_1 _6779_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net17),
    .D(\generated._889[6] ),
    .Q_N(_0021_),
    .Q(\generated._66[6] ));
 sg13g2_dfrbp_1 _6780_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net18),
    .D(\generated._889[7] ),
    .Q_N(_0028_),
    .Q(\generated._66[7] ));
 sg13g2_dfrbp_1 _6781_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net19),
    .D(\generated._889[8] ),
    .Q_N(_0030_),
    .Q(\generated._66[8] ));
 sg13g2_dfrbp_1 _6782_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net20),
    .D(\generated._889[9] ),
    .Q_N(_0032_),
    .Q(\generated._66[9] ));
 sg13g2_dfrbp_1 _6783_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net21),
    .D(\generated._938[3] ),
    .Q_N(_0018_),
    .Q(\generated._69[3] ));
 sg13g2_dfrbp_1 _6784_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net22),
    .D(\generated._938[4] ),
    .Q_N(_0027_),
    .Q(\generated._69[4] ));
 sg13g2_dfrbp_1 _6785_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net23),
    .D(\generated._938[5] ),
    .Q_N(_0029_),
    .Q(\generated._69[5] ));
 sg13g2_dfrbp_1 _6786_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net24),
    .D(\generated._938[6] ),
    .Q_N(_0031_),
    .Q(\generated._69[6] ));
 sg13g2_dfrbp_1 _6787_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net25),
    .D(net535),
    .Q_N(_0033_),
    .Q(\generated._69[7] ));
 sg13g2_dfrbp_1 _6788_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net29),
    .D(net426),
    .Q_N(_0034_),
    .Q(\generated._69[8] ));
 sg13g2_dfrbp_1 _6789_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net243),
    .D(net484),
    .Q_N(_0023_),
    .Q(\generated._69[9] ));
 sg13g2_dfrbp_1 _6790_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net222),
    .D(_0116_),
    .Q_N(_3335_),
    .Q(_0013_));
 sg13g2_dfrbp_1 _6791_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net221),
    .D(_0117_),
    .Q_N(_3334_),
    .Q(_0014_));
 sg13g2_dfrbp_1 _6792_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net30),
    .D(_0118_),
    .Q_N(_3336_),
    .Q(_0015_));
 sg13g2_dfrbp_1 _6793_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net31),
    .D(_0004_),
    .Q_N(_3337_),
    .Q(_0010_));
 sg13g2_dfrbp_1 _6794_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net32),
    .D(_0005_),
    .Q_N(_3338_),
    .Q(_0011_));
 sg13g2_dfrbp_1 _6795_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net33),
    .D(_0006_),
    .Q_N(_3339_),
    .Q(_0012_));
 sg13g2_dfrbp_1 _6796_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net34),
    .D(_0000_),
    .Q_N(_3340_),
    .Q(_0007_));
 sg13g2_dfrbp_1 _6797_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net36),
    .D(_0001_),
    .Q_N(_3341_),
    .Q(_0008_));
 sg13g2_dfrbp_1 _6798_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net220),
    .D(_0002_),
    .Q_N(_3333_),
    .Q(_0009_));
 sg13g2_dfrbp_1 _6799_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net107),
    .D(_0119_),
    .Q_N(_3342_),
    .Q(audio));
 sg13g2_dfrbp_1 _6800_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net219),
    .D(_0003_),
    .Q_N(_3332_),
    .Q(\generated._1148[0] ));
 sg13g2_dfrbp_1 _6801_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net218),
    .D(_0120_),
    .Q_N(_3331_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _6802_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net217),
    .D(_0121_),
    .Q_N(_3330_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _6803_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net216),
    .D(_0122_),
    .Q_N(_3329_),
    .Q(\generated._614[0] ));
 sg13g2_dfrbp_1 _6804_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net214),
    .D(net380),
    .Q_N(_3328_),
    .Q(\generated._614[1] ));
 sg13g2_dfrbp_1 _6805_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net212),
    .D(net352),
    .Q_N(_3327_),
    .Q(\generated._614[2] ));
 sg13g2_dfrbp_1 _6806_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net210),
    .D(net414),
    .Q_N(_3326_),
    .Q(\generated._614[3] ));
 sg13g2_dfrbp_1 _6807_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net208),
    .D(net268),
    .Q_N(_3325_),
    .Q(\generated._614[4] ));
 sg13g2_dfrbp_1 _6808_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net206),
    .D(_0127_),
    .Q_N(_3324_),
    .Q(\generated._614[5] ));
 sg13g2_dfrbp_1 _6809_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net204),
    .D(_0128_),
    .Q_N(_0099_),
    .Q(\generated._221[0] ));
 sg13g2_dfrbp_1 _6810_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net202),
    .D(_0129_),
    .Q_N(_3323_),
    .Q(\generated._221[1] ));
 sg13g2_dfrbp_1 _6811_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net200),
    .D(_0130_),
    .Q_N(_0100_),
    .Q(\generated._221[2] ));
 sg13g2_dfrbp_1 _6812_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net198),
    .D(_0131_),
    .Q_N(_0101_),
    .Q(\generated._221[3] ));
 sg13g2_dfrbp_1 _6813_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net196),
    .D(_0132_),
    .Q_N(_3322_),
    .Q(\generated._1024[0] ));
 sg13g2_dfrbp_1 _6814_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net195),
    .D(_0133_),
    .Q_N(_0106_),
    .Q(\generated._1024[1] ));
 sg13g2_dfrbp_1 _6815_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net194),
    .D(_0134_),
    .Q_N(_0091_),
    .Q(\generated._1024[2] ));
 sg13g2_dfrbp_1 _6816_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net193),
    .D(_0135_),
    .Q_N(_0035_),
    .Q(\generated._434[10] ));
 sg13g2_dfrbp_1 _6817_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net192),
    .D(_0136_),
    .Q_N(_0043_),
    .Q(\generated._434[11] ));
 sg13g2_dfrbp_1 _6818_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net191),
    .D(net500),
    .Q_N(_0042_),
    .Q(\generated._434[12] ));
 sg13g2_dfrbp_1 _6819_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net190),
    .D(net488),
    .Q_N(_0045_),
    .Q(\generated._434[13] ));
 sg13g2_dfrbp_1 _6820_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net189),
    .D(_0139_),
    .Q_N(_0041_),
    .Q(\generated._434[14] ));
 sg13g2_dfrbp_1 _6821_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net188),
    .D(_0140_),
    .Q_N(_0040_),
    .Q(\generated._434[15] ));
 sg13g2_dfrbp_1 _6822_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net187),
    .D(_0141_),
    .Q_N(_0039_),
    .Q(\generated._434[16] ));
 sg13g2_dfrbp_1 _6823_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net186),
    .D(_0142_),
    .Q_N(_0047_),
    .Q(\generated._434[17] ));
 sg13g2_dfrbp_1 _6824_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net185),
    .D(net482),
    .Q_N(_0038_),
    .Q(\generated._434[18] ));
 sg13g2_dfrbp_1 _6825_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net184),
    .D(net332),
    .Q_N(_0037_),
    .Q(\generated._434[19] ));
 sg13g2_dfrbp_1 _6826_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net183),
    .D(net255),
    .Q_N(\generated._1118[0] ),
    .Q(\generated._100[0] ));
 sg13g2_dfrbp_1 _6827_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net182),
    .D(_0146_),
    .Q_N(_3321_),
    .Q(\generated._100[1] ));
 sg13g2_dfrbp_1 _6828_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net181),
    .D(net287),
    .Q_N(_3320_),
    .Q(\generated._100[2] ));
 sg13g2_dfrbp_1 _6829_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net163),
    .D(_0148_),
    .Q_N(_3319_),
    .Q(\generated._100[3] ));
 sg13g2_dfrbp_1 _6830_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net162),
    .D(_0149_),
    .Q_N(_3318_),
    .Q(\generated._100[4] ));
 sg13g2_dfrbp_1 _6831_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net161),
    .D(net389),
    .Q_N(_0026_),
    .Q(\generated._100[5] ));
 sg13g2_dfrbp_1 _6832_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net160),
    .D(_0151_),
    .Q_N(_3317_),
    .Q(\generated._100[6] ));
 sg13g2_dfrbp_1 _6833_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net159),
    .D(_0152_),
    .Q_N(_3316_),
    .Q(\generated._100[7] ));
 sg13g2_dfrbp_1 _6834_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net158),
    .D(_0153_),
    .Q_N(_3315_),
    .Q(\generated._100[8] ));
 sg13g2_dfrbp_1 _6835_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net157),
    .D(_0154_),
    .Q_N(_3314_),
    .Q(\generated._100[9] ));
 sg13g2_dfrbp_1 _6836_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net156),
    .D(_0155_),
    .Q_N(_0075_),
    .Q(\generated._1084[0] ));
 sg13g2_dfrbp_1 _6837_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net155),
    .D(_0156_),
    .Q_N(_3313_),
    .Q(\generated._1084[1] ));
 sg13g2_dfrbp_1 _6838_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net154),
    .D(_0157_),
    .Q_N(_3312_),
    .Q(\generated._1084[2] ));
 sg13g2_dfrbp_1 _6839_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net153),
    .D(net423),
    .Q_N(_3311_),
    .Q(\generated._1084[3] ));
 sg13g2_dfrbp_1 _6840_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net152),
    .D(_0159_),
    .Q_N(_3310_),
    .Q(\generated._1084[4] ));
 sg13g2_dfrbp_1 _6841_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net141),
    .D(_0160_),
    .Q_N(_3309_),
    .Q(\generated._1084[5] ));
 sg13g2_dfrbp_1 _6842_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net140),
    .D(_0161_),
    .Q_N(_3308_),
    .Q(\generated._1084[6] ));
 sg13g2_dfrbp_1 _6843_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net139),
    .D(net528),
    .Q_N(_3307_),
    .Q(\generated._1084[7] ));
 sg13g2_dfrbp_1 _6844_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net138),
    .D(_0163_),
    .Q_N(_3306_),
    .Q(\generated._1084[8] ));
 sg13g2_dfrbp_1 _6845_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net137),
    .D(_0164_),
    .Q_N(_3305_),
    .Q(\generated._1084[9] ));
 sg13g2_dfrbp_1 _6846_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net136),
    .D(net263),
    .Q_N(\generated._1076[0] ),
    .Q(\generated._1078[0] ));
 sg13g2_dfrbp_1 _6847_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net135),
    .D(net334),
    .Q_N(_3304_),
    .Q(\generated._1078[1] ));
 sg13g2_dfrbp_1 _6848_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net134),
    .D(net458),
    .Q_N(_3303_),
    .Q(\generated._1078[2] ));
 sg13g2_dfrbp_1 _6849_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net133),
    .D(net393),
    .Q_N(_3302_),
    .Q(\generated._1078[3] ));
 sg13g2_dfrbp_1 _6850_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net132),
    .D(_0169_),
    .Q_N(_3301_),
    .Q(\generated._1074[0] ));
 sg13g2_dfrbp_1 _6851_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(net477),
    .Q_N(_0109_),
    .Q(\generated._1074[1] ));
 sg13g2_dfrbp_1 _6852_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net130),
    .D(_0171_),
    .Q_N(_0108_),
    .Q(\generated._1074[2] ));
 sg13g2_dfrbp_1 _6853_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net129),
    .D(_0172_),
    .Q_N(\generated._1025[0] ),
    .Q(\generated._970 ));
 sg13g2_dfrbp_1 _6854_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net128),
    .D(_0173_),
    .Q_N(_3300_),
    .Q(\generated._969 ));
 sg13g2_dfrbp_1 _6855_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net127),
    .D(net266),
    .Q_N(\generated._77[0] ),
    .Q(\generated._1000[0] ));
 sg13g2_dfrbp_1 _6856_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net125),
    .D(net305),
    .Q_N(_3299_),
    .Q(\generated._406[1] ));
 sg13g2_dfrbp_1 _6857_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net123),
    .D(_0176_),
    .Q_N(_3298_),
    .Q(\generated._406[2] ));
 sg13g2_dfrbp_1 _6858_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net121),
    .D(_0177_),
    .Q_N(_3297_),
    .Q(\generated._406[3] ));
 sg13g2_dfrbp_1 _6859_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net119),
    .D(_0178_),
    .Q_N(_3296_),
    .Q(\generated._406[4] ));
 sg13g2_dfrbp_1 _6860_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net117),
    .D(net312),
    .Q_N(_3295_),
    .Q(\generated._406[5] ));
 sg13g2_dfrbp_1 _6861_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net105),
    .D(net330),
    .Q_N(_3294_),
    .Q(\generated._406[6] ));
 sg13g2_dfrbp_1 _6862_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net103),
    .D(net319),
    .Q_N(_3293_),
    .Q(\generated._406[7] ));
 sg13g2_dfrbp_1 _6863_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net101),
    .D(net257),
    .Q_N(\generated._941[0] ),
    .Q(\generated._71[0] ));
 sg13g2_dfrbp_1 _6864_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net100),
    .D(net307),
    .Q_N(_3292_),
    .Q(\generated._71[1] ));
 sg13g2_dfrbp_1 _6865_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net99),
    .D(net454),
    .Q_N(_3291_),
    .Q(\generated._71[2] ));
 sg13g2_dfrbp_1 _6866_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net98),
    .D(net402),
    .Q_N(_3290_),
    .Q(\generated._71[3] ));
 sg13g2_dfrbp_1 _6867_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net97),
    .D(net259),
    .Q_N(\generated._698[0] ),
    .Q(\generated._63[0] ));
 sg13g2_dfrbp_1 _6868_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net96),
    .D(net301),
    .Q_N(_3289_),
    .Q(\generated._63[1] ));
 sg13g2_dfrbp_1 _6869_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net95),
    .D(_0188_),
    .Q_N(_3288_),
    .Q(\generated._63[2] ));
 sg13g2_dfrbp_1 _6870_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net108),
    .D(net405),
    .Q_N(_3343_),
    .Q(\generated._63[3] ));
 sg13g2_dfrbp_1 _6871_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net109),
    .D(\generated._561[0] ),
    .Q_N(_0079_),
    .Q(\generated._562[0] ));
 sg13g2_dfrbp_1 _6872_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net110),
    .D(\generated._561[1] ),
    .Q_N(_0057_),
    .Q(\generated._562[1] ));
 sg13g2_dfrbp_1 _6873_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net111),
    .D(\generated._561[2] ),
    .Q_N(_0061_),
    .Q(\generated._562[2] ));
 sg13g2_dfrbp_1 _6874_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net112),
    .D(\generated._561[3] ),
    .Q_N(_0064_),
    .Q(\generated._562[3] ));
 sg13g2_dfrbp_1 _6875_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net113),
    .D(\generated._561[4] ),
    .Q_N(_0066_),
    .Q(\generated._562[4] ));
 sg13g2_dfrbp_1 _6876_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net114),
    .D(\generated._561[5] ),
    .Q_N(_0068_),
    .Q(\generated._562[5] ));
 sg13g2_dfrbp_1 _6877_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net115),
    .D(\generated._561[6] ),
    .Q_N(_0070_),
    .Q(\generated._562[6] ));
 sg13g2_dfrbp_1 _6878_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net116),
    .D(\generated._561[7] ),
    .Q_N(_0072_),
    .Q(\generated._562[7] ));
 sg13g2_dfrbp_1 _6879_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net142),
    .D(\generated._561[8] ),
    .Q_N(_0073_),
    .Q(\generated._562[8] ));
 sg13g2_dfrbp_1 _6880_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net94),
    .D(\generated._561[9] ),
    .Q_N(_0074_),
    .Q(\generated._562[9] ));
 sg13g2_dfrbp_1 _6881_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net93),
    .D(net365),
    .Q_N(_3287_),
    .Q(\generated._69[0] ));
 sg13g2_dfrbp_1 _6882_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net92),
    .D(net508),
    .Q_N(_0025_),
    .Q(\generated._69[1] ));
 sg13g2_dfrbp_1 _6883_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net91),
    .D(net435),
    .Q_N(_0024_),
    .Q(\generated._69[2] ));
 sg13g2_dfrbp_1 _6884_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net90),
    .D(_0193_),
    .Q_N(\generated._891[0] ),
    .Q(\generated._844 ));
 sg13g2_dfrbp_1 _6885_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net89),
    .D(_0194_),
    .Q_N(_3286_),
    .Q(\generated._843 ));
 sg13g2_dfrbp_1 _6886_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net88),
    .D(_0195_),
    .Q_N(_3285_),
    .Q(\generated._425[1] ));
 sg13g2_dfrbp_1 _6887_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net87),
    .D(_0196_),
    .Q_N(_0022_),
    .Q(\generated._66[1] ));
 sg13g2_dfrbp_1 _6888_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net86),
    .D(_0197_),
    .Q_N(_0089_),
    .Q(\generated._66[2] ));
 sg13g2_dfrbp_1 _6889_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net85),
    .D(_0198_),
    .Q_N(_3284_),
    .Q(\generated._1087[0] ));
 sg13g2_dfrbp_1 _6890_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net84),
    .D(_0199_),
    .Q_N(_3283_),
    .Q(\generated._165[4] ));
 sg13g2_dfrbp_1 _6891_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net83),
    .D(_0200_),
    .Q_N(_3282_),
    .Q(\generated._65[2] ));
 sg13g2_dfrbp_1 _6892_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net82),
    .D(_0201_),
    .Q_N(_3281_),
    .Q(\generated._65[3] ));
 sg13g2_dfrbp_1 _6893_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net81),
    .D(_0202_),
    .Q_N(_3280_),
    .Q(\generated._65[4] ));
 sg13g2_dfrbp_1 _6894_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net80),
    .D(_0203_),
    .Q_N(_3279_),
    .Q(\generated._65[5] ));
 sg13g2_dfrbp_1 _6895_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net79),
    .D(_0204_),
    .Q_N(_3278_),
    .Q(\generated._65[6] ));
 sg13g2_dfrbp_1 _6896_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net78),
    .D(_0205_),
    .Q_N(_0080_),
    .Q(\generated._64[0] ));
 sg13g2_dfrbp_1 _6897_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net77),
    .D(net438),
    .Q_N(_0058_),
    .Q(\generated._512[0] ));
 sg13g2_dfrbp_1 _6898_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net76),
    .D(_0207_),
    .Q_N(_0054_),
    .Q(\generated._512[1] ));
 sg13g2_dfrbp_1 _6899_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net75),
    .D(net494),
    .Q_N(_0055_),
    .Q(\generated._512[2] ));
 sg13g2_dfrbp_1 _6900_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net74),
    .D(_0209_),
    .Q_N(_0059_),
    .Q(\generated._512[3] ));
 sg13g2_dfrbp_1 _6901_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net73),
    .D(_0210_),
    .Q_N(_0062_),
    .Q(\generated._512[4] ));
 sg13g2_dfrbp_1 _6902_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net72),
    .D(_0211_),
    .Q_N(_0065_),
    .Q(\generated._512[5] ));
 sg13g2_dfrbp_1 _6903_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net71),
    .D(_0212_),
    .Q_N(_0067_),
    .Q(\generated._512[6] ));
 sg13g2_dfrbp_1 _6904_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net70),
    .D(_0213_),
    .Q_N(_0069_),
    .Q(\generated._512[7] ));
 sg13g2_dfrbp_1 _6905_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net143),
    .D(net490),
    .Q_N(_0071_),
    .Q(\generated._511 ));
 sg13g2_dfrbp_1 _6906_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net144),
    .D(\generated._695[0] ),
    .Q_N(_0036_),
    .Q(\generated._505[0] ));
 sg13g2_dfrbp_1 _6907_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net145),
    .D(\generated._695[1] ),
    .Q_N(_0044_),
    .Q(\generated._505[1] ));
 sg13g2_dfrbp_1 _6908_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net146),
    .D(\generated._695[2] ),
    .Q_N(_3344_),
    .Q(\generated._505[2] ));
 sg13g2_dfrbp_1 _6909_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net147),
    .D(net451),
    .Q_N(_0046_),
    .Q(\generated._505[3] ));
 sg13g2_dfrbp_1 _6910_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net148),
    .D(\generated._695[4] ),
    .Q_N(_3345_),
    .Q(\generated._505[4] ));
 sg13g2_dfrbp_1 _6911_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net149),
    .D(\generated._695[5] ),
    .Q_N(_3346_),
    .Q(\generated._505[5] ));
 sg13g2_dfrbp_1 _6912_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net150),
    .D(net515),
    .Q_N(_3347_),
    .Q(\generated._505[6] ));
 sg13g2_dfrbp_1 _6913_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net151),
    .D(\generated._695[7] ),
    .Q_N(_3348_),
    .Q(\generated._505[7] ));
 sg13g2_dfrbp_1 _6914_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net164),
    .D(\generated._695[8] ),
    .Q_N(_3349_),
    .Q(\generated._505[8] ));
 sg13g2_dfrbp_1 _6915_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net69),
    .D(\generated._695[9] ),
    .Q_N(_3277_),
    .Q(\generated._503 ));
 sg13g2_dfrbp_1 _6916_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net68),
    .D(net250),
    .Q_N(\generated._563[0] ),
    .Q(\generated._510 ));
 sg13g2_dfrbp_1 _6917_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net67),
    .D(_0216_),
    .Q_N(_3276_),
    .Q(\generated._509 ));
 sg13g2_dfrbp_1 _6918_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net66),
    .D(net340),
    .Q_N(_0088_),
    .Q(\generated._501[0] ));
 sg13g2_dfrbp_1 _6919_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net65),
    .D(net408),
    .Q_N(_0087_),
    .Q(\generated._381[0] ));
 sg13g2_dfrbp_1 _6920_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net64),
    .D(_0219_),
    .Q_N(_0093_),
    .Q(\generated._381[1] ));
 sg13g2_dfrbp_1 _6921_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net63),
    .D(net521),
    .Q_N(_0094_),
    .Q(\generated._381[2] ));
 sg13g2_dfrbp_1 _6922_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net62),
    .D(_0221_),
    .Q_N(_0086_),
    .Q(\generated._381[3] ));
 sg13g2_dfrbp_1 _6923_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net61),
    .D(_0222_),
    .Q_N(_0085_),
    .Q(\generated._381[4] ));
 sg13g2_dfrbp_1 _6924_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net60),
    .D(_0223_),
    .Q_N(_0084_),
    .Q(\generated._381[5] ));
 sg13g2_dfrbp_1 _6925_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net59),
    .D(_0224_),
    .Q_N(_0083_),
    .Q(\generated._381[6] ));
 sg13g2_dfrbp_1 _6926_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net58),
    .D(_0225_),
    .Q_N(_0082_),
    .Q(\generated._381[7] ));
 sg13g2_dfrbp_1 _6927_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net165),
    .D(net448),
    .Q_N(_0081_),
    .Q(\generated._380 ));
 sg13g2_dfrbp_1 _6928_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net166),
    .D(\generated._1023[3] ),
    .Q_N(_0092_),
    .Q(\generated._1024[3] ));
 sg13g2_dfrbp_1 _6929_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net167),
    .D(\generated._1023[4] ),
    .Q_N(_0103_),
    .Q(\generated._1024[4] ));
 sg13g2_dfrbp_1 _6930_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net168),
    .D(\generated._1023[5] ),
    .Q_N(_0104_),
    .Q(\generated._1024[5] ));
 sg13g2_dfrbp_1 _6931_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net169),
    .D(\generated._1023[6] ),
    .Q_N(_0105_),
    .Q(\generated._1024[6] ));
 sg13g2_dfrbp_1 _6932_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net170),
    .D(\generated._1023[7] ),
    .Q_N(_0111_),
    .Q(\generated._1024[7] ));
 sg13g2_dfrbp_1 _6933_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net171),
    .D(net518),
    .Q_N(_0113_),
    .Q(\generated._1024[8] ));
 sg13g2_dfrbp_1 _6934_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net172),
    .D(net543),
    .Q_N(_0115_),
    .Q(\generated._1024[9] ));
 sg13g2_dfrbp_1 _6935_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net173),
    .D(net298),
    .Q_N(_0076_),
    .Q(\generated._373[0] ));
 sg13g2_dfrbp_1 _6936_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net174),
    .D(net399),
    .Q_N(_0077_),
    .Q(\generated._373[1] ));
 sg13g2_dfrbp_1 _6937_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net175),
    .D(\generated._481[2] ),
    .Q_N(_3350_),
    .Q(\generated._373[2] ));
 sg13g2_dfrbp_1 _6938_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net176),
    .D(net469),
    .Q_N(_0078_),
    .Q(\generated._373[3] ));
 sg13g2_dfrbp_1 _6939_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net177),
    .D(\generated._481[4] ),
    .Q_N(_3351_),
    .Q(\generated._373[4] ));
 sg13g2_dfrbp_1 _6940_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net178),
    .D(\generated._481[5] ),
    .Q_N(_3352_),
    .Q(\generated._373[5] ));
 sg13g2_dfrbp_1 _6941_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net179),
    .D(\generated._481[6] ),
    .Q_N(_3353_),
    .Q(\generated._373[6] ));
 sg13g2_dfrbp_1 _6942_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net180),
    .D(\generated._481[7] ),
    .Q_N(_3354_),
    .Q(\generated._373[7] ));
 sg13g2_dfrbp_1 _6943_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net229),
    .D(\generated._481[8] ),
    .Q_N(_3355_),
    .Q(\generated._373[8] ));
 sg13g2_dfrbp_1 _6944_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net57),
    .D(net417),
    .Q_N(_3275_),
    .Q(\generated._371 ));
 sg13g2_dfrbp_1 _6945_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net56),
    .D(_0227_),
    .Q_N(_3274_),
    .Q(\generated._16[0] ));
 sg13g2_dfrbp_1 _6946_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net54),
    .D(_0228_),
    .Q_N(_3273_),
    .Q(\generated._16[1] ));
 sg13g2_dfrbp_1 _6947_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net52),
    .D(net279),
    .Q_N(_3272_),
    .Q(\generated._16[2] ));
 sg13g2_dfrbp_1 _6948_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net50),
    .D(_0230_),
    .Q_N(_3271_),
    .Q(\generated._16[3] ));
 sg13g2_dfrbp_1 _6949_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net48),
    .D(net277),
    .Q_N(_0095_),
    .Q(\generated._16[4] ));
 sg13g2_dfrbp_1 _6950_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net46),
    .D(_0232_),
    .Q_N(\generated._328[0] ),
    .Q(\generated._33[0] ));
 sg13g2_dfrbp_1 _6951_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net45),
    .D(net290),
    .Q_N(_3270_),
    .Q(\generated._33[1] ));
 sg13g2_dfrbp_1 _6952_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net44),
    .D(net284),
    .Q_N(_3269_),
    .Q(\generated._33[2] ));
 sg13g2_dfrbp_1 _6953_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net43),
    .D(_0235_),
    .Q_N(_3268_),
    .Q(\generated._33[3] ));
 sg13g2_dfrbp_1 _6954_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net42),
    .D(_0236_),
    .Q_N(_3267_),
    .Q(\generated._33[4] ));
 sg13g2_dfrbp_1 _6955_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net41),
    .D(_0237_),
    .Q_N(_3266_),
    .Q(\generated._33[5] ));
 sg13g2_dfrbp_1 _6956_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net40),
    .D(net270),
    .Q_N(_3265_),
    .Q(\generated._33[6] ));
 sg13g2_dfrbp_1 _6957_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net39),
    .D(net261),
    .Q_N(\generated._485[0] ),
    .Q(\generated._487[0] ));
 sg13g2_dfrbp_1 _6958_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net38),
    .D(net325),
    .Q_N(_3264_),
    .Q(\generated._487[1] ));
 sg13g2_dfrbp_1 _6959_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net37),
    .D(net441),
    .Q_N(_3263_),
    .Q(\generated._487[2] ));
 sg13g2_dfrbp_1 _6960_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net35),
    .D(net397),
    .Q_N(_3262_),
    .Q(\generated._487[3] ));
 sg13g2_dfrbp_1 _6961_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net28),
    .D(_0243_),
    .Q_N(\generated._395[0] ),
    .Q(\generated._379 ));
 sg13g2_dfrbp_1 _6962_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net27),
    .D(_0244_),
    .Q_N(_3261_),
    .Q(\generated._378 ));
 sg13g2_dfrbp_1 _6963_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net26),
    .D(_0245_),
    .Q_N(_3260_),
    .Q(\generated._346[0] ));
 sg13g2_dfrbp_1 _6964_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net241),
    .D(_0246_),
    .Q_N(_0098_),
    .Q(\generated._346[1] ));
 sg13g2_dfrbp_1 _6965_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net239),
    .D(_0247_),
    .Q_N(_0097_),
    .Q(\generated._346[2] ));
 sg13g2_dfrbp_1 _6966_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net237),
    .D(_0248_),
    .Q_N(_0096_),
    .Q(\generated._346[3] ));
 sg13g2_dfrbp_1 _6967_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net228),
    .D(_0249_),
    .Q_N(_3259_),
    .Q(\generated._346[4] ));
 sg13g2_dfrbp_1 _6968_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net226),
    .D(net387),
    .Q_N(_3258_),
    .Q(\generated._346[5] ));
 sg13g2_dfrbp_1 _6969_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net224),
    .D(net421),
    .Q_N(_3257_),
    .Q(\generated._394[0] ));
 sg13g2_dfrbp_1 _6970_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net223),
    .D(_0252_),
    .Q_N(_0052_),
    .Q(\generated._394[1] ));
 sg13g2_dfrbp_1 _6971_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net215),
    .D(_0253_),
    .Q_N(_0053_),
    .Q(\generated._394[2] ));
 sg13g2_dfrbp_1 _6972_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net213),
    .D(_0254_),
    .Q_N(_0050_),
    .Q(\generated._394[3] ));
 sg13g2_dfrbp_1 _6973_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net211),
    .D(_0255_),
    .Q_N(_0048_),
    .Q(\generated._394[4] ));
 sg13g2_dfrbp_1 _6974_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net209),
    .D(net502),
    .Q_N(_0049_),
    .Q(\generated._394[5] ));
 sg13g2_dfrbp_1 _6975_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net207),
    .D(net546),
    .Q_N(_0051_),
    .Q(\generated._394[6] ));
 sg13g2_dfrbp_1 _6976_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net205),
    .D(_0258_),
    .Q_N(_0056_),
    .Q(\generated._394[7] ));
 sg13g2_dfrbp_1 _6977_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net203),
    .D(_0259_),
    .Q_N(_0060_),
    .Q(\generated._394[8] ));
 sg13g2_dfrbp_1 _6978_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net201),
    .D(_0260_),
    .Q_N(_0063_),
    .Q(\generated._394[9] ));
 sg13g2_dfrbp_1 _6979_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net199),
    .D(_0261_),
    .Q_N(_3256_),
    .Q(\generated._28[0] ));
 sg13g2_dfrbp_1 _6980_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net126),
    .D(_0262_),
    .Q_N(_3255_),
    .Q(\generated._28[1] ));
 sg13g2_dfrbp_1 _6981_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net122),
    .D(_0263_),
    .Q_N(_3254_),
    .Q(\generated._28[2] ));
 sg13g2_dfrbp_1 _6982_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net118),
    .D(net378),
    .Q_N(_3253_),
    .Q(\generated._28[3] ));
 sg13g2_dfrbp_1 _6983_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net104),
    .D(_0265_),
    .Q_N(\generated._353[0] ),
    .Q(\generated._357[0] ));
 sg13g2_dfrbp_1 _6984_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net102),
    .D(net273),
    .Q_N(_3252_),
    .Q(\generated._357[1] ));
 sg13g2_dfrbp_1 _6985_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net55),
    .D(_0267_),
    .Q_N(_3251_),
    .Q(\generated._357[2] ));
 sg13g2_dfrbp_1 _6986_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net53),
    .D(_0268_),
    .Q_N(_3250_),
    .Q(\generated._357[3] ));
 sg13g2_dfrbp_1 _6987_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net51),
    .D(_0269_),
    .Q_N(_3249_),
    .Q(\generated._357[4] ));
 sg13g2_dfrbp_1 _6988_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net49),
    .D(_0270_),
    .Q_N(\generated._301[0] ),
    .Q(\generated._21[0] ));
 sg13g2_dfrbp_1 _6989_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net47),
    .D(_0271_),
    .Q_N(_3248_),
    .Q(\generated._21[1] ));
 sg13g2_dfrbp_1 _6990_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net242),
    .D(net293),
    .Q_N(_3247_),
    .Q(\generated._21[2] ));
 sg13g2_dfrbp_1 _6991_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net240),
    .D(_0273_),
    .Q_N(_3246_),
    .Q(\generated._21[3] ));
 sg13g2_dfrbp_1 _6992_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net230),
    .D(_0274_),
    .Q_N(_3356_),
    .Q(\generated._21[4] ));
 sg13g2_dfrbp_1 _6993_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net231),
    .D(\generated._1073[3] ),
    .Q_N(_0102_),
    .Q(\generated._1074[3] ));
 sg13g2_dfrbp_1 _6994_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net232),
    .D(\generated._1073[4] ),
    .Q_N(_0110_),
    .Q(\generated._1074[4] ));
 sg13g2_dfrbp_1 _6995_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net233),
    .D(\generated._1073[5] ),
    .Q_N(_0112_),
    .Q(\generated._1074[5] ));
 sg13g2_dfrbp_1 _6996_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net234),
    .D(\generated._1073[6] ),
    .Q_N(_0114_),
    .Q(\generated._1074[6] ));
 sg13g2_dfrbp_1 _6997_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net235),
    .D(\generated._1073[7] ),
    .Q_N(_0016_),
    .Q(\generated._1074[7] ));
 sg13g2_dfrbp_1 _6998_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net106),
    .D(\generated._1073[8] ),
    .Q_N(_0017_),
    .Q(\generated._1074[8] ));
 sg13g2_dfrbp_1 _6999_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net238),
    .D(net460),
    .Q_N(_0107_),
    .Q(\generated._1074[9] ));
 sg13g2_dfrbp_1 _7000_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net236),
    .D(_0275_),
    .Q_N(_3245_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _7001_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net227),
    .D(_0276_),
    .Q_N(_3244_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _7002_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net225),
    .D(_0277_),
    .Q_N(_3243_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _7003_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net197),
    .D(_0278_),
    .Q_N(_3242_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _7004_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net124),
    .D(_0279_),
    .Q_N(_3241_),
    .Q(\generated._123 ));
 sg13g2_dfrbp_1 _7005_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net120),
    .D(_0280_),
    .Q_N(_3240_),
    .Q(\generated._115 ));
 sg13g2_tiehi _6779__17 (.L_HI(net17));
 sg13g2_tiehi _6780__18 (.L_HI(net18));
 sg13g2_tiehi _6781__19 (.L_HI(net19));
 sg13g2_tiehi _6782__20 (.L_HI(net20));
 sg13g2_tiehi _6783__21 (.L_HI(net21));
 sg13g2_tiehi _6784__22 (.L_HI(net22));
 sg13g2_tiehi _6785__23 (.L_HI(net23));
 sg13g2_tiehi _6786__24 (.L_HI(net24));
 sg13g2_tiehi _6787__25 (.L_HI(net25));
 sg13g2_tiehi _6963__26 (.L_HI(net26));
 sg13g2_tiehi _6962__27 (.L_HI(net27));
 sg13g2_tiehi _6961__28 (.L_HI(net28));
 sg13g2_tiehi _6788__29 (.L_HI(net29));
 sg13g2_tiehi _6792__30 (.L_HI(net30));
 sg13g2_tiehi _6793__31 (.L_HI(net31));
 sg13g2_tiehi _6794__32 (.L_HI(net32));
 sg13g2_tiehi _6795__33 (.L_HI(net33));
 sg13g2_tiehi _6796__34 (.L_HI(net34));
 sg13g2_tiehi _6960__35 (.L_HI(net35));
 sg13g2_tiehi _6797__36 (.L_HI(net36));
 sg13g2_tiehi _6959__37 (.L_HI(net37));
 sg13g2_tiehi _6958__38 (.L_HI(net38));
 sg13g2_tiehi _6957__39 (.L_HI(net39));
 sg13g2_tiehi _6956__40 (.L_HI(net40));
 sg13g2_tiehi _6955__41 (.L_HI(net41));
 sg13g2_tiehi _6954__42 (.L_HI(net42));
 sg13g2_tiehi _6953__43 (.L_HI(net43));
 sg13g2_tiehi _6952__44 (.L_HI(net44));
 sg13g2_tiehi _6951__45 (.L_HI(net45));
 sg13g2_tiehi _6950__46 (.L_HI(net46));
 sg13g2_tiehi _6989__47 (.L_HI(net47));
 sg13g2_tiehi _6949__48 (.L_HI(net48));
 sg13g2_tiehi _6988__49 (.L_HI(net49));
 sg13g2_tiehi _6948__50 (.L_HI(net50));
 sg13g2_tiehi _6987__51 (.L_HI(net51));
 sg13g2_tiehi _6947__52 (.L_HI(net52));
 sg13g2_tiehi _6986__53 (.L_HI(net53));
 sg13g2_tiehi _6946__54 (.L_HI(net54));
 sg13g2_tiehi _6985__55 (.L_HI(net55));
 sg13g2_tiehi _6945__56 (.L_HI(net56));
 sg13g2_tiehi _6944__57 (.L_HI(net57));
 sg13g2_tiehi _6926__58 (.L_HI(net58));
 sg13g2_tiehi _6925__59 (.L_HI(net59));
 sg13g2_tiehi _6924__60 (.L_HI(net60));
 sg13g2_tiehi _6923__61 (.L_HI(net61));
 sg13g2_tiehi _6922__62 (.L_HI(net62));
 sg13g2_tiehi _6921__63 (.L_HI(net63));
 sg13g2_tiehi _6920__64 (.L_HI(net64));
 sg13g2_tiehi _6919__65 (.L_HI(net65));
 sg13g2_tiehi _6918__66 (.L_HI(net66));
 sg13g2_tiehi _6917__67 (.L_HI(net67));
 sg13g2_tiehi _6916__68 (.L_HI(net68));
 sg13g2_tiehi _6915__69 (.L_HI(net69));
 sg13g2_tiehi _6904__70 (.L_HI(net70));
 sg13g2_tiehi _6903__71 (.L_HI(net71));
 sg13g2_tiehi _6902__72 (.L_HI(net72));
 sg13g2_tiehi _6901__73 (.L_HI(net73));
 sg13g2_tiehi _6900__74 (.L_HI(net74));
 sg13g2_tiehi _6899__75 (.L_HI(net75));
 sg13g2_tiehi _6898__76 (.L_HI(net76));
 sg13g2_tiehi _6897__77 (.L_HI(net77));
 sg13g2_tiehi _6896__78 (.L_HI(net78));
 sg13g2_tiehi _6895__79 (.L_HI(net79));
 sg13g2_tiehi _6894__80 (.L_HI(net80));
 sg13g2_tiehi _6893__81 (.L_HI(net81));
 sg13g2_tiehi _6892__82 (.L_HI(net82));
 sg13g2_tiehi _6891__83 (.L_HI(net83));
 sg13g2_tiehi _6890__84 (.L_HI(net84));
 sg13g2_tiehi _6889__85 (.L_HI(net85));
 sg13g2_tiehi _6888__86 (.L_HI(net86));
 sg13g2_tiehi _6887__87 (.L_HI(net87));
 sg13g2_tiehi _6886__88 (.L_HI(net88));
 sg13g2_tiehi _6885__89 (.L_HI(net89));
 sg13g2_tiehi _6884__90 (.L_HI(net90));
 sg13g2_tiehi _6883__91 (.L_HI(net91));
 sg13g2_tiehi _6882__92 (.L_HI(net92));
 sg13g2_tiehi _6881__93 (.L_HI(net93));
 sg13g2_tiehi _6880__94 (.L_HI(net94));
 sg13g2_tiehi _6869__95 (.L_HI(net95));
 sg13g2_tiehi _6868__96 (.L_HI(net96));
 sg13g2_tiehi _6867__97 (.L_HI(net97));
 sg13g2_tiehi _6866__98 (.L_HI(net98));
 sg13g2_tiehi _6865__99 (.L_HI(net99));
 sg13g2_tiehi _6864__100 (.L_HI(net100));
 sg13g2_tiehi _6863__101 (.L_HI(net101));
 sg13g2_tiehi _6984__102 (.L_HI(net102));
 sg13g2_tiehi _6862__103 (.L_HI(net103));
 sg13g2_tiehi _6983__104 (.L_HI(net104));
 sg13g2_tiehi _6861__105 (.L_HI(net105));
 sg13g2_tiehi _6998__106 (.L_HI(net106));
 sg13g2_tiehi _6799__107 (.L_HI(net107));
 sg13g2_tiehi _6870__108 (.L_HI(net108));
 sg13g2_tiehi _6871__109 (.L_HI(net109));
 sg13g2_tiehi _6872__110 (.L_HI(net110));
 sg13g2_tiehi _6873__111 (.L_HI(net111));
 sg13g2_tiehi _6874__112 (.L_HI(net112));
 sg13g2_tiehi _6875__113 (.L_HI(net113));
 sg13g2_tiehi _6876__114 (.L_HI(net114));
 sg13g2_tiehi _6877__115 (.L_HI(net115));
 sg13g2_tiehi _6878__116 (.L_HI(net116));
 sg13g2_tiehi _6860__117 (.L_HI(net117));
 sg13g2_tiehi _6982__118 (.L_HI(net118));
 sg13g2_tiehi _6859__119 (.L_HI(net119));
 sg13g2_tiehi _7005__120 (.L_HI(net120));
 sg13g2_tiehi _6858__121 (.L_HI(net121));
 sg13g2_tiehi _6981__122 (.L_HI(net122));
 sg13g2_tiehi _6857__123 (.L_HI(net123));
 sg13g2_tiehi _7004__124 (.L_HI(net124));
 sg13g2_tiehi _6856__125 (.L_HI(net125));
 sg13g2_tiehi _6980__126 (.L_HI(net126));
 sg13g2_tiehi _6855__127 (.L_HI(net127));
 sg13g2_tiehi _6854__128 (.L_HI(net128));
 sg13g2_tiehi _6853__129 (.L_HI(net129));
 sg13g2_tiehi _6852__130 (.L_HI(net130));
 sg13g2_tiehi _6851__131 (.L_HI(net131));
 sg13g2_tiehi _6850__132 (.L_HI(net132));
 sg13g2_tiehi _6849__133 (.L_HI(net133));
 sg13g2_tiehi _6848__134 (.L_HI(net134));
 sg13g2_tiehi _6847__135 (.L_HI(net135));
 sg13g2_tiehi _6846__136 (.L_HI(net136));
 sg13g2_tiehi _6845__137 (.L_HI(net137));
 sg13g2_tiehi _6844__138 (.L_HI(net138));
 sg13g2_tiehi _6843__139 (.L_HI(net139));
 sg13g2_tiehi _6842__140 (.L_HI(net140));
 sg13g2_tiehi _6841__141 (.L_HI(net141));
 sg13g2_tiehi _6879__142 (.L_HI(net142));
 sg13g2_tiehi _6905__143 (.L_HI(net143));
 sg13g2_tiehi _6906__144 (.L_HI(net144));
 sg13g2_tiehi _6907__145 (.L_HI(net145));
 sg13g2_tiehi _6908__146 (.L_HI(net146));
 sg13g2_tiehi _6909__147 (.L_HI(net147));
 sg13g2_tiehi _6910__148 (.L_HI(net148));
 sg13g2_tiehi _6911__149 (.L_HI(net149));
 sg13g2_tiehi _6912__150 (.L_HI(net150));
 sg13g2_tiehi _6913__151 (.L_HI(net151));
 sg13g2_tiehi _6840__152 (.L_HI(net152));
 sg13g2_tiehi _6839__153 (.L_HI(net153));
 sg13g2_tiehi _6838__154 (.L_HI(net154));
 sg13g2_tiehi _6837__155 (.L_HI(net155));
 sg13g2_tiehi _6836__156 (.L_HI(net156));
 sg13g2_tiehi _6835__157 (.L_HI(net157));
 sg13g2_tiehi _6834__158 (.L_HI(net158));
 sg13g2_tiehi _6833__159 (.L_HI(net159));
 sg13g2_tiehi _6832__160 (.L_HI(net160));
 sg13g2_tiehi _6831__161 (.L_HI(net161));
 sg13g2_tiehi _6830__162 (.L_HI(net162));
 sg13g2_tiehi _6829__163 (.L_HI(net163));
 sg13g2_tiehi _6914__164 (.L_HI(net164));
 sg13g2_tiehi _6927__165 (.L_HI(net165));
 sg13g2_tiehi _6928__166 (.L_HI(net166));
 sg13g2_tiehi _6929__167 (.L_HI(net167));
 sg13g2_tiehi _6930__168 (.L_HI(net168));
 sg13g2_tiehi _6931__169 (.L_HI(net169));
 sg13g2_tiehi _6932__170 (.L_HI(net170));
 sg13g2_tiehi _6933__171 (.L_HI(net171));
 sg13g2_tiehi _6934__172 (.L_HI(net172));
 sg13g2_tiehi _6935__173 (.L_HI(net173));
 sg13g2_tiehi _6936__174 (.L_HI(net174));
 sg13g2_tiehi _6937__175 (.L_HI(net175));
 sg13g2_tiehi _6938__176 (.L_HI(net176));
 sg13g2_tiehi _6939__177 (.L_HI(net177));
 sg13g2_tiehi _6940__178 (.L_HI(net178));
 sg13g2_tiehi _6941__179 (.L_HI(net179));
 sg13g2_tiehi _6942__180 (.L_HI(net180));
 sg13g2_tiehi _6828__181 (.L_HI(net181));
 sg13g2_tiehi _6827__182 (.L_HI(net182));
 sg13g2_tiehi _6826__183 (.L_HI(net183));
 sg13g2_tiehi _6825__184 (.L_HI(net184));
 sg13g2_tiehi _6824__185 (.L_HI(net185));
 sg13g2_tiehi _6823__186 (.L_HI(net186));
 sg13g2_tiehi _6822__187 (.L_HI(net187));
 sg13g2_tiehi _6821__188 (.L_HI(net188));
 sg13g2_tiehi _6820__189 (.L_HI(net189));
 sg13g2_tiehi _6819__190 (.L_HI(net190));
 sg13g2_tiehi _6818__191 (.L_HI(net191));
 sg13g2_tiehi _6817__192 (.L_HI(net192));
 sg13g2_tiehi _6816__193 (.L_HI(net193));
 sg13g2_tiehi _6815__194 (.L_HI(net194));
 sg13g2_tiehi _6814__195 (.L_HI(net195));
 sg13g2_tiehi _6813__196 (.L_HI(net196));
 sg13g2_tiehi _7003__197 (.L_HI(net197));
 sg13g2_tiehi _6812__198 (.L_HI(net198));
 sg13g2_tiehi _6979__199 (.L_HI(net199));
 sg13g2_tiehi _6811__200 (.L_HI(net200));
 sg13g2_tiehi _6978__201 (.L_HI(net201));
 sg13g2_tiehi _6810__202 (.L_HI(net202));
 sg13g2_tiehi _6977__203 (.L_HI(net203));
 sg13g2_tiehi _6809__204 (.L_HI(net204));
 sg13g2_tiehi _6976__205 (.L_HI(net205));
 sg13g2_tiehi _6808__206 (.L_HI(net206));
 sg13g2_tiehi _6975__207 (.L_HI(net207));
 sg13g2_tiehi _6807__208 (.L_HI(net208));
 sg13g2_tiehi _6974__209 (.L_HI(net209));
 sg13g2_tiehi _6806__210 (.L_HI(net210));
 sg13g2_tiehi _6973__211 (.L_HI(net211));
 sg13g2_tiehi _6805__212 (.L_HI(net212));
 sg13g2_tiehi _6972__213 (.L_HI(net213));
 sg13g2_tiehi _6804__214 (.L_HI(net214));
 sg13g2_tiehi _6971__215 (.L_HI(net215));
 sg13g2_tiehi _6803__216 (.L_HI(net216));
 sg13g2_tiehi _6802__217 (.L_HI(net217));
 sg13g2_tiehi _6801__218 (.L_HI(net218));
 sg13g2_tiehi _6800__219 (.L_HI(net219));
 sg13g2_tiehi _6798__220 (.L_HI(net220));
 sg13g2_tiehi _6791__221 (.L_HI(net221));
 sg13g2_tiehi _6790__222 (.L_HI(net222));
 sg13g2_tiehi _6970__223 (.L_HI(net223));
 sg13g2_tiehi _6969__224 (.L_HI(net224));
 sg13g2_tiehi _7002__225 (.L_HI(net225));
 sg13g2_tiehi _6968__226 (.L_HI(net226));
 sg13g2_tiehi _7001__227 (.L_HI(net227));
 sg13g2_tiehi _6967__228 (.L_HI(net228));
 sg13g2_tiehi _6943__229 (.L_HI(net229));
 sg13g2_tiehi _6992__230 (.L_HI(net230));
 sg13g2_tiehi _6993__231 (.L_HI(net231));
 sg13g2_tiehi _6994__232 (.L_HI(net232));
 sg13g2_tiehi _6995__233 (.L_HI(net233));
 sg13g2_tiehi _6996__234 (.L_HI(net234));
 sg13g2_tiehi _6997__235 (.L_HI(net235));
 sg13g2_tiehi _7000__236 (.L_HI(net236));
 sg13g2_tiehi _6966__237 (.L_HI(net237));
 sg13g2_tiehi _6999__238 (.L_HI(net238));
 sg13g2_tiehi _6965__239 (.L_HI(net239));
 sg13g2_tiehi _6991__240 (.L_HI(net240));
 sg13g2_tiehi _6964__241 (.L_HI(net241));
 sg13g2_tiehi _6990__242 (.L_HI(net242));
 sg13g2_tiehi _6789__243 (.L_HI(net243));
 sg13g2_tiehi _6776__244 (.L_HI(net244));
 sg13g2_tiehi _6777__245 (.L_HI(net245));
 sg13g2_tiehi tt_um_edwintorok_246 (.L_HI(net246));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_edwintorok_3 (.L_LO(net3));
 sg13g2_tielo tt_um_edwintorok_4 (.L_LO(net4));
 sg13g2_tielo tt_um_edwintorok_5 (.L_LO(net5));
 sg13g2_tielo tt_um_edwintorok_6 (.L_LO(net6));
 sg13g2_tielo tt_um_edwintorok_7 (.L_LO(net7));
 sg13g2_tielo tt_um_edwintorok_8 (.L_LO(net8));
 sg13g2_tielo tt_um_edwintorok_9 (.L_LO(net9));
 sg13g2_tielo tt_um_edwintorok_10 (.L_LO(net10));
 sg13g2_tielo tt_um_edwintorok_11 (.L_LO(net11));
 sg13g2_tielo tt_um_edwintorok_12 (.L_LO(net12));
 sg13g2_tielo tt_um_edwintorok_13 (.L_LO(net13));
 sg13g2_tielo tt_um_edwintorok_14 (.L_LO(net14));
 sg13g2_tielo tt_um_edwintorok_15 (.L_LO(net15));
 sg13g2_tiehi _6778__16 (.L_HI(net16));
 sg13g2_buf_2 _7251_ (.A(audio),
    .X(uio_out[7]));
 sg13g2_buf_1 _7252_ (.A(\generated._115 ),
    .X(uo_out[3]));
 sg13g2_buf_1 _7253_ (.A(\generated._123 ),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout567 (.X(net567),
    .A(_1742_));
 sg13g2_buf_4 fanout568 (.X(net568),
    .A(_1515_));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(_0639_));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(_2153_));
 sg13g2_buf_4 fanout571 (.X(net571),
    .A(net572));
 sg13g2_buf_2 fanout572 (.A(_0638_),
    .X(net572));
 sg13g2_buf_4 fanout573 (.X(net573),
    .A(net574));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(_0637_));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(_2148_));
 sg13g2_buf_2 fanout576 (.A(_1661_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_0900_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_1669_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_0870_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_1682_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_1459_),
    .X(net581));
 sg13g2_buf_1 fanout582 (.A(_1459_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_0807_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_1985_),
    .X(net584));
 sg13g2_buf_1 fanout585 (.A(_1985_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_1979_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_1978_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(net589),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_1445_),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_0762_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(net593),
    .X(net592));
 sg13g2_buf_1 fanout593 (.A(_0557_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_0454_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_1995_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_0664_),
    .X(net596));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(_0663_));
 sg13g2_buf_2 fanout598 (.A(net600),
    .X(net598));
 sg13g2_buf_1 fanout599 (.A(net600),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_0437_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_0328_),
    .X(net601));
 sg13g2_buf_4 fanout602 (.X(net602),
    .A(_0322_));
 sg13g2_buf_1 fanout603 (.A(_0322_),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_1966_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_1222_),
    .X(net605));
 sg13g2_buf_4 fanout606 (.X(net606),
    .A(_0343_));
 sg13g2_buf_1 fanout607 (.A(_0343_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(net609),
    .X(net608));
 sg13g2_buf_4 fanout609 (.X(net609),
    .A(_0342_));
 sg13g2_buf_2 fanout610 (.A(net611),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_0331_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(net613),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_0331_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_1 fanout615 (.A(net617),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_0321_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(net619),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_3018_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(net622),
    .X(net620));
 sg13g2_buf_1 fanout621 (.A(net622),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_3018_),
    .X(net622));
 sg13g2_buf_4 fanout623 (.X(net623),
    .A(net625));
 sg13g2_buf_2 fanout624 (.A(net625),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_2883_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(net627),
    .X(net626));
 sg13g2_buf_4 fanout627 (.X(net627),
    .A(_1044_));
 sg13g2_buf_4 fanout628 (.X(net628),
    .A(net631));
 sg13g2_buf_2 fanout629 (.A(net630),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(net631),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_1043_),
    .X(net631));
 sg13g2_buf_4 fanout632 (.X(net632),
    .A(net633));
 sg13g2_buf_4 fanout633 (.X(net633),
    .A(_0592_));
 sg13g2_buf_2 fanout634 (.A(net635),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(net639),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(net639),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(net639),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(net639),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_0591_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(net641),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(net642),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_0335_),
    .X(net642));
 sg13g2_buf_4 fanout643 (.X(net643),
    .A(_0335_));
 sg13g2_buf_2 fanout644 (.A(_0335_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(net647),
    .X(net645));
 sg13g2_buf_1 fanout646 (.A(net647),
    .X(net646));
 sg13g2_buf_4 fanout647 (.X(net647),
    .A(_0334_));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(net651));
 sg13g2_buf_2 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(net651),
    .X(net650));
 sg13g2_buf_4 fanout651 (.X(net651),
    .A(_3013_));
 sg13g2_buf_4 fanout652 (.X(net652),
    .A(net653));
 sg13g2_buf_2 fanout653 (.A(net654),
    .X(net653));
 sg13g2_buf_4 fanout654 (.X(net654),
    .A(_3012_));
 sg13g2_buf_2 fanout655 (.A(_0395_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_2854_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_2854_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(\generated._394[0] ),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(net660),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_1 fanout661 (.A(net663),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(net663),
    .X(net662));
 sg13g2_buf_1 fanout663 (.A(net664),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(\generated._378 ),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(net668),
    .X(net665));
 sg13g2_buf_1 fanout666 (.A(net668),
    .X(net666));
 sg13g2_buf_4 fanout667 (.X(net667),
    .A(net668));
 sg13g2_buf_2 fanout668 (.A(\generated._379 ),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(net670),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(net671),
    .X(net670));
 sg13g2_buf_4 fanout671 (.X(net671),
    .A(\generated._371 ));
 sg13g2_buf_2 fanout672 (.A(\generated._501[0] ),
    .X(net672));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(\generated._509 ));
 sg13g2_buf_1 fanout674 (.A(\generated._509 ),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(net678),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(net677),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_1 fanout678 (.A(\generated._509 ),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(net683),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(net682),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(net683),
    .X(net681));
 sg13g2_buf_1 fanout682 (.A(net683),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(\generated._510 ),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(net685),
    .X(net684));
 sg13g2_buf_4 fanout685 (.X(net685),
    .A(\generated._503 ));
 sg13g2_buf_4 fanout686 (.X(net686),
    .A(net548));
 sg13g2_buf_2 fanout687 (.A(\generated._65[3] ),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(\generated._66[2] ),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(\generated._66[1] ),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(\generated._843 ),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(net694),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(net694),
    .X(net693));
 sg13g2_buf_4 fanout694 (.X(net694),
    .A(\generated._843 ));
 sg13g2_buf_4 fanout695 (.X(net695),
    .A(net699));
 sg13g2_buf_2 fanout696 (.A(net699),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(net699),
    .X(net697));
 sg13g2_buf_1 fanout698 (.A(net699),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(\generated._844 ),
    .X(net699));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(\generated._562[0] ));
 sg13g2_buf_2 fanout701 (.A(net703),
    .X(net701));
 sg13g2_buf_1 fanout702 (.A(net703),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(net353),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(net706),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(net706),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(\generated._969 ),
    .X(net706));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(net710));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(net710));
 sg13g2_buf_2 fanout709 (.A(net710),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(\generated._970 ),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(net716),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(net713),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(net716),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(net715),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(net716),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(\generated._1084[9] ),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(net719),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(net719),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(\generated._1084[9] ),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(\generated._100[9] ),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(net537),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(\generated._100[7] ),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(net724),
    .X(net723));
 sg13g2_buf_1 fanout724 (.A(\generated._100[4] ),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(net726),
    .X(net725));
 sg13g2_buf_4 fanout726 (.X(net726),
    .A(net563));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(net411));
 sg13g2_buf_1 fanout728 (.A(\generated._614[5] ),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(net267),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(net413),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(net459),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(\generated._66[9] ),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(\generated._66[8] ),
    .X(net733));
 sg13g2_buf_4 fanout734 (.X(net734),
    .A(\generated._66[7] ));
 sg13g2_buf_2 fanout735 (.A(\generated._66[6] ),
    .X(net735));
 sg13g2_buf_1 fanout736 (.A(\generated._66[6] ),
    .X(net736));
 sg13g2_buf_4 fanout737 (.X(net737),
    .A(\generated._66[5] ));
 sg13g2_buf_4 fanout738 (.X(net738),
    .A(\generated._66[4] ));
 sg13g2_buf_2 fanout739 (.A(\generated._66[4] ),
    .X(net739));
 sg13g2_buf_4 fanout740 (.X(net740),
    .A(\generated._66[3] ));
 sg13g2_buf_2 fanout741 (.A(net742),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(net743),
    .X(net742));
 sg13g2_buf_4 fanout743 (.X(net743),
    .A(_2844_));
 sg13g2_buf_2 fanout744 (.A(net1),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(net747),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(net747),
    .X(net746));
 sg13g2_buf_4 fanout747 (.X(net747),
    .A(net749));
 sg13g2_buf_2 fanout748 (.A(net749),
    .X(net748));
 sg13g2_buf_4 fanout749 (.X(net749),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(uio_in[0]),
    .X(net1));
 sg13g2_tielo tt_um_edwintorok_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_0_clk));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_32_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_34_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_1_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_30_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_31_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_25_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_29_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_22_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_23_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_24_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_3_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_4_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_8_clk));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_5_clk));
 sg13g2_inv_8 clkload20 (.A(clknet_leaf_6_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_7_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_18_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_10_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\generated._301[0] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold2 (.A(\generated._328[0] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold3 (.A(\generated._563[0] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0215_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold5 (.A(\generated._1025[0] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold6 (.A(\generated._891[0] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold7 (.A(\generated._395[0] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold8 (.A(\generated._1118[0] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0145_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold10 (.A(\generated._941[0] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0182_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold12 (.A(\generated._698[0] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0186_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold14 (.A(\generated._485[0] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0239_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold16 (.A(\generated._1076[0] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0165_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold18 (.A(\generated._353[0] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold19 (.A(\generated._77[0] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0174_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold21 (.A(\generated._614[4] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0126_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold23 (.A(\generated._33[6] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0238_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold25 (.A(\generated._357[0] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold26 (.A(_2780_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0266_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold28 (.A(\generated._33[3] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold29 (.A(_2664_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold30 (.A(\generated._16[4] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0231_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold32 (.A(\generated._16[2] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0229_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold34 (.A(\generated._100[8] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold35 (.A(_1313_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold36 (.A(\generated._33[2] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold37 (.A(_2663_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0234_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold39 (.A(\generated._100[2] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold40 (.A(_1305_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0147_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold42 (.A(\generated._33[0] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold43 (.A(_2662_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0233_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold45 (.A(\generated._21[2] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold46 (.A(_2788_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0272_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0100_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold49 (.A(_1247_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0075_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold51 (.A(_1045_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold52 (.A(\generated._481[0] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0098_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold54 (.A(\generated._63[1] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0187_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold56 (.A(\generated._100[7] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold57 (.A(\generated._406[1] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold58 (.A(_1374_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0175_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold60 (.A(\generated._71[0] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0183_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold62 (.A(\generated._33[5] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold63 (.A(_2667_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold64 (.A(\generated._406[5] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold65 (.A(_1382_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0179_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold67 (.A(\generated._346[1] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0101_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold69 (.A(_1249_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold70 (.A(\generated._346[3] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold71 (.A(_2905_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold72 (.A(\generated._406[7] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0181_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold74 (.A(\generated._357[4] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold75 (.A(_2785_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold76 (.A(\generated._28[0] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold77 (.A(_2771_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold78 (.A(\generated._487[1] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0240_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0035_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold81 (.A(\generated._357[2] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold82 (.A(_2781_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold83 (.A(\generated._406[6] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0180_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold85 (.A(\generated._434[19] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0144_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold87 (.A(\generated._1078[0] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0166_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold89 (.A(\generated._1084[0] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold90 (.A(_1324_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold91 (.A(\generated._16[1] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold92 (.A(_2652_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold93 (.A(\generated._501[0] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0217_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold95 (.A(\generated._346[4] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold96 (.A(\generated._221[1] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold97 (.A(_1243_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold98 (.A(\generated._21[0] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold99 (.A(_2786_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold100 (.A(\generated._21[3] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold101 (.A(_2790_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold102 (.A(\generated._16[3] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold103 (.A(\generated._21[4] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold104 (.A(\generated._614[2] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold105 (.A(_1230_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0124_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold107 (.A(\generated._969 ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold108 (.A(\generated._100[0] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold109 (.A(_1304_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold110 (.A(\generated._33[4] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold111 (.A(\generated._1024[0] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold112 (.A(\generated._357[3] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold113 (.A(\generated._16[0] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold114 (.A(\generated._221[0] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold115 (.A(_1240_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold116 (.A(\generated._406[4] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold117 (.A(_1381_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold118 (.A(\generated._69[0] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0190_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold120 (.A(\generated._100[9] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold121 (.A(\generated._28[2] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold122 (.A(_2777_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold123 (.A(\generated._434[10] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold124 (.A(_1259_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold125 (.A(\generated._406[3] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold126 (.A(_1380_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold127 (.A(\generated._28[1] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0036_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0605_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold130 (.A(\generated._63[2] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold131 (.A(\generated._28[3] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0264_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold133 (.A(\generated._614[1] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0123_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold135 (.A(\generated._100[6] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold136 (.A(_1309_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold137 (.A(\generated._505[8] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold138 (.A(\generated._346[2] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold139 (.A(_2914_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold140 (.A(\generated._346[5] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0250_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold142 (.A(\generated._100[5] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0150_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold144 (.A(\generated._1074[0] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold145 (.A(\generated._1078[3] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold146 (.A(_1367_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0168_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold148 (.A(\generated._16[0] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold149 (.A(\generated._487[3] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold150 (.A(_2674_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0242_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0076_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold153 (.A(\generated._481[1] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold154 (.A(\generated._71[3] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold155 (.A(_1392_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0185_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold157 (.A(\generated._63[3] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold158 (.A(_1397_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0189_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0088_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold161 (.A(_2574_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0218_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0030_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0106_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold165 (.A(\generated._614[5] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold166 (.A(_1236_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold167 (.A(\generated._614[3] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0125_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold169 (.A(\generated._373[8] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold170 (.A(_1138_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold171 (.A(\generated._481[9] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold172 (.A(\generated._406[2] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold173 (.A(_1377_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold174 (.A(\generated._394[0] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0251_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold176 (.A(\generated._1084[2] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0158_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0034_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0471_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold180 (.A(\generated._938[8] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold181 (.A(\generated._614[0] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold182 (.A(\generated._1084[8] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold183 (.A(\generated._1024[2] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold184 (.A(_1252_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold185 (.A(\generated._425[1] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0110_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0024_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold188 (.A(_1400_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0192_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0080_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold191 (.A(_2478_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0206_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold193 (.A(\generated._487[2] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold194 (.A(_2673_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0241_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold196 (.A(\generated._100[3] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold197 (.A(_1306_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0022_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold199 (.A(\generated._63[0] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold200 (.A(\generated._434[14] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0082_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0226_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0046_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0680_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold205 (.A(\generated._695[3] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold206 (.A(\generated._71[2] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold207 (.A(_1391_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0184_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold209 (.A(\generated._381[3] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold210 (.A(\generated._1078[2] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold211 (.A(_1366_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0167_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold213 (.A(\generated._66[9] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold214 (.A(\generated._1073[9] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0108_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold216 (.A(_1370_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold217 (.A(\generated._434[16] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold218 (.A(_1286_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold219 (.A(\generated._1084[5] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0067_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold221 (.A(_2548_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0078_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold223 (.A(\generated._481[3] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold224 (.A(\generated._434[15] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold225 (.A(_1283_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold226 (.A(\generated._346[0] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold227 (.A(\generated._512[5] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold228 (.A(_2529_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0109_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold230 (.A(_1369_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0170_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold232 (.A(\generated._1024[7] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0299_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0047_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold235 (.A(_1294_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0143_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold237 (.A(\generated._69[8] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold238 (.A(\generated._938[9] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold239 (.A(\generated._394[7] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold240 (.A(\generated._221[2] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold241 (.A(\generated._434[13] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0138_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0069_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0214_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold245 (.A(\generated._381[1] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold246 (.A(_2581_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold247 (.A(\generated._512[2] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0208_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold249 (.A(\generated._394[8] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold250 (.A(\generated._373[7] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold251 (.A(_1122_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold252 (.A(\generated._434[12] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold253 (.A(_1265_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0137_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold255 (.A(\generated._394[4] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0256_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0065_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold258 (.A(_2539_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold259 (.A(\generated._1084[4] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0025_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold261 (.A(_1399_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0191_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0044_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold264 (.A(\generated._1024[6] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0103_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold266 (.A(_3234_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold267 (.A(\generated._394[2] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold268 (.A(\generated._505[6] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold269 (.A(\generated._695[6] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0111_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0310_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold272 (.A(\generated._1023[8] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0027_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold274 (.A(\generated._381[2] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0220_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0086_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0083_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold278 (.A(_2643_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0084_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold280 (.A(_2635_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold281 (.A(\generated._1084[7] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0162_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold283 (.A(\generated._373[7] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold284 (.A(\generated._1074[7] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold285 (.A(\generated._512[1] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0096_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold287 (.A(\generated._69[6] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0451_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold289 (.A(\generated._938[7] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0048_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold291 (.A(\generated._100[8] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0052_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold293 (.A(\generated._1024[4] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold294 (.A(\generated._505[7] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold295 (.A(\generated._512[3] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0113_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold297 (.A(\generated._1023[9] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold298 (.A(\generated._1084[4] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0051_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0257_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0028_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold302 (.A(\generated._64[0] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0018_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0381_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0029_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0422_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0423_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold308 (.A(\generated._434[17] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold309 (.A(_1291_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0053_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0008_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0059_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold313 (.A(\generated._381[5] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold314 (.A(\generated._373[4] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0057_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold316 (.A(\generated._562[8] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0099_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold318 (.A(\generated._100[9] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold319 (.A(\generated._434[13] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0046_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold321 (.A(\generated._406[1] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold322 (.A(_3169_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold323 (.A(\generated._434[15] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold324 (.A(\generated._373[4] ),
    .X(net753));
 sg13g2_antennanp ANTENNA_1 (.A(_0269_));
 sg13g2_antennanp ANTENNA_2 (.A(_0269_));
 sg13g2_antennanp ANTENNA_3 (.A(_2781_));
 sg13g2_antennanp ANTENNA_4 (.A(_0269_));
 sg13g2_antennanp ANTENNA_5 (.A(_2781_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_4 FILLER_0_28 ();
 sg13g2_fill_2 FILLER_0_48 ();
 sg13g2_fill_1 FILLER_0_55 ();
 sg13g2_fill_2 FILLER_0_68 ();
 sg13g2_fill_1 FILLER_0_70 ();
 sg13g2_fill_1 FILLER_0_84 ();
 sg13g2_fill_2 FILLER_0_95 ();
 sg13g2_decap_8 FILLER_0_102 ();
 sg13g2_decap_4 FILLER_0_109 ();
 sg13g2_fill_2 FILLER_0_117 ();
 sg13g2_fill_1 FILLER_0_119 ();
 sg13g2_decap_4 FILLER_0_130 ();
 sg13g2_fill_1 FILLER_0_151 ();
 sg13g2_fill_1 FILLER_0_161 ();
 sg13g2_decap_4 FILLER_0_166 ();
 sg13g2_fill_1 FILLER_0_170 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_fill_1 FILLER_0_189 ();
 sg13g2_fill_2 FILLER_0_194 ();
 sg13g2_fill_1 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_fill_1 FILLER_0_208 ();
 sg13g2_decap_4 FILLER_0_214 ();
 sg13g2_fill_1 FILLER_0_218 ();
 sg13g2_fill_2 FILLER_0_224 ();
 sg13g2_fill_1 FILLER_0_226 ();
 sg13g2_fill_1 FILLER_0_247 ();
 sg13g2_fill_2 FILLER_0_252 ();
 sg13g2_fill_2 FILLER_0_259 ();
 sg13g2_fill_2 FILLER_0_271 ();
 sg13g2_decap_4 FILLER_0_304 ();
 sg13g2_fill_2 FILLER_0_308 ();
 sg13g2_decap_4 FILLER_0_324 ();
 sg13g2_fill_2 FILLER_0_328 ();
 sg13g2_fill_2 FILLER_0_346 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_4 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_4 FILLER_1_21 ();
 sg13g2_fill_2 FILLER_1_25 ();
 sg13g2_fill_1 FILLER_1_53 ();
 sg13g2_fill_1 FILLER_1_75 ();
 sg13g2_fill_2 FILLER_1_95 ();
 sg13g2_fill_1 FILLER_1_110 ();
 sg13g2_fill_2 FILLER_1_177 ();
 sg13g2_fill_1 FILLER_1_222 ();
 sg13g2_fill_2 FILLER_1_258 ();
 sg13g2_fill_2 FILLER_1_281 ();
 sg13g2_fill_1 FILLER_1_283 ();
 sg13g2_fill_2 FILLER_1_317 ();
 sg13g2_decap_4 FILLER_1_383 ();
 sg13g2_fill_1 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_41 ();
 sg13g2_fill_1 FILLER_2_43 ();
 sg13g2_fill_1 FILLER_2_100 ();
 sg13g2_fill_2 FILLER_2_124 ();
 sg13g2_fill_1 FILLER_2_126 ();
 sg13g2_fill_2 FILLER_2_179 ();
 sg13g2_fill_2 FILLER_2_268 ();
 sg13g2_fill_2 FILLER_2_296 ();
 sg13g2_fill_1 FILLER_2_320 ();
 sg13g2_fill_2 FILLER_2_352 ();
 sg13g2_fill_1 FILLER_2_354 ();
 sg13g2_fill_2 FILLER_2_393 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_4 FILLER_3_14 ();
 sg13g2_fill_2 FILLER_3_44 ();
 sg13g2_fill_2 FILLER_3_65 ();
 sg13g2_fill_1 FILLER_3_83 ();
 sg13g2_fill_2 FILLER_3_112 ();
 sg13g2_fill_1 FILLER_3_122 ();
 sg13g2_fill_2 FILLER_3_172 ();
 sg13g2_fill_1 FILLER_3_174 ();
 sg13g2_fill_2 FILLER_3_217 ();
 sg13g2_fill_1 FILLER_3_219 ();
 sg13g2_fill_1 FILLER_3_242 ();
 sg13g2_fill_2 FILLER_3_255 ();
 sg13g2_fill_1 FILLER_3_309 ();
 sg13g2_fill_1 FILLER_3_336 ();
 sg13g2_fill_1 FILLER_3_355 ();
 sg13g2_fill_2 FILLER_3_370 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_fill_1 FILLER_4_14 ();
 sg13g2_fill_2 FILLER_4_68 ();
 sg13g2_fill_1 FILLER_4_80 ();
 sg13g2_fill_1 FILLER_4_96 ();
 sg13g2_decap_8 FILLER_4_106 ();
 sg13g2_fill_2 FILLER_4_113 ();
 sg13g2_decap_8 FILLER_4_188 ();
 sg13g2_fill_1 FILLER_4_195 ();
 sg13g2_decap_8 FILLER_4_200 ();
 sg13g2_fill_2 FILLER_4_212 ();
 sg13g2_fill_1 FILLER_4_214 ();
 sg13g2_fill_1 FILLER_4_262 ();
 sg13g2_fill_1 FILLER_4_281 ();
 sg13g2_fill_2 FILLER_4_299 ();
 sg13g2_fill_1 FILLER_4_301 ();
 sg13g2_fill_1 FILLER_4_402 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_7 ();
 sg13g2_fill_2 FILLER_5_23 ();
 sg13g2_fill_1 FILLER_5_25 ();
 sg13g2_decap_8 FILLER_5_62 ();
 sg13g2_decap_4 FILLER_5_69 ();
 sg13g2_fill_1 FILLER_5_73 ();
 sg13g2_decap_4 FILLER_5_92 ();
 sg13g2_fill_1 FILLER_5_96 ();
 sg13g2_decap_4 FILLER_5_111 ();
 sg13g2_fill_1 FILLER_5_115 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_4 FILLER_5_182 ();
 sg13g2_fill_2 FILLER_5_186 ();
 sg13g2_fill_2 FILLER_5_212 ();
 sg13g2_fill_1 FILLER_5_214 ();
 sg13g2_fill_1 FILLER_5_401 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_6_54 ();
 sg13g2_fill_1 FILLER_6_56 ();
 sg13g2_decap_4 FILLER_6_61 ();
 sg13g2_fill_2 FILLER_6_77 ();
 sg13g2_fill_2 FILLER_6_142 ();
 sg13g2_fill_1 FILLER_6_166 ();
 sg13g2_fill_2 FILLER_6_183 ();
 sg13g2_fill_1 FILLER_6_237 ();
 sg13g2_fill_1 FILLER_6_269 ();
 sg13g2_fill_1 FILLER_6_275 ();
 sg13g2_fill_2 FILLER_6_285 ();
 sg13g2_fill_1 FILLER_6_363 ();
 sg13g2_fill_1 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_25 ();
 sg13g2_fill_1 FILLER_7_40 ();
 sg13g2_decap_8 FILLER_7_68 ();
 sg13g2_fill_2 FILLER_7_111 ();
 sg13g2_decap_4 FILLER_7_123 ();
 sg13g2_fill_1 FILLER_7_127 ();
 sg13g2_fill_1 FILLER_7_193 ();
 sg13g2_fill_2 FILLER_7_233 ();
 sg13g2_fill_2 FILLER_7_248 ();
 sg13g2_fill_1 FILLER_7_250 ();
 sg13g2_fill_2 FILLER_7_256 ();
 sg13g2_fill_1 FILLER_7_281 ();
 sg13g2_fill_1 FILLER_7_297 ();
 sg13g2_fill_2 FILLER_7_311 ();
 sg13g2_fill_1 FILLER_7_341 ();
 sg13g2_fill_2 FILLER_7_395 ();
 sg13g2_fill_1 FILLER_7_397 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_66 ();
 sg13g2_fill_1 FILLER_8_68 ();
 sg13g2_fill_1 FILLER_8_90 ();
 sg13g2_fill_2 FILLER_8_96 ();
 sg13g2_fill_1 FILLER_8_98 ();
 sg13g2_fill_2 FILLER_8_125 ();
 sg13g2_fill_1 FILLER_8_127 ();
 sg13g2_fill_1 FILLER_8_143 ();
 sg13g2_fill_2 FILLER_8_158 ();
 sg13g2_fill_1 FILLER_8_160 ();
 sg13g2_fill_2 FILLER_8_195 ();
 sg13g2_fill_1 FILLER_8_201 ();
 sg13g2_decap_4 FILLER_8_214 ();
 sg13g2_fill_2 FILLER_8_226 ();
 sg13g2_fill_1 FILLER_8_228 ();
 sg13g2_fill_2 FILLER_8_234 ();
 sg13g2_decap_4 FILLER_8_282 ();
 sg13g2_fill_2 FILLER_8_303 ();
 sg13g2_fill_1 FILLER_8_305 ();
 sg13g2_fill_1 FILLER_8_324 ();
 sg13g2_fill_1 FILLER_8_342 ();
 sg13g2_fill_1 FILLER_8_360 ();
 sg13g2_fill_2 FILLER_8_366 ();
 sg13g2_fill_1 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_9 ();
 sg13g2_decap_4 FILLER_9_23 ();
 sg13g2_fill_1 FILLER_9_27 ();
 sg13g2_fill_2 FILLER_9_84 ();
 sg13g2_fill_2 FILLER_9_96 ();
 sg13g2_fill_1 FILLER_9_98 ();
 sg13g2_fill_2 FILLER_9_103 ();
 sg13g2_fill_1 FILLER_9_113 ();
 sg13g2_fill_1 FILLER_9_124 ();
 sg13g2_decap_8 FILLER_9_173 ();
 sg13g2_decap_4 FILLER_9_183 ();
 sg13g2_fill_1 FILLER_9_187 ();
 sg13g2_decap_4 FILLER_9_192 ();
 sg13g2_decap_8 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_207 ();
 sg13g2_decap_8 FILLER_9_214 ();
 sg13g2_decap_4 FILLER_9_221 ();
 sg13g2_fill_2 FILLER_9_233 ();
 sg13g2_fill_1 FILLER_9_239 ();
 sg13g2_fill_2 FILLER_9_259 ();
 sg13g2_fill_1 FILLER_9_266 ();
 sg13g2_fill_2 FILLER_9_275 ();
 sg13g2_fill_1 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_50 ();
 sg13g2_fill_2 FILLER_10_96 ();
 sg13g2_fill_1 FILLER_10_98 ();
 sg13g2_fill_2 FILLER_10_104 ();
 sg13g2_fill_2 FILLER_10_141 ();
 sg13g2_fill_2 FILLER_10_157 ();
 sg13g2_fill_1 FILLER_10_159 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_4 FILLER_10_175 ();
 sg13g2_fill_1 FILLER_10_179 ();
 sg13g2_fill_2 FILLER_10_201 ();
 sg13g2_fill_1 FILLER_10_203 ();
 sg13g2_fill_2 FILLER_10_215 ();
 sg13g2_fill_1 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_222 ();
 sg13g2_fill_1 FILLER_10_229 ();
 sg13g2_fill_2 FILLER_10_264 ();
 sg13g2_fill_1 FILLER_10_296 ();
 sg13g2_fill_2 FILLER_10_337 ();
 sg13g2_fill_1 FILLER_10_339 ();
 sg13g2_fill_2 FILLER_10_345 ();
 sg13g2_fill_2 FILLER_10_352 ();
 sg13g2_fill_2 FILLER_10_367 ();
 sg13g2_fill_2 FILLER_10_387 ();
 sg13g2_fill_1 FILLER_10_389 ();
 sg13g2_fill_1 FILLER_10_399 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_31 ();
 sg13g2_fill_2 FILLER_11_62 ();
 sg13g2_fill_2 FILLER_11_90 ();
 sg13g2_fill_1 FILLER_11_92 ();
 sg13g2_fill_2 FILLER_11_103 ();
 sg13g2_fill_2 FILLER_11_137 ();
 sg13g2_fill_1 FILLER_11_139 ();
 sg13g2_fill_1 FILLER_11_168 ();
 sg13g2_fill_2 FILLER_11_191 ();
 sg13g2_fill_2 FILLER_11_223 ();
 sg13g2_fill_1 FILLER_11_287 ();
 sg13g2_fill_1 FILLER_11_354 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_33 ();
 sg13g2_fill_2 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_64 ();
 sg13g2_fill_1 FILLER_12_66 ();
 sg13g2_fill_2 FILLER_12_89 ();
 sg13g2_fill_1 FILLER_12_91 ();
 sg13g2_fill_2 FILLER_12_159 ();
 sg13g2_fill_1 FILLER_12_161 ();
 sg13g2_decap_4 FILLER_12_205 ();
 sg13g2_decap_4 FILLER_12_231 ();
 sg13g2_decap_4 FILLER_12_251 ();
 sg13g2_fill_2 FILLER_12_255 ();
 sg13g2_fill_2 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_282 ();
 sg13g2_fill_1 FILLER_12_292 ();
 sg13g2_fill_1 FILLER_12_313 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_22 ();
 sg13g2_decap_8 FILLER_13_29 ();
 sg13g2_fill_1 FILLER_13_41 ();
 sg13g2_fill_1 FILLER_13_67 ();
 sg13g2_fill_2 FILLER_13_81 ();
 sg13g2_fill_1 FILLER_13_83 ();
 sg13g2_fill_1 FILLER_13_148 ();
 sg13g2_decap_4 FILLER_13_153 ();
 sg13g2_fill_2 FILLER_13_157 ();
 sg13g2_fill_1 FILLER_13_173 ();
 sg13g2_decap_4 FILLER_13_191 ();
 sg13g2_fill_1 FILLER_13_195 ();
 sg13g2_fill_1 FILLER_13_201 ();
 sg13g2_decap_8 FILLER_13_234 ();
 sg13g2_fill_2 FILLER_13_241 ();
 sg13g2_fill_1 FILLER_13_303 ();
 sg13g2_fill_2 FILLER_13_321 ();
 sg13g2_fill_2 FILLER_13_349 ();
 sg13g2_fill_2 FILLER_13_373 ();
 sg13g2_fill_1 FILLER_13_375 ();
 sg13g2_fill_2 FILLER_13_388 ();
 sg13g2_fill_1 FILLER_13_390 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_15 ();
 sg13g2_decap_8 FILLER_14_25 ();
 sg13g2_decap_8 FILLER_14_32 ();
 sg13g2_fill_1 FILLER_14_104 ();
 sg13g2_fill_2 FILLER_14_114 ();
 sg13g2_fill_2 FILLER_14_150 ();
 sg13g2_decap_4 FILLER_14_183 ();
 sg13g2_fill_2 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_201 ();
 sg13g2_fill_2 FILLER_14_239 ();
 sg13g2_fill_1 FILLER_14_293 ();
 sg13g2_fill_1 FILLER_14_299 ();
 sg13g2_fill_1 FILLER_14_367 ();
 sg13g2_fill_2 FILLER_14_398 ();
 sg13g2_fill_1 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_7 ();
 sg13g2_decap_4 FILLER_15_25 ();
 sg13g2_fill_1 FILLER_15_29 ();
 sg13g2_decap_8 FILLER_15_38 ();
 sg13g2_fill_2 FILLER_15_45 ();
 sg13g2_fill_1 FILLER_15_47 ();
 sg13g2_fill_2 FILLER_15_89 ();
 sg13g2_fill_1 FILLER_15_158 ();
 sg13g2_fill_1 FILLER_15_163 ();
 sg13g2_fill_2 FILLER_15_168 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_198 ();
 sg13g2_fill_2 FILLER_15_218 ();
 sg13g2_fill_1 FILLER_15_220 ();
 sg13g2_fill_1 FILLER_15_227 ();
 sg13g2_fill_2 FILLER_15_260 ();
 sg13g2_fill_2 FILLER_15_289 ();
 sg13g2_fill_1 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_305 ();
 sg13g2_fill_1 FILLER_15_333 ();
 sg13g2_fill_2 FILLER_15_364 ();
 sg13g2_fill_2 FILLER_15_371 ();
 sg13g2_fill_2 FILLER_15_382 ();
 sg13g2_fill_1 FILLER_15_393 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_fill_1 FILLER_16_17 ();
 sg13g2_decap_4 FILLER_16_49 ();
 sg13g2_fill_1 FILLER_16_57 ();
 sg13g2_fill_2 FILLER_16_71 ();
 sg13g2_fill_1 FILLER_16_73 ();
 sg13g2_fill_2 FILLER_16_81 ();
 sg13g2_fill_2 FILLER_16_147 ();
 sg13g2_fill_1 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_fill_2 FILLER_16_172 ();
 sg13g2_fill_1 FILLER_16_174 ();
 sg13g2_decap_8 FILLER_16_191 ();
 sg13g2_fill_1 FILLER_16_198 ();
 sg13g2_fill_1 FILLER_16_210 ();
 sg13g2_fill_2 FILLER_16_216 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_fill_2 FILLER_16_277 ();
 sg13g2_fill_1 FILLER_16_279 ();
 sg13g2_fill_1 FILLER_16_295 ();
 sg13g2_fill_1 FILLER_16_353 ();
 sg13g2_fill_2 FILLER_16_372 ();
 sg13g2_fill_1 FILLER_16_394 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_70 ();
 sg13g2_fill_1 FILLER_17_141 ();
 sg13g2_fill_2 FILLER_17_164 ();
 sg13g2_decap_4 FILLER_17_187 ();
 sg13g2_fill_2 FILLER_17_191 ();
 sg13g2_fill_1 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_233 ();
 sg13g2_fill_2 FILLER_17_239 ();
 sg13g2_fill_2 FILLER_17_251 ();
 sg13g2_fill_1 FILLER_17_374 ();
 sg13g2_fill_2 FILLER_18_58 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_fill_1 FILLER_18_102 ();
 sg13g2_fill_2 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_117 ();
 sg13g2_fill_2 FILLER_18_140 ();
 sg13g2_fill_2 FILLER_18_180 ();
 sg13g2_fill_2 FILLER_18_186 ();
 sg13g2_decap_4 FILLER_18_196 ();
 sg13g2_fill_2 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_4 FILLER_18_217 ();
 sg13g2_fill_1 FILLER_18_221 ();
 sg13g2_fill_2 FILLER_18_239 ();
 sg13g2_fill_1 FILLER_18_241 ();
 sg13g2_fill_2 FILLER_18_246 ();
 sg13g2_fill_2 FILLER_18_256 ();
 sg13g2_fill_2 FILLER_18_266 ();
 sg13g2_fill_1 FILLER_18_268 ();
 sg13g2_fill_1 FILLER_18_351 ();
 sg13g2_fill_2 FILLER_18_394 ();
 sg13g2_fill_1 FILLER_18_396 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_15 ();
 sg13g2_fill_1 FILLER_19_17 ();
 sg13g2_fill_2 FILLER_19_26 ();
 sg13g2_fill_1 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_53 ();
 sg13g2_fill_1 FILLER_19_65 ();
 sg13g2_fill_1 FILLER_19_92 ();
 sg13g2_fill_1 FILLER_19_158 ();
 sg13g2_fill_2 FILLER_19_177 ();
 sg13g2_fill_1 FILLER_19_179 ();
 sg13g2_fill_2 FILLER_19_194 ();
 sg13g2_fill_1 FILLER_19_196 ();
 sg13g2_decap_4 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_fill_2 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_237 ();
 sg13g2_fill_2 FILLER_19_242 ();
 sg13g2_fill_2 FILLER_19_334 ();
 sg13g2_fill_2 FILLER_19_344 ();
 sg13g2_fill_1 FILLER_19_372 ();
 sg13g2_fill_1 FILLER_19_377 ();
 sg13g2_fill_2 FILLER_19_402 ();
 sg13g2_fill_1 FILLER_19_404 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_20 ();
 sg13g2_fill_1 FILLER_20_27 ();
 sg13g2_fill_2 FILLER_20_111 ();
 sg13g2_fill_1 FILLER_20_127 ();
 sg13g2_fill_1 FILLER_20_165 ();
 sg13g2_fill_2 FILLER_20_188 ();
 sg13g2_fill_1 FILLER_20_190 ();
 sg13g2_fill_1 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_238 ();
 sg13g2_fill_1 FILLER_20_240 ();
 sg13g2_fill_1 FILLER_20_251 ();
 sg13g2_fill_1 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_352 ();
 sg13g2_fill_2 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_17 ();
 sg13g2_fill_1 FILLER_21_19 ();
 sg13g2_fill_1 FILLER_21_33 ();
 sg13g2_fill_1 FILLER_21_67 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_96 ();
 sg13g2_fill_1 FILLER_21_148 ();
 sg13g2_fill_1 FILLER_21_156 ();
 sg13g2_fill_1 FILLER_21_167 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_fill_1 FILLER_21_223 ();
 sg13g2_fill_1 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_259 ();
 sg13g2_fill_2 FILLER_21_287 ();
 sg13g2_fill_2 FILLER_21_355 ();
 sg13g2_fill_2 FILLER_21_366 ();
 sg13g2_fill_2 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_11 ();
 sg13g2_fill_2 FILLER_22_18 ();
 sg13g2_fill_1 FILLER_22_20 ();
 sg13g2_decap_4 FILLER_22_34 ();
 sg13g2_fill_2 FILLER_22_38 ();
 sg13g2_fill_2 FILLER_22_47 ();
 sg13g2_fill_1 FILLER_22_49 ();
 sg13g2_fill_2 FILLER_22_80 ();
 sg13g2_decap_8 FILLER_22_86 ();
 sg13g2_decap_8 FILLER_22_93 ();
 sg13g2_fill_1 FILLER_22_100 ();
 sg13g2_fill_1 FILLER_22_114 ();
 sg13g2_fill_1 FILLER_22_120 ();
 sg13g2_fill_2 FILLER_22_129 ();
 sg13g2_fill_1 FILLER_22_131 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_fill_2 FILLER_22_167 ();
 sg13g2_fill_2 FILLER_22_173 ();
 sg13g2_fill_1 FILLER_22_175 ();
 sg13g2_fill_2 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_188 ();
 sg13g2_decap_4 FILLER_22_210 ();
 sg13g2_fill_2 FILLER_22_214 ();
 sg13g2_fill_2 FILLER_22_225 ();
 sg13g2_fill_1 FILLER_22_227 ();
 sg13g2_fill_1 FILLER_22_292 ();
 sg13g2_fill_2 FILLER_22_337 ();
 sg13g2_fill_1 FILLER_22_339 ();
 sg13g2_fill_1 FILLER_22_367 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_4 FILLER_23_35 ();
 sg13g2_decap_4 FILLER_23_51 ();
 sg13g2_decap_4 FILLER_23_59 ();
 sg13g2_fill_2 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_69 ();
 sg13g2_fill_2 FILLER_23_82 ();
 sg13g2_fill_2 FILLER_23_123 ();
 sg13g2_decap_4 FILLER_23_136 ();
 sg13g2_fill_1 FILLER_23_167 ();
 sg13g2_decap_8 FILLER_23_171 ();
 sg13g2_fill_2 FILLER_23_178 ();
 sg13g2_decap_4 FILLER_23_208 ();
 sg13g2_fill_2 FILLER_23_212 ();
 sg13g2_fill_2 FILLER_23_232 ();
 sg13g2_fill_1 FILLER_23_234 ();
 sg13g2_fill_2 FILLER_23_287 ();
 sg13g2_fill_2 FILLER_23_320 ();
 sg13g2_fill_2 FILLER_23_381 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_13 ();
 sg13g2_decap_8 FILLER_24_26 ();
 sg13g2_decap_4 FILLER_24_33 ();
 sg13g2_decap_8 FILLER_24_54 ();
 sg13g2_fill_1 FILLER_24_96 ();
 sg13g2_decap_8 FILLER_24_137 ();
 sg13g2_decap_4 FILLER_24_144 ();
 sg13g2_fill_1 FILLER_24_178 ();
 sg13g2_fill_2 FILLER_24_187 ();
 sg13g2_fill_1 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_201 ();
 sg13g2_decap_4 FILLER_24_208 ();
 sg13g2_fill_2 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_227 ();
 sg13g2_fill_2 FILLER_24_240 ();
 sg13g2_fill_1 FILLER_24_259 ();
 sg13g2_fill_1 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_307 ();
 sg13g2_fill_2 FILLER_24_326 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_fill_1 FILLER_24_387 ();
 sg13g2_fill_2 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_21 ();
 sg13g2_fill_2 FILLER_25_35 ();
 sg13g2_fill_1 FILLER_25_37 ();
 sg13g2_decap_8 FILLER_25_50 ();
 sg13g2_fill_2 FILLER_25_81 ();
 sg13g2_fill_1 FILLER_25_83 ();
 sg13g2_fill_2 FILLER_25_116 ();
 sg13g2_fill_1 FILLER_25_144 ();
 sg13g2_fill_1 FILLER_25_177 ();
 sg13g2_fill_2 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_199 ();
 sg13g2_decap_8 FILLER_25_204 ();
 sg13g2_fill_2 FILLER_25_287 ();
 sg13g2_fill_1 FILLER_25_289 ();
 sg13g2_fill_2 FILLER_25_352 ();
 sg13g2_fill_1 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_394 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_2 FILLER_26_25 ();
 sg13g2_fill_1 FILLER_26_27 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_fill_2 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_92 ();
 sg13g2_decap_8 FILLER_26_141 ();
 sg13g2_decap_4 FILLER_26_148 ();
 sg13g2_fill_1 FILLER_26_164 ();
 sg13g2_fill_2 FILLER_26_190 ();
 sg13g2_fill_1 FILLER_26_192 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_fill_2 FILLER_26_225 ();
 sg13g2_fill_1 FILLER_26_227 ();
 sg13g2_fill_2 FILLER_26_242 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_fill_1 FILLER_26_378 ();
 sg13g2_fill_2 FILLER_26_388 ();
 sg13g2_fill_2 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_27_13 ();
 sg13g2_decap_4 FILLER_27_48 ();
 sg13g2_fill_1 FILLER_27_52 ();
 sg13g2_fill_2 FILLER_27_65 ();
 sg13g2_fill_1 FILLER_27_75 ();
 sg13g2_fill_1 FILLER_27_84 ();
 sg13g2_fill_1 FILLER_27_100 ();
 sg13g2_fill_1 FILLER_27_123 ();
 sg13g2_decap_8 FILLER_27_150 ();
 sg13g2_fill_2 FILLER_27_157 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_fill_1 FILLER_27_165 ();
 sg13g2_decap_8 FILLER_27_170 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_fill_1 FILLER_27_239 ();
 sg13g2_fill_2 FILLER_27_247 ();
 sg13g2_fill_1 FILLER_27_249 ();
 sg13g2_fill_1 FILLER_27_337 ();
 sg13g2_fill_2 FILLER_27_364 ();
 sg13g2_fill_2 FILLER_27_371 ();
 sg13g2_fill_2 FILLER_27_391 ();
 sg13g2_fill_1 FILLER_27_393 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_27 ();
 sg13g2_fill_2 FILLER_28_41 ();
 sg13g2_fill_2 FILLER_28_69 ();
 sg13g2_fill_1 FILLER_28_85 ();
 sg13g2_fill_1 FILLER_28_96 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_206 ();
 sg13g2_fill_1 FILLER_28_212 ();
 sg13g2_decap_4 FILLER_28_221 ();
 sg13g2_fill_2 FILLER_28_265 ();
 sg13g2_fill_1 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_378 ();
 sg13g2_fill_2 FILLER_28_392 ();
 sg13g2_fill_1 FILLER_28_394 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_17 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_42 ();
 sg13g2_fill_2 FILLER_29_52 ();
 sg13g2_fill_1 FILLER_29_72 ();
 sg13g2_decap_8 FILLER_29_167 ();
 sg13g2_decap_8 FILLER_29_174 ();
 sg13g2_decap_4 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_fill_2 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_29_202 ();
 sg13g2_decap_8 FILLER_29_211 ();
 sg13g2_fill_2 FILLER_29_218 ();
 sg13g2_fill_2 FILLER_29_229 ();
 sg13g2_fill_1 FILLER_29_231 ();
 sg13g2_fill_2 FILLER_29_250 ();
 sg13g2_fill_2 FILLER_29_261 ();
 sg13g2_fill_1 FILLER_29_263 ();
 sg13g2_fill_1 FILLER_29_291 ();
 sg13g2_fill_2 FILLER_29_332 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_4 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_32 ();
 sg13g2_fill_2 FILLER_30_54 ();
 sg13g2_fill_1 FILLER_30_56 ();
 sg13g2_fill_2 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_101 ();
 sg13g2_fill_2 FILLER_30_145 ();
 sg13g2_fill_1 FILLER_30_178 ();
 sg13g2_decap_8 FILLER_30_187 ();
 sg13g2_decap_8 FILLER_30_194 ();
 sg13g2_decap_8 FILLER_30_201 ();
 sg13g2_fill_1 FILLER_30_208 ();
 sg13g2_fill_1 FILLER_30_239 ();
 sg13g2_fill_1 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_18 ();
 sg13g2_fill_1 FILLER_31_20 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_fill_2 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_80 ();
 sg13g2_fill_1 FILLER_31_309 ();
 sg13g2_fill_2 FILLER_31_366 ();
 sg13g2_fill_1 FILLER_31_368 ();
 sg13g2_fill_1 FILLER_31_395 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_39 ();
 sg13g2_fill_1 FILLER_32_46 ();
 sg13g2_fill_1 FILLER_32_76 ();
 sg13g2_fill_2 FILLER_32_99 ();
 sg13g2_fill_1 FILLER_32_176 ();
 sg13g2_decap_4 FILLER_32_220 ();
 sg13g2_fill_1 FILLER_32_238 ();
 sg13g2_fill_2 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_fill_2 FILLER_32_377 ();
 sg13g2_fill_1 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_16 ();
 sg13g2_fill_1 FILLER_33_23 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_107 ();
 sg13g2_fill_1 FILLER_33_129 ();
 sg13g2_decap_4 FILLER_33_190 ();
 sg13g2_fill_1 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_306 ();
 sg13g2_fill_1 FILLER_33_313 ();
 sg13g2_fill_2 FILLER_33_367 ();
 sg13g2_fill_1 FILLER_33_369 ();
 sg13g2_fill_2 FILLER_33_375 ();
 sg13g2_fill_1 FILLER_33_377 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_4 ();
 sg13g2_fill_2 FILLER_34_27 ();
 sg13g2_fill_2 FILLER_34_59 ();
 sg13g2_fill_1 FILLER_34_61 ();
 sg13g2_fill_2 FILLER_34_80 ();
 sg13g2_decap_4 FILLER_34_98 ();
 sg13g2_fill_2 FILLER_34_107 ();
 sg13g2_fill_1 FILLER_34_109 ();
 sg13g2_fill_1 FILLER_34_118 ();
 sg13g2_fill_2 FILLER_34_135 ();
 sg13g2_fill_1 FILLER_34_137 ();
 sg13g2_fill_2 FILLER_34_178 ();
 sg13g2_fill_1 FILLER_34_180 ();
 sg13g2_fill_2 FILLER_34_223 ();
 sg13g2_fill_2 FILLER_34_297 ();
 sg13g2_fill_1 FILLER_34_299 ();
 sg13g2_fill_2 FILLER_34_353 ();
 sg13g2_fill_2 FILLER_34_371 ();
 sg13g2_fill_2 FILLER_34_381 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_42 ();
 sg13g2_fill_1 FILLER_35_47 ();
 sg13g2_decap_8 FILLER_35_69 ();
 sg13g2_decap_8 FILLER_35_76 ();
 sg13g2_fill_2 FILLER_35_87 ();
 sg13g2_fill_1 FILLER_35_89 ();
 sg13g2_fill_1 FILLER_35_111 ();
 sg13g2_fill_2 FILLER_35_126 ();
 sg13g2_fill_1 FILLER_35_128 ();
 sg13g2_fill_2 FILLER_35_150 ();
 sg13g2_fill_1 FILLER_35_152 ();
 sg13g2_fill_2 FILLER_35_169 ();
 sg13g2_fill_1 FILLER_35_171 ();
 sg13g2_fill_1 FILLER_35_180 ();
 sg13g2_decap_4 FILLER_35_230 ();
 sg13g2_fill_2 FILLER_35_257 ();
 sg13g2_fill_1 FILLER_35_305 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_4 ();
 sg13g2_fill_2 FILLER_36_36 ();
 sg13g2_fill_1 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_69 ();
 sg13g2_fill_2 FILLER_36_104 ();
 sg13g2_fill_1 FILLER_36_106 ();
 sg13g2_fill_1 FILLER_36_127 ();
 sg13g2_fill_2 FILLER_36_165 ();
 sg13g2_fill_1 FILLER_36_171 ();
 sg13g2_fill_2 FILLER_36_212 ();
 sg13g2_fill_1 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_395 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_15 ();
 sg13g2_decap_4 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_25 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_51 ();
 sg13g2_fill_1 FILLER_37_68 ();
 sg13g2_fill_1 FILLER_37_87 ();
 sg13g2_fill_2 FILLER_37_107 ();
 sg13g2_fill_1 FILLER_37_109 ();
 sg13g2_fill_1 FILLER_37_124 ();
 sg13g2_fill_2 FILLER_37_141 ();
 sg13g2_decap_8 FILLER_37_151 ();
 sg13g2_fill_2 FILLER_37_158 ();
 sg13g2_fill_2 FILLER_37_192 ();
 sg13g2_fill_2 FILLER_37_205 ();
 sg13g2_fill_1 FILLER_37_207 ();
 sg13g2_fill_1 FILLER_37_264 ();
 sg13g2_fill_2 FILLER_37_327 ();
 sg13g2_fill_2 FILLER_37_338 ();
 sg13g2_fill_1 FILLER_37_365 ();
 sg13g2_fill_2 FILLER_37_375 ();
 sg13g2_fill_1 FILLER_37_377 ();
 sg13g2_fill_2 FILLER_37_383 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_fill_2 FILLER_38_48 ();
 sg13g2_fill_1 FILLER_38_50 ();
 sg13g2_decap_8 FILLER_38_134 ();
 sg13g2_decap_8 FILLER_38_141 ();
 sg13g2_fill_2 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_172 ();
 sg13g2_fill_2 FILLER_38_223 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_276 ();
 sg13g2_fill_1 FILLER_38_340 ();
 sg13g2_fill_2 FILLER_38_345 ();
 sg13g2_fill_1 FILLER_38_347 ();
 sg13g2_fill_2 FILLER_38_364 ();
 sg13g2_fill_2 FILLER_38_380 ();
 sg13g2_fill_1 FILLER_38_382 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_14 ();
 sg13g2_fill_2 FILLER_39_23 ();
 sg13g2_fill_1 FILLER_39_25 ();
 sg13g2_decap_8 FILLER_39_43 ();
 sg13g2_decap_4 FILLER_39_50 ();
 sg13g2_fill_1 FILLER_39_54 ();
 sg13g2_fill_2 FILLER_39_59 ();
 sg13g2_fill_1 FILLER_39_61 ();
 sg13g2_decap_8 FILLER_39_106 ();
 sg13g2_decap_4 FILLER_39_113 ();
 sg13g2_fill_2 FILLER_39_117 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_fill_1 FILLER_39_133 ();
 sg13g2_fill_1 FILLER_39_144 ();
 sg13g2_fill_2 FILLER_39_162 ();
 sg13g2_fill_1 FILLER_39_177 ();
 sg13g2_fill_1 FILLER_39_200 ();
 sg13g2_fill_1 FILLER_39_244 ();
 sg13g2_fill_1 FILLER_39_254 ();
 sg13g2_fill_2 FILLER_39_265 ();
 sg13g2_fill_1 FILLER_39_267 ();
 sg13g2_fill_2 FILLER_39_286 ();
 sg13g2_fill_1 FILLER_39_288 ();
 sg13g2_fill_2 FILLER_39_298 ();
 sg13g2_fill_1 FILLER_39_300 ();
 sg13g2_fill_1 FILLER_39_319 ();
 sg13g2_decap_4 FILLER_39_334 ();
 sg13g2_fill_2 FILLER_39_338 ();
 sg13g2_fill_1 FILLER_39_348 ();
 sg13g2_fill_2 FILLER_39_375 ();
 sg13g2_fill_1 FILLER_39_377 ();
 sg13g2_fill_1 FILLER_39_385 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_40 ();
 sg13g2_fill_1 FILLER_40_60 ();
 sg13g2_fill_2 FILLER_40_88 ();
 sg13g2_fill_1 FILLER_40_90 ();
 sg13g2_decap_4 FILLER_40_103 ();
 sg13g2_fill_1 FILLER_40_107 ();
 sg13g2_decap_8 FILLER_40_114 ();
 sg13g2_decap_4 FILLER_40_133 ();
 sg13g2_fill_2 FILLER_40_141 ();
 sg13g2_fill_1 FILLER_40_143 ();
 sg13g2_fill_1 FILLER_40_179 ();
 sg13g2_decap_4 FILLER_40_219 ();
 sg13g2_fill_1 FILLER_40_266 ();
 sg13g2_fill_2 FILLER_40_303 ();
 sg13g2_fill_1 FILLER_40_305 ();
 sg13g2_fill_2 FILLER_40_315 ();
 sg13g2_fill_2 FILLER_40_322 ();
 sg13g2_decap_4 FILLER_40_332 ();
 sg13g2_fill_2 FILLER_40_336 ();
 sg13g2_fill_2 FILLER_40_343 ();
 sg13g2_fill_1 FILLER_40_345 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_7 ();
 sg13g2_decap_4 FILLER_41_24 ();
 sg13g2_fill_2 FILLER_41_28 ();
 sg13g2_fill_1 FILLER_41_35 ();
 sg13g2_fill_2 FILLER_41_65 ();
 sg13g2_fill_2 FILLER_41_72 ();
 sg13g2_fill_1 FILLER_41_74 ();
 sg13g2_fill_2 FILLER_41_96 ();
 sg13g2_fill_1 FILLER_41_98 ();
 sg13g2_decap_4 FILLER_41_120 ();
 sg13g2_fill_1 FILLER_41_124 ();
 sg13g2_fill_2 FILLER_41_132 ();
 sg13g2_fill_1 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_172 ();
 sg13g2_fill_1 FILLER_41_217 ();
 sg13g2_fill_2 FILLER_41_235 ();
 sg13g2_fill_1 FILLER_41_237 ();
 sg13g2_fill_2 FILLER_41_315 ();
 sg13g2_fill_1 FILLER_41_317 ();
 sg13g2_decap_4 FILLER_41_339 ();
 sg13g2_fill_1 FILLER_41_343 ();
 sg13g2_decap_4 FILLER_41_348 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_29 ();
 sg13g2_fill_2 FILLER_42_44 ();
 sg13g2_fill_1 FILLER_42_46 ();
 sg13g2_fill_2 FILLER_42_56 ();
 sg13g2_fill_1 FILLER_42_58 ();
 sg13g2_fill_2 FILLER_42_99 ();
 sg13g2_fill_2 FILLER_42_112 ();
 sg13g2_fill_1 FILLER_42_122 ();
 sg13g2_decap_4 FILLER_42_169 ();
 sg13g2_fill_1 FILLER_42_177 ();
 sg13g2_fill_1 FILLER_42_234 ();
 sg13g2_fill_1 FILLER_42_279 ();
 sg13g2_fill_2 FILLER_42_334 ();
 sg13g2_decap_4 FILLER_42_352 ();
 sg13g2_fill_2 FILLER_42_376 ();
 sg13g2_fill_2 FILLER_43_34 ();
 sg13g2_fill_1 FILLER_43_51 ();
 sg13g2_fill_2 FILLER_43_62 ();
 sg13g2_fill_1 FILLER_43_64 ();
 sg13g2_fill_1 FILLER_43_84 ();
 sg13g2_fill_1 FILLER_43_94 ();
 sg13g2_fill_2 FILLER_43_120 ();
 sg13g2_fill_1 FILLER_43_122 ();
 sg13g2_decap_4 FILLER_43_197 ();
 sg13g2_fill_1 FILLER_43_224 ();
 sg13g2_fill_1 FILLER_43_230 ();
 sg13g2_fill_1 FILLER_43_244 ();
 sg13g2_fill_2 FILLER_43_280 ();
 sg13g2_decap_4 FILLER_43_297 ();
 sg13g2_fill_1 FILLER_43_306 ();
 sg13g2_fill_2 FILLER_43_324 ();
 sg13g2_fill_1 FILLER_43_326 ();
 sg13g2_fill_1 FILLER_43_344 ();
 sg13g2_decap_4 FILLER_44_26 ();
 sg13g2_fill_2 FILLER_44_35 ();
 sg13g2_fill_2 FILLER_44_65 ();
 sg13g2_fill_2 FILLER_44_106 ();
 sg13g2_decap_8 FILLER_44_128 ();
 sg13g2_decap_8 FILLER_44_135 ();
 sg13g2_decap_8 FILLER_44_142 ();
 sg13g2_fill_2 FILLER_44_149 ();
 sg13g2_fill_1 FILLER_44_151 ();
 sg13g2_fill_2 FILLER_44_162 ();
 sg13g2_fill_1 FILLER_44_164 ();
 sg13g2_fill_2 FILLER_44_216 ();
 sg13g2_decap_8 FILLER_44_274 ();
 sg13g2_fill_2 FILLER_44_285 ();
 sg13g2_decap_8 FILLER_44_297 ();
 sg13g2_decap_4 FILLER_44_316 ();
 sg13g2_fill_1 FILLER_44_320 ();
 sg13g2_fill_1 FILLER_44_324 ();
 sg13g2_decap_4 FILLER_44_333 ();
 sg13g2_fill_1 FILLER_44_337 ();
 sg13g2_fill_1 FILLER_44_370 ();
 sg13g2_fill_2 FILLER_44_397 ();
 sg13g2_fill_1 FILLER_44_399 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_decap_4 FILLER_45_38 ();
 sg13g2_fill_1 FILLER_45_47 ();
 sg13g2_fill_1 FILLER_45_53 ();
 sg13g2_fill_1 FILLER_45_66 ();
 sg13g2_fill_1 FILLER_45_71 ();
 sg13g2_fill_1 FILLER_45_93 ();
 sg13g2_fill_1 FILLER_45_99 ();
 sg13g2_decap_8 FILLER_45_124 ();
 sg13g2_fill_2 FILLER_45_136 ();
 sg13g2_fill_1 FILLER_45_138 ();
 sg13g2_fill_1 FILLER_45_144 ();
 sg13g2_fill_2 FILLER_45_155 ();
 sg13g2_fill_2 FILLER_45_161 ();
 sg13g2_fill_1 FILLER_45_163 ();
 sg13g2_fill_2 FILLER_45_208 ();
 sg13g2_fill_2 FILLER_45_225 ();
 sg13g2_decap_8 FILLER_45_271 ();
 sg13g2_fill_1 FILLER_45_308 ();
 sg13g2_fill_1 FILLER_45_335 ();
 sg13g2_fill_1 FILLER_45_341 ();
 sg13g2_fill_2 FILLER_45_346 ();
 sg13g2_fill_2 FILLER_45_372 ();
 sg13g2_fill_1 FILLER_45_374 ();
 sg13g2_fill_2 FILLER_45_384 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_22 ();
 sg13g2_fill_1 FILLER_46_41 ();
 sg13g2_fill_1 FILLER_46_59 ();
 sg13g2_fill_2 FILLER_46_108 ();
 sg13g2_fill_1 FILLER_46_110 ();
 sg13g2_fill_2 FILLER_46_153 ();
 sg13g2_fill_1 FILLER_46_155 ();
 sg13g2_fill_2 FILLER_46_169 ();
 sg13g2_fill_1 FILLER_46_171 ();
 sg13g2_fill_1 FILLER_46_199 ();
 sg13g2_fill_2 FILLER_46_217 ();
 sg13g2_fill_2 FILLER_46_230 ();
 sg13g2_fill_2 FILLER_46_250 ();
 sg13g2_decap_8 FILLER_46_257 ();
 sg13g2_decap_4 FILLER_46_264 ();
 sg13g2_fill_1 FILLER_46_268 ();
 sg13g2_fill_1 FILLER_46_291 ();
 sg13g2_fill_2 FILLER_46_297 ();
 sg13g2_decap_4 FILLER_46_311 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_fill_2 FILLER_46_343 ();
 sg13g2_fill_2 FILLER_46_363 ();
 sg13g2_fill_1 FILLER_46_373 ();
 sg13g2_fill_2 FILLER_47_35 ();
 sg13g2_fill_1 FILLER_47_37 ();
 sg13g2_fill_2 FILLER_47_43 ();
 sg13g2_fill_1 FILLER_47_55 ();
 sg13g2_fill_2 FILLER_47_76 ();
 sg13g2_fill_2 FILLER_47_113 ();
 sg13g2_fill_1 FILLER_47_115 ();
 sg13g2_fill_2 FILLER_47_133 ();
 sg13g2_fill_1 FILLER_47_140 ();
 sg13g2_decap_4 FILLER_47_180 ();
 sg13g2_fill_1 FILLER_47_210 ();
 sg13g2_fill_2 FILLER_47_215 ();
 sg13g2_fill_1 FILLER_47_225 ();
 sg13g2_decap_4 FILLER_47_239 ();
 sg13g2_fill_2 FILLER_47_243 ();
 sg13g2_fill_1 FILLER_47_253 ();
 sg13g2_fill_1 FILLER_47_271 ();
 sg13g2_fill_1 FILLER_47_278 ();
 sg13g2_fill_2 FILLER_47_311 ();
 sg13g2_fill_1 FILLER_47_313 ();
 sg13g2_fill_2 FILLER_47_348 ();
 sg13g2_fill_2 FILLER_47_367 ();
 sg13g2_fill_1 FILLER_47_369 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_21 ();
 sg13g2_fill_1 FILLER_48_23 ();
 sg13g2_fill_1 FILLER_48_42 ();
 sg13g2_fill_2 FILLER_48_53 ();
 sg13g2_fill_1 FILLER_48_55 ();
 sg13g2_decap_4 FILLER_48_119 ();
 sg13g2_fill_2 FILLER_48_128 ();
 sg13g2_fill_1 FILLER_48_149 ();
 sg13g2_decap_4 FILLER_48_168 ();
 sg13g2_decap_4 FILLER_48_188 ();
 sg13g2_decap_8 FILLER_48_197 ();
 sg13g2_fill_1 FILLER_48_204 ();
 sg13g2_fill_1 FILLER_48_210 ();
 sg13g2_fill_1 FILLER_48_230 ();
 sg13g2_fill_1 FILLER_48_285 ();
 sg13g2_fill_1 FILLER_48_297 ();
 sg13g2_decap_4 FILLER_48_307 ();
 sg13g2_fill_1 FILLER_48_311 ();
 sg13g2_fill_1 FILLER_48_324 ();
 sg13g2_fill_2 FILLER_48_338 ();
 sg13g2_fill_2 FILLER_48_352 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_14 ();
 sg13g2_fill_1 FILLER_49_25 ();
 sg13g2_fill_1 FILLER_49_35 ();
 sg13g2_fill_2 FILLER_49_69 ();
 sg13g2_fill_1 FILLER_49_105 ();
 sg13g2_fill_2 FILLER_49_114 ();
 sg13g2_fill_1 FILLER_49_116 ();
 sg13g2_decap_4 FILLER_49_122 ();
 sg13g2_fill_1 FILLER_49_136 ();
 sg13g2_decap_4 FILLER_49_142 ();
 sg13g2_fill_2 FILLER_49_154 ();
 sg13g2_fill_1 FILLER_49_156 ();
 sg13g2_decap_4 FILLER_49_161 ();
 sg13g2_fill_1 FILLER_49_165 ();
 sg13g2_decap_8 FILLER_49_191 ();
 sg13g2_fill_1 FILLER_49_198 ();
 sg13g2_fill_2 FILLER_49_212 ();
 sg13g2_fill_2 FILLER_49_300 ();
 sg13g2_fill_1 FILLER_49_302 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_fill_2 FILLER_49_361 ();
 sg13g2_fill_1 FILLER_49_363 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_11 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_4 FILLER_50_28 ();
 sg13g2_fill_2 FILLER_50_32 ();
 sg13g2_fill_2 FILLER_50_51 ();
 sg13g2_fill_2 FILLER_50_65 ();
 sg13g2_fill_2 FILLER_50_71 ();
 sg13g2_fill_1 FILLER_50_73 ();
 sg13g2_fill_1 FILLER_50_83 ();
 sg13g2_fill_2 FILLER_50_96 ();
 sg13g2_fill_1 FILLER_50_98 ();
 sg13g2_fill_1 FILLER_50_104 ();
 sg13g2_fill_2 FILLER_50_145 ();
 sg13g2_fill_1 FILLER_50_147 ();
 sg13g2_fill_2 FILLER_50_163 ();
 sg13g2_decap_4 FILLER_50_169 ();
 sg13g2_fill_1 FILLER_50_173 ();
 sg13g2_decap_8 FILLER_50_186 ();
 sg13g2_decap_4 FILLER_50_193 ();
 sg13g2_fill_2 FILLER_50_218 ();
 sg13g2_fill_1 FILLER_50_220 ();
 sg13g2_fill_2 FILLER_50_244 ();
 sg13g2_fill_1 FILLER_50_246 ();
 sg13g2_fill_1 FILLER_50_265 ();
 sg13g2_fill_2 FILLER_50_297 ();
 sg13g2_fill_2 FILLER_50_321 ();
 sg13g2_fill_1 FILLER_50_323 ();
 sg13g2_fill_2 FILLER_50_345 ();
 sg13g2_fill_2 FILLER_50_351 ();
 sg13g2_fill_2 FILLER_50_366 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_55 ();
 sg13g2_fill_2 FILLER_51_81 ();
 sg13g2_fill_1 FILLER_51_104 ();
 sg13g2_fill_1 FILLER_51_123 ();
 sg13g2_fill_2 FILLER_51_141 ();
 sg13g2_fill_2 FILLER_51_159 ();
 sg13g2_fill_1 FILLER_51_161 ();
 sg13g2_decap_8 FILLER_51_175 ();
 sg13g2_decap_4 FILLER_51_182 ();
 sg13g2_fill_1 FILLER_51_186 ();
 sg13g2_decap_8 FILLER_51_192 ();
 sg13g2_decap_8 FILLER_51_199 ();
 sg13g2_fill_2 FILLER_51_236 ();
 sg13g2_fill_1 FILLER_51_238 ();
 sg13g2_fill_2 FILLER_51_250 ();
 sg13g2_fill_1 FILLER_51_252 ();
 sg13g2_fill_1 FILLER_51_258 ();
 sg13g2_fill_2 FILLER_51_356 ();
 sg13g2_fill_1 FILLER_51_371 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_fill_1 FILLER_52_26 ();
 sg13g2_fill_2 FILLER_52_60 ();
 sg13g2_fill_1 FILLER_52_98 ();
 sg13g2_decap_4 FILLER_52_104 ();
 sg13g2_fill_1 FILLER_52_119 ();
 sg13g2_fill_2 FILLER_52_125 ();
 sg13g2_fill_1 FILLER_52_127 ();
 sg13g2_fill_2 FILLER_52_137 ();
 sg13g2_fill_2 FILLER_52_162 ();
 sg13g2_fill_1 FILLER_52_173 ();
 sg13g2_fill_2 FILLER_52_187 ();
 sg13g2_fill_2 FILLER_52_212 ();
 sg13g2_decap_4 FILLER_52_221 ();
 sg13g2_fill_1 FILLER_52_225 ();
 sg13g2_fill_1 FILLER_52_242 ();
 sg13g2_fill_1 FILLER_52_320 ();
 sg13g2_fill_2 FILLER_52_348 ();
 sg13g2_fill_1 FILLER_52_360 ();
 sg13g2_fill_2 FILLER_52_366 ();
 sg13g2_fill_1 FILLER_52_368 ();
 sg13g2_fill_1 FILLER_53_10 ();
 sg13g2_fill_2 FILLER_53_30 ();
 sg13g2_fill_1 FILLER_53_32 ();
 sg13g2_fill_2 FILLER_53_38 ();
 sg13g2_fill_1 FILLER_53_40 ();
 sg13g2_fill_2 FILLER_53_77 ();
 sg13g2_fill_1 FILLER_53_79 ();
 sg13g2_fill_2 FILLER_53_89 ();
 sg13g2_fill_1 FILLER_53_91 ();
 sg13g2_fill_2 FILLER_53_113 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_fill_2 FILLER_53_142 ();
 sg13g2_fill_1 FILLER_53_160 ();
 sg13g2_fill_2 FILLER_53_180 ();
 sg13g2_fill_1 FILLER_53_182 ();
 sg13g2_fill_1 FILLER_53_212 ();
 sg13g2_decap_4 FILLER_53_222 ();
 sg13g2_fill_1 FILLER_53_226 ();
 sg13g2_fill_1 FILLER_53_238 ();
 sg13g2_fill_2 FILLER_53_244 ();
 sg13g2_fill_1 FILLER_53_246 ();
 sg13g2_fill_2 FILLER_53_301 ();
 sg13g2_fill_1 FILLER_53_303 ();
 sg13g2_fill_2 FILLER_53_354 ();
 sg13g2_fill_1 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_6 ();
 sg13g2_fill_1 FILLER_54_27 ();
 sg13g2_fill_1 FILLER_54_51 ();
 sg13g2_decap_4 FILLER_54_101 ();
 sg13g2_fill_1 FILLER_54_105 ();
 sg13g2_fill_1 FILLER_54_125 ();
 sg13g2_fill_2 FILLER_54_145 ();
 sg13g2_fill_2 FILLER_54_258 ();
 sg13g2_fill_1 FILLER_54_260 ();
 sg13g2_fill_2 FILLER_54_306 ();
 sg13g2_fill_2 FILLER_54_320 ();
 sg13g2_fill_2 FILLER_54_339 ();
 sg13g2_fill_1 FILLER_54_360 ();
 sg13g2_fill_1 FILLER_54_399 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_4 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_32 ();
 sg13g2_fill_2 FILLER_55_60 ();
 sg13g2_fill_1 FILLER_55_70 ();
 sg13g2_fill_1 FILLER_55_105 ();
 sg13g2_fill_1 FILLER_55_125 ();
 sg13g2_fill_2 FILLER_55_175 ();
 sg13g2_fill_1 FILLER_55_177 ();
 sg13g2_fill_1 FILLER_55_188 ();
 sg13g2_fill_2 FILLER_55_210 ();
 sg13g2_fill_1 FILLER_55_212 ();
 sg13g2_fill_2 FILLER_55_218 ();
 sg13g2_fill_2 FILLER_55_296 ();
 sg13g2_fill_1 FILLER_55_315 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_36 ();
 sg13g2_fill_2 FILLER_56_43 ();
 sg13g2_fill_1 FILLER_56_100 ();
 sg13g2_fill_1 FILLER_56_135 ();
 sg13g2_fill_1 FILLER_56_144 ();
 sg13g2_fill_2 FILLER_56_159 ();
 sg13g2_fill_1 FILLER_56_161 ();
 sg13g2_fill_1 FILLER_56_168 ();
 sg13g2_fill_2 FILLER_56_174 ();
 sg13g2_fill_2 FILLER_56_181 ();
 sg13g2_decap_8 FILLER_56_193 ();
 sg13g2_decap_8 FILLER_56_200 ();
 sg13g2_decap_8 FILLER_56_207 ();
 sg13g2_decap_8 FILLER_56_214 ();
 sg13g2_decap_8 FILLER_56_221 ();
 sg13g2_decap_4 FILLER_56_228 ();
 sg13g2_fill_2 FILLER_56_232 ();
 sg13g2_fill_2 FILLER_56_241 ();
 sg13g2_fill_2 FILLER_56_252 ();
 sg13g2_fill_1 FILLER_56_254 ();
 sg13g2_fill_2 FILLER_56_260 ();
 sg13g2_fill_1 FILLER_56_262 ();
 sg13g2_fill_1 FILLER_56_382 ();
 sg13g2_fill_2 FILLER_57_35 ();
 sg13g2_fill_2 FILLER_57_47 ();
 sg13g2_fill_2 FILLER_57_87 ();
 sg13g2_decap_4 FILLER_57_97 ();
 sg13g2_fill_1 FILLER_57_101 ();
 sg13g2_fill_1 FILLER_57_110 ();
 sg13g2_fill_1 FILLER_57_124 ();
 sg13g2_fill_2 FILLER_57_133 ();
 sg13g2_fill_1 FILLER_57_155 ();
 sg13g2_fill_1 FILLER_57_161 ();
 sg13g2_fill_1 FILLER_57_166 ();
 sg13g2_fill_1 FILLER_57_183 ();
 sg13g2_decap_4 FILLER_57_194 ();
 sg13g2_fill_2 FILLER_57_198 ();
 sg13g2_fill_1 FILLER_57_242 ();
 sg13g2_fill_2 FILLER_57_282 ();
 sg13g2_fill_1 FILLER_57_284 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_4 FILLER_58_7 ();
 sg13g2_decap_4 FILLER_58_15 ();
 sg13g2_fill_2 FILLER_58_45 ();
 sg13g2_decap_8 FILLER_58_57 ();
 sg13g2_decap_8 FILLER_58_64 ();
 sg13g2_fill_2 FILLER_58_71 ();
 sg13g2_decap_8 FILLER_58_90 ();
 sg13g2_decap_8 FILLER_58_113 ();
 sg13g2_fill_2 FILLER_58_120 ();
 sg13g2_fill_2 FILLER_58_132 ();
 sg13g2_fill_1 FILLER_58_134 ();
 sg13g2_fill_2 FILLER_58_159 ();
 sg13g2_fill_1 FILLER_58_161 ();
 sg13g2_fill_2 FILLER_58_191 ();
 sg13g2_fill_1 FILLER_58_193 ();
 sg13g2_fill_2 FILLER_58_219 ();
 sg13g2_fill_2 FILLER_58_241 ();
 sg13g2_fill_2 FILLER_58_257 ();
 sg13g2_fill_2 FILLER_58_321 ();
 sg13g2_fill_2 FILLER_58_327 ();
 sg13g2_fill_2 FILLER_58_341 ();
 sg13g2_fill_1 FILLER_58_343 ();
 sg13g2_fill_1 FILLER_58_399 ();
 sg13g2_fill_2 FILLER_59_26 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_4 FILLER_59_70 ();
 sg13g2_fill_2 FILLER_59_74 ();
 sg13g2_fill_2 FILLER_59_85 ();
 sg13g2_fill_1 FILLER_59_87 ();
 sg13g2_fill_1 FILLER_59_107 ();
 sg13g2_fill_2 FILLER_59_127 ();
 sg13g2_fill_1 FILLER_59_129 ();
 sg13g2_fill_2 FILLER_59_154 ();
 sg13g2_fill_1 FILLER_59_156 ();
 sg13g2_fill_2 FILLER_59_194 ();
 sg13g2_decap_4 FILLER_59_216 ();
 sg13g2_fill_2 FILLER_59_220 ();
 sg13g2_fill_2 FILLER_59_265 ();
 sg13g2_fill_1 FILLER_59_267 ();
 sg13g2_fill_2 FILLER_59_294 ();
 sg13g2_fill_2 FILLER_59_322 ();
 sg13g2_fill_2 FILLER_59_380 ();
 sg13g2_fill_1 FILLER_59_382 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_7 ();
 sg13g2_decap_4 FILLER_60_23 ();
 sg13g2_fill_1 FILLER_60_27 ();
 sg13g2_fill_2 FILLER_60_38 ();
 sg13g2_fill_1 FILLER_60_40 ();
 sg13g2_decap_4 FILLER_60_46 ();
 sg13g2_fill_2 FILLER_60_50 ();
 sg13g2_fill_1 FILLER_60_58 ();
 sg13g2_decap_8 FILLER_60_85 ();
 sg13g2_decap_8 FILLER_60_92 ();
 sg13g2_fill_1 FILLER_60_99 ();
 sg13g2_fill_2 FILLER_60_124 ();
 sg13g2_fill_1 FILLER_60_147 ();
 sg13g2_decap_8 FILLER_60_171 ();
 sg13g2_fill_2 FILLER_60_178 ();
 sg13g2_fill_1 FILLER_60_180 ();
 sg13g2_decap_8 FILLER_60_189 ();
 sg13g2_decap_4 FILLER_60_208 ();
 sg13g2_fill_1 FILLER_60_256 ();
 sg13g2_fill_2 FILLER_60_264 ();
 sg13g2_fill_1 FILLER_60_266 ();
 sg13g2_fill_2 FILLER_60_276 ();
 sg13g2_fill_1 FILLER_60_287 ();
 sg13g2_fill_1 FILLER_60_322 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_4 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_4 ();
 sg13g2_fill_1 FILLER_61_20 ();
 sg13g2_decap_4 FILLER_61_32 ();
 sg13g2_fill_2 FILLER_61_41 ();
 sg13g2_decap_4 FILLER_61_92 ();
 sg13g2_fill_1 FILLER_61_96 ();
 sg13g2_fill_2 FILLER_61_106 ();
 sg13g2_fill_1 FILLER_61_132 ();
 sg13g2_fill_1 FILLER_61_151 ();
 sg13g2_fill_2 FILLER_61_168 ();
 sg13g2_fill_1 FILLER_61_170 ();
 sg13g2_decap_4 FILLER_61_176 ();
 sg13g2_fill_1 FILLER_61_180 ();
 sg13g2_decap_8 FILLER_61_186 ();
 sg13g2_decap_8 FILLER_61_193 ();
 sg13g2_decap_8 FILLER_61_200 ();
 sg13g2_fill_1 FILLER_61_207 ();
 sg13g2_fill_1 FILLER_61_226 ();
 sg13g2_fill_1 FILLER_61_235 ();
 sg13g2_fill_1 FILLER_61_245 ();
 sg13g2_fill_2 FILLER_61_325 ();
 sg13g2_fill_1 FILLER_61_337 ();
 sg13g2_fill_1 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_31 ();
 sg13g2_fill_2 FILLER_62_37 ();
 sg13g2_fill_2 FILLER_62_54 ();
 sg13g2_fill_2 FILLER_62_61 ();
 sg13g2_fill_2 FILLER_62_102 ();
 sg13g2_fill_2 FILLER_62_113 ();
 sg13g2_fill_1 FILLER_62_138 ();
 sg13g2_fill_2 FILLER_62_143 ();
 sg13g2_decap_4 FILLER_62_161 ();
 sg13g2_decap_4 FILLER_62_192 ();
 sg13g2_fill_2 FILLER_62_250 ();
 sg13g2_fill_1 FILLER_62_252 ();
 sg13g2_fill_2 FILLER_62_265 ();
 sg13g2_fill_2 FILLER_62_360 ();
 sg13g2_fill_1 FILLER_62_362 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_fill_2 FILLER_63_26 ();
 sg13g2_fill_1 FILLER_63_65 ();
 sg13g2_decap_4 FILLER_63_92 ();
 sg13g2_fill_1 FILLER_63_96 ();
 sg13g2_decap_4 FILLER_63_109 ();
 sg13g2_fill_2 FILLER_63_117 ();
 sg13g2_fill_1 FILLER_63_119 ();
 sg13g2_decap_4 FILLER_63_135 ();
 sg13g2_fill_1 FILLER_63_139 ();
 sg13g2_decap_4 FILLER_63_144 ();
 sg13g2_fill_1 FILLER_63_180 ();
 sg13g2_fill_1 FILLER_63_185 ();
 sg13g2_fill_2 FILLER_63_234 ();
 sg13g2_fill_2 FILLER_63_242 ();
 sg13g2_fill_1 FILLER_63_244 ();
 sg13g2_fill_2 FILLER_63_262 ();
 sg13g2_fill_1 FILLER_63_324 ();
 sg13g2_decap_4 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_36 ();
 sg13g2_decap_4 FILLER_64_43 ();
 sg13g2_fill_1 FILLER_64_57 ();
 sg13g2_fill_1 FILLER_64_66 ();
 sg13g2_fill_2 FILLER_64_71 ();
 sg13g2_fill_1 FILLER_64_73 ();
 sg13g2_decap_4 FILLER_64_143 ();
 sg13g2_decap_4 FILLER_64_151 ();
 sg13g2_fill_2 FILLER_64_155 ();
 sg13g2_fill_1 FILLER_64_225 ();
 sg13g2_fill_1 FILLER_64_294 ();
 sg13g2_fill_1 FILLER_64_345 ();
 sg13g2_fill_2 FILLER_64_372 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_22 ();
 sg13g2_fill_2 FILLER_65_41 ();
 sg13g2_fill_1 FILLER_65_43 ();
 sg13g2_decap_8 FILLER_65_83 ();
 sg13g2_decap_8 FILLER_65_90 ();
 sg13g2_decap_4 FILLER_65_109 ();
 sg13g2_fill_1 FILLER_65_142 ();
 sg13g2_fill_1 FILLER_65_165 ();
 sg13g2_decap_8 FILLER_65_179 ();
 sg13g2_fill_1 FILLER_65_203 ();
 sg13g2_fill_1 FILLER_65_250 ();
 sg13g2_fill_1 FILLER_65_270 ();
 sg13g2_fill_1 FILLER_65_375 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_22 ();
 sg13g2_fill_1 FILLER_66_48 ();
 sg13g2_decap_4 FILLER_66_59 ();
 sg13g2_fill_1 FILLER_66_63 ();
 sg13g2_fill_2 FILLER_66_69 ();
 sg13g2_decap_8 FILLER_66_79 ();
 sg13g2_decap_8 FILLER_66_86 ();
 sg13g2_fill_2 FILLER_66_93 ();
 sg13g2_fill_1 FILLER_66_95 ();
 sg13g2_fill_2 FILLER_66_104 ();
 sg13g2_decap_4 FILLER_66_157 ();
 sg13g2_fill_1 FILLER_66_161 ();
 sg13g2_fill_1 FILLER_66_170 ();
 sg13g2_fill_2 FILLER_66_175 ();
 sg13g2_fill_1 FILLER_66_177 ();
 sg13g2_fill_1 FILLER_66_233 ();
 sg13g2_fill_2 FILLER_66_250 ();
 sg13g2_fill_1 FILLER_66_297 ();
 sg13g2_fill_2 FILLER_66_329 ();
 sg13g2_fill_1 FILLER_66_349 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_fill_1 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_18 ();
 sg13g2_fill_2 FILLER_67_51 ();
 sg13g2_fill_1 FILLER_67_94 ();
 sg13g2_fill_2 FILLER_67_124 ();
 sg13g2_fill_2 FILLER_67_136 ();
 sg13g2_fill_2 FILLER_67_172 ();
 sg13g2_fill_1 FILLER_67_181 ();
 sg13g2_fill_1 FILLER_67_223 ();
 sg13g2_fill_1 FILLER_67_274 ();
 sg13g2_fill_1 FILLER_67_288 ();
 sg13g2_fill_2 FILLER_67_324 ();
 sg13g2_fill_2 FILLER_67_330 ();
 sg13g2_fill_1 FILLER_67_350 ();
 sg13g2_fill_2 FILLER_67_363 ();
 sg13g2_fill_1 FILLER_67_365 ();
 sg13g2_fill_2 FILLER_67_372 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_fill_2 FILLER_68_33 ();
 sg13g2_fill_2 FILLER_68_43 ();
 sg13g2_decap_8 FILLER_68_57 ();
 sg13g2_decap_8 FILLER_68_85 ();
 sg13g2_fill_2 FILLER_68_117 ();
 sg13g2_fill_1 FILLER_68_119 ();
 sg13g2_decap_4 FILLER_68_141 ();
 sg13g2_fill_2 FILLER_68_145 ();
 sg13g2_decap_8 FILLER_68_151 ();
 sg13g2_fill_1 FILLER_68_158 ();
 sg13g2_fill_1 FILLER_68_225 ();
 sg13g2_fill_2 FILLER_68_248 ();
 sg13g2_fill_2 FILLER_68_351 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_29 ();
 sg13g2_fill_2 FILLER_69_48 ();
 sg13g2_fill_2 FILLER_69_70 ();
 sg13g2_fill_2 FILLER_69_90 ();
 sg13g2_fill_2 FILLER_69_105 ();
 sg13g2_fill_1 FILLER_69_107 ();
 sg13g2_fill_2 FILLER_69_129 ();
 sg13g2_decap_8 FILLER_69_136 ();
 sg13g2_decap_8 FILLER_69_155 ();
 sg13g2_decap_4 FILLER_69_162 ();
 sg13g2_fill_2 FILLER_69_211 ();
 sg13g2_fill_1 FILLER_69_243 ();
 sg13g2_fill_2 FILLER_69_292 ();
 sg13g2_fill_1 FILLER_69_294 ();
 sg13g2_fill_2 FILLER_69_313 ();
 sg13g2_fill_1 FILLER_69_315 ();
 sg13g2_fill_2 FILLER_69_356 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_22 ();
 sg13g2_fill_2 FILLER_70_29 ();
 sg13g2_fill_1 FILLER_70_31 ();
 sg13g2_fill_2 FILLER_70_47 ();
 sg13g2_fill_1 FILLER_70_49 ();
 sg13g2_fill_1 FILLER_70_69 ();
 sg13g2_fill_2 FILLER_70_118 ();
 sg13g2_fill_2 FILLER_70_125 ();
 sg13g2_decap_8 FILLER_70_139 ();
 sg13g2_fill_1 FILLER_70_146 ();
 sg13g2_decap_8 FILLER_70_165 ();
 sg13g2_fill_2 FILLER_70_172 ();
 sg13g2_fill_2 FILLER_70_241 ();
 sg13g2_fill_1 FILLER_70_252 ();
 sg13g2_fill_1 FILLER_70_279 ();
 sg13g2_fill_1 FILLER_70_295 ();
 sg13g2_fill_1 FILLER_70_307 ();
 sg13g2_fill_2 FILLER_70_318 ();
 sg13g2_fill_1 FILLER_70_320 ();
 sg13g2_fill_2 FILLER_70_338 ();
 sg13g2_fill_1 FILLER_70_340 ();
 sg13g2_fill_2 FILLER_70_393 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_decap_4 FILLER_71_20 ();
 sg13g2_decap_4 FILLER_71_29 ();
 sg13g2_fill_2 FILLER_71_33 ();
 sg13g2_decap_4 FILLER_71_40 ();
 sg13g2_fill_1 FILLER_71_44 ();
 sg13g2_fill_2 FILLER_71_49 ();
 sg13g2_fill_1 FILLER_71_51 ();
 sg13g2_fill_1 FILLER_71_60 ();
 sg13g2_fill_2 FILLER_71_70 ();
 sg13g2_fill_1 FILLER_71_72 ();
 sg13g2_fill_2 FILLER_71_79 ();
 sg13g2_decap_8 FILLER_71_93 ();
 sg13g2_decap_4 FILLER_71_114 ();
 sg13g2_fill_2 FILLER_71_123 ();
 sg13g2_decap_4 FILLER_71_135 ();
 sg13g2_fill_2 FILLER_71_139 ();
 sg13g2_decap_4 FILLER_71_174 ();
 sg13g2_fill_2 FILLER_71_178 ();
 sg13g2_fill_1 FILLER_71_275 ();
 sg13g2_fill_2 FILLER_71_333 ();
 sg13g2_fill_2 FILLER_71_361 ();
 sg13g2_fill_2 FILLER_71_398 ();
 sg13g2_fill_1 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_46 ();
 sg13g2_decap_4 FILLER_72_53 ();
 sg13g2_fill_2 FILLER_72_57 ();
 sg13g2_decap_8 FILLER_72_92 ();
 sg13g2_fill_1 FILLER_72_99 ();
 sg13g2_fill_2 FILLER_72_136 ();
 sg13g2_fill_1 FILLER_72_138 ();
 sg13g2_decap_4 FILLER_72_144 ();
 sg13g2_fill_1 FILLER_72_148 ();
 sg13g2_decap_4 FILLER_72_170 ();
 sg13g2_fill_1 FILLER_72_174 ();
 sg13g2_fill_1 FILLER_72_237 ();
 sg13g2_fill_2 FILLER_72_345 ();
 sg13g2_fill_2 FILLER_73_22 ();
 sg13g2_fill_2 FILLER_73_32 ();
 sg13g2_fill_1 FILLER_73_34 ();
 sg13g2_decap_8 FILLER_73_39 ();
 sg13g2_fill_2 FILLER_73_59 ();
 sg13g2_fill_1 FILLER_73_61 ();
 sg13g2_decap_8 FILLER_73_74 ();
 sg13g2_fill_2 FILLER_73_81 ();
 sg13g2_fill_2 FILLER_73_104 ();
 sg13g2_fill_1 FILLER_73_146 ();
 sg13g2_fill_2 FILLER_73_163 ();
 sg13g2_fill_1 FILLER_73_165 ();
 sg13g2_fill_1 FILLER_73_171 ();
 sg13g2_fill_1 FILLER_73_199 ();
 sg13g2_fill_2 FILLER_73_217 ();
 sg13g2_fill_1 FILLER_73_219 ();
 sg13g2_fill_1 FILLER_73_264 ();
 sg13g2_fill_2 FILLER_73_278 ();
 sg13g2_decap_4 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_4 ();
 sg13g2_fill_2 FILLER_74_14 ();
 sg13g2_fill_1 FILLER_74_16 ();
 sg13g2_fill_2 FILLER_74_38 ();
 sg13g2_decap_8 FILLER_74_74 ();
 sg13g2_decap_4 FILLER_74_81 ();
 sg13g2_fill_2 FILLER_74_173 ();
 sg13g2_fill_1 FILLER_74_175 ();
 sg13g2_fill_2 FILLER_74_192 ();
 sg13g2_fill_1 FILLER_74_209 ();
 sg13g2_fill_1 FILLER_74_250 ();
 sg13g2_fill_2 FILLER_74_267 ();
 sg13g2_fill_2 FILLER_74_292 ();
 sg13g2_fill_2 FILLER_74_324 ();
 sg13g2_fill_2 FILLER_74_358 ();
 sg13g2_fill_1 FILLER_74_366 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_4 FILLER_75_29 ();
 sg13g2_decap_4 FILLER_75_61 ();
 sg13g2_fill_2 FILLER_75_65 ();
 sg13g2_fill_1 FILLER_75_88 ();
 sg13g2_decap_8 FILLER_75_110 ();
 sg13g2_decap_8 FILLER_75_117 ();
 sg13g2_fill_2 FILLER_75_124 ();
 sg13g2_fill_1 FILLER_75_126 ();
 sg13g2_decap_4 FILLER_75_132 ();
 sg13g2_fill_1 FILLER_75_136 ();
 sg13g2_fill_2 FILLER_75_147 ();
 sg13g2_fill_1 FILLER_75_149 ();
 sg13g2_fill_2 FILLER_75_163 ();
 sg13g2_fill_2 FILLER_75_245 ();
 sg13g2_fill_1 FILLER_75_247 ();
 sg13g2_fill_2 FILLER_75_253 ();
 sg13g2_fill_1 FILLER_75_255 ();
 sg13g2_fill_1 FILLER_75_266 ();
 sg13g2_fill_2 FILLER_75_276 ();
 sg13g2_fill_1 FILLER_75_292 ();
 sg13g2_fill_1 FILLER_75_317 ();
 sg13g2_fill_1 FILLER_75_382 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_7 ();
 sg13g2_fill_1 FILLER_76_12 ();
 sg13g2_fill_2 FILLER_76_23 ();
 sg13g2_fill_1 FILLER_76_25 ();
 sg13g2_fill_1 FILLER_76_38 ();
 sg13g2_decap_4 FILLER_76_44 ();
 sg13g2_fill_1 FILLER_76_58 ();
 sg13g2_fill_1 FILLER_76_97 ();
 sg13g2_fill_2 FILLER_76_103 ();
 sg13g2_decap_8 FILLER_76_115 ();
 sg13g2_decap_8 FILLER_76_122 ();
 sg13g2_fill_2 FILLER_76_129 ();
 sg13g2_fill_1 FILLER_76_131 ();
 sg13g2_fill_2 FILLER_76_152 ();
 sg13g2_fill_1 FILLER_76_154 ();
 sg13g2_fill_1 FILLER_76_173 ();
 sg13g2_fill_2 FILLER_76_239 ();
 sg13g2_fill_1 FILLER_76_269 ();
 sg13g2_fill_2 FILLER_76_306 ();
 sg13g2_fill_2 FILLER_76_318 ();
 sg13g2_fill_2 FILLER_76_333 ();
 sg13g2_fill_1 FILLER_76_379 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_fill_1 FILLER_77_36 ();
 sg13g2_fill_2 FILLER_77_61 ();
 sg13g2_fill_2 FILLER_77_84 ();
 sg13g2_fill_1 FILLER_77_107 ();
 sg13g2_fill_1 FILLER_77_113 ();
 sg13g2_fill_2 FILLER_77_122 ();
 sg13g2_fill_2 FILLER_77_173 ();
 sg13g2_fill_1 FILLER_77_199 ();
 sg13g2_fill_2 FILLER_77_205 ();
 sg13g2_fill_1 FILLER_77_207 ();
 sg13g2_fill_1 FILLER_77_272 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_7 ();
 sg13g2_fill_1 FILLER_78_9 ();
 sg13g2_fill_2 FILLER_78_44 ();
 sg13g2_fill_1 FILLER_78_46 ();
 sg13g2_fill_2 FILLER_78_150 ();
 sg13g2_fill_2 FILLER_78_171 ();
 sg13g2_fill_2 FILLER_78_237 ();
 sg13g2_fill_1 FILLER_78_239 ();
 sg13g2_fill_2 FILLER_78_274 ();
 sg13g2_fill_1 FILLER_78_276 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_fill_1 FILLER_79_34 ();
 sg13g2_fill_1 FILLER_79_44 ();
 sg13g2_decap_4 FILLER_79_73 ();
 sg13g2_fill_2 FILLER_79_80 ();
 sg13g2_fill_1 FILLER_79_82 ();
 sg13g2_fill_2 FILLER_79_157 ();
 sg13g2_fill_1 FILLER_79_159 ();
 sg13g2_fill_2 FILLER_79_184 ();
 sg13g2_fill_2 FILLER_79_212 ();
 sg13g2_fill_2 FILLER_79_218 ();
 sg13g2_fill_1 FILLER_79_220 ();
 sg13g2_fill_1 FILLER_79_252 ();
 sg13g2_fill_2 FILLER_79_265 ();
 sg13g2_fill_1 FILLER_79_267 ();
 sg13g2_fill_2 FILLER_79_317 ();
 sg13g2_fill_1 FILLER_79_364 ();
 sg13g2_fill_2 FILLER_79_391 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_4 FILLER_80_28 ();
 sg13g2_fill_1 FILLER_80_32 ();
 sg13g2_decap_8 FILLER_80_37 ();
 sg13g2_decap_8 FILLER_80_44 ();
 sg13g2_fill_1 FILLER_80_51 ();
 sg13g2_fill_1 FILLER_80_55 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_fill_1 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_fill_1 FILLER_80_111 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_fill_1 FILLER_80_123 ();
 sg13g2_fill_2 FILLER_80_140 ();
 sg13g2_fill_2 FILLER_80_187 ();
 sg13g2_fill_2 FILLER_80_201 ();
 sg13g2_fill_2 FILLER_80_229 ();
 sg13g2_fill_1 FILLER_80_231 ();
 sg13g2_fill_1 FILLER_80_236 ();
 sg13g2_fill_1 FILLER_80_265 ();
 sg13g2_fill_2 FILLER_80_274 ();
 sg13g2_fill_2 FILLER_80_288 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net246;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
endmodule

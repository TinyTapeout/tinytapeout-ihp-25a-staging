module tt_um_pdm_pitch_filter_arghunter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire net27;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire \u_top_module.addr[0] ;
 wire \u_top_module.addr[1] ;
 wire \u_top_module.addr[2] ;
 wire \u_top_module.addr[3] ;
 wire \u_top_module.addr[4] ;
 wire \u_top_module.addr[5] ;
 wire \u_top_module.addr[6] ;
 wire \u_top_module.addr[7] ;
 wire \u_top_module.capture_reg[0] ;
 wire \u_top_module.capture_reg[1] ;
 wire \u_top_module.capture_reg[2] ;
 wire \u_top_module.capture_reg[3] ;
 wire \u_top_module.capture_reg[4] ;
 wire \u_top_module.capture_reg[5] ;
 wire \u_top_module.capture_reg[6] ;
 wire \u_top_module.capture_reg[7] ;
 wire \u_top_module.dec_clk ;
 wire \u_top_module.dec_data ;
 wire \u_top_module.decimation_ratio[0] ;
 wire \u_top_module.decimation_ratio[1] ;
 wire \u_top_module.decimation_ratio[2] ;
 wire \u_top_module.decimation_ratio[3] ;
 wire \u_top_module.decimation_ratio[4] ;
 wire \u_top_module.decimation_ratio[5] ;
 wire \u_top_module.decimation_ratio[6] ;
 wire \u_top_module.decimation_ratio[7] ;
 wire \u_top_module.filter_length[0] ;
 wire \u_top_module.filter_length[1] ;
 wire \u_top_module.filter_length[2] ;
 wire \u_top_module.filter_length[3] ;
 wire \u_top_module.filter_length[4] ;
 wire \u_top_module.filter_length[5] ;
 wire \u_top_module.filter_length[6] ;
 wire \u_top_module.filter_length[7] ;
 wire \u_top_module.mem_out[0] ;
 wire \u_top_module.mem_out[1] ;
 wire \u_top_module.mem_out[2] ;
 wire \u_top_module.mem_out[3] ;
 wire \u_top_module.mem_out[4] ;
 wire \u_top_module.mem_out[5] ;
 wire \u_top_module.mem_out[6] ;
 wire \u_top_module.mem_out[7] ;
 wire \u_top_module.out ;
 wire \u_top_module.u_decimator.counter[0] ;
 wire \u_top_module.u_decimator.counter[1] ;
 wire \u_top_module.u_decimator.counter[2] ;
 wire \u_top_module.u_decimator.counter[3] ;
 wire \u_top_module.u_decimator.counter[4] ;
 wire \u_top_module.u_decimator.counter[5] ;
 wire \u_top_module.u_decimator.counter[6] ;
 wire \u_top_module.u_decimator.counter[7] ;
 wire \u_top_module.u_filter.shift_reg[0] ;
 wire \u_top_module.u_filter.shift_reg[100] ;
 wire \u_top_module.u_filter.shift_reg[101] ;
 wire \u_top_module.u_filter.shift_reg[102] ;
 wire \u_top_module.u_filter.shift_reg[103] ;
 wire \u_top_module.u_filter.shift_reg[104] ;
 wire \u_top_module.u_filter.shift_reg[105] ;
 wire \u_top_module.u_filter.shift_reg[106] ;
 wire \u_top_module.u_filter.shift_reg[107] ;
 wire \u_top_module.u_filter.shift_reg[108] ;
 wire \u_top_module.u_filter.shift_reg[109] ;
 wire \u_top_module.u_filter.shift_reg[10] ;
 wire \u_top_module.u_filter.shift_reg[110] ;
 wire \u_top_module.u_filter.shift_reg[111] ;
 wire \u_top_module.u_filter.shift_reg[112] ;
 wire \u_top_module.u_filter.shift_reg[113] ;
 wire \u_top_module.u_filter.shift_reg[114] ;
 wire \u_top_module.u_filter.shift_reg[115] ;
 wire \u_top_module.u_filter.shift_reg[116] ;
 wire \u_top_module.u_filter.shift_reg[117] ;
 wire \u_top_module.u_filter.shift_reg[118] ;
 wire \u_top_module.u_filter.shift_reg[119] ;
 wire \u_top_module.u_filter.shift_reg[11] ;
 wire \u_top_module.u_filter.shift_reg[120] ;
 wire \u_top_module.u_filter.shift_reg[121] ;
 wire \u_top_module.u_filter.shift_reg[122] ;
 wire \u_top_module.u_filter.shift_reg[123] ;
 wire \u_top_module.u_filter.shift_reg[124] ;
 wire \u_top_module.u_filter.shift_reg[125] ;
 wire \u_top_module.u_filter.shift_reg[126] ;
 wire \u_top_module.u_filter.shift_reg[127] ;
 wire \u_top_module.u_filter.shift_reg[128] ;
 wire \u_top_module.u_filter.shift_reg[129] ;
 wire \u_top_module.u_filter.shift_reg[12] ;
 wire \u_top_module.u_filter.shift_reg[130] ;
 wire \u_top_module.u_filter.shift_reg[131] ;
 wire \u_top_module.u_filter.shift_reg[132] ;
 wire \u_top_module.u_filter.shift_reg[133] ;
 wire \u_top_module.u_filter.shift_reg[134] ;
 wire \u_top_module.u_filter.shift_reg[135] ;
 wire \u_top_module.u_filter.shift_reg[136] ;
 wire \u_top_module.u_filter.shift_reg[137] ;
 wire \u_top_module.u_filter.shift_reg[138] ;
 wire \u_top_module.u_filter.shift_reg[139] ;
 wire \u_top_module.u_filter.shift_reg[13] ;
 wire \u_top_module.u_filter.shift_reg[140] ;
 wire \u_top_module.u_filter.shift_reg[141] ;
 wire \u_top_module.u_filter.shift_reg[142] ;
 wire \u_top_module.u_filter.shift_reg[143] ;
 wire \u_top_module.u_filter.shift_reg[144] ;
 wire \u_top_module.u_filter.shift_reg[145] ;
 wire \u_top_module.u_filter.shift_reg[146] ;
 wire \u_top_module.u_filter.shift_reg[147] ;
 wire \u_top_module.u_filter.shift_reg[148] ;
 wire \u_top_module.u_filter.shift_reg[149] ;
 wire \u_top_module.u_filter.shift_reg[14] ;
 wire \u_top_module.u_filter.shift_reg[150] ;
 wire \u_top_module.u_filter.shift_reg[151] ;
 wire \u_top_module.u_filter.shift_reg[152] ;
 wire \u_top_module.u_filter.shift_reg[153] ;
 wire \u_top_module.u_filter.shift_reg[154] ;
 wire \u_top_module.u_filter.shift_reg[155] ;
 wire \u_top_module.u_filter.shift_reg[156] ;
 wire \u_top_module.u_filter.shift_reg[157] ;
 wire \u_top_module.u_filter.shift_reg[158] ;
 wire \u_top_module.u_filter.shift_reg[159] ;
 wire \u_top_module.u_filter.shift_reg[15] ;
 wire \u_top_module.u_filter.shift_reg[160] ;
 wire \u_top_module.u_filter.shift_reg[161] ;
 wire \u_top_module.u_filter.shift_reg[162] ;
 wire \u_top_module.u_filter.shift_reg[163] ;
 wire \u_top_module.u_filter.shift_reg[164] ;
 wire \u_top_module.u_filter.shift_reg[165] ;
 wire \u_top_module.u_filter.shift_reg[166] ;
 wire \u_top_module.u_filter.shift_reg[167] ;
 wire \u_top_module.u_filter.shift_reg[168] ;
 wire \u_top_module.u_filter.shift_reg[169] ;
 wire \u_top_module.u_filter.shift_reg[16] ;
 wire \u_top_module.u_filter.shift_reg[170] ;
 wire \u_top_module.u_filter.shift_reg[171] ;
 wire \u_top_module.u_filter.shift_reg[172] ;
 wire \u_top_module.u_filter.shift_reg[173] ;
 wire \u_top_module.u_filter.shift_reg[174] ;
 wire \u_top_module.u_filter.shift_reg[175] ;
 wire \u_top_module.u_filter.shift_reg[176] ;
 wire \u_top_module.u_filter.shift_reg[177] ;
 wire \u_top_module.u_filter.shift_reg[178] ;
 wire \u_top_module.u_filter.shift_reg[179] ;
 wire \u_top_module.u_filter.shift_reg[17] ;
 wire \u_top_module.u_filter.shift_reg[180] ;
 wire \u_top_module.u_filter.shift_reg[181] ;
 wire \u_top_module.u_filter.shift_reg[182] ;
 wire \u_top_module.u_filter.shift_reg[183] ;
 wire \u_top_module.u_filter.shift_reg[184] ;
 wire \u_top_module.u_filter.shift_reg[185] ;
 wire \u_top_module.u_filter.shift_reg[186] ;
 wire \u_top_module.u_filter.shift_reg[187] ;
 wire \u_top_module.u_filter.shift_reg[188] ;
 wire \u_top_module.u_filter.shift_reg[189] ;
 wire \u_top_module.u_filter.shift_reg[18] ;
 wire \u_top_module.u_filter.shift_reg[190] ;
 wire \u_top_module.u_filter.shift_reg[191] ;
 wire \u_top_module.u_filter.shift_reg[192] ;
 wire \u_top_module.u_filter.shift_reg[193] ;
 wire \u_top_module.u_filter.shift_reg[194] ;
 wire \u_top_module.u_filter.shift_reg[195] ;
 wire \u_top_module.u_filter.shift_reg[196] ;
 wire \u_top_module.u_filter.shift_reg[197] ;
 wire \u_top_module.u_filter.shift_reg[198] ;
 wire \u_top_module.u_filter.shift_reg[199] ;
 wire \u_top_module.u_filter.shift_reg[19] ;
 wire \u_top_module.u_filter.shift_reg[1] ;
 wire \u_top_module.u_filter.shift_reg[200] ;
 wire \u_top_module.u_filter.shift_reg[201] ;
 wire \u_top_module.u_filter.shift_reg[202] ;
 wire \u_top_module.u_filter.shift_reg[203] ;
 wire \u_top_module.u_filter.shift_reg[204] ;
 wire \u_top_module.u_filter.shift_reg[205] ;
 wire \u_top_module.u_filter.shift_reg[206] ;
 wire \u_top_module.u_filter.shift_reg[207] ;
 wire \u_top_module.u_filter.shift_reg[208] ;
 wire \u_top_module.u_filter.shift_reg[209] ;
 wire \u_top_module.u_filter.shift_reg[20] ;
 wire \u_top_module.u_filter.shift_reg[210] ;
 wire \u_top_module.u_filter.shift_reg[211] ;
 wire \u_top_module.u_filter.shift_reg[212] ;
 wire \u_top_module.u_filter.shift_reg[213] ;
 wire \u_top_module.u_filter.shift_reg[214] ;
 wire \u_top_module.u_filter.shift_reg[215] ;
 wire \u_top_module.u_filter.shift_reg[216] ;
 wire \u_top_module.u_filter.shift_reg[217] ;
 wire \u_top_module.u_filter.shift_reg[218] ;
 wire \u_top_module.u_filter.shift_reg[219] ;
 wire \u_top_module.u_filter.shift_reg[21] ;
 wire \u_top_module.u_filter.shift_reg[220] ;
 wire \u_top_module.u_filter.shift_reg[221] ;
 wire \u_top_module.u_filter.shift_reg[222] ;
 wire \u_top_module.u_filter.shift_reg[223] ;
 wire \u_top_module.u_filter.shift_reg[224] ;
 wire \u_top_module.u_filter.shift_reg[225] ;
 wire \u_top_module.u_filter.shift_reg[226] ;
 wire \u_top_module.u_filter.shift_reg[227] ;
 wire \u_top_module.u_filter.shift_reg[228] ;
 wire \u_top_module.u_filter.shift_reg[229] ;
 wire \u_top_module.u_filter.shift_reg[22] ;
 wire \u_top_module.u_filter.shift_reg[230] ;
 wire \u_top_module.u_filter.shift_reg[231] ;
 wire \u_top_module.u_filter.shift_reg[232] ;
 wire \u_top_module.u_filter.shift_reg[233] ;
 wire \u_top_module.u_filter.shift_reg[234] ;
 wire \u_top_module.u_filter.shift_reg[235] ;
 wire \u_top_module.u_filter.shift_reg[236] ;
 wire \u_top_module.u_filter.shift_reg[237] ;
 wire \u_top_module.u_filter.shift_reg[238] ;
 wire \u_top_module.u_filter.shift_reg[239] ;
 wire \u_top_module.u_filter.shift_reg[23] ;
 wire \u_top_module.u_filter.shift_reg[240] ;
 wire \u_top_module.u_filter.shift_reg[241] ;
 wire \u_top_module.u_filter.shift_reg[242] ;
 wire \u_top_module.u_filter.shift_reg[243] ;
 wire \u_top_module.u_filter.shift_reg[244] ;
 wire \u_top_module.u_filter.shift_reg[245] ;
 wire \u_top_module.u_filter.shift_reg[246] ;
 wire \u_top_module.u_filter.shift_reg[247] ;
 wire \u_top_module.u_filter.shift_reg[248] ;
 wire \u_top_module.u_filter.shift_reg[249] ;
 wire \u_top_module.u_filter.shift_reg[24] ;
 wire \u_top_module.u_filter.shift_reg[250] ;
 wire \u_top_module.u_filter.shift_reg[251] ;
 wire \u_top_module.u_filter.shift_reg[252] ;
 wire \u_top_module.u_filter.shift_reg[253] ;
 wire \u_top_module.u_filter.shift_reg[254] ;
 wire \u_top_module.u_filter.shift_reg[25] ;
 wire \u_top_module.u_filter.shift_reg[26] ;
 wire \u_top_module.u_filter.shift_reg[27] ;
 wire \u_top_module.u_filter.shift_reg[28] ;
 wire \u_top_module.u_filter.shift_reg[29] ;
 wire \u_top_module.u_filter.shift_reg[2] ;
 wire \u_top_module.u_filter.shift_reg[30] ;
 wire \u_top_module.u_filter.shift_reg[31] ;
 wire \u_top_module.u_filter.shift_reg[32] ;
 wire \u_top_module.u_filter.shift_reg[33] ;
 wire \u_top_module.u_filter.shift_reg[34] ;
 wire \u_top_module.u_filter.shift_reg[35] ;
 wire \u_top_module.u_filter.shift_reg[36] ;
 wire \u_top_module.u_filter.shift_reg[37] ;
 wire \u_top_module.u_filter.shift_reg[38] ;
 wire \u_top_module.u_filter.shift_reg[39] ;
 wire \u_top_module.u_filter.shift_reg[3] ;
 wire \u_top_module.u_filter.shift_reg[40] ;
 wire \u_top_module.u_filter.shift_reg[41] ;
 wire \u_top_module.u_filter.shift_reg[42] ;
 wire \u_top_module.u_filter.shift_reg[43] ;
 wire \u_top_module.u_filter.shift_reg[44] ;
 wire \u_top_module.u_filter.shift_reg[45] ;
 wire \u_top_module.u_filter.shift_reg[46] ;
 wire \u_top_module.u_filter.shift_reg[47] ;
 wire \u_top_module.u_filter.shift_reg[48] ;
 wire \u_top_module.u_filter.shift_reg[49] ;
 wire \u_top_module.u_filter.shift_reg[4] ;
 wire \u_top_module.u_filter.shift_reg[50] ;
 wire \u_top_module.u_filter.shift_reg[51] ;
 wire \u_top_module.u_filter.shift_reg[52] ;
 wire \u_top_module.u_filter.shift_reg[53] ;
 wire \u_top_module.u_filter.shift_reg[54] ;
 wire \u_top_module.u_filter.shift_reg[55] ;
 wire \u_top_module.u_filter.shift_reg[56] ;
 wire \u_top_module.u_filter.shift_reg[57] ;
 wire \u_top_module.u_filter.shift_reg[58] ;
 wire \u_top_module.u_filter.shift_reg[59] ;
 wire \u_top_module.u_filter.shift_reg[5] ;
 wire \u_top_module.u_filter.shift_reg[60] ;
 wire \u_top_module.u_filter.shift_reg[61] ;
 wire \u_top_module.u_filter.shift_reg[62] ;
 wire \u_top_module.u_filter.shift_reg[63] ;
 wire \u_top_module.u_filter.shift_reg[64] ;
 wire \u_top_module.u_filter.shift_reg[65] ;
 wire \u_top_module.u_filter.shift_reg[66] ;
 wire \u_top_module.u_filter.shift_reg[67] ;
 wire \u_top_module.u_filter.shift_reg[68] ;
 wire \u_top_module.u_filter.shift_reg[69] ;
 wire \u_top_module.u_filter.shift_reg[6] ;
 wire \u_top_module.u_filter.shift_reg[70] ;
 wire \u_top_module.u_filter.shift_reg[71] ;
 wire \u_top_module.u_filter.shift_reg[72] ;
 wire \u_top_module.u_filter.shift_reg[73] ;
 wire \u_top_module.u_filter.shift_reg[74] ;
 wire \u_top_module.u_filter.shift_reg[75] ;
 wire \u_top_module.u_filter.shift_reg[76] ;
 wire \u_top_module.u_filter.shift_reg[77] ;
 wire \u_top_module.u_filter.shift_reg[78] ;
 wire \u_top_module.u_filter.shift_reg[79] ;
 wire \u_top_module.u_filter.shift_reg[7] ;
 wire \u_top_module.u_filter.shift_reg[80] ;
 wire \u_top_module.u_filter.shift_reg[81] ;
 wire \u_top_module.u_filter.shift_reg[82] ;
 wire \u_top_module.u_filter.shift_reg[83] ;
 wire \u_top_module.u_filter.shift_reg[84] ;
 wire \u_top_module.u_filter.shift_reg[85] ;
 wire \u_top_module.u_filter.shift_reg[86] ;
 wire \u_top_module.u_filter.shift_reg[87] ;
 wire \u_top_module.u_filter.shift_reg[88] ;
 wire \u_top_module.u_filter.shift_reg[89] ;
 wire \u_top_module.u_filter.shift_reg[8] ;
 wire \u_top_module.u_filter.shift_reg[90] ;
 wire \u_top_module.u_filter.shift_reg[91] ;
 wire \u_top_module.u_filter.shift_reg[92] ;
 wire \u_top_module.u_filter.shift_reg[93] ;
 wire \u_top_module.u_filter.shift_reg[94] ;
 wire \u_top_module.u_filter.shift_reg[95] ;
 wire \u_top_module.u_filter.shift_reg[96] ;
 wire \u_top_module.u_filter.shift_reg[97] ;
 wire \u_top_module.u_filter.shift_reg[98] ;
 wire \u_top_module.u_filter.shift_reg[99] ;
 wire \u_top_module.u_filter.shift_reg[9] ;
 wire \u_top_module.u_i2s_bus.counter[0] ;
 wire \u_top_module.u_i2s_bus.counter[1] ;
 wire \u_top_module.u_i2s_bus.counter[2] ;
 wire \u_top_module.u_i2s_bus.counter[3] ;
 wire \u_top_module.u_i2s_bus.counter[4] ;
 wire \u_top_module.u_i2s_bus.counter[5] ;
 wire \u_top_module.u_i2s_bus.counter[6] ;
 wire \u_top_module.u_i2s_bus.counter[7] ;
 wire \u_top_module.u_i2s_bus.dec_clk ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.prev_lr_clk ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[9].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.u_mux_shift.sum_res ;
 wire \u_top_module.u_memory.memory[0][0] ;
 wire \u_top_module.u_memory.memory[0][1] ;
 wire \u_top_module.u_memory.memory[0][2] ;
 wire \u_top_module.u_memory.memory[0][3] ;
 wire \u_top_module.u_memory.memory[0][4] ;
 wire \u_top_module.u_memory.memory[0][5] ;
 wire \u_top_module.u_memory.memory[0][6] ;
 wire \u_top_module.u_memory.memory[0][7] ;
 wire \u_top_module.u_memory.memory[1][0] ;
 wire \u_top_module.u_memory.memory[1][1] ;
 wire \u_top_module.u_memory.memory[1][2] ;
 wire \u_top_module.u_memory.memory[1][3] ;
 wire \u_top_module.u_memory.memory[1][4] ;
 wire \u_top_module.u_memory.memory[1][5] ;
 wire \u_top_module.u_memory.memory[1][6] ;
 wire \u_top_module.u_memory.memory[1][7] ;
 wire \u_top_module.u_memory.memory[2][0] ;
 wire \u_top_module.u_memory.memory[2][1] ;
 wire \u_top_module.u_memory.memory[2][2] ;
 wire \u_top_module.u_memory.memory[2][3] ;
 wire \u_top_module.u_memory.memory[2][4] ;
 wire \u_top_module.u_memory.memory[2][5] ;
 wire \u_top_module.u_memory.memory[2][6] ;
 wire \u_top_module.u_memory.memory[2][7] ;
 wire \u_top_module.u_memory.memory[3][0] ;
 wire \u_top_module.u_memory.memory[3][1] ;
 wire \u_top_module.u_memory.memory[3][2] ;
 wire \u_top_module.u_memory.memory[3][3] ;
 wire \u_top_module.u_memory.memory[3][4] ;
 wire \u_top_module.u_memory.memory[3][5] ;
 wire \u_top_module.u_memory.memory[3][6] ;
 wire \u_top_module.u_memory.memory[3][7] ;
 wire \u_top_module.u_memory.memory[4][0] ;
 wire \u_top_module.u_memory.memory[4][1] ;
 wire \u_top_module.u_memory.memory[4][2] ;
 wire \u_top_module.u_memory.memory[4][3] ;
 wire \u_top_module.u_memory.memory[4][4] ;
 wire \u_top_module.u_memory.memory[4][5] ;
 wire \u_top_module.u_memory.memory[4][6] ;
 wire \u_top_module.u_memory.memory[4][7] ;
 wire \u_top_module.u_memory.memory[5][0] ;
 wire \u_top_module.u_memory.memory[5][1] ;
 wire \u_top_module.u_memory.memory[5][2] ;
 wire \u_top_module.u_memory.memory[5][3] ;
 wire \u_top_module.u_memory.memory[5][4] ;
 wire \u_top_module.u_memory.memory[5][5] ;
 wire \u_top_module.u_memory.memory[5][6] ;
 wire \u_top_module.u_memory.memory[5][7] ;
 wire \u_top_module.u_memory.memory[6][0] ;
 wire \u_top_module.u_memory.memory[6][1] ;
 wire \u_top_module.u_memory.memory[6][2] ;
 wire \u_top_module.u_memory.memory[6][3] ;
 wire \u_top_module.u_memory.memory[6][4] ;
 wire \u_top_module.u_memory.memory[6][5] ;
 wire \u_top_module.u_memory.memory[6][6] ;
 wire \u_top_module.u_memory.memory[6][7] ;
 wire \u_top_module.u_memory.memory[7][0] ;
 wire \u_top_module.u_memory.memory[7][1] ;
 wire \u_top_module.u_memory.memory[7][2] ;
 wire \u_top_module.u_memory.memory[7][3] ;
 wire \u_top_module.u_memory.memory[7][4] ;
 wire \u_top_module.u_memory.memory[7][5] ;
 wire \u_top_module.u_memory.memory[7][6] ;
 wire \u_top_module.u_memory.memory[7][7] ;
 wire \u_top_module.u_spi_port.cs_n_prev ;
 wire \u_top_module.u_spi_port.shift_reg[0] ;
 wire \u_top_module.u_spi_port.shift_reg[10] ;
 wire \u_top_module.u_spi_port.shift_reg[11] ;
 wire \u_top_module.u_spi_port.shift_reg[12] ;
 wire \u_top_module.u_spi_port.shift_reg[13] ;
 wire \u_top_module.u_spi_port.shift_reg[14] ;
 wire \u_top_module.u_spi_port.shift_reg[15] ;
 wire \u_top_module.u_spi_port.shift_reg[1] ;
 wire \u_top_module.u_spi_port.shift_reg[2] ;
 wire \u_top_module.u_spi_port.shift_reg[3] ;
 wire \u_top_module.u_spi_port.shift_reg[4] ;
 wire \u_top_module.u_spi_port.shift_reg[5] ;
 wire \u_top_module.u_spi_port.shift_reg[6] ;
 wire \u_top_module.u_spi_port.shift_reg[7] ;
 wire \u_top_module.u_spi_port.shift_reg[8] ;
 wire \u_top_module.u_spi_port.shift_reg[9] ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1;
 wire net2;
 wire net3;
 wire net4;

 sg13g2_inv_1 _1311_ (.Y(_0030_),
    .A(net2));
 sg13g2_inv_1 _1312_ (.Y(_0546_),
    .A(\u_top_module.addr[1] ));
 sg13g2_inv_1 _1313_ (.Y(_0031_),
    .A(net980));
 sg13g2_inv_1 _1314_ (.Y(_0547_),
    .A(\u_top_module.u_decimator.counter[0] ));
 sg13g2_inv_1 _1315_ (.Y(_0548_),
    .A(\u_top_module.u_decimator.counter[1] ));
 sg13g2_inv_1 _1316_ (.Y(_0549_),
    .A(\u_top_module.decimation_ratio[1] ));
 sg13g2_inv_1 _1317_ (.Y(_0550_),
    .A(\u_top_module.decimation_ratio[3] ));
 sg13g2_inv_1 _1318_ (.Y(_0551_),
    .A(\u_top_module.decimation_ratio[2] ));
 sg13g2_inv_1 _1319_ (.Y(_0552_),
    .A(\u_top_module.decimation_ratio[6] ));
 sg13g2_inv_1 _1320_ (.Y(_0553_),
    .A(\u_top_module.u_decimator.counter[5] ));
 sg13g2_inv_1 _1321_ (.Y(_0554_),
    .A(\u_top_module.u_decimator.counter[4] ));
 sg13g2_inv_1 _1322_ (.Y(_0555_),
    .A(\u_top_module.decimation_ratio[4] ));
 sg13g2_inv_1 _1323_ (.Y(_0556_),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ));
 sg13g2_inv_1 _1324_ (.Y(_0557_),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ));
 sg13g2_inv_2 _1325_ (.Y(_0558_),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ));
 sg13g2_inv_1 _1326_ (.Y(_0559_),
    .A(\u_top_module.filter_length[4] ));
 sg13g2_inv_1 _1327_ (.Y(_0560_),
    .A(net834));
 sg13g2_inv_1 _1328_ (.Y(_0561_),
    .A(net865));
 sg13g2_inv_1 _1329_ (.Y(_0562_),
    .A(\u_top_module.u_filter.shift_reg[42] ));
 sg13g2_inv_1 _1330_ (.Y(_0563_),
    .A(\u_top_module.u_filter.shift_reg[151] ));
 sg13g2_inv_1 _1331_ (.Y(_0564_),
    .A(\u_top_module.u_filter.shift_reg[215] ));
 sg13g2_inv_1 _1332_ (.Y(_0565_),
    .A(\u_top_module.u_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_and2_1 _1333_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.out ),
    .B(net1018),
    .X(_0170_));
 sg13g2_nor2_1 _1334_ (.A(\u_top_module.addr[3] ),
    .B(\u_top_module.addr[2] ),
    .Y(_0566_));
 sg13g2_nor4_2 _1335_ (.A(\u_top_module.addr[5] ),
    .B(\u_top_module.addr[4] ),
    .C(\u_top_module.addr[7] ),
    .Y(_0567_),
    .D(\u_top_module.addr[6] ));
 sg13g2_nand2_1 _1336_ (.Y(_0568_),
    .A(\u_top_module.addr[0] ),
    .B(_0546_));
 sg13g2_nand4_1 _1337_ (.B(_0546_),
    .C(_0566_),
    .A(\u_top_module.addr[0] ),
    .Y(_0001_),
    .D(_0567_));
 sg13g2_nor2_1 _1338_ (.A(\u_top_module.addr[0] ),
    .B(\u_top_module.addr[1] ),
    .Y(_0569_));
 sg13g2_nand3_1 _1339_ (.B(_0567_),
    .C(_0569_),
    .A(_0566_),
    .Y(_0000_));
 sg13g2_nor2_1 _1340_ (.A(\u_top_module.addr[2] ),
    .B(_0568_),
    .Y(_0570_));
 sg13g2_nor2_1 _1341_ (.A(_0027_),
    .B(_0568_),
    .Y(_0571_));
 sg13g2_nand2_1 _1342_ (.Y(_0572_),
    .A(\u_top_module.addr[0] ),
    .B(\u_top_module.addr[1] ));
 sg13g2_nor2_1 _1343_ (.A(\u_top_module.addr[2] ),
    .B(_0572_),
    .Y(_0573_));
 sg13g2_nor2_1 _1344_ (.A(_0027_),
    .B(_0572_),
    .Y(_0574_));
 sg13g2_nand2b_1 _1345_ (.Y(_0575_),
    .B(\u_top_module.addr[1] ),
    .A_N(\u_top_module.addr[0] ));
 sg13g2_nor2_1 _1346_ (.A(_0027_),
    .B(_0575_),
    .Y(_0576_));
 sg13g2_nor3_1 _1347_ (.A(\u_top_module.addr[2] ),
    .B(\u_top_module.addr[0] ),
    .C(\u_top_module.addr[1] ),
    .Y(_0577_));
 sg13g2_nand2b_2 _1348_ (.Y(_0578_),
    .B(_0569_),
    .A_N(\u_top_module.addr[2] ));
 sg13g2_a21oi_1 _1349_ (.A1(\u_top_module.u_memory.memory[6][0] ),
    .A2(net878),
    .Y(_0579_),
    .B1(_0577_));
 sg13g2_nor3_1 _1350_ (.A(\u_top_module.addr[0] ),
    .B(\u_top_module.addr[1] ),
    .C(_0027_),
    .Y(_0580_));
 sg13g2_nor2_1 _1351_ (.A(\u_top_module.addr[2] ),
    .B(_0575_),
    .Y(_0581_));
 sg13g2_a22oi_1 _1352_ (.Y(_0582_),
    .B1(net882),
    .B2(\u_top_module.u_memory.memory[3][0] ),
    .A2(net872),
    .A1(\u_top_module.u_memory.memory[5][0] ));
 sg13g2_a22oi_1 _1353_ (.Y(_0583_),
    .B1(net876),
    .B2(\u_top_module.u_memory.memory[2][0] ),
    .A2(net880),
    .A1(\u_top_module.u_memory.memory[7][0] ));
 sg13g2_a22oi_1 _1354_ (.Y(_0584_),
    .B1(net894),
    .B2(\u_top_module.u_memory.memory[4][0] ),
    .A2(net874),
    .A1(\u_top_module.u_memory.memory[1][0] ));
 sg13g2_nand4_1 _1355_ (.B(_0582_),
    .C(_0583_),
    .A(_0579_),
    .Y(_0585_),
    .D(_0584_));
 sg13g2_o21ai_1 _1356_ (.B1(_0585_),
    .Y(_0586_),
    .A1(\u_top_module.u_memory.memory[0][0] ),
    .A2(_0578_));
 sg13g2_inv_1 _1357_ (.Y(_0197_),
    .A(_0586_));
 sg13g2_a21oi_1 _1358_ (.A1(\u_top_module.u_memory.memory[6][1] ),
    .A2(net877),
    .Y(_0587_),
    .B1(net895));
 sg13g2_a22oi_1 _1359_ (.Y(_0588_),
    .B1(net875),
    .B2(\u_top_module.u_memory.memory[2][1] ),
    .A2(net881),
    .A1(\u_top_module.u_memory.memory[3][1] ));
 sg13g2_a22oi_1 _1360_ (.Y(_0589_),
    .B1(net893),
    .B2(\u_top_module.u_memory.memory[4][1] ),
    .A2(net871),
    .A1(\u_top_module.u_memory.memory[5][1] ));
 sg13g2_a22oi_1 _1361_ (.Y(_0590_),
    .B1(net879),
    .B2(\u_top_module.u_memory.memory[7][1] ),
    .A2(net873),
    .A1(\u_top_module.u_memory.memory[1][1] ));
 sg13g2_nand4_1 _1362_ (.B(_0588_),
    .C(_0589_),
    .A(_0587_),
    .Y(_0591_),
    .D(_0590_));
 sg13g2_o21ai_1 _1363_ (.B1(_0591_),
    .Y(_0592_),
    .A1(\u_top_module.u_memory.memory[0][1] ),
    .A2(_0578_));
 sg13g2_inv_1 _1364_ (.Y(_0198_),
    .A(_0592_));
 sg13g2_a21oi_1 _1365_ (.A1(\u_top_module.u_memory.memory[4][2] ),
    .A2(net894),
    .Y(_0593_),
    .B1(net896));
 sg13g2_a22oi_1 _1366_ (.Y(_0594_),
    .B1(net878),
    .B2(\u_top_module.u_memory.memory[6][2] ),
    .A2(net874),
    .A1(\u_top_module.u_memory.memory[1][2] ));
 sg13g2_a22oi_1 _1367_ (.Y(_0595_),
    .B1(net876),
    .B2(\u_top_module.u_memory.memory[2][2] ),
    .A2(net882),
    .A1(\u_top_module.u_memory.memory[3][2] ));
 sg13g2_a22oi_1 _1368_ (.Y(_0596_),
    .B1(net880),
    .B2(\u_top_module.u_memory.memory[7][2] ),
    .A2(net872),
    .A1(\u_top_module.u_memory.memory[5][2] ));
 sg13g2_nand4_1 _1369_ (.B(_0594_),
    .C(_0595_),
    .A(_0593_),
    .Y(_0597_),
    .D(_0596_));
 sg13g2_o21ai_1 _1370_ (.B1(_0597_),
    .Y(_0598_),
    .A1(\u_top_module.u_memory.memory[0][2] ),
    .A2(_0578_));
 sg13g2_inv_1 _1371_ (.Y(_0199_),
    .A(_0598_));
 sg13g2_a22oi_1 _1372_ (.Y(_0599_),
    .B1(net877),
    .B2(\u_top_module.u_memory.memory[6][3] ),
    .A2(net881),
    .A1(\u_top_module.u_memory.memory[3][3] ));
 sg13g2_a22oi_1 _1373_ (.Y(_0600_),
    .B1(net875),
    .B2(\u_top_module.u_memory.memory[2][3] ),
    .A2(net893),
    .A1(\u_top_module.u_memory.memory[4][3] ));
 sg13g2_a22oi_1 _1374_ (.Y(_0601_),
    .B1(net879),
    .B2(\u_top_module.u_memory.memory[7][3] ),
    .A2(net871),
    .A1(\u_top_module.u_memory.memory[5][3] ));
 sg13g2_a21oi_1 _1375_ (.A1(\u_top_module.u_memory.memory[1][3] ),
    .A2(net873),
    .Y(_0602_),
    .B1(net896));
 sg13g2_nand4_1 _1376_ (.B(_0600_),
    .C(_0601_),
    .A(_0599_),
    .Y(_0603_),
    .D(_0602_));
 sg13g2_o21ai_1 _1377_ (.B1(_0603_),
    .Y(_0604_),
    .A1(\u_top_module.u_memory.memory[0][3] ),
    .A2(_0578_));
 sg13g2_inv_1 _1378_ (.Y(_0200_),
    .A(_0604_));
 sg13g2_a22oi_1 _1379_ (.Y(_0605_),
    .B1(net893),
    .B2(\u_top_module.u_memory.memory[4][4] ),
    .A2(net879),
    .A1(\u_top_module.u_memory.memory[7][4] ));
 sg13g2_a22oi_1 _1380_ (.Y(_0606_),
    .B1(net881),
    .B2(\u_top_module.u_memory.memory[3][4] ),
    .A2(net873),
    .A1(\u_top_module.u_memory.memory[1][4] ));
 sg13g2_a22oi_1 _1381_ (.Y(_0607_),
    .B1(net877),
    .B2(\u_top_module.u_memory.memory[6][4] ),
    .A2(net871),
    .A1(\u_top_module.u_memory.memory[5][4] ));
 sg13g2_a21oi_1 _1382_ (.A1(\u_top_module.u_memory.memory[2][4] ),
    .A2(net875),
    .Y(_0608_),
    .B1(net895));
 sg13g2_nand4_1 _1383_ (.B(_0606_),
    .C(_0607_),
    .A(_0605_),
    .Y(_0609_),
    .D(_0608_));
 sg13g2_o21ai_1 _1384_ (.B1(_0609_),
    .Y(_0610_),
    .A1(\u_top_module.u_memory.memory[0][4] ),
    .A2(_0578_));
 sg13g2_inv_1 _1385_ (.Y(_0201_),
    .A(_0610_));
 sg13g2_a22oi_1 _1386_ (.Y(_0611_),
    .B1(net876),
    .B2(\u_top_module.u_memory.memory[2][5] ),
    .A2(net882),
    .A1(\u_top_module.u_memory.memory[3][5] ));
 sg13g2_a22oi_1 _1387_ (.Y(_0612_),
    .B1(net894),
    .B2(\u_top_module.u_memory.memory[4][5] ),
    .A2(net872),
    .A1(\u_top_module.u_memory.memory[5][5] ));
 sg13g2_a22oi_1 _1388_ (.Y(_0613_),
    .B1(net880),
    .B2(\u_top_module.u_memory.memory[7][5] ),
    .A2(net874),
    .A1(\u_top_module.u_memory.memory[1][5] ));
 sg13g2_a21oi_1 _1389_ (.A1(\u_top_module.u_memory.memory[6][5] ),
    .A2(net878),
    .Y(_0614_),
    .B1(net896));
 sg13g2_nand4_1 _1390_ (.B(_0612_),
    .C(_0613_),
    .A(_0611_),
    .Y(_0615_),
    .D(_0614_));
 sg13g2_o21ai_1 _1391_ (.B1(_0615_),
    .Y(_0616_),
    .A1(\u_top_module.u_memory.memory[0][5] ),
    .A2(_0578_));
 sg13g2_inv_1 _1392_ (.Y(_0202_),
    .A(_0616_));
 sg13g2_a22oi_1 _1393_ (.Y(_0617_),
    .B1(net880),
    .B2(\u_top_module.u_memory.memory[7][6] ),
    .A2(net872),
    .A1(\u_top_module.u_memory.memory[5][6] ));
 sg13g2_a22oi_1 _1394_ (.Y(_0618_),
    .B1(net882),
    .B2(\u_top_module.u_memory.memory[3][6] ),
    .A2(net874),
    .A1(\u_top_module.u_memory.memory[1][6] ));
 sg13g2_a22oi_1 _1395_ (.Y(_0619_),
    .B1(net876),
    .B2(\u_top_module.u_memory.memory[2][6] ),
    .A2(net878),
    .A1(\u_top_module.u_memory.memory[6][6] ));
 sg13g2_a21oi_1 _1396_ (.A1(\u_top_module.u_memory.memory[4][6] ),
    .A2(net894),
    .Y(_0620_),
    .B1(net895));
 sg13g2_nand4_1 _1397_ (.B(_0618_),
    .C(_0619_),
    .A(_0617_),
    .Y(_0621_),
    .D(_0620_));
 sg13g2_o21ai_1 _1398_ (.B1(_0621_),
    .Y(_0622_),
    .A1(\u_top_module.u_memory.memory[0][6] ),
    .A2(_0578_));
 sg13g2_inv_1 _1399_ (.Y(_0203_),
    .A(_0622_));
 sg13g2_a22oi_1 _1400_ (.Y(_0623_),
    .B1(net893),
    .B2(\u_top_module.u_memory.memory[4][7] ),
    .A2(net877),
    .A1(\u_top_module.u_memory.memory[6][7] ));
 sg13g2_a22oi_1 _1401_ (.Y(_0624_),
    .B1(net875),
    .B2(\u_top_module.u_memory.memory[2][7] ),
    .A2(net881),
    .A1(\u_top_module.u_memory.memory[3][7] ));
 sg13g2_a22oi_1 _1402_ (.Y(_0625_),
    .B1(net879),
    .B2(\u_top_module.u_memory.memory[7][7] ),
    .A2(net871),
    .A1(\u_top_module.u_memory.memory[5][7] ));
 sg13g2_a21oi_1 _1403_ (.A1(\u_top_module.u_memory.memory[1][7] ),
    .A2(net873),
    .Y(_0626_),
    .B1(net895));
 sg13g2_nand4_1 _1404_ (.B(_0624_),
    .C(_0625_),
    .A(_0623_),
    .Y(_0627_),
    .D(_0626_));
 sg13g2_o21ai_1 _1405_ (.B1(_0627_),
    .Y(_0628_),
    .A1(\u_top_module.u_memory.memory[0][7] ),
    .A2(_0578_));
 sg13g2_inv_1 _1406_ (.Y(_0204_),
    .A(_0628_));
 sg13g2_or2_2 _1407_ (.X(_0629_),
    .B(\u_top_module.u_i2s_bus.counter[6] ),
    .A(\u_top_module.u_i2s_bus.counter[7] ));
 sg13g2_nor2_1 _1408_ (.A(\u_top_module.u_i2s_bus.counter[0] ),
    .B(_0629_),
    .Y(_0011_));
 sg13g2_nor2_1 _1409_ (.A(\u_top_module.u_i2s_bus.counter[0] ),
    .B(\u_top_module.u_i2s_bus.counter[1] ),
    .Y(_0630_));
 sg13g2_and2_1 _1410_ (.A(\u_top_module.u_i2s_bus.counter[0] ),
    .B(\u_top_module.u_i2s_bus.counter[1] ),
    .X(_0631_));
 sg13g2_nor3_1 _1411_ (.A(_0629_),
    .B(_0630_),
    .C(_0631_),
    .Y(_0012_));
 sg13g2_nor2_1 _1412_ (.A(\u_top_module.u_i2s_bus.counter[2] ),
    .B(_0631_),
    .Y(_0632_));
 sg13g2_and2_1 _1413_ (.A(\u_top_module.u_i2s_bus.counter[2] ),
    .B(_0631_),
    .X(_0633_));
 sg13g2_nor3_1 _1414_ (.A(_0629_),
    .B(_0632_),
    .C(_0633_),
    .Y(_0013_));
 sg13g2_nor2_1 _1415_ (.A(\u_top_module.u_i2s_bus.counter[3] ),
    .B(_0633_),
    .Y(_0634_));
 sg13g2_and2_1 _1416_ (.A(\u_top_module.u_i2s_bus.counter[3] ),
    .B(_0633_),
    .X(_0635_));
 sg13g2_nor3_1 _1417_ (.A(_0629_),
    .B(_0634_),
    .C(_0635_),
    .Y(_0014_));
 sg13g2_nor2_1 _1418_ (.A(\u_top_module.u_i2s_bus.counter[4] ),
    .B(_0635_),
    .Y(_0636_));
 sg13g2_and2_1 _1419_ (.A(\u_top_module.u_i2s_bus.counter[4] ),
    .B(_0635_),
    .X(_0637_));
 sg13g2_nor3_1 _1420_ (.A(_0629_),
    .B(_0636_),
    .C(_0637_),
    .Y(_0015_));
 sg13g2_nand2_1 _1421_ (.Y(_0638_),
    .A(\u_top_module.u_i2s_bus.counter[5] ),
    .B(_0637_));
 sg13g2_xnor2_1 _1422_ (.Y(_0639_),
    .A(\u_top_module.u_i2s_bus.counter[5] ),
    .B(_0637_));
 sg13g2_nor2_1 _1423_ (.A(_0629_),
    .B(_0639_),
    .Y(_0016_));
 sg13g2_nor2_1 _1424_ (.A(_0629_),
    .B(_0638_),
    .Y(_0017_));
 sg13g2_nand2b_1 _1425_ (.Y(_0640_),
    .B(\u_top_module.u_i2s_bus.dec_clk ),
    .A_N(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.prev_lr_clk ));
 sg13g2_mux2_1 _1426_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ),
    .S(net891),
    .X(_0020_));
 sg13g2_mux2_1 _1427_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.out ),
    .S(net892),
    .X(_0021_));
 sg13g2_nand2_1 _1428_ (.Y(_0641_),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.out ),
    .B(net891));
 sg13g2_o21ai_1 _1429_ (.B1(_0641_),
    .Y(_0022_),
    .A1(_0556_),
    .A2(net891));
 sg13g2_nand2_1 _1430_ (.Y(_0642_),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.out ),
    .B(net891));
 sg13g2_o21ai_1 _1431_ (.B1(_0642_),
    .Y(_0023_),
    .A1(_0557_),
    .A2(net889));
 sg13g2_nand2_1 _1432_ (.Y(_0643_),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.out ),
    .B(net890));
 sg13g2_o21ai_1 _1433_ (.B1(_0643_),
    .Y(_0024_),
    .A1(_0558_),
    .A2(net889));
 sg13g2_mux2_1 _1434_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.out ),
    .S(net889),
    .X(_0025_));
 sg13g2_mux2_1 _1435_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.out ),
    .S(net889),
    .X(_0026_));
 sg13g2_nand2b_1 _1436_ (.Y(_0644_),
    .B(\u_top_module.u_decimator.counter[7] ),
    .A_N(\u_top_module.decimation_ratio[7] ));
 sg13g2_a22oi_1 _1437_ (.Y(_0645_),
    .B1(_0548_),
    .B2(\u_top_module.decimation_ratio[1] ),
    .A2(\u_top_module.decimation_ratio[0] ),
    .A1(_0547_));
 sg13g2_a221oi_1 _1438_ (.B2(_0551_),
    .C1(_0645_),
    .B1(\u_top_module.u_decimator.counter[2] ),
    .A1(\u_top_module.u_decimator.counter[1] ),
    .Y(_0646_),
    .A2(_0549_));
 sg13g2_nand2b_1 _1439_ (.Y(_0647_),
    .B(\u_top_module.decimation_ratio[3] ),
    .A_N(\u_top_module.u_decimator.counter[3] ));
 sg13g2_o21ai_1 _1440_ (.B1(_0647_),
    .Y(_0648_),
    .A1(\u_top_module.u_decimator.counter[2] ),
    .A2(_0551_));
 sg13g2_a22oi_1 _1441_ (.Y(_0649_),
    .B1(\u_top_module.u_decimator.counter[4] ),
    .B2(_0555_),
    .A2(_0550_),
    .A1(\u_top_module.u_decimator.counter[3] ));
 sg13g2_o21ai_1 _1442_ (.B1(_0649_),
    .Y(_0650_),
    .A1(_0646_),
    .A2(_0648_));
 sg13g2_a22oi_1 _1443_ (.Y(_0651_),
    .B1(_0554_),
    .B2(\u_top_module.decimation_ratio[4] ),
    .A2(\u_top_module.decimation_ratio[5] ),
    .A1(_0553_));
 sg13g2_nor2_1 _1444_ (.A(_0553_),
    .B(\u_top_module.decimation_ratio[5] ),
    .Y(_0652_));
 sg13g2_a221oi_1 _1445_ (.B2(_0651_),
    .C1(_0652_),
    .B1(_0650_),
    .A1(\u_top_module.u_decimator.counter[6] ),
    .Y(_0653_),
    .A2(_0552_));
 sg13g2_nand2b_1 _1446_ (.Y(_0654_),
    .B(\u_top_module.decimation_ratio[7] ),
    .A_N(\u_top_module.u_decimator.counter[7] ));
 sg13g2_o21ai_1 _1447_ (.B1(_0654_),
    .Y(_0655_),
    .A1(\u_top_module.u_decimator.counter[6] ),
    .A2(_0552_));
 sg13g2_o21ai_1 _1448_ (.B1(_0644_),
    .Y(_0656_),
    .A1(_0653_),
    .A2(_0655_));
 sg13g2_nor2_1 _1449_ (.A(\u_top_module.u_decimator.counter[0] ),
    .B(_0656_),
    .Y(_0002_));
 sg13g2_xnor2_1 _1450_ (.Y(_0657_),
    .A(\u_top_module.u_decimator.counter[0] ),
    .B(\u_top_module.u_decimator.counter[1] ));
 sg13g2_nor2_1 _1451_ (.A(_0656_),
    .B(_0657_),
    .Y(_0003_));
 sg13g2_and3_1 _1452_ (.X(_0658_),
    .A(\u_top_module.u_decimator.counter[0] ),
    .B(\u_top_module.u_decimator.counter[1] ),
    .C(\u_top_module.u_decimator.counter[2] ));
 sg13g2_a21oi_1 _1453_ (.A1(\u_top_module.u_decimator.counter[0] ),
    .A2(\u_top_module.u_decimator.counter[1] ),
    .Y(_0659_),
    .B1(\u_top_module.u_decimator.counter[2] ));
 sg13g2_nor3_1 _1454_ (.A(net792),
    .B(_0658_),
    .C(_0659_),
    .Y(_0004_));
 sg13g2_nor2_1 _1455_ (.A(\u_top_module.u_decimator.counter[3] ),
    .B(_0658_),
    .Y(_0660_));
 sg13g2_and2_1 _1456_ (.A(\u_top_module.u_decimator.counter[3] ),
    .B(_0658_),
    .X(_0661_));
 sg13g2_nor3_1 _1457_ (.A(net792),
    .B(_0660_),
    .C(_0661_),
    .Y(_0005_));
 sg13g2_nor2_1 _1458_ (.A(\u_top_module.u_decimator.counter[4] ),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_and2_1 _1459_ (.A(\u_top_module.u_decimator.counter[4] ),
    .B(_0661_),
    .X(_0663_));
 sg13g2_nor3_1 _1460_ (.A(net792),
    .B(_0662_),
    .C(_0663_),
    .Y(_0006_));
 sg13g2_xnor2_1 _1461_ (.Y(_0664_),
    .A(\u_top_module.u_decimator.counter[5] ),
    .B(_0663_));
 sg13g2_nor2_1 _1462_ (.A(net792),
    .B(_0664_),
    .Y(_0007_));
 sg13g2_a21oi_1 _1463_ (.A1(\u_top_module.u_decimator.counter[5] ),
    .A2(_0663_),
    .Y(_0665_),
    .B1(\u_top_module.u_decimator.counter[6] ));
 sg13g2_nand3_1 _1464_ (.B(\u_top_module.u_decimator.counter[5] ),
    .C(_0663_),
    .A(\u_top_module.u_decimator.counter[6] ),
    .Y(_0666_));
 sg13g2_nand2b_1 _1465_ (.Y(_0667_),
    .B(_0666_),
    .A_N(_0665_));
 sg13g2_nor2_1 _1466_ (.A(net792),
    .B(_0667_),
    .Y(_0008_));
 sg13g2_xor2_1 _1467_ (.B(_0666_),
    .A(\u_top_module.u_decimator.counter[7] ),
    .X(_0668_));
 sg13g2_nor2_1 _1468_ (.A(net792),
    .B(_0668_),
    .Y(_0009_));
 sg13g2_mux2_1 _1469_ (.A0(\u_top_module.dec_data ),
    .A1(net3),
    .S(net792),
    .X(_0064_));
 sg13g2_nor2_1 _1470_ (.A(_0565_),
    .B(net891),
    .Y(_0065_));
 sg13g2_mux2_1 _1471_ (.A0(\u_top_module.u_memory.memory[0][0] ),
    .A1(net950),
    .S(net896),
    .X(_0066_));
 sg13g2_mux2_1 _1472_ (.A0(\u_top_module.u_memory.memory[0][1] ),
    .A1(net949),
    .S(net895),
    .X(_0067_));
 sg13g2_mux2_1 _1473_ (.A0(\u_top_module.u_memory.memory[0][2] ),
    .A1(net948),
    .S(net896),
    .X(_0068_));
 sg13g2_mux2_1 _1474_ (.A0(\u_top_module.u_memory.memory[0][3] ),
    .A1(net947),
    .S(net896),
    .X(_0069_));
 sg13g2_mux2_1 _1475_ (.A0(\u_top_module.u_memory.memory[0][4] ),
    .A1(net946),
    .S(net895),
    .X(_0070_));
 sg13g2_mux2_1 _1476_ (.A0(\u_top_module.u_memory.memory[0][5] ),
    .A1(net945),
    .S(net896),
    .X(_0071_));
 sg13g2_mux2_1 _1477_ (.A0(\u_top_module.u_memory.memory[0][6] ),
    .A1(net944),
    .S(net895),
    .X(_0072_));
 sg13g2_mux2_1 _1478_ (.A0(\u_top_module.u_memory.memory[0][7] ),
    .A1(net943),
    .S(net895),
    .X(_0073_));
 sg13g2_mux2_1 _1479_ (.A0(\u_top_module.u_memory.memory[1][0] ),
    .A1(net950),
    .S(net874),
    .X(_0074_));
 sg13g2_mux2_1 _1480_ (.A0(\u_top_module.u_memory.memory[1][1] ),
    .A1(net949),
    .S(net873),
    .X(_0075_));
 sg13g2_mux2_1 _1481_ (.A0(\u_top_module.u_memory.memory[1][2] ),
    .A1(net948),
    .S(net874),
    .X(_0076_));
 sg13g2_mux2_1 _1482_ (.A0(\u_top_module.u_memory.memory[1][3] ),
    .A1(net947),
    .S(net873),
    .X(_0077_));
 sg13g2_mux2_1 _1483_ (.A0(\u_top_module.u_memory.memory[1][4] ),
    .A1(net946),
    .S(net873),
    .X(_0078_));
 sg13g2_mux2_1 _1484_ (.A0(\u_top_module.u_memory.memory[1][5] ),
    .A1(net945),
    .S(net874),
    .X(_0079_));
 sg13g2_mux2_1 _1485_ (.A0(\u_top_module.u_memory.memory[1][6] ),
    .A1(net944),
    .S(net874),
    .X(_0080_));
 sg13g2_mux2_1 _1486_ (.A0(\u_top_module.u_memory.memory[1][7] ),
    .A1(net943),
    .S(net873),
    .X(_0081_));
 sg13g2_mux2_1 _1487_ (.A0(\u_top_module.u_memory.memory[5][0] ),
    .A1(net950),
    .S(net872),
    .X(_0082_));
 sg13g2_mux2_1 _1488_ (.A0(\u_top_module.u_memory.memory[5][1] ),
    .A1(net949),
    .S(net871),
    .X(_0083_));
 sg13g2_mux2_1 _1489_ (.A0(\u_top_module.u_memory.memory[5][2] ),
    .A1(net948),
    .S(net872),
    .X(_0084_));
 sg13g2_mux2_1 _1490_ (.A0(\u_top_module.u_memory.memory[5][3] ),
    .A1(net947),
    .S(net871),
    .X(_0085_));
 sg13g2_mux2_1 _1491_ (.A0(\u_top_module.u_memory.memory[5][4] ),
    .A1(net946),
    .S(net871),
    .X(_0086_));
 sg13g2_mux2_1 _1492_ (.A0(\u_top_module.u_memory.memory[5][5] ),
    .A1(net945),
    .S(net872),
    .X(_0087_));
 sg13g2_mux2_1 _1493_ (.A0(\u_top_module.u_memory.memory[5][6] ),
    .A1(net944),
    .S(net872),
    .X(_0088_));
 sg13g2_mux2_1 _1494_ (.A0(\u_top_module.u_memory.memory[5][7] ),
    .A1(net943),
    .S(net871),
    .X(_0089_));
 sg13g2_mux2_1 _1495_ (.A0(\u_top_module.u_memory.memory[2][0] ),
    .A1(net950),
    .S(net876),
    .X(_0090_));
 sg13g2_mux2_1 _1496_ (.A0(\u_top_module.u_memory.memory[2][1] ),
    .A1(net949),
    .S(net875),
    .X(_0091_));
 sg13g2_mux2_1 _1497_ (.A0(\u_top_module.u_memory.memory[2][2] ),
    .A1(net948),
    .S(net876),
    .X(_0092_));
 sg13g2_mux2_1 _1498_ (.A0(\u_top_module.u_memory.memory[2][3] ),
    .A1(net947),
    .S(net875),
    .X(_0093_));
 sg13g2_mux2_1 _1499_ (.A0(\u_top_module.u_memory.memory[2][4] ),
    .A1(net946),
    .S(net875),
    .X(_0094_));
 sg13g2_mux2_1 _1500_ (.A0(\u_top_module.u_memory.memory[2][5] ),
    .A1(net945),
    .S(net876),
    .X(_0095_));
 sg13g2_mux2_1 _1501_ (.A0(\u_top_module.u_memory.memory[2][6] ),
    .A1(net944),
    .S(net876),
    .X(_0096_));
 sg13g2_mux2_1 _1502_ (.A0(\u_top_module.u_memory.memory[2][7] ),
    .A1(net943),
    .S(net875),
    .X(_0097_));
 sg13g2_mux2_1 _1503_ (.A0(\u_top_module.u_memory.memory[3][0] ),
    .A1(net950),
    .S(net882),
    .X(_0098_));
 sg13g2_mux2_1 _1504_ (.A0(\u_top_module.u_memory.memory[3][1] ),
    .A1(net949),
    .S(net881),
    .X(_0099_));
 sg13g2_mux2_1 _1505_ (.A0(\u_top_module.u_memory.memory[3][2] ),
    .A1(net948),
    .S(net882),
    .X(_0100_));
 sg13g2_mux2_1 _1506_ (.A0(\u_top_module.u_memory.memory[3][3] ),
    .A1(net947),
    .S(net881),
    .X(_0101_));
 sg13g2_mux2_1 _1507_ (.A0(\u_top_module.u_memory.memory[3][4] ),
    .A1(net946),
    .S(net881),
    .X(_0102_));
 sg13g2_mux2_1 _1508_ (.A0(\u_top_module.u_memory.memory[3][5] ),
    .A1(net945),
    .S(net882),
    .X(_0103_));
 sg13g2_mux2_1 _1509_ (.A0(\u_top_module.u_memory.memory[3][6] ),
    .A1(net944),
    .S(net882),
    .X(_0104_));
 sg13g2_mux2_1 _1510_ (.A0(\u_top_module.u_memory.memory[3][7] ),
    .A1(net943),
    .S(net881),
    .X(_0105_));
 sg13g2_mux2_1 _1511_ (.A0(\u_top_module.u_memory.memory[6][0] ),
    .A1(net950),
    .S(net878),
    .X(_0106_));
 sg13g2_mux2_1 _1512_ (.A0(\u_top_module.u_memory.memory[6][1] ),
    .A1(net949),
    .S(net877),
    .X(_0107_));
 sg13g2_mux2_1 _1513_ (.A0(\u_top_module.u_memory.memory[6][2] ),
    .A1(net948),
    .S(net878),
    .X(_0108_));
 sg13g2_mux2_1 _1514_ (.A0(\u_top_module.u_memory.memory[6][3] ),
    .A1(net947),
    .S(net877),
    .X(_0109_));
 sg13g2_mux2_1 _1515_ (.A0(\u_top_module.u_memory.memory[6][4] ),
    .A1(net946),
    .S(net877),
    .X(_0110_));
 sg13g2_mux2_1 _1516_ (.A0(\u_top_module.u_memory.memory[6][5] ),
    .A1(net945),
    .S(net878),
    .X(_0111_));
 sg13g2_mux2_1 _1517_ (.A0(\u_top_module.u_memory.memory[6][6] ),
    .A1(net944),
    .S(net878),
    .X(_0112_));
 sg13g2_mux2_1 _1518_ (.A0(\u_top_module.u_memory.memory[6][7] ),
    .A1(net943),
    .S(net877),
    .X(_0113_));
 sg13g2_mux2_1 _1519_ (.A0(\u_top_module.u_memory.memory[4][0] ),
    .A1(net950),
    .S(net894),
    .X(_0114_));
 sg13g2_mux2_1 _1520_ (.A0(\u_top_module.u_memory.memory[4][1] ),
    .A1(net949),
    .S(net893),
    .X(_0115_));
 sg13g2_mux2_1 _1521_ (.A0(\u_top_module.u_memory.memory[4][2] ),
    .A1(net948),
    .S(net894),
    .X(_0116_));
 sg13g2_mux2_1 _1522_ (.A0(\u_top_module.u_memory.memory[4][3] ),
    .A1(net947),
    .S(net893),
    .X(_0117_));
 sg13g2_mux2_1 _1523_ (.A0(\u_top_module.u_memory.memory[4][4] ),
    .A1(net946),
    .S(net893),
    .X(_0118_));
 sg13g2_mux2_1 _1524_ (.A0(\u_top_module.u_memory.memory[4][5] ),
    .A1(net945),
    .S(net894),
    .X(_0119_));
 sg13g2_mux2_1 _1525_ (.A0(\u_top_module.u_memory.memory[4][6] ),
    .A1(net944),
    .S(net894),
    .X(_0120_));
 sg13g2_mux2_1 _1526_ (.A0(\u_top_module.u_memory.memory[4][7] ),
    .A1(net943),
    .S(net893),
    .X(_0121_));
 sg13g2_nor2_2 _1527_ (.A(_0030_),
    .B(\u_top_module.u_spi_port.cs_n_prev ),
    .Y(_0669_));
 sg13g2_mux2_1 _1528_ (.A0(\u_top_module.capture_reg[0] ),
    .A1(\u_top_module.u_spi_port.shift_reg[0] ),
    .S(net885),
    .X(_0122_));
 sg13g2_mux2_1 _1529_ (.A0(\u_top_module.capture_reg[1] ),
    .A1(\u_top_module.u_spi_port.shift_reg[1] ),
    .S(net886),
    .X(_0123_));
 sg13g2_mux2_1 _1530_ (.A0(\u_top_module.capture_reg[2] ),
    .A1(\u_top_module.u_spi_port.shift_reg[2] ),
    .S(net886),
    .X(_0124_));
 sg13g2_mux2_1 _1531_ (.A0(\u_top_module.capture_reg[3] ),
    .A1(\u_top_module.u_spi_port.shift_reg[3] ),
    .S(net886),
    .X(_0125_));
 sg13g2_mux2_1 _1532_ (.A0(\u_top_module.capture_reg[4] ),
    .A1(\u_top_module.u_spi_port.shift_reg[4] ),
    .S(net886),
    .X(_0126_));
 sg13g2_mux2_1 _1533_ (.A0(\u_top_module.capture_reg[5] ),
    .A1(\u_top_module.u_spi_port.shift_reg[5] ),
    .S(net886),
    .X(_0127_));
 sg13g2_mux2_1 _1534_ (.A0(\u_top_module.capture_reg[6] ),
    .A1(\u_top_module.u_spi_port.shift_reg[6] ),
    .S(net886),
    .X(_0128_));
 sg13g2_mux2_1 _1535_ (.A0(\u_top_module.capture_reg[7] ),
    .A1(\u_top_module.u_spi_port.shift_reg[7] ),
    .S(net886),
    .X(_0129_));
 sg13g2_mux2_1 _1536_ (.A0(\u_top_module.addr[0] ),
    .A1(\u_top_module.u_spi_port.shift_reg[8] ),
    .S(net885),
    .X(_0130_));
 sg13g2_nand2_1 _1537_ (.Y(_0670_),
    .A(\u_top_module.u_spi_port.shift_reg[9] ),
    .B(net885));
 sg13g2_o21ai_1 _1538_ (.B1(_0670_),
    .Y(_0131_),
    .A1(_0546_),
    .A2(net885));
 sg13g2_mux2_1 _1539_ (.A0(\u_top_module.addr[2] ),
    .A1(\u_top_module.u_spi_port.shift_reg[10] ),
    .S(net885),
    .X(_0132_));
 sg13g2_mux2_1 _1540_ (.A0(\u_top_module.addr[3] ),
    .A1(\u_top_module.u_spi_port.shift_reg[11] ),
    .S(_0669_),
    .X(_0133_));
 sg13g2_mux2_1 _1541_ (.A0(\u_top_module.addr[4] ),
    .A1(\u_top_module.u_spi_port.shift_reg[12] ),
    .S(_0669_),
    .X(_0134_));
 sg13g2_mux2_1 _1542_ (.A0(\u_top_module.addr[5] ),
    .A1(\u_top_module.u_spi_port.shift_reg[13] ),
    .S(net885),
    .X(_0135_));
 sg13g2_mux2_1 _1543_ (.A0(\u_top_module.addr[6] ),
    .A1(\u_top_module.u_spi_port.shift_reg[14] ),
    .S(net885),
    .X(_0136_));
 sg13g2_mux2_1 _1544_ (.A0(\u_top_module.addr[7] ),
    .A1(\u_top_module.u_spi_port.shift_reg[15] ),
    .S(net885),
    .X(_0137_));
 sg13g2_mux2_1 _1545_ (.A0(\u_top_module.u_memory.memory[7][0] ),
    .A1(net950),
    .S(net880),
    .X(_0138_));
 sg13g2_mux2_1 _1546_ (.A0(\u_top_module.u_memory.memory[7][1] ),
    .A1(net949),
    .S(net879),
    .X(_0139_));
 sg13g2_mux2_1 _1547_ (.A0(\u_top_module.u_memory.memory[7][2] ),
    .A1(net948),
    .S(net880),
    .X(_0140_));
 sg13g2_mux2_1 _1548_ (.A0(\u_top_module.u_memory.memory[7][3] ),
    .A1(net947),
    .S(net879),
    .X(_0141_));
 sg13g2_mux2_1 _1549_ (.A0(\u_top_module.u_memory.memory[7][4] ),
    .A1(net946),
    .S(net879),
    .X(_0142_));
 sg13g2_mux2_1 _1550_ (.A0(\u_top_module.u_memory.memory[7][5] ),
    .A1(net945),
    .S(net880),
    .X(_0143_));
 sg13g2_mux2_1 _1551_ (.A0(\u_top_module.u_memory.memory[7][6] ),
    .A1(net944),
    .S(net880),
    .X(_0144_));
 sg13g2_mux2_1 _1552_ (.A0(\u_top_module.u_memory.memory[7][7] ),
    .A1(net943),
    .S(net879),
    .X(_0145_));
 sg13g2_nand2_1 _1553_ (.Y(_0671_),
    .A(_0030_),
    .B(net979));
 sg13g2_mux2_1 _1554_ (.A0(net1),
    .A1(\u_top_module.u_spi_port.shift_reg[0] ),
    .S(net884),
    .X(_0146_));
 sg13g2_mux2_1 _1555_ (.A0(\u_top_module.u_spi_port.shift_reg[0] ),
    .A1(\u_top_module.u_spi_port.shift_reg[1] ),
    .S(net883),
    .X(_0147_));
 sg13g2_mux2_1 _1556_ (.A0(\u_top_module.u_spi_port.shift_reg[1] ),
    .A1(\u_top_module.u_spi_port.shift_reg[2] ),
    .S(net883),
    .X(_0148_));
 sg13g2_mux2_1 _1557_ (.A0(\u_top_module.u_spi_port.shift_reg[2] ),
    .A1(\u_top_module.u_spi_port.shift_reg[3] ),
    .S(net883),
    .X(_0149_));
 sg13g2_mux2_1 _1558_ (.A0(\u_top_module.u_spi_port.shift_reg[3] ),
    .A1(\u_top_module.u_spi_port.shift_reg[4] ),
    .S(net883),
    .X(_0150_));
 sg13g2_mux2_1 _1559_ (.A0(\u_top_module.u_spi_port.shift_reg[4] ),
    .A1(\u_top_module.u_spi_port.shift_reg[5] ),
    .S(net883),
    .X(_0151_));
 sg13g2_mux2_1 _1560_ (.A0(\u_top_module.u_spi_port.shift_reg[5] ),
    .A1(\u_top_module.u_spi_port.shift_reg[6] ),
    .S(net883),
    .X(_0152_));
 sg13g2_mux2_1 _1561_ (.A0(\u_top_module.u_spi_port.shift_reg[6] ),
    .A1(\u_top_module.u_spi_port.shift_reg[7] ),
    .S(net883),
    .X(_0153_));
 sg13g2_mux2_1 _1562_ (.A0(\u_top_module.u_spi_port.shift_reg[7] ),
    .A1(\u_top_module.u_spi_port.shift_reg[8] ),
    .S(net883),
    .X(_0154_));
 sg13g2_mux2_1 _1563_ (.A0(\u_top_module.u_spi_port.shift_reg[8] ),
    .A1(\u_top_module.u_spi_port.shift_reg[9] ),
    .S(net884),
    .X(_0155_));
 sg13g2_mux2_1 _1564_ (.A0(\u_top_module.u_spi_port.shift_reg[9] ),
    .A1(\u_top_module.u_spi_port.shift_reg[10] ),
    .S(net884),
    .X(_0156_));
 sg13g2_mux2_1 _1565_ (.A0(\u_top_module.u_spi_port.shift_reg[10] ),
    .A1(\u_top_module.u_spi_port.shift_reg[11] ),
    .S(net884),
    .X(_0157_));
 sg13g2_mux2_1 _1566_ (.A0(\u_top_module.u_spi_port.shift_reg[11] ),
    .A1(\u_top_module.u_spi_port.shift_reg[12] ),
    .S(net884),
    .X(_0158_));
 sg13g2_mux2_1 _1567_ (.A0(\u_top_module.u_spi_port.shift_reg[12] ),
    .A1(\u_top_module.u_spi_port.shift_reg[13] ),
    .S(net884),
    .X(_0159_));
 sg13g2_mux2_1 _1568_ (.A0(\u_top_module.u_spi_port.shift_reg[13] ),
    .A1(\u_top_module.u_spi_port.shift_reg[14] ),
    .S(net884),
    .X(_0160_));
 sg13g2_mux2_1 _1569_ (.A0(\u_top_module.u_spi_port.shift_reg[14] ),
    .A1(\u_top_module.u_spi_port.shift_reg[15] ),
    .S(net884),
    .X(_0161_));
 sg13g2_nor2_1 _1570_ (.A(net845),
    .B(net861),
    .Y(_0672_));
 sg13g2_or2_2 _1571_ (.X(_0673_),
    .B(net865),
    .A(net849));
 sg13g2_nor3_2 _1572_ (.A(net836),
    .B(net849),
    .C(net863),
    .Y(_0674_));
 sg13g2_or3_1 _1573_ (.A(net836),
    .B(net848),
    .C(net863),
    .X(_0675_));
 sg13g2_nor4_2 _1574_ (.A(\u_top_module.filter_length[3] ),
    .B(net836),
    .C(net850),
    .Y(_0676_),
    .D(net864));
 sg13g2_and2_1 _1575_ (.A(_0559_),
    .B(_0676_),
    .X(_0677_));
 sg13g2_nor3_1 _1576_ (.A(\u_top_module.filter_length[7] ),
    .B(\u_top_module.filter_length[6] ),
    .C(\u_top_module.filter_length[5] ),
    .Y(_0678_));
 sg13g2_and3_2 _1577_ (.X(_0679_),
    .A(_0559_),
    .B(_0676_),
    .C(_0678_));
 sg13g2_nand3_1 _1578_ (.B(_0676_),
    .C(_0678_),
    .A(_0559_),
    .Y(_0680_));
 sg13g2_nand3_1 _1579_ (.B(\u_top_module.u_filter.shift_reg[159] ),
    .C(net805),
    .A(net830),
    .Y(_0681_));
 sg13g2_and2_1 _1580_ (.A(net845),
    .B(net861),
    .X(_0682_));
 sg13g2_nand2_1 _1581_ (.Y(_0683_),
    .A(net844),
    .B(net861));
 sg13g2_o21ai_1 _1582_ (.B1(net823),
    .Y(_0684_),
    .A1(\u_top_module.u_filter.shift_reg[158] ),
    .A2(net812));
 sg13g2_o21ai_1 _1583_ (.B1(net835),
    .Y(_0685_),
    .A1(net844),
    .A2(net861));
 sg13g2_or2_1 _1584_ (.X(_0686_),
    .B(\u_top_module.u_filter.shift_reg[157] ),
    .A(net858));
 sg13g2_o21ai_1 _1585_ (.B1(_0686_),
    .Y(_0687_),
    .A1(net841),
    .A2(\u_top_module.u_filter.shift_reg[156] ));
 sg13g2_and2_2 _1586_ (.A(net820),
    .B(net809),
    .X(_0688_));
 sg13g2_nand2_1 _1587_ (.Y(_0689_),
    .A(net820),
    .B(net809));
 sg13g2_a221oi_1 _1588_ (.B2(net819),
    .C1(net800),
    .B1(_0687_),
    .A1(_0681_),
    .Y(_0690_),
    .A2(_0684_));
 sg13g2_xnor2_1 _1589_ (.Y(_0691_),
    .A(\u_top_module.filter_length[4] ),
    .B(_0676_));
 sg13g2_xnor2_1 _1590_ (.Y(_0692_),
    .A(_0559_),
    .B(_0676_));
 sg13g2_nor2_1 _1591_ (.A(net858),
    .B(\u_top_module.u_filter.shift_reg[153] ),
    .Y(_0693_));
 sg13g2_nor2_1 _1592_ (.A(net841),
    .B(\u_top_module.u_filter.shift_reg[152] ),
    .Y(_0694_));
 sg13g2_o21ai_1 _1593_ (.B1(net824),
    .Y(_0695_),
    .A1(_0693_),
    .A2(_0694_));
 sg13g2_o21ai_1 _1594_ (.B1(net800),
    .Y(_0696_),
    .A1(net832),
    .A2(\u_top_module.u_filter.shift_reg[155] ));
 sg13g2_o21ai_1 _1595_ (.B1(_0695_),
    .Y(_0697_),
    .A1(\u_top_module.u_filter.shift_reg[154] ),
    .A2(net812));
 sg13g2_o21ai_1 _1596_ (.B1(net797),
    .Y(_0698_),
    .A1(_0696_),
    .A2(_0697_));
 sg13g2_xnor2_1 _1597_ (.Y(_0699_),
    .A(\u_top_module.filter_length[3] ),
    .B(_0674_));
 sg13g2_xnor2_1 _1598_ (.Y(_0700_),
    .A(\u_top_module.filter_length[3] ),
    .B(net822));
 sg13g2_a21o_1 _1599_ (.A2(\u_top_module.u_filter.shift_reg[141] ),
    .A1(net840),
    .B1(net857),
    .X(_0701_));
 sg13g2_or2_1 _1600_ (.X(_0702_),
    .B(\u_top_module.u_filter.shift_reg[140] ),
    .A(net841));
 sg13g2_a22oi_1 _1601_ (.Y(_0703_),
    .B1(_0701_),
    .B2(_0702_),
    .A2(net829),
    .A1(\u_top_module.u_filter.shift_reg[143] ));
 sg13g2_nor2_1 _1602_ (.A(\u_top_module.u_filter.shift_reg[142] ),
    .B(net812),
    .Y(_0704_));
 sg13g2_or3_1 _1603_ (.A(net800),
    .B(_0703_),
    .C(_0704_),
    .X(_0705_));
 sg13g2_nor2_1 _1604_ (.A(net857),
    .B(\u_top_module.u_filter.shift_reg[137] ),
    .Y(_0706_));
 sg13g2_nor2_1 _1605_ (.A(net840),
    .B(\u_top_module.u_filter.shift_reg[136] ),
    .Y(_0707_));
 sg13g2_o21ai_1 _1606_ (.B1(net824),
    .Y(_0708_),
    .A1(_0706_),
    .A2(_0707_));
 sg13g2_nand3b_1 _1607_ (.B(net857),
    .C(net840),
    .Y(_0709_),
    .A_N(\u_top_module.u_filter.shift_reg[138] ));
 sg13g2_nand2b_1 _1608_ (.Y(_0710_),
    .B(net834),
    .A_N(\u_top_module.u_filter.shift_reg[139] ));
 sg13g2_and4_1 _1609_ (.A(net819),
    .B(net809),
    .C(_0709_),
    .D(_0710_),
    .X(_0711_));
 sg13g2_a21oi_1 _1610_ (.A1(_0708_),
    .A2(_0711_),
    .Y(_0712_),
    .B1(net797));
 sg13g2_a21oi_1 _1611_ (.A1(_0705_),
    .A2(_0712_),
    .Y(_0713_),
    .B1(_0699_));
 sg13g2_o21ai_1 _1612_ (.B1(_0713_),
    .Y(_0714_),
    .A1(_0690_),
    .A2(_0698_));
 sg13g2_nor2b_1 _1613_ (.A(\u_top_module.filter_length[5] ),
    .B_N(_0677_),
    .Y(_0715_));
 sg13g2_xnor2_1 _1614_ (.Y(_0716_),
    .A(\u_top_module.filter_length[5] ),
    .B(_0677_));
 sg13g2_xor2_1 _1615_ (.B(_0677_),
    .A(\u_top_module.filter_length[5] ),
    .X(_0717_));
 sg13g2_mux4_1 _1616_ (.S0(net857),
    .A0(\u_top_module.u_filter.shift_reg[135] ),
    .A1(\u_top_module.u_filter.shift_reg[132] ),
    .A2(\u_top_module.u_filter.shift_reg[133] ),
    .A3(\u_top_module.u_filter.shift_reg[134] ),
    .S1(net840),
    .X(_0718_));
 sg13g2_nand3_1 _1617_ (.B(net798),
    .C(_0718_),
    .A(net806),
    .Y(_0719_));
 sg13g2_nor2_1 _1618_ (.A(net857),
    .B(\u_top_module.u_filter.shift_reg[129] ),
    .Y(_0720_));
 sg13g2_nor2_1 _1619_ (.A(net840),
    .B(\u_top_module.u_filter.shift_reg[128] ),
    .Y(_0721_));
 sg13g2_o21ai_1 _1620_ (.B1(net824),
    .Y(_0722_),
    .A1(_0720_),
    .A2(_0721_));
 sg13g2_nand2b_1 _1621_ (.Y(_0723_),
    .B(net834),
    .A_N(\u_top_module.u_filter.shift_reg[131] ));
 sg13g2_nand2b_1 _1622_ (.Y(_0724_),
    .B(net818),
    .A_N(\u_top_module.u_filter.shift_reg[130] ));
 sg13g2_nand4_1 _1623_ (.B(_0722_),
    .C(_0723_),
    .A(net800),
    .Y(_0725_),
    .D(_0724_));
 sg13g2_nand3_1 _1624_ (.B(_0719_),
    .C(_0725_),
    .A(_0691_),
    .Y(_0726_));
 sg13g2_nor2_1 _1625_ (.A(net857),
    .B(\u_top_module.u_filter.shift_reg[145] ),
    .Y(_0727_));
 sg13g2_nor2_1 _1626_ (.A(net840),
    .B(\u_top_module.u_filter.shift_reg[144] ),
    .Y(_0728_));
 sg13g2_o21ai_1 _1627_ (.B1(net824),
    .Y(_0729_),
    .A1(_0727_),
    .A2(_0728_));
 sg13g2_nand2b_1 _1628_ (.Y(_0730_),
    .B(net834),
    .A_N(\u_top_module.u_filter.shift_reg[147] ));
 sg13g2_nand2b_1 _1629_ (.Y(_0731_),
    .B(net818),
    .A_N(\u_top_module.u_filter.shift_reg[146] ));
 sg13g2_nand4_1 _1630_ (.B(_0729_),
    .C(_0730_),
    .A(net800),
    .Y(_0732_),
    .D(_0731_));
 sg13g2_nand3_1 _1631_ (.B(net857),
    .C(\u_top_module.u_filter.shift_reg[150] ),
    .A(net840),
    .Y(_0733_));
 sg13g2_nand2b_1 _1632_ (.Y(_0734_),
    .B(\u_top_module.u_filter.shift_reg[149] ),
    .A_N(net857));
 sg13g2_nand2b_1 _1633_ (.Y(_0735_),
    .B(\u_top_module.u_filter.shift_reg[148] ),
    .A_N(net840));
 sg13g2_nand4_1 _1634_ (.B(_0733_),
    .C(_0734_),
    .A(net824),
    .Y(_0736_),
    .D(_0735_));
 sg13g2_o21ai_1 _1635_ (.B1(net809),
    .Y(_0737_),
    .A1(_0563_),
    .A2(net819));
 sg13g2_a21oi_1 _1636_ (.A1(_0736_),
    .A2(_0737_),
    .Y(_0738_),
    .B1(_0691_));
 sg13g2_a21oi_2 _1637_ (.B1(net793),
    .Y(_0739_),
    .A2(_0738_),
    .A1(_0732_));
 sg13g2_a21oi_1 _1638_ (.A1(_0726_),
    .A2(_0739_),
    .Y(_0740_),
    .B1(_0717_));
 sg13g2_nand2b_1 _1639_ (.Y(_0741_),
    .B(_0715_),
    .A_N(\u_top_module.filter_length[6] ));
 sg13g2_nand2b_1 _1640_ (.Y(_0742_),
    .B(\u_top_module.filter_length[6] ),
    .A_N(_0715_));
 sg13g2_nand2_2 _1641_ (.Y(_0743_),
    .A(_0741_),
    .B(_0742_));
 sg13g2_nand3_1 _1642_ (.B(\u_top_module.u_filter.shift_reg[191] ),
    .C(net805),
    .A(net830),
    .Y(_0744_));
 sg13g2_o21ai_1 _1643_ (.B1(net825),
    .Y(_0745_),
    .A1(\u_top_module.u_filter.shift_reg[190] ),
    .A2(net813));
 sg13g2_or2_1 _1644_ (.X(_0746_),
    .B(\u_top_module.u_filter.shift_reg[189] ),
    .A(net859));
 sg13g2_o21ai_1 _1645_ (.B1(_0746_),
    .Y(_0747_),
    .A1(net843),
    .A2(\u_top_module.u_filter.shift_reg[188] ));
 sg13g2_a221oi_1 _1646_ (.B2(net819),
    .C1(net802),
    .B1(_0747_),
    .A1(_0744_),
    .Y(_0748_),
    .A2(_0745_));
 sg13g2_nor2_1 _1647_ (.A(net856),
    .B(\u_top_module.u_filter.shift_reg[185] ),
    .Y(_0749_));
 sg13g2_nor2_1 _1648_ (.A(net842),
    .B(\u_top_module.u_filter.shift_reg[184] ),
    .Y(_0750_));
 sg13g2_o21ai_1 _1649_ (.B1(net823),
    .Y(_0751_),
    .A1(_0749_),
    .A2(_0750_));
 sg13g2_o21ai_1 _1650_ (.B1(net801),
    .Y(_0752_),
    .A1(net832),
    .A2(\u_top_module.u_filter.shift_reg[187] ));
 sg13g2_o21ai_1 _1651_ (.B1(_0751_),
    .Y(_0753_),
    .A1(\u_top_module.u_filter.shift_reg[186] ),
    .A2(net812));
 sg13g2_o21ai_1 _1652_ (.B1(net793),
    .Y(_0754_),
    .A1(_0752_),
    .A2(_0753_));
 sg13g2_nor2_1 _1653_ (.A(net856),
    .B(\u_top_module.u_filter.shift_reg[177] ),
    .Y(_0755_));
 sg13g2_nor2_1 _1654_ (.A(net839),
    .B(\u_top_module.u_filter.shift_reg[176] ),
    .Y(_0756_));
 sg13g2_o21ai_1 _1655_ (.B1(net823),
    .Y(_0757_),
    .A1(_0755_),
    .A2(_0756_));
 sg13g2_nand2b_1 _1656_ (.Y(_0758_),
    .B(net834),
    .A_N(\u_top_module.u_filter.shift_reg[179] ));
 sg13g2_nand3b_1 _1657_ (.B(net856),
    .C(net839),
    .Y(_0759_),
    .A_N(\u_top_module.u_filter.shift_reg[178] ));
 sg13g2_and4_1 _1658_ (.A(net819),
    .B(net809),
    .C(_0758_),
    .D(_0759_),
    .X(_0760_));
 sg13g2_a21oi_1 _1659_ (.A1(_0757_),
    .A2(_0760_),
    .Y(_0761_),
    .B1(net793));
 sg13g2_mux4_1 _1660_ (.S0(net856),
    .A0(\u_top_module.u_filter.shift_reg[183] ),
    .A1(\u_top_module.u_filter.shift_reg[180] ),
    .A2(\u_top_module.u_filter.shift_reg[181] ),
    .A3(\u_top_module.u_filter.shift_reg[182] ),
    .S1(net839),
    .X(_0762_));
 sg13g2_nand3_1 _1661_ (.B(net798),
    .C(_0762_),
    .A(net805),
    .Y(_0763_));
 sg13g2_a21oi_1 _1662_ (.A1(_0761_),
    .A2(_0763_),
    .Y(_0764_),
    .B1(_0691_));
 sg13g2_o21ai_1 _1663_ (.B1(_0764_),
    .Y(_0765_),
    .A1(_0748_),
    .A2(_0754_));
 sg13g2_nor2_1 _1664_ (.A(net860),
    .B(\u_top_module.u_filter.shift_reg[161] ),
    .Y(_0766_));
 sg13g2_nor2_1 _1665_ (.A(net844),
    .B(\u_top_module.u_filter.shift_reg[160] ),
    .Y(_0767_));
 sg13g2_o21ai_1 _1666_ (.B1(net825),
    .Y(_0768_),
    .A1(_0766_),
    .A2(_0767_));
 sg13g2_nand2b_1 _1667_ (.Y(_0769_),
    .B(net835),
    .A_N(\u_top_module.u_filter.shift_reg[163] ));
 sg13g2_nand3b_1 _1668_ (.B(net860),
    .C(net844),
    .Y(_0770_),
    .A_N(\u_top_module.u_filter.shift_reg[162] ));
 sg13g2_and4_1 _1669_ (.A(net820),
    .B(net811),
    .C(_0769_),
    .D(_0770_),
    .X(_0771_));
 sg13g2_and2_1 _1670_ (.A(\u_top_module.u_filter.shift_reg[167] ),
    .B(_0674_),
    .X(_0772_));
 sg13g2_nor2_1 _1671_ (.A(net845),
    .B(\u_top_module.u_filter.shift_reg[164] ),
    .Y(_0205_));
 sg13g2_nor2_1 _1672_ (.A(net861),
    .B(\u_top_module.u_filter.shift_reg[165] ),
    .Y(_0206_));
 sg13g2_nor3_1 _1673_ (.A(net809),
    .B(_0205_),
    .C(_0206_),
    .Y(_0207_));
 sg13g2_nand2b_1 _1674_ (.Y(_0208_),
    .B(net818),
    .A_N(\u_top_module.u_filter.shift_reg[166] ));
 sg13g2_o21ai_1 _1675_ (.B1(_0208_),
    .Y(_0209_),
    .A1(_0772_),
    .A2(_0207_));
 sg13g2_a21oi_1 _1676_ (.A1(_0768_),
    .A2(_0771_),
    .Y(_0210_),
    .B1(net796));
 sg13g2_nor2_1 _1677_ (.A(net860),
    .B(\u_top_module.u_filter.shift_reg[169] ),
    .Y(_0211_));
 sg13g2_nor2_1 _1678_ (.A(net843),
    .B(\u_top_module.u_filter.shift_reg[168] ),
    .Y(_0212_));
 sg13g2_o21ai_1 _1679_ (.B1(net832),
    .Y(_0213_),
    .A1(_0211_),
    .A2(_0212_));
 sg13g2_nand2b_1 _1680_ (.Y(_0214_),
    .B(net818),
    .A_N(\u_top_module.u_filter.shift_reg[170] ));
 sg13g2_nand2b_1 _1681_ (.Y(_0215_),
    .B(net834),
    .A_N(\u_top_module.u_filter.shift_reg[171] ));
 sg13g2_nand4_1 _1682_ (.B(_0213_),
    .C(_0214_),
    .A(net802),
    .Y(_0216_),
    .D(_0215_));
 sg13g2_mux4_1 _1683_ (.S0(net858),
    .A0(\u_top_module.u_filter.shift_reg[175] ),
    .A1(\u_top_module.u_filter.shift_reg[172] ),
    .A2(\u_top_module.u_filter.shift_reg[173] ),
    .A3(\u_top_module.u_filter.shift_reg[174] ),
    .S1(net841),
    .X(_0217_));
 sg13g2_a21oi_1 _1684_ (.A1(net798),
    .A2(_0217_),
    .Y(_0218_),
    .B1(_0699_));
 sg13g2_a221oi_1 _1685_ (.B2(_0218_),
    .C1(net797),
    .B1(_0216_),
    .A1(_0209_),
    .Y(_0219_),
    .A2(_0210_));
 sg13g2_nor2_1 _1686_ (.A(_0716_),
    .B(_0219_),
    .Y(_0220_));
 sg13g2_a221oi_1 _1687_ (.B2(_0220_),
    .C1(_0743_),
    .B1(_0765_),
    .A1(_0714_),
    .Y(_0221_),
    .A2(_0740_));
 sg13g2_nand3_1 _1688_ (.B(\u_top_module.u_filter.shift_reg[223] ),
    .C(net808),
    .A(net831),
    .Y(_0222_));
 sg13g2_o21ai_1 _1689_ (.B1(net828),
    .Y(_0223_),
    .A1(\u_top_module.u_filter.shift_reg[222] ),
    .A2(net815));
 sg13g2_or2_1 _1690_ (.X(_0224_),
    .B(\u_top_module.u_filter.shift_reg[221] ),
    .A(net868));
 sg13g2_o21ai_1 _1691_ (.B1(_0224_),
    .Y(_0225_),
    .A1(net853),
    .A2(\u_top_module.u_filter.shift_reg[220] ));
 sg13g2_a221oi_1 _1692_ (.B2(net822),
    .C1(net804),
    .B1(_0225_),
    .A1(_0222_),
    .Y(_0226_),
    .A2(_0223_));
 sg13g2_nor2_1 _1693_ (.A(net869),
    .B(\u_top_module.u_filter.shift_reg[217] ),
    .Y(_0227_));
 sg13g2_nor2_1 _1694_ (.A(net853),
    .B(\u_top_module.u_filter.shift_reg[216] ),
    .Y(_0228_));
 sg13g2_o21ai_1 _1695_ (.B1(net828),
    .Y(_0229_),
    .A1(_0227_),
    .A2(_0228_));
 sg13g2_o21ai_1 _1696_ (.B1(net804),
    .Y(_0230_),
    .A1(net833),
    .A2(\u_top_module.u_filter.shift_reg[219] ));
 sg13g2_o21ai_1 _1697_ (.B1(_0229_),
    .Y(_0231_),
    .A1(\u_top_module.u_filter.shift_reg[218] ),
    .A2(net815));
 sg13g2_o21ai_1 _1698_ (.B1(net795),
    .Y(_0232_),
    .A1(_0230_),
    .A2(_0231_));
 sg13g2_a21o_1 _1699_ (.A2(\u_top_module.u_filter.shift_reg[213] ),
    .A1(net830),
    .B1(net829),
    .X(_0233_));
 sg13g2_nor2b_1 _1700_ (.A(net854),
    .B_N(\u_top_module.u_filter.shift_reg[212] ),
    .Y(_0234_));
 sg13g2_a21o_1 _1701_ (.A2(net818),
    .A1(\u_top_module.u_filter.shift_reg[214] ),
    .B1(_0234_),
    .X(_0235_));
 sg13g2_o21ai_1 _1702_ (.B1(net811),
    .Y(_0236_),
    .A1(_0564_),
    .A2(net821));
 sg13g2_o21ai_1 _1703_ (.B1(_0236_),
    .Y(_0237_),
    .A1(_0233_),
    .A2(_0235_));
 sg13g2_nor2_1 _1704_ (.A(net868),
    .B(\u_top_module.u_filter.shift_reg[209] ),
    .Y(_0238_));
 sg13g2_nor2_1 _1705_ (.A(net854),
    .B(\u_top_module.u_filter.shift_reg[208] ),
    .Y(_0239_));
 sg13g2_o21ai_1 _1706_ (.B1(net833),
    .Y(_0240_),
    .A1(_0238_),
    .A2(_0239_));
 sg13g2_nand2b_1 _1707_ (.Y(_0241_),
    .B(net837),
    .A_N(\u_top_module.u_filter.shift_reg[211] ));
 sg13g2_nand3b_1 _1708_ (.B(net868),
    .C(net854),
    .Y(_0242_),
    .A_N(\u_top_module.u_filter.shift_reg[210] ));
 sg13g2_and4_1 _1709_ (.A(net821),
    .B(net810),
    .C(_0241_),
    .D(_0242_),
    .X(_0243_));
 sg13g2_a21oi_1 _1710_ (.A1(_0240_),
    .A2(_0243_),
    .Y(_0244_),
    .B1(net794));
 sg13g2_a21oi_1 _1711_ (.A1(_0237_),
    .A2(_0244_),
    .Y(_0245_),
    .B1(_0691_));
 sg13g2_o21ai_1 _1712_ (.B1(_0245_),
    .Y(_0246_),
    .A1(_0226_),
    .A2(_0232_));
 sg13g2_nand2b_1 _1713_ (.Y(_0247_),
    .B(net847),
    .A_N(\u_top_module.u_filter.shift_reg[205] ));
 sg13g2_nor2b_1 _1714_ (.A(net847),
    .B_N(\u_top_module.u_filter.shift_reg[204] ),
    .Y(_0248_));
 sg13g2_a221oi_1 _1715_ (.B2(net831),
    .C1(_0248_),
    .B1(_0247_),
    .A1(\u_top_module.u_filter.shift_reg[206] ),
    .Y(_0249_),
    .A2(net817));
 sg13g2_nor2_1 _1716_ (.A(\u_top_module.u_filter.shift_reg[207] ),
    .B(net827),
    .Y(_0250_));
 sg13g2_nor2_1 _1717_ (.A(net866),
    .B(\u_top_module.u_filter.shift_reg[201] ),
    .Y(_0251_));
 sg13g2_nor2_1 _1718_ (.A(net851),
    .B(\u_top_module.u_filter.shift_reg[200] ),
    .Y(_0252_));
 sg13g2_o21ai_1 _1719_ (.B1(net833),
    .Y(_0253_),
    .A1(_0251_),
    .A2(_0252_));
 sg13g2_nand2b_1 _1720_ (.Y(_0254_),
    .B(net837),
    .A_N(\u_top_module.u_filter.shift_reg[203] ));
 sg13g2_nand3b_1 _1721_ (.B(net866),
    .C(net851),
    .Y(_0255_),
    .A_N(\u_top_module.u_filter.shift_reg[202] ));
 sg13g2_nor2_1 _1722_ (.A(net864),
    .B(\u_top_module.u_filter.shift_reg[193] ),
    .Y(_0256_));
 sg13g2_nor2_1 _1723_ (.A(net850),
    .B(\u_top_module.u_filter.shift_reg[192] ),
    .Y(_0257_));
 sg13g2_o21ai_1 _1724_ (.B1(net827),
    .Y(_0258_),
    .A1(_0256_),
    .A2(_0257_));
 sg13g2_nand2b_1 _1725_ (.Y(_0259_),
    .B(net817),
    .A_N(\u_top_module.u_filter.shift_reg[194] ));
 sg13g2_nand2b_1 _1726_ (.Y(_0260_),
    .B(net836),
    .A_N(\u_top_module.u_filter.shift_reg[195] ));
 sg13g2_or4_1 _1727_ (.A(_0679_),
    .B(net803),
    .C(_0249_),
    .D(_0250_),
    .X(_0261_));
 sg13g2_and4_1 _1728_ (.A(net821),
    .B(net811),
    .C(_0254_),
    .D(_0255_),
    .X(_0262_));
 sg13g2_a21oi_1 _1729_ (.A1(_0253_),
    .A2(_0262_),
    .Y(_0263_),
    .B1(_0699_));
 sg13g2_nand4_1 _1730_ (.B(_0258_),
    .C(_0259_),
    .A(net803),
    .Y(_0264_),
    .D(_0260_));
 sg13g2_mux4_1 _1731_ (.S0(net864),
    .A0(\u_top_module.u_filter.shift_reg[199] ),
    .A1(\u_top_module.u_filter.shift_reg[196] ),
    .A2(\u_top_module.u_filter.shift_reg[197] ),
    .A3(\u_top_module.u_filter.shift_reg[198] ),
    .S1(net847),
    .X(_0265_));
 sg13g2_nand3_1 _1732_ (.B(net799),
    .C(_0265_),
    .A(net807),
    .Y(_0266_));
 sg13g2_nand3_1 _1733_ (.B(_0264_),
    .C(_0266_),
    .A(_0699_),
    .Y(_0267_));
 sg13g2_a21oi_1 _1734_ (.A1(_0261_),
    .A2(_0263_),
    .Y(_0268_),
    .B1(net797));
 sg13g2_a21oi_1 _1735_ (.A1(_0267_),
    .A2(_0268_),
    .Y(_0269_),
    .B1(_0717_));
 sg13g2_nand3_1 _1736_ (.B(\u_top_module.u_filter.shift_reg[239] ),
    .C(net808),
    .A(net830),
    .Y(_0270_));
 sg13g2_o21ai_1 _1737_ (.B1(net828),
    .Y(_0271_),
    .A1(\u_top_module.u_filter.shift_reg[238] ),
    .A2(net814));
 sg13g2_or2_1 _1738_ (.X(_0272_),
    .B(\u_top_module.u_filter.shift_reg[237] ),
    .A(net868));
 sg13g2_o21ai_1 _1739_ (.B1(_0272_),
    .Y(_0273_),
    .A1(net853),
    .A2(\u_top_module.u_filter.shift_reg[236] ));
 sg13g2_a221oi_1 _1740_ (.B2(net837),
    .C1(net804),
    .B1(_0273_),
    .A1(_0270_),
    .Y(_0274_),
    .A2(_0271_));
 sg13g2_nor2_1 _1741_ (.A(net869),
    .B(\u_top_module.u_filter.shift_reg[233] ),
    .Y(_0275_));
 sg13g2_nor2_1 _1742_ (.A(net853),
    .B(\u_top_module.u_filter.shift_reg[232] ),
    .Y(_0276_));
 sg13g2_o21ai_1 _1743_ (.B1(net826),
    .Y(_0277_),
    .A1(_0275_),
    .A2(_0276_));
 sg13g2_o21ai_1 _1744_ (.B1(net804),
    .Y(_0278_),
    .A1(net832),
    .A2(\u_top_module.u_filter.shift_reg[235] ));
 sg13g2_o21ai_1 _1745_ (.B1(_0277_),
    .Y(_0279_),
    .A1(\u_top_module.u_filter.shift_reg[234] ),
    .A2(net814));
 sg13g2_o21ai_1 _1746_ (.B1(net794),
    .Y(_0280_),
    .A1(_0278_),
    .A2(_0279_));
 sg13g2_nand2b_1 _1747_ (.Y(_0281_),
    .B(net854),
    .A_N(\u_top_module.u_filter.shift_reg[229] ));
 sg13g2_nor2b_1 _1748_ (.A(net853),
    .B_N(\u_top_module.u_filter.shift_reg[228] ),
    .Y(_0282_));
 sg13g2_a221oi_1 _1749_ (.B2(net830),
    .C1(_0282_),
    .B1(_0281_),
    .A1(\u_top_module.u_filter.shift_reg[230] ),
    .Y(_0283_),
    .A2(net817));
 sg13g2_nand2_1 _1750_ (.Y(_0284_),
    .A(\u_top_module.u_filter.shift_reg[231] ),
    .B(_0674_));
 sg13g2_a21o_1 _1751_ (.A2(_0284_),
    .A1(net810),
    .B1(_0283_),
    .X(_0285_));
 sg13g2_nor2_1 _1752_ (.A(net868),
    .B(\u_top_module.u_filter.shift_reg[225] ),
    .Y(_0286_));
 sg13g2_nor2_1 _1753_ (.A(net853),
    .B(\u_top_module.u_filter.shift_reg[224] ),
    .Y(_0287_));
 sg13g2_o21ai_1 _1754_ (.B1(net826),
    .Y(_0288_),
    .A1(_0286_),
    .A2(_0287_));
 sg13g2_nand2b_1 _1755_ (.Y(_0289_),
    .B(net837),
    .A_N(\u_top_module.u_filter.shift_reg[227] ));
 sg13g2_nand3b_1 _1756_ (.B(net868),
    .C(net853),
    .Y(_0290_),
    .A_N(\u_top_module.u_filter.shift_reg[226] ));
 sg13g2_and4_1 _1757_ (.A(net821),
    .B(net810),
    .C(_0289_),
    .D(_0290_),
    .X(_0291_));
 sg13g2_a21oi_1 _1758_ (.A1(_0288_),
    .A2(_0291_),
    .Y(_0292_),
    .B1(net794));
 sg13g2_a21oi_1 _1759_ (.A1(_0285_),
    .A2(_0292_),
    .Y(_0293_),
    .B1(net797));
 sg13g2_o21ai_1 _1760_ (.B1(_0293_),
    .Y(_0294_),
    .A1(_0274_),
    .A2(_0280_));
 sg13g2_nor2_1 _1761_ (.A(net849),
    .B(\u_top_module.u_filter.shift_reg[252] ),
    .Y(_0295_));
 sg13g2_nor2_1 _1762_ (.A(net865),
    .B(\u_top_module.u_filter.shift_reg[253] ),
    .Y(_0296_));
 sg13g2_nor4_1 _1763_ (.A(net829),
    .B(net817),
    .C(_0295_),
    .D(_0296_),
    .Y(_0297_));
 sg13g2_and2_1 _1764_ (.A(\u_top_module.u_filter.shift_reg[254] ),
    .B(net817),
    .X(_0298_));
 sg13g2_o21ai_1 _1765_ (.B1(net799),
    .Y(_0299_),
    .A1(_0297_),
    .A2(_0298_));
 sg13g2_nand2b_1 _1766_ (.Y(_0300_),
    .B(net817),
    .A_N(\u_top_module.u_filter.shift_reg[250] ));
 sg13g2_nor2_1 _1767_ (.A(net863),
    .B(\u_top_module.u_filter.shift_reg[249] ),
    .Y(_0301_));
 sg13g2_nor2_1 _1768_ (.A(net848),
    .B(\u_top_module.u_filter.shift_reg[248] ),
    .Y(_0302_));
 sg13g2_o21ai_1 _1769_ (.B1(net827),
    .Y(_0303_),
    .A1(_0301_),
    .A2(_0302_));
 sg13g2_nand2b_1 _1770_ (.Y(_0304_),
    .B(net836),
    .A_N(\u_top_module.u_filter.shift_reg[251] ));
 sg13g2_nand4_1 _1771_ (.B(_0300_),
    .C(_0303_),
    .A(net803),
    .Y(_0305_),
    .D(_0304_));
 sg13g2_nand3_1 _1772_ (.B(_0299_),
    .C(_0305_),
    .A(net795),
    .Y(_0306_));
 sg13g2_and2_1 _1773_ (.A(\u_top_module.u_filter.shift_reg[247] ),
    .B(_0674_),
    .X(_0307_));
 sg13g2_nor2_1 _1774_ (.A(net863),
    .B(\u_top_module.u_filter.shift_reg[245] ),
    .Y(_0308_));
 sg13g2_nor2_1 _1775_ (.A(net849),
    .B(\u_top_module.u_filter.shift_reg[244] ),
    .Y(_0309_));
 sg13g2_nor3_1 _1776_ (.A(net810),
    .B(_0308_),
    .C(_0309_),
    .Y(_0310_));
 sg13g2_nand2b_1 _1777_ (.Y(_0311_),
    .B(net817),
    .A_N(\u_top_module.u_filter.shift_reg[246] ));
 sg13g2_o21ai_1 _1778_ (.B1(_0311_),
    .Y(_0312_),
    .A1(_0307_),
    .A2(_0310_));
 sg13g2_nor2_1 _1779_ (.A(net868),
    .B(\u_top_module.u_filter.shift_reg[241] ),
    .Y(_0313_));
 sg13g2_nor2_1 _1780_ (.A(net854),
    .B(\u_top_module.u_filter.shift_reg[240] ),
    .Y(_0314_));
 sg13g2_o21ai_1 _1781_ (.B1(net826),
    .Y(_0315_),
    .A1(_0313_),
    .A2(_0314_));
 sg13g2_nand2b_1 _1782_ (.Y(_0316_),
    .B(net837),
    .A_N(\u_top_module.u_filter.shift_reg[243] ));
 sg13g2_nand3b_1 _1783_ (.B(net868),
    .C(net854),
    .Y(_0317_),
    .A_N(\u_top_module.u_filter.shift_reg[242] ));
 sg13g2_and4_1 _1784_ (.A(net821),
    .B(net810),
    .C(_0316_),
    .D(_0317_),
    .X(_0318_));
 sg13g2_a21oi_1 _1785_ (.A1(_0315_),
    .A2(_0318_),
    .Y(_0319_),
    .B1(net794));
 sg13g2_a21oi_1 _1786_ (.A1(_0312_),
    .A2(_0319_),
    .Y(_0320_),
    .B1(_0691_));
 sg13g2_a21oi_1 _1787_ (.A1(_0306_),
    .A2(_0320_),
    .Y(_0321_),
    .B1(_0716_));
 sg13g2_a22oi_1 _1788_ (.Y(_0322_),
    .B1(_0294_),
    .B2(_0321_),
    .A2(_0269_),
    .A1(_0246_));
 sg13g2_nand2_1 _1789_ (.Y(_0323_),
    .A(\u_top_module.filter_length[7] ),
    .B(_0741_));
 sg13g2_nand2_1 _1790_ (.Y(_0324_),
    .A(net807),
    .B(_0323_));
 sg13g2_a221oi_1 _1791_ (.B2(net807),
    .C1(_0221_),
    .B1(_0323_),
    .A1(_0743_),
    .Y(_0325_),
    .A2(_0322_));
 sg13g2_nand3_1 _1792_ (.B(\u_top_module.u_filter.shift_reg[79] ),
    .C(net806),
    .A(net830),
    .Y(_0326_));
 sg13g2_o21ai_1 _1793_ (.B1(net825),
    .Y(_0327_),
    .A1(\u_top_module.u_filter.shift_reg[78] ),
    .A2(net813));
 sg13g2_or2_1 _1794_ (.X(_0328_),
    .B(\u_top_module.u_filter.shift_reg[76] ),
    .A(net845));
 sg13g2_o21ai_1 _1795_ (.B1(_0328_),
    .Y(_0329_),
    .A1(net861),
    .A2(\u_top_module.u_filter.shift_reg[77] ));
 sg13g2_a221oi_1 _1796_ (.B2(net820),
    .C1(net802),
    .B1(_0329_),
    .A1(_0326_),
    .Y(_0330_),
    .A2(_0327_));
 sg13g2_nor2_1 _1797_ (.A(net860),
    .B(\u_top_module.u_filter.shift_reg[73] ),
    .Y(_0331_));
 sg13g2_nor2_1 _1798_ (.A(net848),
    .B(\u_top_module.u_filter.shift_reg[72] ),
    .Y(_0332_));
 sg13g2_o21ai_1 _1799_ (.B1(net825),
    .Y(_0333_),
    .A1(_0331_),
    .A2(_0332_));
 sg13g2_o21ai_1 _1800_ (.B1(_0333_),
    .Y(_0334_),
    .A1(\u_top_module.u_filter.shift_reg[74] ),
    .A2(net814));
 sg13g2_o21ai_1 _1801_ (.B1(net802),
    .Y(_0335_),
    .A1(net832),
    .A2(\u_top_module.u_filter.shift_reg[75] ));
 sg13g2_o21ai_1 _1802_ (.B1(net793),
    .Y(_0336_),
    .A1(_0334_),
    .A2(_0335_));
 sg13g2_a21o_1 _1803_ (.A2(\u_top_module.u_filter.shift_reg[69] ),
    .A1(net848),
    .B1(net863),
    .X(_0337_));
 sg13g2_or2_1 _1804_ (.X(_0338_),
    .B(\u_top_module.u_filter.shift_reg[68] ),
    .A(net848));
 sg13g2_a22oi_1 _1805_ (.Y(_0339_),
    .B1(_0337_),
    .B2(_0338_),
    .A2(net829),
    .A1(\u_top_module.u_filter.shift_reg[71] ));
 sg13g2_nor2_1 _1806_ (.A(\u_top_module.u_filter.shift_reg[70] ),
    .B(net814),
    .Y(_0340_));
 sg13g2_or3_1 _1807_ (.A(net803),
    .B(_0339_),
    .C(_0340_),
    .X(_0341_));
 sg13g2_nor2_1 _1808_ (.A(net863),
    .B(\u_top_module.u_filter.shift_reg[65] ),
    .Y(_0342_));
 sg13g2_nor2_1 _1809_ (.A(net848),
    .B(\u_top_module.u_filter.shift_reg[64] ),
    .Y(_0343_));
 sg13g2_o21ai_1 _1810_ (.B1(net827),
    .Y(_0344_),
    .A1(_0342_),
    .A2(_0343_));
 sg13g2_nand3b_1 _1811_ (.B(net863),
    .C(net848),
    .Y(_0345_),
    .A_N(\u_top_module.u_filter.shift_reg[66] ));
 sg13g2_nand2b_1 _1812_ (.Y(_0346_),
    .B(net836),
    .A_N(\u_top_module.u_filter.shift_reg[67] ));
 sg13g2_and4_1 _1813_ (.A(net822),
    .B(net810),
    .C(_0345_),
    .D(_0346_),
    .X(_0347_));
 sg13g2_a21oi_1 _1814_ (.A1(_0344_),
    .A2(_0347_),
    .Y(_0348_),
    .B1(net795));
 sg13g2_a21oi_1 _1815_ (.A1(_0341_),
    .A2(_0348_),
    .Y(_0349_),
    .B1(_0692_));
 sg13g2_o21ai_1 _1816_ (.B1(_0349_),
    .Y(_0350_),
    .A1(_0330_),
    .A2(_0336_));
 sg13g2_nand3_1 _1817_ (.B(\u_top_module.u_filter.shift_reg[95] ),
    .C(net805),
    .A(net830),
    .Y(_0351_));
 sg13g2_o21ai_1 _1818_ (.B1(net823),
    .Y(_0352_),
    .A1(\u_top_module.u_filter.shift_reg[94] ),
    .A2(net813));
 sg13g2_or2_1 _1819_ (.X(_0353_),
    .B(\u_top_module.u_filter.shift_reg[93] ),
    .A(net860));
 sg13g2_o21ai_1 _1820_ (.B1(_0353_),
    .Y(_0354_),
    .A1(net844),
    .A2(\u_top_module.u_filter.shift_reg[92] ));
 sg13g2_a221oi_1 _1821_ (.B2(net819),
    .C1(net801),
    .B1(_0354_),
    .A1(_0351_),
    .Y(_0355_),
    .A2(_0352_));
 sg13g2_nor2_1 _1822_ (.A(net858),
    .B(\u_top_module.u_filter.shift_reg[89] ),
    .Y(_0356_));
 sg13g2_nor2_1 _1823_ (.A(net841),
    .B(\u_top_module.u_filter.shift_reg[88] ),
    .Y(_0357_));
 sg13g2_o21ai_1 _1824_ (.B1(net824),
    .Y(_0358_),
    .A1(_0356_),
    .A2(_0357_));
 sg13g2_o21ai_1 _1825_ (.B1(net801),
    .Y(_0359_),
    .A1(net832),
    .A2(\u_top_module.u_filter.shift_reg[91] ));
 sg13g2_o21ai_1 _1826_ (.B1(_0358_),
    .Y(_0360_),
    .A1(\u_top_module.u_filter.shift_reg[90] ),
    .A2(net812));
 sg13g2_o21ai_1 _1827_ (.B1(net793),
    .Y(_0361_),
    .A1(_0359_),
    .A2(_0360_));
 sg13g2_a21o_1 _1828_ (.A2(\u_top_module.u_filter.shift_reg[85] ),
    .A1(net844),
    .B1(net860),
    .X(_0362_));
 sg13g2_or2_1 _1829_ (.X(_0363_),
    .B(\u_top_module.u_filter.shift_reg[84] ),
    .A(net844));
 sg13g2_a22oi_1 _1830_ (.Y(_0364_),
    .B1(_0362_),
    .B2(_0363_),
    .A2(net829),
    .A1(\u_top_module.u_filter.shift_reg[87] ));
 sg13g2_nor2_1 _1831_ (.A(\u_top_module.u_filter.shift_reg[86] ),
    .B(net813),
    .Y(_0365_));
 sg13g2_or3_1 _1832_ (.A(net802),
    .B(_0364_),
    .C(_0365_),
    .X(_0366_));
 sg13g2_nor2_1 _1833_ (.A(net860),
    .B(\u_top_module.u_filter.shift_reg[81] ),
    .Y(_0367_));
 sg13g2_nor2_1 _1834_ (.A(net845),
    .B(\u_top_module.u_filter.shift_reg[80] ),
    .Y(_0368_));
 sg13g2_o21ai_1 _1835_ (.B1(net825),
    .Y(_0369_),
    .A1(_0367_),
    .A2(_0368_));
 sg13g2_nand3b_1 _1836_ (.B(net860),
    .C(net844),
    .Y(_0370_),
    .A_N(\u_top_module.u_filter.shift_reg[82] ));
 sg13g2_nand2b_1 _1837_ (.Y(_0371_),
    .B(net835),
    .A_N(\u_top_module.u_filter.shift_reg[83] ));
 sg13g2_and4_1 _1838_ (.A(net820),
    .B(net811),
    .C(_0370_),
    .D(_0371_),
    .X(_0372_));
 sg13g2_a21oi_1 _1839_ (.A1(_0369_),
    .A2(_0372_),
    .Y(_0373_),
    .B1(net796));
 sg13g2_a21oi_1 _1840_ (.A1(_0366_),
    .A2(_0373_),
    .Y(_0374_),
    .B1(_0691_));
 sg13g2_o21ai_1 _1841_ (.B1(_0374_),
    .Y(_0375_),
    .A1(_0355_),
    .A2(_0361_));
 sg13g2_nand3_1 _1842_ (.B(_0350_),
    .C(_0375_),
    .A(_0716_),
    .Y(_0376_));
 sg13g2_nand3_1 _1843_ (.B(\u_top_module.u_filter.shift_reg[127] ),
    .C(net805),
    .A(net830),
    .Y(_0377_));
 sg13g2_o21ai_1 _1844_ (.B1(net823),
    .Y(_0378_),
    .A1(\u_top_module.u_filter.shift_reg[126] ),
    .A2(net812));
 sg13g2_or2_1 _1845_ (.X(_0379_),
    .B(\u_top_module.u_filter.shift_reg[125] ),
    .A(net858));
 sg13g2_o21ai_1 _1846_ (.B1(_0379_),
    .Y(_0380_),
    .A1(net842),
    .A2(\u_top_module.u_filter.shift_reg[124] ));
 sg13g2_a221oi_1 _1847_ (.B2(net819),
    .C1(net800),
    .B1(_0380_),
    .A1(_0377_),
    .Y(_0381_),
    .A2(_0378_));
 sg13g2_nor2_1 _1848_ (.A(net856),
    .B(\u_top_module.u_filter.shift_reg[121] ),
    .Y(_0382_));
 sg13g2_nor2_1 _1849_ (.A(net839),
    .B(\u_top_module.u_filter.shift_reg[120] ),
    .Y(_0383_));
 sg13g2_o21ai_1 _1850_ (.B1(net823),
    .Y(_0384_),
    .A1(_0382_),
    .A2(_0383_));
 sg13g2_o21ai_1 _1851_ (.B1(net800),
    .Y(_0385_),
    .A1(net832),
    .A2(\u_top_module.u_filter.shift_reg[123] ));
 sg13g2_o21ai_1 _1852_ (.B1(_0384_),
    .Y(_0386_),
    .A1(\u_top_module.u_filter.shift_reg[122] ),
    .A2(net812));
 sg13g2_o21ai_1 _1853_ (.B1(net793),
    .Y(_0387_),
    .A1(_0385_),
    .A2(_0386_));
 sg13g2_a21o_1 _1854_ (.A2(\u_top_module.u_filter.shift_reg[117] ),
    .A1(net839),
    .B1(net856),
    .X(_0388_));
 sg13g2_or2_1 _1855_ (.X(_0389_),
    .B(\u_top_module.u_filter.shift_reg[116] ),
    .A(net839));
 sg13g2_a22oi_1 _1856_ (.Y(_0390_),
    .B1(_0388_),
    .B2(_0389_),
    .A2(net829),
    .A1(\u_top_module.u_filter.shift_reg[119] ));
 sg13g2_nor2_1 _1857_ (.A(\u_top_module.u_filter.shift_reg[118] ),
    .B(net812),
    .Y(_0391_));
 sg13g2_or3_1 _1858_ (.A(net800),
    .B(_0390_),
    .C(_0391_),
    .X(_0392_));
 sg13g2_nor2_1 _1859_ (.A(net856),
    .B(\u_top_module.u_filter.shift_reg[113] ),
    .Y(_0393_));
 sg13g2_nor2_1 _1860_ (.A(net839),
    .B(\u_top_module.u_filter.shift_reg[112] ),
    .Y(_0394_));
 sg13g2_o21ai_1 _1861_ (.B1(net823),
    .Y(_0395_),
    .A1(_0393_),
    .A2(_0394_));
 sg13g2_nand3b_1 _1862_ (.B(net856),
    .C(net839),
    .Y(_0396_),
    .A_N(\u_top_module.u_filter.shift_reg[114] ));
 sg13g2_nand2b_1 _1863_ (.Y(_0397_),
    .B(net834),
    .A_N(\u_top_module.u_filter.shift_reg[115] ));
 sg13g2_and4_1 _1864_ (.A(net819),
    .B(net809),
    .C(_0396_),
    .D(_0397_),
    .X(_0398_));
 sg13g2_a21oi_1 _1865_ (.A1(_0395_),
    .A2(_0398_),
    .Y(_0399_),
    .B1(net793));
 sg13g2_a21oi_1 _1866_ (.A1(_0392_),
    .A2(_0399_),
    .Y(_0400_),
    .B1(_0691_));
 sg13g2_o21ai_1 _1867_ (.B1(_0400_),
    .Y(_0401_),
    .A1(_0381_),
    .A2(_0387_));
 sg13g2_nor2_1 _1868_ (.A(net859),
    .B(\u_top_module.u_filter.shift_reg[97] ),
    .Y(_0402_));
 sg13g2_nor2_1 _1869_ (.A(net843),
    .B(\u_top_module.u_filter.shift_reg[96] ),
    .Y(_0403_));
 sg13g2_o21ai_1 _1870_ (.B1(net825),
    .Y(_0404_),
    .A1(_0402_),
    .A2(_0403_));
 sg13g2_nand3b_1 _1871_ (.B(net859),
    .C(net843),
    .Y(_0405_),
    .A_N(\u_top_module.u_filter.shift_reg[98] ));
 sg13g2_nand2b_1 _1872_ (.Y(_0406_),
    .B(net835),
    .A_N(\u_top_module.u_filter.shift_reg[99] ));
 sg13g2_and4_1 _1873_ (.A(net820),
    .B(net809),
    .C(_0405_),
    .D(_0406_),
    .X(_0407_));
 sg13g2_a21oi_1 _1874_ (.A1(_0404_),
    .A2(_0407_),
    .Y(_0408_),
    .B1(net796));
 sg13g2_mux4_1 _1875_ (.S0(net859),
    .A0(\u_top_module.u_filter.shift_reg[103] ),
    .A1(\u_top_module.u_filter.shift_reg[100] ),
    .A2(\u_top_module.u_filter.shift_reg[101] ),
    .A3(\u_top_module.u_filter.shift_reg[102] ),
    .S1(net843),
    .X(_0409_));
 sg13g2_nand3_1 _1876_ (.B(net798),
    .C(_0409_),
    .A(net805),
    .Y(_0410_));
 sg13g2_nor2_1 _1877_ (.A(net859),
    .B(\u_top_module.u_filter.shift_reg[105] ),
    .Y(_0411_));
 sg13g2_nor2_1 _1878_ (.A(net843),
    .B(\u_top_module.u_filter.shift_reg[104] ),
    .Y(_0412_));
 sg13g2_o21ai_1 _1879_ (.B1(net823),
    .Y(_0413_),
    .A1(_0411_),
    .A2(_0412_));
 sg13g2_nand2b_1 _1880_ (.Y(_0414_),
    .B(net834),
    .A_N(\u_top_module.u_filter.shift_reg[107] ));
 sg13g2_nand2b_1 _1881_ (.Y(_0415_),
    .B(net818),
    .A_N(\u_top_module.u_filter.shift_reg[106] ));
 sg13g2_nand4_1 _1882_ (.B(_0413_),
    .C(_0414_),
    .A(net801),
    .Y(_0416_),
    .D(_0415_));
 sg13g2_mux4_1 _1883_ (.S0(net858),
    .A0(\u_top_module.u_filter.shift_reg[111] ),
    .A1(\u_top_module.u_filter.shift_reg[108] ),
    .A2(\u_top_module.u_filter.shift_reg[109] ),
    .A3(\u_top_module.u_filter.shift_reg[110] ),
    .S1(net842),
    .X(_0417_));
 sg13g2_nand3_1 _1884_ (.B(net798),
    .C(_0417_),
    .A(net805),
    .Y(_0418_));
 sg13g2_nand3_1 _1885_ (.B(_0416_),
    .C(_0418_),
    .A(net793),
    .Y(_0419_));
 sg13g2_a21oi_1 _1886_ (.A1(_0408_),
    .A2(_0410_),
    .Y(_0420_),
    .B1(net797));
 sg13g2_a21oi_2 _1887_ (.B1(_0716_),
    .Y(_0421_),
    .A2(_0420_),
    .A1(_0419_));
 sg13g2_a22oi_1 _1888_ (.Y(_0422_),
    .B1(_0401_),
    .B2(_0421_),
    .A2(_0742_),
    .A1(_0741_));
 sg13g2_nand3_1 _1889_ (.B(\u_top_module.u_filter.shift_reg[31] ),
    .C(net808),
    .A(net831),
    .Y(_0423_));
 sg13g2_o21ai_1 _1890_ (.B1(net826),
    .Y(_0424_),
    .A1(\u_top_module.u_filter.shift_reg[30] ),
    .A2(net814));
 sg13g2_or2_1 _1891_ (.X(_0425_),
    .B(\u_top_module.u_filter.shift_reg[29] ),
    .A(net866));
 sg13g2_o21ai_1 _1892_ (.B1(_0425_),
    .Y(_0426_),
    .A1(net851),
    .A2(\u_top_module.u_filter.shift_reg[28] ));
 sg13g2_a221oi_1 _1893_ (.B2(net821),
    .C1(net804),
    .B1(_0426_),
    .A1(_0423_),
    .Y(_0427_),
    .A2(_0424_));
 sg13g2_nor2_1 _1894_ (.A(net866),
    .B(\u_top_module.u_filter.shift_reg[25] ),
    .Y(_0428_));
 sg13g2_nor2_1 _1895_ (.A(net851),
    .B(\u_top_module.u_filter.shift_reg[24] ),
    .Y(_0429_));
 sg13g2_o21ai_1 _1896_ (.B1(net826),
    .Y(_0430_),
    .A1(_0428_),
    .A2(_0429_));
 sg13g2_o21ai_1 _1897_ (.B1(net804),
    .Y(_0431_),
    .A1(net832),
    .A2(\u_top_module.u_filter.shift_reg[27] ));
 sg13g2_o21ai_1 _1898_ (.B1(_0430_),
    .Y(_0432_),
    .A1(\u_top_module.u_filter.shift_reg[26] ),
    .A2(net815));
 sg13g2_o21ai_1 _1899_ (.B1(net794),
    .Y(_0433_),
    .A1(_0431_),
    .A2(_0432_));
 sg13g2_a21o_1 _1900_ (.A2(\u_top_module.u_filter.shift_reg[21] ),
    .A1(net852),
    .B1(net867),
    .X(_0434_));
 sg13g2_or2_1 _1901_ (.X(_0435_),
    .B(\u_top_module.u_filter.shift_reg[20] ),
    .A(net852));
 sg13g2_a22oi_1 _1902_ (.Y(_0436_),
    .B1(_0434_),
    .B2(_0435_),
    .A2(net829),
    .A1(\u_top_module.u_filter.shift_reg[23] ));
 sg13g2_nor2_1 _1903_ (.A(\u_top_module.u_filter.shift_reg[22] ),
    .B(net815),
    .Y(_0437_));
 sg13g2_or3_1 _1904_ (.A(net804),
    .B(_0436_),
    .C(_0437_),
    .X(_0438_));
 sg13g2_nor2_1 _1905_ (.A(net867),
    .B(\u_top_module.u_filter.shift_reg[17] ),
    .Y(_0439_));
 sg13g2_nor2_1 _1906_ (.A(net852),
    .B(\u_top_module.u_filter.shift_reg[16] ),
    .Y(_0440_));
 sg13g2_o21ai_1 _1907_ (.B1(net826),
    .Y(_0441_),
    .A1(_0439_),
    .A2(_0440_));
 sg13g2_nand3b_1 _1908_ (.B(net867),
    .C(net852),
    .Y(_0442_),
    .A_N(\u_top_module.u_filter.shift_reg[18] ));
 sg13g2_nand2b_1 _1909_ (.Y(_0443_),
    .B(net837),
    .A_N(\u_top_module.u_filter.shift_reg[19] ));
 sg13g2_and4_1 _1910_ (.A(net821),
    .B(net810),
    .C(_0442_),
    .D(_0443_),
    .X(_0444_));
 sg13g2_a21oi_1 _1911_ (.A1(_0441_),
    .A2(_0444_),
    .Y(_0445_),
    .B1(net794));
 sg13g2_a21oi_1 _1912_ (.A1(_0438_),
    .A2(_0445_),
    .Y(_0446_),
    .B1(_0691_));
 sg13g2_o21ai_1 _1913_ (.B1(_0446_),
    .Y(_0447_),
    .A1(_0427_),
    .A2(_0433_));
 sg13g2_nor2_1 _1914_ (.A(net866),
    .B(\u_top_module.u_filter.shift_reg[1] ),
    .Y(_0448_));
 sg13g2_nor2_1 _1915_ (.A(net851),
    .B(\u_top_module.u_filter.shift_reg[0] ),
    .Y(_0449_));
 sg13g2_o21ai_1 _1916_ (.B1(net826),
    .Y(_0450_),
    .A1(_0448_),
    .A2(_0449_));
 sg13g2_nand3b_1 _1917_ (.B(net866),
    .C(net851),
    .Y(_0451_),
    .A_N(\u_top_module.u_filter.shift_reg[2] ));
 sg13g2_nand2b_1 _1918_ (.Y(_0452_),
    .B(net837),
    .A_N(\u_top_module.u_filter.shift_reg[3] ));
 sg13g2_and4_1 _1919_ (.A(net821),
    .B(net811),
    .C(_0451_),
    .D(_0452_),
    .X(_0453_));
 sg13g2_a21oi_2 _1920_ (.B1(net794),
    .Y(_0454_),
    .A2(_0453_),
    .A1(_0450_));
 sg13g2_mux4_1 _1921_ (.S0(net866),
    .A0(\u_top_module.u_filter.shift_reg[7] ),
    .A1(\u_top_module.u_filter.shift_reg[4] ),
    .A2(\u_top_module.u_filter.shift_reg[5] ),
    .A3(\u_top_module.u_filter.shift_reg[6] ),
    .S1(net851),
    .X(_0455_));
 sg13g2_nand3_1 _1922_ (.B(net799),
    .C(_0455_),
    .A(net807),
    .Y(_0456_));
 sg13g2_a21oi_1 _1923_ (.A1(_0454_),
    .A2(_0456_),
    .Y(_0457_),
    .B1(net797));
 sg13g2_nand2b_1 _1924_ (.Y(_0458_),
    .B(net817),
    .A_N(\u_top_module.u_filter.shift_reg[10] ));
 sg13g2_nand2b_1 _1925_ (.Y(_0459_),
    .B(net836),
    .A_N(\u_top_module.u_filter.shift_reg[11] ));
 sg13g2_nor2_1 _1926_ (.A(net866),
    .B(\u_top_module.u_filter.shift_reg[9] ),
    .Y(_0460_));
 sg13g2_nor2_1 _1927_ (.A(net851),
    .B(\u_top_module.u_filter.shift_reg[8] ),
    .Y(_0461_));
 sg13g2_o21ai_1 _1928_ (.B1(net826),
    .Y(_0462_),
    .A1(_0460_),
    .A2(_0461_));
 sg13g2_nand4_1 _1929_ (.B(_0458_),
    .C(_0459_),
    .A(net803),
    .Y(_0463_),
    .D(_0462_));
 sg13g2_mux4_1 _1930_ (.S0(net867),
    .A0(\u_top_module.u_filter.shift_reg[15] ),
    .A1(\u_top_module.u_filter.shift_reg[12] ),
    .A2(\u_top_module.u_filter.shift_reg[13] ),
    .A3(\u_top_module.u_filter.shift_reg[14] ),
    .S1(net853),
    .X(_0464_));
 sg13g2_nand3_1 _1931_ (.B(net798),
    .C(_0464_),
    .A(net808),
    .Y(_0465_));
 sg13g2_nand3_1 _1932_ (.B(_0463_),
    .C(_0465_),
    .A(net794),
    .Y(_0466_));
 sg13g2_a21oi_1 _1933_ (.A1(_0457_),
    .A2(_0466_),
    .Y(_0467_),
    .B1(_0717_));
 sg13g2_nand3_1 _1934_ (.B(\u_top_module.u_filter.shift_reg[63] ),
    .C(net807),
    .A(net831),
    .Y(_0468_));
 sg13g2_o21ai_1 _1935_ (.B1(net827),
    .Y(_0469_),
    .A1(\u_top_module.u_filter.shift_reg[62] ),
    .A2(net814));
 sg13g2_or2_1 _1936_ (.X(_0470_),
    .B(\u_top_module.u_filter.shift_reg[61] ),
    .A(net863));
 sg13g2_o21ai_1 _1937_ (.B1(_0470_),
    .Y(_0471_),
    .A1(net848),
    .A2(\u_top_module.u_filter.shift_reg[60] ));
 sg13g2_a221oi_1 _1938_ (.B2(net822),
    .C1(net803),
    .B1(_0471_),
    .A1(_0468_),
    .Y(_0472_),
    .A2(_0469_));
 sg13g2_nor2_1 _1939_ (.A(net864),
    .B(\u_top_module.u_filter.shift_reg[57] ),
    .Y(_0473_));
 sg13g2_nor2_1 _1940_ (.A(net847),
    .B(\u_top_module.u_filter.shift_reg[56] ),
    .Y(_0474_));
 sg13g2_o21ai_1 _1941_ (.B1(net827),
    .Y(_0475_),
    .A1(_0473_),
    .A2(_0474_));
 sg13g2_o21ai_1 _1942_ (.B1(net803),
    .Y(_0476_),
    .A1(net833),
    .A2(\u_top_module.u_filter.shift_reg[59] ));
 sg13g2_o21ai_1 _1943_ (.B1(_0475_),
    .Y(_0477_),
    .A1(\u_top_module.u_filter.shift_reg[58] ),
    .A2(net814));
 sg13g2_o21ai_1 _1944_ (.B1(net795),
    .Y(_0478_),
    .A1(_0476_),
    .A2(_0477_));
 sg13g2_nor2_1 _1945_ (.A(_0472_),
    .B(_0478_),
    .Y(_0479_));
 sg13g2_nor2_1 _1946_ (.A(net864),
    .B(\u_top_module.u_filter.shift_reg[49] ),
    .Y(_0480_));
 sg13g2_nor2_1 _1947_ (.A(net847),
    .B(\u_top_module.u_filter.shift_reg[48] ),
    .Y(_0481_));
 sg13g2_o21ai_1 _1948_ (.B1(net827),
    .Y(_0482_),
    .A1(_0480_),
    .A2(_0481_));
 sg13g2_o21ai_1 _1949_ (.B1(_0482_),
    .Y(_0483_),
    .A1(\u_top_module.u_filter.shift_reg[50] ),
    .A2(net814));
 sg13g2_o21ai_1 _1950_ (.B1(net803),
    .Y(_0484_),
    .A1(net833),
    .A2(\u_top_module.u_filter.shift_reg[51] ));
 sg13g2_mux4_1 _1951_ (.S0(net864),
    .A0(\u_top_module.u_filter.shift_reg[55] ),
    .A1(\u_top_module.u_filter.shift_reg[52] ),
    .A2(\u_top_module.u_filter.shift_reg[53] ),
    .A3(\u_top_module.u_filter.shift_reg[54] ),
    .S1(net847),
    .X(_0485_));
 sg13g2_nand3_1 _1952_ (.B(net799),
    .C(_0485_),
    .A(net807),
    .Y(_0486_));
 sg13g2_o21ai_1 _1953_ (.B1(_0486_),
    .Y(_0487_),
    .A1(_0483_),
    .A2(_0484_));
 sg13g2_o21ai_1 _1954_ (.B1(net797),
    .Y(_0488_),
    .A1(net795),
    .A2(_0487_));
 sg13g2_nor2_1 _1955_ (.A(net864),
    .B(\u_top_module.u_filter.shift_reg[33] ),
    .Y(_0489_));
 sg13g2_nor2_1 _1956_ (.A(net847),
    .B(\u_top_module.u_filter.shift_reg[32] ),
    .Y(_0490_));
 sg13g2_o21ai_1 _1957_ (.B1(net827),
    .Y(_0491_),
    .A1(_0489_),
    .A2(_0490_));
 sg13g2_nand3b_1 _1958_ (.B(net864),
    .C(net847),
    .Y(_0492_),
    .A_N(\u_top_module.u_filter.shift_reg[34] ));
 sg13g2_nand2b_1 _1959_ (.Y(_0493_),
    .B(net836),
    .A_N(\u_top_module.u_filter.shift_reg[35] ));
 sg13g2_and4_1 _1960_ (.A(net822),
    .B(net810),
    .C(_0492_),
    .D(_0493_),
    .X(_0494_));
 sg13g2_a21oi_1 _1961_ (.A1(_0491_),
    .A2(_0494_),
    .Y(_0495_),
    .B1(net795));
 sg13g2_mux4_1 _1962_ (.S0(net859),
    .A0(\u_top_module.u_filter.shift_reg[39] ),
    .A1(\u_top_module.u_filter.shift_reg[36] ),
    .A2(\u_top_module.u_filter.shift_reg[37] ),
    .A3(\u_top_module.u_filter.shift_reg[38] ),
    .S1(net843),
    .X(_0496_));
 sg13g2_nand3_1 _1963_ (.B(net798),
    .C(_0496_),
    .A(net806),
    .Y(_0497_));
 sg13g2_a21oi_1 _1964_ (.A1(_0495_),
    .A2(_0497_),
    .Y(_0498_),
    .B1(_0692_));
 sg13g2_nor2_1 _1965_ (.A(\u_top_module.u_filter.shift_reg[46] ),
    .B(net813),
    .Y(_0499_));
 sg13g2_a21o_1 _1966_ (.A2(\u_top_module.u_filter.shift_reg[45] ),
    .A1(net843),
    .B1(net859),
    .X(_0500_));
 sg13g2_or2_1 _1967_ (.X(_0501_),
    .B(\u_top_module.u_filter.shift_reg[44] ),
    .A(net846));
 sg13g2_a22oi_1 _1968_ (.Y(_0502_),
    .B1(_0500_),
    .B2(_0501_),
    .A2(_0672_),
    .A1(\u_top_module.u_filter.shift_reg[47] ));
 sg13g2_o21ai_1 _1969_ (.B1(net846),
    .Y(_0503_),
    .A1(net859),
    .A2(\u_top_module.u_filter.shift_reg[41] ));
 sg13g2_a22oi_1 _1970_ (.Y(_0504_),
    .B1(\u_top_module.u_filter.shift_reg[43] ),
    .B2(net829),
    .A2(\u_top_module.u_filter.shift_reg[40] ),
    .A1(net862));
 sg13g2_a221oi_1 _1971_ (.B2(_0504_),
    .C1(net798),
    .B1(_0503_),
    .A1(_0562_),
    .Y(_0505_),
    .A2(net818));
 sg13g2_nor4_1 _1972_ (.A(_0679_),
    .B(net802),
    .C(_0499_),
    .D(_0502_),
    .Y(_0506_));
 sg13g2_or3_1 _1973_ (.A(_0699_),
    .B(_0505_),
    .C(_0506_),
    .X(_0507_));
 sg13g2_a21oi_1 _1974_ (.A1(_0498_),
    .A2(_0507_),
    .Y(_0508_),
    .B1(_0716_));
 sg13g2_o21ai_1 _1975_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_0479_),
    .A2(_0488_));
 sg13g2_a21oi_1 _1976_ (.A1(_0447_),
    .A2(_0467_),
    .Y(_0510_),
    .B1(_0743_));
 sg13g2_a221oi_1 _1977_ (.B2(_0510_),
    .C1(_0324_),
    .B1(_0509_),
    .A1(_0376_),
    .Y(_0511_),
    .A2(_0422_));
 sg13g2_or3_2 _1978_ (.A(\u_top_module.u_i2s_bus.u_mux_shift.sum_res ),
    .B(_0325_),
    .C(_0511_),
    .X(_0512_));
 sg13g2_o21ai_1 _1979_ (.B1(\u_top_module.u_i2s_bus.u_mux_shift.sum_res ),
    .Y(_0513_),
    .A1(_0325_),
    .A2(_0511_));
 sg13g2_a21o_1 _1980_ (.A2(_0513_),
    .A1(_0512_),
    .B1(_0028_),
    .X(_0514_));
 sg13g2_nand3_1 _1981_ (.B(_0512_),
    .C(_0513_),
    .A(_0028_),
    .Y(_0515_));
 sg13g2_nand3_1 _1982_ (.B(_0514_),
    .C(_0515_),
    .A(net807),
    .Y(_0516_));
 sg13g2_o21ai_1 _1983_ (.B1(_0516_),
    .Y(_0162_),
    .A1(_0565_),
    .A2(net807));
 sg13g2_nand2_1 _1984_ (.Y(_0517_),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .B(_0679_));
 sg13g2_nand2b_1 _1985_ (.Y(_0518_),
    .B(_0512_),
    .A_N(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ));
 sg13g2_xor2_1 _1986_ (.B(_0512_),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .X(_0519_));
 sg13g2_xnor2_1 _1987_ (.Y(_0520_),
    .A(_0514_),
    .B(_0519_));
 sg13g2_o21ai_1 _1988_ (.B1(_0517_),
    .Y(_0163_),
    .A1(_0679_),
    .A2(_0520_));
 sg13g2_nor2_1 _1989_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .B(net806),
    .Y(_0521_));
 sg13g2_o21ai_1 _1990_ (.B1(_0518_),
    .Y(_0522_),
    .A1(_0514_),
    .A2(_0519_));
 sg13g2_nor2b_1 _1991_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .B_N(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .Y(_0523_));
 sg13g2_xnor2_1 _1992_ (.Y(_0524_),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .B(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ));
 sg13g2_xnor2_1 _1993_ (.Y(_0525_),
    .A(_0522_),
    .B(_0524_));
 sg13g2_a21oi_1 _1994_ (.A1(net806),
    .A2(_0525_),
    .Y(_0164_),
    .B1(_0521_));
 sg13g2_nand2_1 _1995_ (.Y(_0526_),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .B(_0679_));
 sg13g2_xnor2_1 _1996_ (.Y(_0527_),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .B(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ));
 sg13g2_a21o_1 _1997_ (.A2(_0524_),
    .A1(_0522_),
    .B1(_0523_),
    .X(_0528_));
 sg13g2_xnor2_1 _1998_ (.Y(_0529_),
    .A(_0527_),
    .B(_0528_));
 sg13g2_o21ai_1 _1999_ (.B1(_0526_),
    .Y(_0165_),
    .A1(_0679_),
    .A2(_0529_));
 sg13g2_xor2_1 _2000_ (.B(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .X(_0530_));
 sg13g2_nand3_1 _2001_ (.B(_0524_),
    .C(_0527_),
    .A(_0522_),
    .Y(_0531_));
 sg13g2_o21ai_1 _2002_ (.B1(_0556_),
    .Y(_0532_),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .A2(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ));
 sg13g2_nand3_1 _2003_ (.B(_0531_),
    .C(_0532_),
    .A(_0530_),
    .Y(_0533_));
 sg13g2_a21o_1 _2004_ (.A2(_0532_),
    .A1(_0531_),
    .B1(_0530_),
    .X(_0534_));
 sg13g2_nand3_1 _2005_ (.B(_0533_),
    .C(_0534_),
    .A(net806),
    .Y(_0535_));
 sg13g2_o21ai_1 _2006_ (.B1(_0535_),
    .Y(_0166_),
    .A1(_0557_),
    .A2(net806));
 sg13g2_xor2_1 _2007_ (.B(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .X(_0536_));
 sg13g2_o21ai_1 _2008_ (.B1(_0534_),
    .Y(_0537_),
    .A1(_0556_),
    .A2(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ));
 sg13g2_xnor2_1 _2009_ (.Y(_0538_),
    .A(_0536_),
    .B(_0537_));
 sg13g2_nor2_1 _2010_ (.A(_0679_),
    .B(_0538_),
    .Y(_0539_));
 sg13g2_a21oi_1 _2011_ (.A1(_0558_),
    .A2(_0679_),
    .Y(_0167_),
    .B1(_0539_));
 sg13g2_o21ai_1 _2012_ (.B1(_0558_),
    .Y(_0540_),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .A2(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ));
 sg13g2_o21ai_1 _2013_ (.B1(_0540_),
    .Y(_0541_),
    .A1(_0534_),
    .A2(_0536_));
 sg13g2_o21ai_1 _2014_ (.B1(net805),
    .Y(_0542_),
    .A1(_0558_),
    .A2(_0541_));
 sg13g2_a21oi_1 _2015_ (.A1(_0558_),
    .A2(_0541_),
    .Y(_0543_),
    .B1(_0542_));
 sg13g2_xor2_1 _2016_ (.B(_0543_),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .X(_0168_));
 sg13g2_mux2_1 _2017_ (.A0(_0541_),
    .A1(_0558_),
    .S(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .X(_0544_));
 sg13g2_nor2_1 _2018_ (.A(_0542_),
    .B(_0544_),
    .Y(_0545_));
 sg13g2_xor2_1 _2019_ (.B(_0545_),
    .A(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .X(_0169_));
 sg13g2_and2_1 _2020_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.out ),
    .B(net889),
    .X(_0171_));
 sg13g2_and2_1 _2021_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.out ),
    .B(net892),
    .X(_0172_));
 sg13g2_and2_1 _2022_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.out ),
    .B(net889),
    .X(_0173_));
 sg13g2_mux2_1 _2023_ (.A0(\u_top_module.u_i2s_bus.dec_clk ),
    .A1(_0019_),
    .S(_0629_),
    .X(_0174_));
 sg13g2_and2_1 _2024_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ),
    .B(net889),
    .X(_0175_));
 sg13g2_and2_1 _2025_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.out ),
    .B(net890),
    .X(_0176_));
 sg13g2_and2_1 _2026_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.out ),
    .B(net890),
    .X(_0177_));
 sg13g2_and2_1 _2027_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.out ),
    .B(net889),
    .X(_0178_));
 sg13g2_and2_1 _2028_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.out ),
    .B(net888),
    .X(_0179_));
 sg13g2_and2_1 _2029_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.out ),
    .B(net888),
    .X(_0180_));
 sg13g2_and2_1 _2030_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.out ),
    .B(net888),
    .X(_0181_));
 sg13g2_and2_1 _2031_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.out ),
    .B(net887),
    .X(_0182_));
 sg13g2_and2_1 _2032_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.out ),
    .B(net887),
    .X(_0183_));
 sg13g2_and2_1 _2033_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.out ),
    .B(net887),
    .X(_0184_));
 sg13g2_and2_1 _2034_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.out ),
    .B(net887),
    .X(_0185_));
 sg13g2_and2_1 _2035_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.out ),
    .B(net887),
    .X(_0186_));
 sg13g2_and2_1 _2036_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.out ),
    .B(net887),
    .X(_0187_));
 sg13g2_and2_1 _2037_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.out ),
    .B(net887),
    .X(_0188_));
 sg13g2_and2_1 _2038_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.out ),
    .B(net887),
    .X(_0189_));
 sg13g2_and2_1 _2039_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.out ),
    .B(net888),
    .X(_0190_));
 sg13g2_and2_1 _2040_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.out ),
    .B(net888),
    .X(_0191_));
 sg13g2_and2_1 _2041_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.out ),
    .B(net888),
    .X(_0192_));
 sg13g2_and2_1 _2042_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.out ),
    .B(net891),
    .X(_0193_));
 sg13g2_and2_1 _2043_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.out ),
    .B(net891),
    .X(_0194_));
 sg13g2_and2_1 _2044_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.out ),
    .B(net891),
    .X(_0195_));
 sg13g2_mux2_1 _2045_ (.A0(net931),
    .A1(_0010_),
    .S(net792),
    .X(_0196_));
 sg13g2_inv_1 _2046_ (.Y(_0032_),
    .A(net964));
 sg13g2_inv_1 _2047_ (.Y(_0033_),
    .A(net965));
 sg13g2_inv_1 _2048_ (.Y(_0034_),
    .A(net965));
 sg13g2_inv_1 _2049_ (.Y(_0035_),
    .A(net958));
 sg13g2_inv_1 _2050_ (.Y(_0036_),
    .A(net958));
 sg13g2_inv_1 _2051_ (.Y(_0037_),
    .A(net957));
 sg13g2_inv_1 _2052_ (.Y(_0038_),
    .A(net957));
 sg13g2_inv_1 _2053_ (.Y(_0039_),
    .A(net956));
 sg13g2_inv_1 _2054_ (.Y(_0040_),
    .A(net956));
 sg13g2_inv_1 _2055_ (.Y(_0041_),
    .A(net956));
 sg13g2_inv_1 _2056_ (.Y(_0042_),
    .A(net957));
 sg13g2_inv_1 _2057_ (.Y(_0043_),
    .A(net958));
 sg13g2_inv_1 _2058_ (.Y(_0044_),
    .A(net958));
 sg13g2_inv_1 _2059_ (.Y(_0045_),
    .A(net953));
 sg13g2_inv_1 _2060_ (.Y(_0046_),
    .A(net953));
 sg13g2_inv_1 _2061_ (.Y(_0047_),
    .A(net953));
 sg13g2_inv_1 _2062_ (.Y(_0048_),
    .A(net952));
 sg13g2_inv_1 _2063_ (.Y(_0049_),
    .A(net955));
 sg13g2_inv_1 _2064_ (.Y(_0050_),
    .A(net955));
 sg13g2_inv_1 _2065_ (.Y(_0051_),
    .A(net955));
 sg13g2_inv_1 _2066_ (.Y(_0052_),
    .A(net951));
 sg13g2_inv_1 _2067_ (.Y(_0053_),
    .A(net951));
 sg13g2_inv_1 _2068_ (.Y(_0054_),
    .A(net951));
 sg13g2_inv_1 _2069_ (.Y(_0055_),
    .A(net952));
 sg13g2_inv_1 _2070_ (.Y(_0056_),
    .A(net952));
 sg13g2_inv_1 _2071_ (.Y(_0057_),
    .A(net954));
 sg13g2_inv_1 _2072_ (.Y(_0058_),
    .A(net953));
 sg13g2_inv_1 _2073_ (.Y(_0059_),
    .A(net955));
 sg13g2_inv_1 _2074_ (.Y(_0060_),
    .A(net965));
 sg13g2_inv_1 _2075_ (.Y(_0061_),
    .A(net965));
 sg13g2_inv_1 _2076_ (.Y(_0062_),
    .A(net963));
 sg13g2_inv_1 _2077_ (.Y(_0063_),
    .A(net971));
 sg13g2_dfrbp_1 _2078_ (.CLK(net981),
    .RESET_B(net1026),
    .D(_0005_),
    .Q_N(_0937_),
    .Q(\u_top_module.u_decimator.counter[3] ));
 sg13g2_dfrbp_1 _2079_ (.CLK(net978),
    .RESET_B(net1026),
    .D(_0006_),
    .Q_N(_0938_),
    .Q(\u_top_module.u_decimator.counter[4] ));
 sg13g2_dfrbp_1 _2080_ (.CLK(net978),
    .RESET_B(net1038),
    .D(_0007_),
    .Q_N(_0939_),
    .Q(\u_top_module.u_decimator.counter[5] ));
 sg13g2_dfrbp_1 _2081_ (.CLK(net972),
    .RESET_B(net1038),
    .D(_0008_),
    .Q_N(_0940_),
    .Q(\u_top_module.u_decimator.counter[6] ));
 sg13g2_dfrbp_1 _2082_ (.CLK(net971),
    .RESET_B(net1038),
    .D(_0009_),
    .Q_N(_0936_),
    .Q(\u_top_module.u_decimator.counter[7] ));
 sg13g2_dfrbp_1 _2083_ (.CLK(net980),
    .RESET_B(net1039),
    .D(_0064_),
    .Q_N(_0028_),
    .Q(\u_top_module.dec_data ));
 sg13g2_dllrq_1 _2084_ (.D(\u_top_module.mem_out[0] ),
    .GATE_N(_0001_),
    .RESET_B(net27),
    .Q(\u_top_module.filter_length[0] ));
 sg13g2_dllrq_1 _2085_ (.D(\u_top_module.mem_out[1] ),
    .GATE_N(_0001_),
    .RESET_B(net28),
    .Q(\u_top_module.filter_length[1] ));
 sg13g2_dllrq_1 _2086_ (.D(\u_top_module.mem_out[2] ),
    .GATE_N(_0001_),
    .RESET_B(net29),
    .Q(\u_top_module.filter_length[2] ));
 sg13g2_dllrq_1 _2087_ (.D(\u_top_module.mem_out[3] ),
    .GATE_N(_0001_),
    .RESET_B(net30),
    .Q(\u_top_module.filter_length[3] ));
 sg13g2_dllrq_1 _2088_ (.D(\u_top_module.mem_out[4] ),
    .GATE_N(_0001_),
    .RESET_B(net31),
    .Q(\u_top_module.filter_length[4] ));
 sg13g2_dllrq_1 _2089_ (.D(\u_top_module.mem_out[5] ),
    .GATE_N(_0001_),
    .RESET_B(net32),
    .Q(\u_top_module.filter_length[5] ));
 sg13g2_dllrq_1 _2090_ (.D(\u_top_module.mem_out[6] ),
    .GATE_N(_0001_),
    .RESET_B(net33),
    .Q(\u_top_module.filter_length[6] ));
 sg13g2_dllrq_1 _2091_ (.D(\u_top_module.mem_out[7] ),
    .GATE_N(_0001_),
    .RESET_B(net34),
    .Q(\u_top_module.filter_length[7] ));
 sg13g2_dllrq_1 _2092_ (.D(\u_top_module.mem_out[0] ),
    .GATE_N(_0000_),
    .RESET_B(net35),
    .Q(\u_top_module.decimation_ratio[0] ));
 sg13g2_dllrq_1 _2093_ (.D(\u_top_module.mem_out[1] ),
    .GATE_N(_0000_),
    .RESET_B(net36),
    .Q(\u_top_module.decimation_ratio[1] ));
 sg13g2_dllrq_1 _2094_ (.D(\u_top_module.mem_out[2] ),
    .GATE_N(_0000_),
    .RESET_B(net37),
    .Q(\u_top_module.decimation_ratio[2] ));
 sg13g2_dllrq_1 _2095_ (.D(\u_top_module.mem_out[3] ),
    .GATE_N(_0000_),
    .RESET_B(net38),
    .Q(\u_top_module.decimation_ratio[3] ));
 sg13g2_dllrq_1 _2096_ (.D(\u_top_module.mem_out[4] ),
    .GATE_N(_0000_),
    .RESET_B(net39),
    .Q(\u_top_module.decimation_ratio[4] ));
 sg13g2_dllrq_1 _2097_ (.D(\u_top_module.mem_out[5] ),
    .GATE_N(_0000_),
    .RESET_B(net40),
    .Q(\u_top_module.decimation_ratio[5] ));
 sg13g2_dllrq_1 _2098_ (.D(\u_top_module.mem_out[6] ),
    .GATE_N(_0000_),
    .RESET_B(net41),
    .Q(\u_top_module.decimation_ratio[6] ));
 sg13g2_dllrq_1 _2099_ (.D(\u_top_module.mem_out[7] ),
    .GATE_N(_0000_),
    .RESET_B(net42),
    .Q(\u_top_module.decimation_ratio[7] ));
 sg13g2_dfrbp_1 _2100_ (.CLK(net972),
    .RESET_B(net43),
    .D(_0197_),
    .Q_N(_0941_),
    .Q(\u_top_module.mem_out[0] ));
 sg13g2_dfrbp_1 _2101_ (.CLK(net971),
    .RESET_B(net44),
    .D(_0198_),
    .Q_N(_0942_),
    .Q(\u_top_module.mem_out[1] ));
 sg13g2_dfrbp_1 _2102_ (.CLK(net978),
    .RESET_B(net45),
    .D(_0199_),
    .Q_N(_0943_),
    .Q(\u_top_module.mem_out[2] ));
 sg13g2_dfrbp_1 _2103_ (.CLK(net971),
    .RESET_B(net46),
    .D(_0200_),
    .Q_N(_0944_),
    .Q(\u_top_module.mem_out[3] ));
 sg13g2_dfrbp_1 _2104_ (.CLK(net971),
    .RESET_B(net47),
    .D(_0201_),
    .Q_N(_0945_),
    .Q(\u_top_module.mem_out[4] ));
 sg13g2_dfrbp_1 _2105_ (.CLK(net972),
    .RESET_B(net48),
    .D(_0202_),
    .Q_N(_0946_),
    .Q(\u_top_module.mem_out[5] ));
 sg13g2_dfrbp_1 _2106_ (.CLK(net971),
    .RESET_B(net107),
    .D(_0203_),
    .Q_N(_0947_),
    .Q(\u_top_module.mem_out[6] ));
 sg13g2_dfrbp_1 _2107_ (.CLK(net971),
    .RESET_B(net50),
    .D(_0204_),
    .Q_N(_0935_),
    .Q(\u_top_module.mem_out[7] ));
 sg13g2_dfrbp_1 _2108_ (.CLK(net964),
    .RESET_B(net49),
    .D(_0065_),
    .Q_N(_0934_),
    .Q(\u_top_module.u_i2s_bus.u_mux_shift.data ));
 sg13g2_dfrbp_1 _2109_ (.CLK(net972),
    .RESET_B(net1026),
    .D(_0066_),
    .Q_N(_0933_),
    .Q(\u_top_module.u_memory.memory[0][0] ));
 sg13g2_dfrbp_1 _2110_ (.CLK(net971),
    .RESET_B(net1017),
    .D(_0067_),
    .Q_N(_0932_),
    .Q(\u_top_module.u_memory.memory[0][1] ));
 sg13g2_dfrbp_1 _2111_ (.CLK(net974),
    .RESET_B(net1019),
    .D(_0068_),
    .Q_N(_0931_),
    .Q(\u_top_module.u_memory.memory[0][2] ));
 sg13g2_dfrbp_1 _2112_ (.CLK(net967),
    .RESET_B(net1013),
    .D(_0069_),
    .Q_N(_0930_),
    .Q(\u_top_module.u_memory.memory[0][3] ));
 sg13g2_dfrbp_1 _2113_ (.CLK(net967),
    .RESET_B(net1013),
    .D(_0070_),
    .Q_N(_0929_),
    .Q(\u_top_module.u_memory.memory[0][4] ));
 sg13g2_dfrbp_1 _2114_ (.CLK(net968),
    .RESET_B(net1019),
    .D(_0071_),
    .Q_N(_0928_),
    .Q(\u_top_module.u_memory.memory[0][5] ));
 sg13g2_dfrbp_1 _2115_ (.CLK(net967),
    .RESET_B(net1016),
    .D(_0072_),
    .Q_N(_0927_),
    .Q(\u_top_module.u_memory.memory[0][6] ));
 sg13g2_dfrbp_1 _2116_ (.CLK(net970),
    .RESET_B(net1014),
    .D(_0073_),
    .Q_N(_0926_),
    .Q(\u_top_module.u_memory.memory[0][7] ));
 sg13g2_dfrbp_1 _2117_ (.CLK(net969),
    .RESET_B(net1018),
    .D(_0074_),
    .Q_N(_0925_),
    .Q(\u_top_module.u_memory.memory[1][0] ));
 sg13g2_dfrbp_1 _2118_ (.CLK(net961),
    .RESET_B(net1017),
    .D(_0075_),
    .Q_N(_0924_),
    .Q(\u_top_module.u_memory.memory[1][1] ));
 sg13g2_dfrbp_1 _2119_ (.CLK(net969),
    .RESET_B(net1019),
    .D(_0076_),
    .Q_N(_0923_),
    .Q(\u_top_module.u_memory.memory[1][2] ));
 sg13g2_dfrbp_1 _2120_ (.CLK(net961),
    .RESET_B(net1013),
    .D(_0077_),
    .Q_N(_0922_),
    .Q(\u_top_module.u_memory.memory[1][3] ));
 sg13g2_dfrbp_1 _2121_ (.CLK(net960),
    .RESET_B(net1012),
    .D(_0078_),
    .Q_N(_0921_),
    .Q(\u_top_module.u_memory.memory[1][4] ));
 sg13g2_dfrbp_1 _2122_ (.CLK(net968),
    .RESET_B(net1020),
    .D(_0079_),
    .Q_N(_0920_),
    .Q(\u_top_module.u_memory.memory[1][5] ));
 sg13g2_dfrbp_1 _2123_ (.CLK(net967),
    .RESET_B(net1015),
    .D(_0080_),
    .Q_N(_0919_),
    .Q(\u_top_module.u_memory.memory[1][6] ));
 sg13g2_dfrbp_1 _2124_ (.CLK(net959),
    .RESET_B(net1014),
    .D(_0081_),
    .Q_N(_0918_),
    .Q(\u_top_module.u_memory.memory[1][7] ));
 sg13g2_dfrbp_1 _2125_ (.CLK(net972),
    .RESET_B(net1018),
    .D(_0082_),
    .Q_N(_0917_),
    .Q(\u_top_module.u_memory.memory[5][0] ));
 sg13g2_dfrbp_1 _2126_ (.CLK(net963),
    .RESET_B(net1017),
    .D(_0083_),
    .Q_N(_0916_),
    .Q(\u_top_module.u_memory.memory[5][1] ));
 sg13g2_dfrbp_1 _2127_ (.CLK(net974),
    .RESET_B(net1019),
    .D(_0084_),
    .Q_N(_0915_),
    .Q(\u_top_module.u_memory.memory[5][2] ));
 sg13g2_dfrbp_1 _2128_ (.CLK(net961),
    .RESET_B(net1013),
    .D(_0085_),
    .Q_N(_0914_),
    .Q(\u_top_module.u_memory.memory[5][3] ));
 sg13g2_dfrbp_1 _2129_ (.CLK(net960),
    .RESET_B(net1012),
    .D(_0086_),
    .Q_N(_0913_),
    .Q(\u_top_module.u_memory.memory[5][4] ));
 sg13g2_dfrbp_1 _2130_ (.CLK(net973),
    .RESET_B(net1020),
    .D(_0087_),
    .Q_N(_0912_),
    .Q(\u_top_module.u_memory.memory[5][5] ));
 sg13g2_dfrbp_1 _2131_ (.CLK(net967),
    .RESET_B(net1015),
    .D(_0088_),
    .Q_N(_0911_),
    .Q(\u_top_module.u_memory.memory[5][6] ));
 sg13g2_dfrbp_1 _2132_ (.CLK(net959),
    .RESET_B(net1011),
    .D(_0089_),
    .Q_N(_0910_),
    .Q(\u_top_module.u_memory.memory[5][7] ));
 sg13g2_dfrbp_1 _2133_ (.CLK(net969),
    .RESET_B(net1015),
    .D(_0090_),
    .Q_N(_0909_),
    .Q(\u_top_module.u_memory.memory[2][0] ));
 sg13g2_dfrbp_1 _2134_ (.CLK(net963),
    .RESET_B(net1017),
    .D(_0091_),
    .Q_N(_0908_),
    .Q(\u_top_module.u_memory.memory[2][1] ));
 sg13g2_dfrbp_1 _2135_ (.CLK(net974),
    .RESET_B(net1019),
    .D(_0092_),
    .Q_N(_0907_),
    .Q(\u_top_module.u_memory.memory[2][2] ));
 sg13g2_dfrbp_1 _2136_ (.CLK(net962),
    .RESET_B(net1013),
    .D(_0093_),
    .Q_N(_0906_),
    .Q(\u_top_module.u_memory.memory[2][3] ));
 sg13g2_dfrbp_1 _2137_ (.CLK(net967),
    .RESET_B(net1012),
    .D(_0094_),
    .Q_N(_0905_),
    .Q(\u_top_module.u_memory.memory[2][4] ));
 sg13g2_dfrbp_1 _2138_ (.CLK(net973),
    .RESET_B(net1020),
    .D(_0095_),
    .Q_N(_0904_),
    .Q(\u_top_module.u_memory.memory[2][5] ));
 sg13g2_dfrbp_1 _2139_ (.CLK(net968),
    .RESET_B(net1015),
    .D(_0096_),
    .Q_N(_0903_),
    .Q(\u_top_module.u_memory.memory[2][6] ));
 sg13g2_dfrbp_1 _2140_ (.CLK(net959),
    .RESET_B(net1011),
    .D(_0097_),
    .Q_N(_0902_),
    .Q(\u_top_module.u_memory.memory[2][7] ));
 sg13g2_dfrbp_1 _2141_ (.CLK(net972),
    .RESET_B(net1018),
    .D(_0098_),
    .Q_N(_0901_),
    .Q(\u_top_module.u_memory.memory[3][0] ));
 sg13g2_dfrbp_1 _2142_ (.CLK(net963),
    .RESET_B(net1017),
    .D(_0099_),
    .Q_N(_0900_),
    .Q(\u_top_module.u_memory.memory[3][1] ));
 sg13g2_dfrbp_1 _2143_ (.CLK(net974),
    .RESET_B(net1023),
    .D(_0100_),
    .Q_N(_0899_),
    .Q(\u_top_module.u_memory.memory[3][2] ));
 sg13g2_dfrbp_1 _2144_ (.CLK(net961),
    .RESET_B(net1013),
    .D(_0101_),
    .Q_N(_0898_),
    .Q(\u_top_module.u_memory.memory[3][3] ));
 sg13g2_dfrbp_1 _2145_ (.CLK(net960),
    .RESET_B(net1012),
    .D(_0102_),
    .Q_N(_0897_),
    .Q(\u_top_module.u_memory.memory[3][4] ));
 sg13g2_dfrbp_1 _2146_ (.CLK(net973),
    .RESET_B(net1020),
    .D(_0103_),
    .Q_N(_0896_),
    .Q(\u_top_module.u_memory.memory[3][5] ));
 sg13g2_dfrbp_1 _2147_ (.CLK(net968),
    .RESET_B(net1015),
    .D(_0104_),
    .Q_N(_0895_),
    .Q(\u_top_module.u_memory.memory[3][6] ));
 sg13g2_dfrbp_1 _2148_ (.CLK(net959),
    .RESET_B(net1011),
    .D(_0105_),
    .Q_N(_0894_),
    .Q(\u_top_module.u_memory.memory[3][7] ));
 sg13g2_dfrbp_1 _2149_ (.CLK(net972),
    .RESET_B(net1018),
    .D(_0106_),
    .Q_N(_0893_),
    .Q(\u_top_module.u_memory.memory[6][0] ));
 sg13g2_dfrbp_1 _2150_ (.CLK(net963),
    .RESET_B(net1017),
    .D(_0107_),
    .Q_N(_0892_),
    .Q(\u_top_module.u_memory.memory[6][1] ));
 sg13g2_dfrbp_1 _2151_ (.CLK(net969),
    .RESET_B(net1019),
    .D(_0108_),
    .Q_N(_0891_),
    .Q(\u_top_module.u_memory.memory[6][2] ));
 sg13g2_dfrbp_1 _2152_ (.CLK(net961),
    .RESET_B(net1013),
    .D(_0109_),
    .Q_N(_0890_),
    .Q(\u_top_module.u_memory.memory[6][3] ));
 sg13g2_dfrbp_1 _2153_ (.CLK(net960),
    .RESET_B(net1011),
    .D(_0110_),
    .Q_N(_0889_),
    .Q(\u_top_module.u_memory.memory[6][4] ));
 sg13g2_dfrbp_1 _2154_ (.CLK(net968),
    .RESET_B(net1020),
    .D(_0111_),
    .Q_N(_0888_),
    .Q(\u_top_module.u_memory.memory[6][5] ));
 sg13g2_dfrbp_1 _2155_ (.CLK(net967),
    .RESET_B(net1015),
    .D(_0112_),
    .Q_N(_0887_),
    .Q(\u_top_module.u_memory.memory[6][6] ));
 sg13g2_dfrbp_1 _2156_ (.CLK(net959),
    .RESET_B(net1011),
    .D(_0113_),
    .Q_N(_0886_),
    .Q(\u_top_module.u_memory.memory[6][7] ));
 sg13g2_dfrbp_1 _2157_ (.CLK(net968),
    .RESET_B(net1018),
    .D(_0114_),
    .Q_N(_0885_),
    .Q(\u_top_module.u_memory.memory[4][0] ));
 sg13g2_dfrbp_1 _2158_ (.CLK(net963),
    .RESET_B(net1017),
    .D(_0115_),
    .Q_N(_0884_),
    .Q(\u_top_module.u_memory.memory[4][1] ));
 sg13g2_dfrbp_1 _2159_ (.CLK(net969),
    .RESET_B(net1019),
    .D(_0116_),
    .Q_N(_0883_),
    .Q(\u_top_module.u_memory.memory[4][2] ));
 sg13g2_dfrbp_1 _2160_ (.CLK(net961),
    .RESET_B(net984),
    .D(_0117_),
    .Q_N(_0882_),
    .Q(\u_top_module.u_memory.memory[4][3] ));
 sg13g2_dfrbp_1 _2161_ (.CLK(net960),
    .RESET_B(net1011),
    .D(_0118_),
    .Q_N(_0881_),
    .Q(\u_top_module.u_memory.memory[4][4] ));
 sg13g2_dfrbp_1 _2162_ (.CLK(net973),
    .RESET_B(net1020),
    .D(_0119_),
    .Q_N(_0880_),
    .Q(\u_top_module.u_memory.memory[4][5] ));
 sg13g2_dfrbp_1 _2163_ (.CLK(net967),
    .RESET_B(net1015),
    .D(_0120_),
    .Q_N(_0879_),
    .Q(\u_top_module.u_memory.memory[4][6] ));
 sg13g2_dfrbp_1 _2164_ (.CLK(net959),
    .RESET_B(net1011),
    .D(_0121_),
    .Q_N(_0878_),
    .Q(\u_top_module.u_memory.memory[4][7] ));
 sg13g2_dfrbp_1 _2165_ (.CLK(net980),
    .RESET_B(net1024),
    .D(_0030_),
    .Q_N(\u_top_module.u_spi_port.cs_n_prev ),
    .Q(_0029_));
 sg13g2_dfrbp_1 _2166_ (.CLK(net976),
    .RESET_B(net1023),
    .D(_0122_),
    .Q_N(_0877_),
    .Q(\u_top_module.capture_reg[0] ));
 sg13g2_dfrbp_1 _2167_ (.CLK(net976),
    .RESET_B(net1022),
    .D(_0123_),
    .Q_N(_0876_),
    .Q(\u_top_module.capture_reg[1] ));
 sg13g2_dfrbp_1 _2168_ (.CLK(net973),
    .RESET_B(net1022),
    .D(_0124_),
    .Q_N(_0875_),
    .Q(\u_top_module.capture_reg[2] ));
 sg13g2_dfrbp_1 _2169_ (.CLK(net976),
    .RESET_B(net1023),
    .D(_0125_),
    .Q_N(_0874_),
    .Q(\u_top_module.capture_reg[3] ));
 sg13g2_dfrbp_1 _2170_ (.CLK(net975),
    .RESET_B(net1021),
    .D(_0126_),
    .Q_N(_0873_),
    .Q(\u_top_module.capture_reg[4] ));
 sg13g2_dfrbp_1 _2171_ (.CLK(net973),
    .RESET_B(net1020),
    .D(_0127_),
    .Q_N(_0872_),
    .Q(\u_top_module.capture_reg[5] ));
 sg13g2_dfrbp_1 _2172_ (.CLK(net973),
    .RESET_B(net1021),
    .D(_0128_),
    .Q_N(_0871_),
    .Q(\u_top_module.capture_reg[6] ));
 sg13g2_dfrbp_1 _2173_ (.CLK(net975),
    .RESET_B(net1021),
    .D(_0129_),
    .Q_N(_0870_),
    .Q(\u_top_module.capture_reg[7] ));
 sg13g2_dfrbp_1 _2174_ (.CLK(net973),
    .RESET_B(net1024),
    .D(_0130_),
    .Q_N(_0869_),
    .Q(\u_top_module.addr[0] ));
 sg13g2_dfrbp_1 _2175_ (.CLK(net978),
    .RESET_B(net1026),
    .D(_0131_),
    .Q_N(_0868_),
    .Q(\u_top_module.addr[1] ));
 sg13g2_dfrbp_1 _2176_ (.CLK(net978),
    .RESET_B(net1026),
    .D(_0132_),
    .Q_N(_0027_),
    .Q(\u_top_module.addr[2] ));
 sg13g2_dfrbp_1 _2177_ (.CLK(net978),
    .RESET_B(net1024),
    .D(_0133_),
    .Q_N(_0867_),
    .Q(\u_top_module.addr[3] ));
 sg13g2_dfrbp_1 _2178_ (.CLK(net979),
    .RESET_B(net1025),
    .D(_0134_),
    .Q_N(_0866_),
    .Q(\u_top_module.addr[4] ));
 sg13g2_dfrbp_1 _2179_ (.CLK(net979),
    .RESET_B(net1025),
    .D(_0135_),
    .Q_N(_0865_),
    .Q(\u_top_module.addr[5] ));
 sg13g2_dfrbp_1 _2180_ (.CLK(net979),
    .RESET_B(net1025),
    .D(_0136_),
    .Q_N(_0864_),
    .Q(\u_top_module.addr[6] ));
 sg13g2_dfrbp_1 _2181_ (.CLK(net979),
    .RESET_B(net1025),
    .D(_0137_),
    .Q_N(_0863_),
    .Q(\u_top_module.addr[7] ));
 sg13g2_dfrbp_1 _2182_ (.CLK(net969),
    .RESET_B(net1016),
    .D(_0138_),
    .Q_N(_0862_),
    .Q(\u_top_module.u_memory.memory[7][0] ));
 sg13g2_dfrbp_1 _2183_ (.CLK(net963),
    .RESET_B(net1017),
    .D(_0139_),
    .Q_N(_0861_),
    .Q(\u_top_module.u_memory.memory[7][1] ));
 sg13g2_dfrbp_1 _2184_ (.CLK(net974),
    .RESET_B(net1019),
    .D(_0140_),
    .Q_N(_0860_),
    .Q(\u_top_module.u_memory.memory[7][2] ));
 sg13g2_dfrbp_1 _2185_ (.CLK(net962),
    .RESET_B(net1013),
    .D(_0141_),
    .Q_N(_0859_),
    .Q(\u_top_module.u_memory.memory[7][3] ));
 sg13g2_dfrbp_1 _2186_ (.CLK(net959),
    .RESET_B(net1012),
    .D(_0142_),
    .Q_N(_0858_),
    .Q(\u_top_module.u_memory.memory[7][4] ));
 sg13g2_dfrbp_1 _2187_ (.CLK(net968),
    .RESET_B(net1020),
    .D(_0143_),
    .Q_N(_0857_),
    .Q(\u_top_module.u_memory.memory[7][5] ));
 sg13g2_dfrbp_1 _2188_ (.CLK(net968),
    .RESET_B(net1015),
    .D(_0144_),
    .Q_N(_0856_),
    .Q(\u_top_module.u_memory.memory[7][6] ));
 sg13g2_dfrbp_1 _2189_ (.CLK(net959),
    .RESET_B(net1011),
    .D(_0145_),
    .Q_N(_0855_),
    .Q(\u_top_module.u_memory.memory[7][7] ));
 sg13g2_dfrbp_1 _2190_ (.CLK(net976),
    .RESET_B(net1022),
    .D(_0146_),
    .Q_N(_0854_),
    .Q(\u_top_module.u_spi_port.shift_reg[0] ));
 sg13g2_dfrbp_1 _2191_ (.CLK(net976),
    .RESET_B(net1022),
    .D(_0147_),
    .Q_N(_0853_),
    .Q(\u_top_module.u_spi_port.shift_reg[1] ));
 sg13g2_dfrbp_1 _2192_ (.CLK(net975),
    .RESET_B(net1022),
    .D(_0148_),
    .Q_N(_0852_),
    .Q(\u_top_module.u_spi_port.shift_reg[2] ));
 sg13g2_dfrbp_1 _2193_ (.CLK(net975),
    .RESET_B(net1021),
    .D(_0149_),
    .Q_N(_0851_),
    .Q(\u_top_module.u_spi_port.shift_reg[3] ));
 sg13g2_dfrbp_1 _2194_ (.CLK(net975),
    .RESET_B(net1021),
    .D(_0150_),
    .Q_N(_0850_),
    .Q(\u_top_module.u_spi_port.shift_reg[4] ));
 sg13g2_dfrbp_1 _2195_ (.CLK(net975),
    .RESET_B(net1021),
    .D(_0151_),
    .Q_N(_0849_),
    .Q(\u_top_module.u_spi_port.shift_reg[5] ));
 sg13g2_dfrbp_1 _2196_ (.CLK(net975),
    .RESET_B(net1021),
    .D(_0152_),
    .Q_N(_0848_),
    .Q(\u_top_module.u_spi_port.shift_reg[6] ));
 sg13g2_dfrbp_1 _2197_ (.CLK(net975),
    .RESET_B(net1021),
    .D(_0153_),
    .Q_N(_0847_),
    .Q(\u_top_module.u_spi_port.shift_reg[7] ));
 sg13g2_dfrbp_1 _2198_ (.CLK(net976),
    .RESET_B(net1022),
    .D(_0154_),
    .Q_N(_0846_),
    .Q(\u_top_module.u_spi_port.shift_reg[8] ));
 sg13g2_dfrbp_1 _2199_ (.CLK(net976),
    .RESET_B(net1022),
    .D(_0155_),
    .Q_N(_0845_),
    .Q(\u_top_module.u_spi_port.shift_reg[9] ));
 sg13g2_dfrbp_1 _2200_ (.CLK(net976),
    .RESET_B(net1024),
    .D(_0156_),
    .Q_N(_0844_),
    .Q(\u_top_module.u_spi_port.shift_reg[10] ));
 sg13g2_dfrbp_1 _2201_ (.CLK(net979),
    .RESET_B(net1024),
    .D(_0157_),
    .Q_N(_0843_),
    .Q(\u_top_module.u_spi_port.shift_reg[11] ));
 sg13g2_dfrbp_1 _2202_ (.CLK(net979),
    .RESET_B(net1024),
    .D(_0158_),
    .Q_N(_0842_),
    .Q(\u_top_module.u_spi_port.shift_reg[12] ));
 sg13g2_dfrbp_1 _2203_ (.CLK(net979),
    .RESET_B(net1024),
    .D(_0159_),
    .Q_N(_0841_),
    .Q(\u_top_module.u_spi_port.shift_reg[13] ));
 sg13g2_dfrbp_1 _2204_ (.CLK(net980),
    .RESET_B(net1024),
    .D(_0160_),
    .Q_N(_0840_),
    .Q(\u_top_module.u_spi_port.shift_reg[14] ));
 sg13g2_dfrbp_1 _2205_ (.CLK(net980),
    .RESET_B(net1025),
    .D(_0161_),
    .Q_N(_0839_),
    .Q(\u_top_module.u_spi_port.shift_reg[15] ));
 sg13g2_dfrbp_1 _2206_ (.CLK(net920),
    .RESET_B(net1029),
    .D(_0162_),
    .Q_N(_0838_),
    .Q(\u_top_module.u_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2207_ (.CLK(net920),
    .RESET_B(net1002),
    .D(_0163_),
    .Q_N(_0837_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2208_ (.CLK(net912),
    .RESET_B(net985),
    .D(_0164_),
    .Q_N(_0836_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2209_ (.CLK(net912),
    .RESET_B(net1002),
    .D(_0165_),
    .Q_N(_0835_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2210_ (.CLK(net910),
    .RESET_B(net985),
    .D(_0166_),
    .Q_N(_0834_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2211_ (.CLK(net910),
    .RESET_B(net985),
    .D(_0167_),
    .Q_N(_0833_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2212_ (.CLK(net910),
    .RESET_B(net985),
    .D(_0168_),
    .Q_N(_0832_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2213_ (.CLK(net900),
    .RESET_B(net1051),
    .D(_0169_),
    .Q_N(_0948_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2214_ (.CLK(net954),
    .RESET_B(net984),
    .D(_0011_),
    .Q_N(_0949_),
    .Q(\u_top_module.u_i2s_bus.counter[0] ));
 sg13g2_dfrbp_1 _2215_ (.CLK(net954),
    .RESET_B(net984),
    .D(_0012_),
    .Q_N(_0950_),
    .Q(\u_top_module.u_i2s_bus.counter[1] ));
 sg13g2_dfrbp_1 _2216_ (.CLK(net954),
    .RESET_B(net984),
    .D(_0013_),
    .Q_N(_0951_),
    .Q(\u_top_module.u_i2s_bus.counter[2] ));
 sg13g2_dfrbp_1 _2217_ (.CLK(net954),
    .RESET_B(net984),
    .D(_0014_),
    .Q_N(_0952_),
    .Q(\u_top_module.u_i2s_bus.counter[3] ));
 sg13g2_dfrbp_1 _2218_ (.CLK(net954),
    .RESET_B(net985),
    .D(_0015_),
    .Q_N(_0953_),
    .Q(\u_top_module.u_i2s_bus.counter[4] ));
 sg13g2_dfrbp_1 _2219_ (.CLK(net962),
    .RESET_B(net985),
    .D(_0016_),
    .Q_N(_0954_),
    .Q(\u_top_module.u_i2s_bus.counter[5] ));
 sg13g2_dfrbp_1 _2220_ (.CLK(net962),
    .RESET_B(net984),
    .D(_0017_),
    .Q_N(_0955_),
    .Q(\u_top_module.u_i2s_bus.counter[6] ));
 sg13g2_dfrbp_1 _2221_ (.CLK(net962),
    .RESET_B(net984),
    .D(net26),
    .Q_N(_0831_),
    .Q(\u_top_module.u_i2s_bus.counter[7] ));
 sg13g2_dfrbp_1 _2222_ (.CLK(_0031_),
    .RESET_B(net106),
    .D(_0170_),
    .Q_N(_0830_),
    .Q(\u_top_module.out ));
 sg13g2_dfrbp_1 _2223_ (.CLK(net956),
    .RESET_B(net105),
    .D(_0171_),
    .Q_N(_0829_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[9].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2224_ (.CLK(_0032_),
    .RESET_B(net108),
    .D(\u_top_module.u_i2s_bus.u_mux_shift.data ),
    .Q_N(_0956_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _2225_ (.CLK(net964),
    .RESET_B(net104),
    .D(_0020_),
    .Q_N(_0828_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2226_ (.CLK(_0033_),
    .RESET_B(net109),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.data ),
    .Q_N(_0957_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2227_ (.CLK(net965),
    .RESET_B(net103),
    .D(_0021_),
    .Q_N(_0827_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2228_ (.CLK(_0034_),
    .RESET_B(net110),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.data ),
    .Q_N(_0958_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2229_ (.CLK(net965),
    .RESET_B(net102),
    .D(_0022_),
    .Q_N(_0826_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2230_ (.CLK(_0035_),
    .RESET_B(net111),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.data ),
    .Q_N(_0959_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2231_ (.CLK(net958),
    .RESET_B(net101),
    .D(_0023_),
    .Q_N(_0825_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2232_ (.CLK(_0036_),
    .RESET_B(net112),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.data ),
    .Q_N(_0960_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2233_ (.CLK(net956),
    .RESET_B(net100),
    .D(_0024_),
    .Q_N(_0824_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2234_ (.CLK(_0037_),
    .RESET_B(net113),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.data ),
    .Q_N(_0961_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2235_ (.CLK(net957),
    .RESET_B(net99),
    .D(_0025_),
    .Q_N(_0823_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2236_ (.CLK(_0038_),
    .RESET_B(net114),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.data ),
    .Q_N(_0962_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2237_ (.CLK(net956),
    .RESET_B(net98),
    .D(_0026_),
    .Q_N(_0822_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2238_ (.CLK(_0039_),
    .RESET_B(net97),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.data ),
    .Q_N(_0821_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2239_ (.CLK(net964),
    .RESET_B(net96),
    .D(_0172_),
    .Q_N(_0820_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2240_ (.CLK(_0040_),
    .RESET_B(net95),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.data ),
    .Q_N(_0819_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2241_ (.CLK(net956),
    .RESET_B(net94),
    .D(_0173_),
    .Q_N(_0818_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2242_ (.CLK(_0041_),
    .RESET_B(net115),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[9].u_mux_shift.data ),
    .Q_N(_0963_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _2243_ (.CLK(net962),
    .RESET_B(net93),
    .D(\u_top_module.u_i2s_bus.dec_clk ),
    .Q_N(_0817_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.prev_lr_clk ));
 sg13g2_dfrbp_1 _2244_ (.CLK(net962),
    .RESET_B(net984),
    .D(_0174_),
    .Q_N(_0019_),
    .Q(\u_top_module.u_i2s_bus.dec_clk ));
 sg13g2_dfrbp_1 _2245_ (.CLK(_0042_),
    .RESET_B(net92),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.data ),
    .Q_N(_0816_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2246_ (.CLK(net956),
    .RESET_B(net91),
    .D(_0175_),
    .Q_N(_0815_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2247_ (.CLK(_0043_),
    .RESET_B(net90),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.data ),
    .Q_N(_0814_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2248_ (.CLK(net958),
    .RESET_B(net89),
    .D(_0176_),
    .Q_N(_0813_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2249_ (.CLK(_0044_),
    .RESET_B(net88),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.data ),
    .Q_N(_0812_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2250_ (.CLK(net958),
    .RESET_B(net87),
    .D(_0177_),
    .Q_N(_0811_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2251_ (.CLK(_0045_),
    .RESET_B(net86),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.data ),
    .Q_N(_0810_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2252_ (.CLK(net953),
    .RESET_B(net85),
    .D(_0178_),
    .Q_N(_0809_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2253_ (.CLK(_0046_),
    .RESET_B(net84),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.data ),
    .Q_N(_0808_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2254_ (.CLK(net953),
    .RESET_B(net83),
    .D(_0179_),
    .Q_N(_0807_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2255_ (.CLK(_0047_),
    .RESET_B(net82),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.data ),
    .Q_N(_0806_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2256_ (.CLK(net953),
    .RESET_B(net81),
    .D(_0180_),
    .Q_N(_0805_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2257_ (.CLK(_0048_),
    .RESET_B(net80),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.data ),
    .Q_N(_0804_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2258_ (.CLK(net952),
    .RESET_B(net79),
    .D(_0181_),
    .Q_N(_0803_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2259_ (.CLK(_0049_),
    .RESET_B(net78),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.data ),
    .Q_N(_0802_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2260_ (.CLK(net952),
    .RESET_B(net77),
    .D(_0182_),
    .Q_N(_0801_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2261_ (.CLK(_0050_),
    .RESET_B(net76),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.data ),
    .Q_N(_0800_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2262_ (.CLK(net952),
    .RESET_B(net75),
    .D(_0183_),
    .Q_N(_0799_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2263_ (.CLK(_0051_),
    .RESET_B(net74),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.data ),
    .Q_N(_0798_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2264_ (.CLK(net952),
    .RESET_B(net73),
    .D(_0184_),
    .Q_N(_0797_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2265_ (.CLK(_0052_),
    .RESET_B(net72),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.data ),
    .Q_N(_0796_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2266_ (.CLK(net951),
    .RESET_B(net71),
    .D(_0185_),
    .Q_N(_0795_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2267_ (.CLK(_0053_),
    .RESET_B(net70),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.data ),
    .Q_N(_0794_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2268_ (.CLK(net951),
    .RESET_B(net69),
    .D(_0186_),
    .Q_N(_0793_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2269_ (.CLK(_0054_),
    .RESET_B(net68),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.data ),
    .Q_N(_0792_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2270_ (.CLK(net951),
    .RESET_B(net67),
    .D(_0187_),
    .Q_N(_0791_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2271_ (.CLK(_0055_),
    .RESET_B(net66),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.data ),
    .Q_N(_0790_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2272_ (.CLK(net951),
    .RESET_B(net65),
    .D(_0188_),
    .Q_N(_0789_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2273_ (.CLK(_0056_),
    .RESET_B(net64),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.data ),
    .Q_N(_0788_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2274_ (.CLK(net951),
    .RESET_B(net63),
    .D(_0189_),
    .Q_N(_0787_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2275_ (.CLK(_0057_),
    .RESET_B(net62),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.data ),
    .Q_N(_0786_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2276_ (.CLK(net954),
    .RESET_B(net61),
    .D(_0190_),
    .Q_N(_0785_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2277_ (.CLK(_0058_),
    .RESET_B(net60),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.data ),
    .Q_N(_0784_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2278_ (.CLK(net954),
    .RESET_B(net59),
    .D(_0191_),
    .Q_N(_0783_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2279_ (.CLK(_0059_),
    .RESET_B(net58),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.data ),
    .Q_N(_0782_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2280_ (.CLK(net953),
    .RESET_B(net57),
    .D(_0192_),
    .Q_N(_0781_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2281_ (.CLK(_0060_),
    .RESET_B(net56),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.data ),
    .Q_N(_0780_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2282_ (.CLK(net965),
    .RESET_B(net55),
    .D(_0193_),
    .Q_N(_0779_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2283_ (.CLK(_0061_),
    .RESET_B(net54),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.data ),
    .Q_N(_0778_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2284_ (.CLK(net965),
    .RESET_B(net53),
    .D(_0194_),
    .Q_N(_0777_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2285_ (.CLK(_0062_),
    .RESET_B(net52),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.data ),
    .Q_N(_0776_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2286_ (.CLK(net963),
    .RESET_B(net51),
    .D(_0195_),
    .Q_N(_0775_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2287_ (.CLK(_0063_),
    .RESET_B(net116),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.data ),
    .Q_N(_0964_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2288_ (.CLK(net931),
    .RESET_B(net1039),
    .D(\u_top_module.dec_data ),
    .Q_N(_0965_),
    .Q(\u_top_module.u_filter.shift_reg[0] ));
 sg13g2_dfrbp_1 _2289_ (.CLK(net931),
    .RESET_B(net1039),
    .D(\u_top_module.u_filter.shift_reg[0] ),
    .Q_N(_0966_),
    .Q(\u_top_module.u_filter.shift_reg[1] ));
 sg13g2_dfrbp_1 _2290_ (.CLK(net931),
    .RESET_B(net1039),
    .D(\u_top_module.u_filter.shift_reg[1] ),
    .Q_N(_0967_),
    .Q(\u_top_module.u_filter.shift_reg[2] ));
 sg13g2_dfrbp_1 _2291_ (.CLK(net931),
    .RESET_B(net1039),
    .D(\u_top_module.u_filter.shift_reg[2] ),
    .Q_N(_0968_),
    .Q(\u_top_module.u_filter.shift_reg[3] ));
 sg13g2_dfrbp_1 _2292_ (.CLK(net931),
    .RESET_B(net1039),
    .D(\u_top_module.u_filter.shift_reg[3] ),
    .Q_N(_0969_),
    .Q(\u_top_module.u_filter.shift_reg[4] ));
 sg13g2_dfrbp_1 _2293_ (.CLK(net931),
    .RESET_B(net1041),
    .D(\u_top_module.u_filter.shift_reg[4] ),
    .Q_N(_0970_),
    .Q(\u_top_module.u_filter.shift_reg[5] ));
 sg13g2_dfrbp_1 _2294_ (.CLK(net931),
    .RESET_B(net1041),
    .D(\u_top_module.u_filter.shift_reg[5] ),
    .Q_N(_0971_),
    .Q(\u_top_module.u_filter.shift_reg[6] ));
 sg13g2_dfrbp_1 _2295_ (.CLK(net932),
    .RESET_B(net1039),
    .D(\u_top_module.u_filter.shift_reg[6] ),
    .Q_N(_0972_),
    .Q(\u_top_module.u_filter.shift_reg[7] ));
 sg13g2_dfrbp_1 _2296_ (.CLK(net932),
    .RESET_B(net1040),
    .D(\u_top_module.u_filter.shift_reg[7] ),
    .Q_N(_0973_),
    .Q(\u_top_module.u_filter.shift_reg[8] ));
 sg13g2_dfrbp_1 _2297_ (.CLK(net932),
    .RESET_B(net1041),
    .D(\u_top_module.u_filter.shift_reg[8] ),
    .Q_N(_0974_),
    .Q(\u_top_module.u_filter.shift_reg[9] ));
 sg13g2_dfrbp_1 _2298_ (.CLK(net930),
    .RESET_B(net1041),
    .D(\u_top_module.u_filter.shift_reg[9] ),
    .Q_N(_0975_),
    .Q(\u_top_module.u_filter.shift_reg[10] ));
 sg13g2_dfrbp_1 _2299_ (.CLK(net937),
    .RESET_B(net1040),
    .D(\u_top_module.u_filter.shift_reg[10] ),
    .Q_N(_0976_),
    .Q(\u_top_module.u_filter.shift_reg[11] ));
 sg13g2_dfrbp_1 _2300_ (.CLK(net937),
    .RESET_B(net1046),
    .D(\u_top_module.u_filter.shift_reg[11] ),
    .Q_N(_0977_),
    .Q(\u_top_module.u_filter.shift_reg[12] ));
 sg13g2_dfrbp_1 _2301_ (.CLK(net936),
    .RESET_B(net1046),
    .D(\u_top_module.u_filter.shift_reg[12] ),
    .Q_N(_0978_),
    .Q(\u_top_module.u_filter.shift_reg[13] ));
 sg13g2_dfrbp_1 _2302_ (.CLK(net937),
    .RESET_B(net1046),
    .D(\u_top_module.u_filter.shift_reg[13] ),
    .Q_N(_0979_),
    .Q(\u_top_module.u_filter.shift_reg[14] ));
 sg13g2_dfrbp_1 _2303_ (.CLK(net936),
    .RESET_B(net1048),
    .D(\u_top_module.u_filter.shift_reg[14] ),
    .Q_N(_0980_),
    .Q(\u_top_module.u_filter.shift_reg[15] ));
 sg13g2_dfrbp_1 _2304_ (.CLK(net936),
    .RESET_B(net1040),
    .D(\u_top_module.u_filter.shift_reg[15] ),
    .Q_N(_0981_),
    .Q(\u_top_module.u_filter.shift_reg[16] ));
 sg13g2_dfrbp_1 _2305_ (.CLK(net930),
    .RESET_B(net1040),
    .D(\u_top_module.u_filter.shift_reg[16] ),
    .Q_N(_0982_),
    .Q(\u_top_module.u_filter.shift_reg[17] ));
 sg13g2_dfrbp_1 _2306_ (.CLK(net930),
    .RESET_B(net1040),
    .D(\u_top_module.u_filter.shift_reg[17] ),
    .Q_N(_0983_),
    .Q(\u_top_module.u_filter.shift_reg[18] ));
 sg13g2_dfrbp_1 _2307_ (.CLK(net930),
    .RESET_B(net1040),
    .D(\u_top_module.u_filter.shift_reg[18] ),
    .Q_N(_0984_),
    .Q(\u_top_module.u_filter.shift_reg[19] ));
 sg13g2_dfrbp_1 _2308_ (.CLK(net930),
    .RESET_B(net1040),
    .D(\u_top_module.u_filter.shift_reg[19] ),
    .Q_N(_0985_),
    .Q(\u_top_module.u_filter.shift_reg[20] ));
 sg13g2_dfrbp_1 _2309_ (.CLK(net930),
    .RESET_B(net1040),
    .D(\u_top_module.u_filter.shift_reg[20] ),
    .Q_N(_0986_),
    .Q(\u_top_module.u_filter.shift_reg[21] ));
 sg13g2_dfrbp_1 _2310_ (.CLK(net930),
    .RESET_B(net1038),
    .D(\u_top_module.u_filter.shift_reg[21] ),
    .Q_N(_0987_),
    .Q(\u_top_module.u_filter.shift_reg[22] ));
 sg13g2_dfrbp_1 _2311_ (.CLK(net930),
    .RESET_B(net1038),
    .D(\u_top_module.u_filter.shift_reg[22] ),
    .Q_N(_0988_),
    .Q(\u_top_module.u_filter.shift_reg[23] ));
 sg13g2_dfrbp_1 _2312_ (.CLK(net933),
    .RESET_B(net1038),
    .D(\u_top_module.u_filter.shift_reg[23] ),
    .Q_N(_0989_),
    .Q(\u_top_module.u_filter.shift_reg[24] ));
 sg13g2_dfrbp_1 _2313_ (.CLK(net933),
    .RESET_B(net1038),
    .D(\u_top_module.u_filter.shift_reg[24] ),
    .Q_N(_0990_),
    .Q(\u_top_module.u_filter.shift_reg[25] ));
 sg13g2_dfrbp_1 _2314_ (.CLK(net933),
    .RESET_B(net1038),
    .D(\u_top_module.u_filter.shift_reg[25] ),
    .Q_N(_0991_),
    .Q(\u_top_module.u_filter.shift_reg[26] ));
 sg13g2_dfrbp_1 _2315_ (.CLK(net933),
    .RESET_B(net1042),
    .D(\u_top_module.u_filter.shift_reg[26] ),
    .Q_N(_0992_),
    .Q(\u_top_module.u_filter.shift_reg[27] ));
 sg13g2_dfrbp_1 _2316_ (.CLK(net933),
    .RESET_B(net1042),
    .D(\u_top_module.u_filter.shift_reg[27] ),
    .Q_N(_0993_),
    .Q(\u_top_module.u_filter.shift_reg[28] ));
 sg13g2_dfrbp_1 _2317_ (.CLK(net935),
    .RESET_B(net1045),
    .D(\u_top_module.u_filter.shift_reg[28] ),
    .Q_N(_0994_),
    .Q(\u_top_module.u_filter.shift_reg[29] ));
 sg13g2_dfrbp_1 _2318_ (.CLK(net935),
    .RESET_B(net1045),
    .D(\u_top_module.u_filter.shift_reg[29] ),
    .Q_N(_0995_),
    .Q(\u_top_module.u_filter.shift_reg[30] ));
 sg13g2_dfrbp_1 _2319_ (.CLK(net935),
    .RESET_B(net1045),
    .D(\u_top_module.u_filter.shift_reg[30] ),
    .Q_N(_0996_),
    .Q(\u_top_module.u_filter.shift_reg[31] ));
 sg13g2_dfrbp_1 _2320_ (.CLK(net927),
    .RESET_B(net1036),
    .D(\u_top_module.u_filter.shift_reg[31] ),
    .Q_N(_0997_),
    .Q(\u_top_module.u_filter.shift_reg[32] ));
 sg13g2_dfrbp_1 _2321_ (.CLK(net923),
    .RESET_B(net1033),
    .D(\u_top_module.u_filter.shift_reg[32] ),
    .Q_N(_0998_),
    .Q(\u_top_module.u_filter.shift_reg[33] ));
 sg13g2_dfrbp_1 _2322_ (.CLK(net923),
    .RESET_B(net1033),
    .D(\u_top_module.u_filter.shift_reg[33] ),
    .Q_N(_0999_),
    .Q(\u_top_module.u_filter.shift_reg[34] ));
 sg13g2_dfrbp_1 _2323_ (.CLK(net923),
    .RESET_B(net1009),
    .D(\u_top_module.u_filter.shift_reg[34] ),
    .Q_N(_1000_),
    .Q(\u_top_module.u_filter.shift_reg[35] ));
 sg13g2_dfrbp_1 _2324_ (.CLK(net920),
    .RESET_B(net1002),
    .D(\u_top_module.u_filter.shift_reg[35] ),
    .Q_N(_1001_),
    .Q(\u_top_module.u_filter.shift_reg[36] ));
 sg13g2_dfrbp_1 _2325_ (.CLK(net912),
    .RESET_B(net1002),
    .D(\u_top_module.u_filter.shift_reg[36] ),
    .Q_N(_1002_),
    .Q(\u_top_module.u_filter.shift_reg[37] ));
 sg13g2_dfrbp_1 _2326_ (.CLK(net912),
    .RESET_B(net1002),
    .D(\u_top_module.u_filter.shift_reg[37] ),
    .Q_N(_1003_),
    .Q(\u_top_module.u_filter.shift_reg[38] ));
 sg13g2_dfrbp_1 _2327_ (.CLK(net912),
    .RESET_B(net1002),
    .D(\u_top_module.u_filter.shift_reg[38] ),
    .Q_N(_1004_),
    .Q(\u_top_module.u_filter.shift_reg[39] ));
 sg13g2_dfrbp_1 _2328_ (.CLK(net912),
    .RESET_B(net1002),
    .D(\u_top_module.u_filter.shift_reg[39] ),
    .Q_N(_1005_),
    .Q(\u_top_module.u_filter.shift_reg[40] ));
 sg13g2_dfrbp_1 _2329_ (.CLK(net913),
    .RESET_B(net1003),
    .D(\u_top_module.u_filter.shift_reg[40] ),
    .Q_N(_1006_),
    .Q(\u_top_module.u_filter.shift_reg[41] ));
 sg13g2_dfrbp_1 _2330_ (.CLK(net913),
    .RESET_B(net1003),
    .D(\u_top_module.u_filter.shift_reg[41] ),
    .Q_N(_1007_),
    .Q(\u_top_module.u_filter.shift_reg[42] ));
 sg13g2_dfrbp_1 _2331_ (.CLK(net913),
    .RESET_B(net1003),
    .D(\u_top_module.u_filter.shift_reg[42] ),
    .Q_N(_1008_),
    .Q(\u_top_module.u_filter.shift_reg[43] ));
 sg13g2_dfrbp_1 _2332_ (.CLK(net913),
    .RESET_B(net1003),
    .D(\u_top_module.u_filter.shift_reg[43] ),
    .Q_N(_1009_),
    .Q(\u_top_module.u_filter.shift_reg[44] ));
 sg13g2_dfrbp_1 _2333_ (.CLK(net913),
    .RESET_B(net1002),
    .D(\u_top_module.u_filter.shift_reg[44] ),
    .Q_N(_1010_),
    .Q(\u_top_module.u_filter.shift_reg[45] ));
 sg13g2_dfrbp_1 _2334_ (.CLK(net912),
    .RESET_B(net1003),
    .D(\u_top_module.u_filter.shift_reg[45] ),
    .Q_N(_1011_),
    .Q(\u_top_module.u_filter.shift_reg[46] ));
 sg13g2_dfrbp_1 _2335_ (.CLK(net912),
    .RESET_B(net1003),
    .D(\u_top_module.u_filter.shift_reg[46] ),
    .Q_N(_1012_),
    .Q(\u_top_module.u_filter.shift_reg[47] ));
 sg13g2_dfrbp_1 _2336_ (.CLK(net921),
    .RESET_B(net1003),
    .D(\u_top_module.u_filter.shift_reg[47] ),
    .Q_N(_1013_),
    .Q(\u_top_module.u_filter.shift_reg[48] ));
 sg13g2_dfrbp_1 _2337_ (.CLK(net921),
    .RESET_B(net1032),
    .D(\u_top_module.u_filter.shift_reg[48] ),
    .Q_N(_1014_),
    .Q(\u_top_module.u_filter.shift_reg[49] ));
 sg13g2_dfrbp_1 _2338_ (.CLK(net921),
    .RESET_B(net1032),
    .D(\u_top_module.u_filter.shift_reg[49] ),
    .Q_N(_1015_),
    .Q(\u_top_module.u_filter.shift_reg[50] ));
 sg13g2_dfrbp_1 _2339_ (.CLK(net921),
    .RESET_B(net1032),
    .D(\u_top_module.u_filter.shift_reg[50] ),
    .Q_N(_1016_),
    .Q(\u_top_module.u_filter.shift_reg[51] ));
 sg13g2_dfrbp_1 _2340_ (.CLK(net920),
    .RESET_B(net1029),
    .D(\u_top_module.u_filter.shift_reg[51] ),
    .Q_N(_1017_),
    .Q(\u_top_module.u_filter.shift_reg[52] ));
 sg13g2_dfrbp_1 _2341_ (.CLK(net920),
    .RESET_B(net1029),
    .D(\u_top_module.u_filter.shift_reg[52] ),
    .Q_N(_1018_),
    .Q(\u_top_module.u_filter.shift_reg[53] ));
 sg13g2_dfrbp_1 _2342_ (.CLK(net920),
    .RESET_B(net1029),
    .D(\u_top_module.u_filter.shift_reg[53] ),
    .Q_N(_1019_),
    .Q(\u_top_module.u_filter.shift_reg[54] ));
 sg13g2_dfrbp_1 _2343_ (.CLK(net920),
    .RESET_B(net1029),
    .D(\u_top_module.u_filter.shift_reg[54] ),
    .Q_N(_1020_),
    .Q(\u_top_module.u_filter.shift_reg[55] ));
 sg13g2_dfrbp_1 _2344_ (.CLK(net921),
    .RESET_B(net1029),
    .D(\u_top_module.u_filter.shift_reg[55] ),
    .Q_N(_1021_),
    .Q(\u_top_module.u_filter.shift_reg[56] ));
 sg13g2_dfrbp_1 _2345_ (.CLK(net920),
    .RESET_B(net1029),
    .D(\u_top_module.u_filter.shift_reg[56] ),
    .Q_N(_1022_),
    .Q(\u_top_module.u_filter.shift_reg[57] ));
 sg13g2_dfrbp_1 _2346_ (.CLK(net925),
    .RESET_B(net1029),
    .D(\u_top_module.u_filter.shift_reg[57] ),
    .Q_N(_1023_),
    .Q(\u_top_module.u_filter.shift_reg[58] ));
 sg13g2_dfrbp_1 _2347_ (.CLK(net925),
    .RESET_B(net1033),
    .D(\u_top_module.u_filter.shift_reg[58] ),
    .Q_N(_1024_),
    .Q(\u_top_module.u_filter.shift_reg[59] ));
 sg13g2_dfrbp_1 _2348_ (.CLK(net923),
    .RESET_B(net1033),
    .D(\u_top_module.u_filter.shift_reg[59] ),
    .Q_N(_1025_),
    .Q(\u_top_module.u_filter.shift_reg[60] ));
 sg13g2_dfrbp_1 _2349_ (.CLK(net923),
    .RESET_B(net1033),
    .D(\u_top_module.u_filter.shift_reg[60] ),
    .Q_N(_1026_),
    .Q(\u_top_module.u_filter.shift_reg[61] ));
 sg13g2_dfrbp_1 _2350_ (.CLK(net923),
    .RESET_B(net1033),
    .D(\u_top_module.u_filter.shift_reg[61] ),
    .Q_N(_1027_),
    .Q(\u_top_module.u_filter.shift_reg[62] ));
 sg13g2_dfrbp_1 _2351_ (.CLK(net923),
    .RESET_B(net1033),
    .D(\u_top_module.u_filter.shift_reg[62] ),
    .Q_N(_1028_),
    .Q(\u_top_module.u_filter.shift_reg[63] ));
 sg13g2_dfrbp_1 _2352_ (.CLK(net923),
    .RESET_B(net1033),
    .D(\u_top_module.u_filter.shift_reg[63] ),
    .Q_N(_1029_),
    .Q(\u_top_module.u_filter.shift_reg[64] ));
 sg13g2_dfrbp_1 _2353_ (.CLK(net924),
    .RESET_B(net1037),
    .D(\u_top_module.u_filter.shift_reg[64] ),
    .Q_N(_1030_),
    .Q(\u_top_module.u_filter.shift_reg[65] ));
 sg13g2_dfrbp_1 _2354_ (.CLK(net924),
    .RESET_B(net1034),
    .D(\u_top_module.u_filter.shift_reg[65] ),
    .Q_N(_1031_),
    .Q(\u_top_module.u_filter.shift_reg[66] ));
 sg13g2_dfrbp_1 _2355_ (.CLK(net924),
    .RESET_B(net1034),
    .D(\u_top_module.u_filter.shift_reg[66] ),
    .Q_N(_1032_),
    .Q(\u_top_module.u_filter.shift_reg[67] ));
 sg13g2_dfrbp_1 _2356_ (.CLK(net925),
    .RESET_B(net1034),
    .D(\u_top_module.u_filter.shift_reg[67] ),
    .Q_N(_1033_),
    .Q(\u_top_module.u_filter.shift_reg[68] ));
 sg13g2_dfrbp_1 _2357_ (.CLK(net924),
    .RESET_B(net1034),
    .D(\u_top_module.u_filter.shift_reg[68] ),
    .Q_N(_1034_),
    .Q(\u_top_module.u_filter.shift_reg[69] ));
 sg13g2_dfrbp_1 _2358_ (.CLK(net924),
    .RESET_B(net1034),
    .D(\u_top_module.u_filter.shift_reg[69] ),
    .Q_N(_1035_),
    .Q(\u_top_module.u_filter.shift_reg[70] ));
 sg13g2_dfrbp_1 _2359_ (.CLK(net924),
    .RESET_B(net1034),
    .D(\u_top_module.u_filter.shift_reg[70] ),
    .Q_N(_1036_),
    .Q(\u_top_module.u_filter.shift_reg[71] ));
 sg13g2_dfrbp_1 _2360_ (.CLK(net924),
    .RESET_B(net1037),
    .D(\u_top_module.u_filter.shift_reg[71] ),
    .Q_N(_1037_),
    .Q(\u_top_module.u_filter.shift_reg[72] ));
 sg13g2_dfrbp_1 _2361_ (.CLK(net924),
    .RESET_B(net1008),
    .D(\u_top_module.u_filter.shift_reg[72] ),
    .Q_N(_1038_),
    .Q(\u_top_module.u_filter.shift_reg[73] ));
 sg13g2_dfrbp_1 _2362_ (.CLK(net917),
    .RESET_B(net1008),
    .D(\u_top_module.u_filter.shift_reg[73] ),
    .Q_N(_1039_),
    .Q(\u_top_module.u_filter.shift_reg[74] ));
 sg13g2_dfrbp_1 _2363_ (.CLK(net917),
    .RESET_B(net1008),
    .D(\u_top_module.u_filter.shift_reg[74] ),
    .Q_N(_1040_),
    .Q(\u_top_module.u_filter.shift_reg[75] ));
 sg13g2_dfrbp_1 _2364_ (.CLK(net918),
    .RESET_B(net1009),
    .D(\u_top_module.u_filter.shift_reg[75] ),
    .Q_N(_1041_),
    .Q(\u_top_module.u_filter.shift_reg[76] ));
 sg13g2_dfrbp_1 _2365_ (.CLK(net917),
    .RESET_B(net1008),
    .D(\u_top_module.u_filter.shift_reg[76] ),
    .Q_N(_1042_),
    .Q(\u_top_module.u_filter.shift_reg[77] ));
 sg13g2_dfrbp_1 _2366_ (.CLK(net917),
    .RESET_B(net1008),
    .D(\u_top_module.u_filter.shift_reg[77] ),
    .Q_N(_1043_),
    .Q(\u_top_module.u_filter.shift_reg[78] ));
 sg13g2_dfrbp_1 _2367_ (.CLK(net917),
    .RESET_B(net1008),
    .D(\u_top_module.u_filter.shift_reg[78] ),
    .Q_N(_1044_),
    .Q(\u_top_module.u_filter.shift_reg[79] ));
 sg13g2_dfrbp_1 _2368_ (.CLK(net917),
    .RESET_B(net1008),
    .D(\u_top_module.u_filter.shift_reg[79] ),
    .Q_N(_1045_),
    .Q(\u_top_module.u_filter.shift_reg[80] ));
 sg13g2_dfrbp_1 _2369_ (.CLK(net917),
    .RESET_B(net1008),
    .D(\u_top_module.u_filter.shift_reg[80] ),
    .Q_N(_1046_),
    .Q(\u_top_module.u_filter.shift_reg[81] ));
 sg13g2_dfrbp_1 _2370_ (.CLK(net917),
    .RESET_B(net1007),
    .D(\u_top_module.u_filter.shift_reg[81] ),
    .Q_N(_1047_),
    .Q(\u_top_module.u_filter.shift_reg[82] ));
 sg13g2_dfrbp_1 _2371_ (.CLK(net919),
    .RESET_B(net1007),
    .D(\u_top_module.u_filter.shift_reg[82] ),
    .Q_N(_1048_),
    .Q(\u_top_module.u_filter.shift_reg[83] ));
 sg13g2_dfrbp_1 _2372_ (.CLK(net915),
    .RESET_B(net1006),
    .D(\u_top_module.u_filter.shift_reg[83] ),
    .Q_N(_1049_),
    .Q(\u_top_module.u_filter.shift_reg[84] ));
 sg13g2_dfrbp_1 _2373_ (.CLK(net915),
    .RESET_B(net1006),
    .D(\u_top_module.u_filter.shift_reg[84] ),
    .Q_N(_1050_),
    .Q(\u_top_module.u_filter.shift_reg[85] ));
 sg13g2_dfrbp_1 _2374_ (.CLK(net915),
    .RESET_B(net1006),
    .D(\u_top_module.u_filter.shift_reg[85] ),
    .Q_N(_1051_),
    .Q(\u_top_module.u_filter.shift_reg[86] ));
 sg13g2_dfrbp_1 _2375_ (.CLK(net915),
    .RESET_B(net1006),
    .D(\u_top_module.u_filter.shift_reg[86] ),
    .Q_N(_1052_),
    .Q(\u_top_module.u_filter.shift_reg[87] ));
 sg13g2_dfrbp_1 _2376_ (.CLK(net915),
    .RESET_B(net1006),
    .D(\u_top_module.u_filter.shift_reg[87] ),
    .Q_N(_1053_),
    .Q(\u_top_module.u_filter.shift_reg[88] ));
 sg13g2_dfrbp_1 _2377_ (.CLK(net907),
    .RESET_B(net998),
    .D(\u_top_module.u_filter.shift_reg[88] ),
    .Q_N(_1054_),
    .Q(\u_top_module.u_filter.shift_reg[89] ));
 sg13g2_dfrbp_1 _2378_ (.CLK(net907),
    .RESET_B(net998),
    .D(\u_top_module.u_filter.shift_reg[89] ),
    .Q_N(_1055_),
    .Q(\u_top_module.u_filter.shift_reg[90] ));
 sg13g2_dfrbp_1 _2379_ (.CLK(net907),
    .RESET_B(net998),
    .D(\u_top_module.u_filter.shift_reg[90] ),
    .Q_N(_1056_),
    .Q(\u_top_module.u_filter.shift_reg[91] ));
 sg13g2_dfrbp_1 _2380_ (.CLK(net907),
    .RESET_B(net998),
    .D(\u_top_module.u_filter.shift_reg[91] ),
    .Q_N(_1057_),
    .Q(\u_top_module.u_filter.shift_reg[92] ));
 sg13g2_dfrbp_1 _2381_ (.CLK(net915),
    .RESET_B(net1006),
    .D(\u_top_module.u_filter.shift_reg[92] ),
    .Q_N(_1058_),
    .Q(\u_top_module.u_filter.shift_reg[93] ));
 sg13g2_dfrbp_1 _2382_ (.CLK(net915),
    .RESET_B(net1006),
    .D(\u_top_module.u_filter.shift_reg[93] ),
    .Q_N(_1059_),
    .Q(\u_top_module.u_filter.shift_reg[94] ));
 sg13g2_dfrbp_1 _2383_ (.CLK(net915),
    .RESET_B(net1006),
    .D(\u_top_module.u_filter.shift_reg[94] ),
    .Q_N(_1060_),
    .Q(\u_top_module.u_filter.shift_reg[95] ));
 sg13g2_dfrbp_1 _2384_ (.CLK(net916),
    .RESET_B(net1005),
    .D(\u_top_module.u_filter.shift_reg[95] ),
    .Q_N(_1061_),
    .Q(\u_top_module.u_filter.shift_reg[96] ));
 sg13g2_dfrbp_1 _2385_ (.CLK(net911),
    .RESET_B(net1001),
    .D(\u_top_module.u_filter.shift_reg[96] ),
    .Q_N(_1062_),
    .Q(\u_top_module.u_filter.shift_reg[97] ));
 sg13g2_dfrbp_1 _2386_ (.CLK(net911),
    .RESET_B(net1001),
    .D(\u_top_module.u_filter.shift_reg[97] ),
    .Q_N(_1063_),
    .Q(\u_top_module.u_filter.shift_reg[98] ));
 sg13g2_dfrbp_1 _2387_ (.CLK(net911),
    .RESET_B(net1001),
    .D(\u_top_module.u_filter.shift_reg[98] ),
    .Q_N(_1064_),
    .Q(\u_top_module.u_filter.shift_reg[99] ));
 sg13g2_dfrbp_1 _2388_ (.CLK(net911),
    .RESET_B(net1000),
    .D(\u_top_module.u_filter.shift_reg[99] ),
    .Q_N(_1065_),
    .Q(\u_top_module.u_filter.shift_reg[100] ));
 sg13g2_dfrbp_1 _2389_ (.CLK(net910),
    .RESET_B(net1000),
    .D(\u_top_module.u_filter.shift_reg[100] ),
    .Q_N(_1066_),
    .Q(\u_top_module.u_filter.shift_reg[101] ));
 sg13g2_dfrbp_1 _2390_ (.CLK(net910),
    .RESET_B(net1000),
    .D(\u_top_module.u_filter.shift_reg[101] ),
    .Q_N(_1067_),
    .Q(\u_top_module.u_filter.shift_reg[102] ));
 sg13g2_dfrbp_1 _2391_ (.CLK(net910),
    .RESET_B(net1000),
    .D(\u_top_module.u_filter.shift_reg[102] ),
    .Q_N(_1068_),
    .Q(\u_top_module.u_filter.shift_reg[103] ));
 sg13g2_dfrbp_1 _2392_ (.CLK(net910),
    .RESET_B(net1000),
    .D(\u_top_module.u_filter.shift_reg[103] ),
    .Q_N(_1069_),
    .Q(\u_top_module.u_filter.shift_reg[104] ));
 sg13g2_dfrbp_1 _2393_ (.CLK(net910),
    .RESET_B(net1000),
    .D(\u_top_module.u_filter.shift_reg[104] ),
    .Q_N(_1070_),
    .Q(\u_top_module.u_filter.shift_reg[105] ));
 sg13g2_dfrbp_1 _2394_ (.CLK(net914),
    .RESET_B(net1000),
    .D(\u_top_module.u_filter.shift_reg[105] ),
    .Q_N(_1071_),
    .Q(\u_top_module.u_filter.shift_reg[106] ));
 sg13g2_dfrbp_1 _2395_ (.CLK(net914),
    .RESET_B(net989),
    .D(\u_top_module.u_filter.shift_reg[106] ),
    .Q_N(_1072_),
    .Q(\u_top_module.u_filter.shift_reg[107] ));
 sg13g2_dfrbp_1 _2396_ (.CLK(net900),
    .RESET_B(net989),
    .D(\u_top_module.u_filter.shift_reg[107] ),
    .Q_N(_1073_),
    .Q(\u_top_module.u_filter.shift_reg[108] ));
 sg13g2_dfrbp_1 _2397_ (.CLK(net900),
    .RESET_B(net989),
    .D(\u_top_module.u_filter.shift_reg[108] ),
    .Q_N(_1074_),
    .Q(\u_top_module.u_filter.shift_reg[109] ));
 sg13g2_dfrbp_1 _2398_ (.CLK(net900),
    .RESET_B(net989),
    .D(\u_top_module.u_filter.shift_reg[109] ),
    .Q_N(_1075_),
    .Q(\u_top_module.u_filter.shift_reg[110] ));
 sg13g2_dfrbp_1 _2399_ (.CLK(net900),
    .RESET_B(net989),
    .D(\u_top_module.u_filter.shift_reg[110] ),
    .Q_N(_1076_),
    .Q(\u_top_module.u_filter.shift_reg[111] ));
 sg13g2_dfrbp_1 _2400_ (.CLK(net900),
    .RESET_B(net989),
    .D(\u_top_module.u_filter.shift_reg[111] ),
    .Q_N(_1077_),
    .Q(\u_top_module.u_filter.shift_reg[112] ));
 sg13g2_dfrbp_1 _2401_ (.CLK(net899),
    .RESET_B(net986),
    .D(\u_top_module.u_filter.shift_reg[112] ),
    .Q_N(_1078_),
    .Q(\u_top_module.u_filter.shift_reg[113] ));
 sg13g2_dfrbp_1 _2402_ (.CLK(net899),
    .RESET_B(net986),
    .D(\u_top_module.u_filter.shift_reg[113] ),
    .Q_N(_1079_),
    .Q(\u_top_module.u_filter.shift_reg[114] ));
 sg13g2_dfrbp_1 _2403_ (.CLK(net898),
    .RESET_B(net986),
    .D(\u_top_module.u_filter.shift_reg[114] ),
    .Q_N(_1080_),
    .Q(\u_top_module.u_filter.shift_reg[115] ));
 sg13g2_dfrbp_1 _2404_ (.CLK(net897),
    .RESET_B(net986),
    .D(\u_top_module.u_filter.shift_reg[115] ),
    .Q_N(_1081_),
    .Q(\u_top_module.u_filter.shift_reg[116] ));
 sg13g2_dfrbp_1 _2405_ (.CLK(net897),
    .RESET_B(net987),
    .D(\u_top_module.u_filter.shift_reg[116] ),
    .Q_N(_1082_),
    .Q(\u_top_module.u_filter.shift_reg[117] ));
 sg13g2_dfrbp_1 _2406_ (.CLK(net897),
    .RESET_B(net987),
    .D(\u_top_module.u_filter.shift_reg[117] ),
    .Q_N(_1083_),
    .Q(\u_top_module.u_filter.shift_reg[118] ));
 sg13g2_dfrbp_1 _2407_ (.CLK(net897),
    .RESET_B(net987),
    .D(\u_top_module.u_filter.shift_reg[118] ),
    .Q_N(_1084_),
    .Q(\u_top_module.u_filter.shift_reg[119] ));
 sg13g2_dfrbp_1 _2408_ (.CLK(net897),
    .RESET_B(net987),
    .D(\u_top_module.u_filter.shift_reg[119] ),
    .Q_N(_1085_),
    .Q(\u_top_module.u_filter.shift_reg[120] ));
 sg13g2_dfrbp_1 _2409_ (.CLK(net897),
    .RESET_B(net987),
    .D(\u_top_module.u_filter.shift_reg[120] ),
    .Q_N(_1086_),
    .Q(\u_top_module.u_filter.shift_reg[121] ));
 sg13g2_dfrbp_1 _2410_ (.CLK(net898),
    .RESET_B(net987),
    .D(\u_top_module.u_filter.shift_reg[121] ),
    .Q_N(_1087_),
    .Q(\u_top_module.u_filter.shift_reg[122] ));
 sg13g2_dfrbp_1 _2411_ (.CLK(net898),
    .RESET_B(net988),
    .D(\u_top_module.u_filter.shift_reg[122] ),
    .Q_N(_1088_),
    .Q(\u_top_module.u_filter.shift_reg[123] ));
 sg13g2_dfrbp_1 _2412_ (.CLK(net901),
    .RESET_B(net990),
    .D(\u_top_module.u_filter.shift_reg[123] ),
    .Q_N(_1089_),
    .Q(\u_top_module.u_filter.shift_reg[124] ));
 sg13g2_dfrbp_1 _2413_ (.CLK(net901),
    .RESET_B(net990),
    .D(\u_top_module.u_filter.shift_reg[124] ),
    .Q_N(_1090_),
    .Q(\u_top_module.u_filter.shift_reg[125] ));
 sg13g2_dfrbp_1 _2414_ (.CLK(net901),
    .RESET_B(net990),
    .D(\u_top_module.u_filter.shift_reg[125] ),
    .Q_N(_1091_),
    .Q(\u_top_module.u_filter.shift_reg[126] ));
 sg13g2_dfrbp_1 _2415_ (.CLK(net901),
    .RESET_B(net989),
    .D(\u_top_module.u_filter.shift_reg[126] ),
    .Q_N(_1092_),
    .Q(\u_top_module.u_filter.shift_reg[127] ));
 sg13g2_dfrbp_1 _2416_ (.CLK(net906),
    .RESET_B(net997),
    .D(\u_top_module.u_filter.shift_reg[127] ),
    .Q_N(_1093_),
    .Q(\u_top_module.u_filter.shift_reg[128] ));
 sg13g2_dfrbp_1 _2417_ (.CLK(net902),
    .RESET_B(net993),
    .D(\u_top_module.u_filter.shift_reg[128] ),
    .Q_N(_1094_),
    .Q(\u_top_module.u_filter.shift_reg[129] ));
 sg13g2_dfrbp_1 _2418_ (.CLK(net905),
    .RESET_B(net993),
    .D(\u_top_module.u_filter.shift_reg[129] ),
    .Q_N(_1095_),
    .Q(\u_top_module.u_filter.shift_reg[130] ));
 sg13g2_dfrbp_1 _2419_ (.CLK(net902),
    .RESET_B(net992),
    .D(\u_top_module.u_filter.shift_reg[130] ),
    .Q_N(_1096_),
    .Q(\u_top_module.u_filter.shift_reg[131] ));
 sg13g2_dfrbp_1 _2420_ (.CLK(net902),
    .RESET_B(net992),
    .D(\u_top_module.u_filter.shift_reg[131] ),
    .Q_N(_1097_),
    .Q(\u_top_module.u_filter.shift_reg[132] ));
 sg13g2_dfrbp_1 _2421_ (.CLK(net902),
    .RESET_B(net992),
    .D(\u_top_module.u_filter.shift_reg[132] ),
    .Q_N(_1098_),
    .Q(\u_top_module.u_filter.shift_reg[133] ));
 sg13g2_dfrbp_1 _2422_ (.CLK(net902),
    .RESET_B(net992),
    .D(\u_top_module.u_filter.shift_reg[133] ),
    .Q_N(_1099_),
    .Q(\u_top_module.u_filter.shift_reg[134] ));
 sg13g2_dfrbp_1 _2423_ (.CLK(net902),
    .RESET_B(net992),
    .D(\u_top_module.u_filter.shift_reg[134] ),
    .Q_N(_1100_),
    .Q(\u_top_module.u_filter.shift_reg[135] ));
 sg13g2_dfrbp_1 _2424_ (.CLK(net902),
    .RESET_B(net992),
    .D(\u_top_module.u_filter.shift_reg[135] ),
    .Q_N(_1101_),
    .Q(\u_top_module.u_filter.shift_reg[136] ));
 sg13g2_dfrbp_1 _2425_ (.CLK(net902),
    .RESET_B(net992),
    .D(\u_top_module.u_filter.shift_reg[136] ),
    .Q_N(_1102_),
    .Q(\u_top_module.u_filter.shift_reg[137] ));
 sg13g2_dfrbp_1 _2426_ (.CLK(net903),
    .RESET_B(net992),
    .D(\u_top_module.u_filter.shift_reg[137] ),
    .Q_N(_1103_),
    .Q(\u_top_module.u_filter.shift_reg[138] ));
 sg13g2_dfrbp_1 _2427_ (.CLK(net903),
    .RESET_B(net994),
    .D(\u_top_module.u_filter.shift_reg[138] ),
    .Q_N(_1104_),
    .Q(\u_top_module.u_filter.shift_reg[139] ));
 sg13g2_dfrbp_1 _2428_ (.CLK(net903),
    .RESET_B(net994),
    .D(\u_top_module.u_filter.shift_reg[139] ),
    .Q_N(_1105_),
    .Q(\u_top_module.u_filter.shift_reg[140] ));
 sg13g2_dfrbp_1 _2429_ (.CLK(net903),
    .RESET_B(net994),
    .D(\u_top_module.u_filter.shift_reg[140] ),
    .Q_N(_1106_),
    .Q(\u_top_module.u_filter.shift_reg[141] ));
 sg13g2_dfrbp_1 _2430_ (.CLK(net903),
    .RESET_B(net994),
    .D(\u_top_module.u_filter.shift_reg[141] ),
    .Q_N(_1107_),
    .Q(\u_top_module.u_filter.shift_reg[142] ));
 sg13g2_dfrbp_1 _2431_ (.CLK(net903),
    .RESET_B(net994),
    .D(\u_top_module.u_filter.shift_reg[142] ),
    .Q_N(_1108_),
    .Q(\u_top_module.u_filter.shift_reg[143] ));
 sg13g2_dfrbp_1 _2432_ (.CLK(net904),
    .RESET_B(net994),
    .D(\u_top_module.u_filter.shift_reg[143] ),
    .Q_N(_1109_),
    .Q(\u_top_module.u_filter.shift_reg[144] ));
 sg13g2_dfrbp_1 _2433_ (.CLK(net903),
    .RESET_B(net994),
    .D(\u_top_module.u_filter.shift_reg[144] ),
    .Q_N(_1110_),
    .Q(\u_top_module.u_filter.shift_reg[145] ));
 sg13g2_dfrbp_1 _2434_ (.CLK(net903),
    .RESET_B(net994),
    .D(\u_top_module.u_filter.shift_reg[145] ),
    .Q_N(_1111_),
    .Q(\u_top_module.u_filter.shift_reg[146] ));
 sg13g2_dfrbp_1 _2435_ (.CLK(net904),
    .RESET_B(net995),
    .D(\u_top_module.u_filter.shift_reg[146] ),
    .Q_N(_1112_),
    .Q(\u_top_module.u_filter.shift_reg[147] ));
 sg13g2_dfrbp_1 _2436_ (.CLK(net904),
    .RESET_B(net995),
    .D(\u_top_module.u_filter.shift_reg[147] ),
    .Q_N(_1113_),
    .Q(\u_top_module.u_filter.shift_reg[148] ));
 sg13g2_dfrbp_1 _2437_ (.CLK(net904),
    .RESET_B(net995),
    .D(\u_top_module.u_filter.shift_reg[148] ),
    .Q_N(_1114_),
    .Q(\u_top_module.u_filter.shift_reg[149] ));
 sg13g2_dfrbp_1 _2438_ (.CLK(net904),
    .RESET_B(net995),
    .D(\u_top_module.u_filter.shift_reg[149] ),
    .Q_N(_1115_),
    .Q(\u_top_module.u_filter.shift_reg[150] ));
 sg13g2_dfrbp_1 _2439_ (.CLK(net904),
    .RESET_B(net995),
    .D(\u_top_module.u_filter.shift_reg[150] ),
    .Q_N(_1116_),
    .Q(\u_top_module.u_filter.shift_reg[151] ));
 sg13g2_dfrbp_1 _2440_ (.CLK(net908),
    .RESET_B(net998),
    .D(\u_top_module.u_filter.shift_reg[151] ),
    .Q_N(_1117_),
    .Q(\u_top_module.u_filter.shift_reg[152] ));
 sg13g2_dfrbp_1 _2441_ (.CLK(net908),
    .RESET_B(net998),
    .D(\u_top_module.u_filter.shift_reg[152] ),
    .Q_N(_1118_),
    .Q(\u_top_module.u_filter.shift_reg[153] ));
 sg13g2_dfrbp_1 _2442_ (.CLK(net907),
    .RESET_B(net998),
    .D(\u_top_module.u_filter.shift_reg[153] ),
    .Q_N(_1119_),
    .Q(\u_top_module.u_filter.shift_reg[154] ));
 sg13g2_dfrbp_1 _2443_ (.CLK(net907),
    .RESET_B(net998),
    .D(\u_top_module.u_filter.shift_reg[154] ),
    .Q_N(_1120_),
    .Q(\u_top_module.u_filter.shift_reg[155] ));
 sg13g2_dfrbp_1 _2444_ (.CLK(net906),
    .RESET_B(net997),
    .D(\u_top_module.u_filter.shift_reg[155] ),
    .Q_N(_1121_),
    .Q(\u_top_module.u_filter.shift_reg[156] ));
 sg13g2_dfrbp_1 _2445_ (.CLK(net906),
    .RESET_B(net997),
    .D(\u_top_module.u_filter.shift_reg[156] ),
    .Q_N(_1122_),
    .Q(\u_top_module.u_filter.shift_reg[157] ));
 sg13g2_dfrbp_1 _2446_ (.CLK(net906),
    .RESET_B(net997),
    .D(\u_top_module.u_filter.shift_reg[157] ),
    .Q_N(_1123_),
    .Q(\u_top_module.u_filter.shift_reg[158] ));
 sg13g2_dfrbp_1 _2447_ (.CLK(net906),
    .RESET_B(net997),
    .D(\u_top_module.u_filter.shift_reg[158] ),
    .Q_N(_1124_),
    .Q(\u_top_module.u_filter.shift_reg[159] ));
 sg13g2_dfrbp_1 _2448_ (.CLK(net906),
    .RESET_B(net997),
    .D(\u_top_module.u_filter.shift_reg[159] ),
    .Q_N(_1125_),
    .Q(\u_top_module.u_filter.shift_reg[160] ));
 sg13g2_dfrbp_1 _2449_ (.CLK(net916),
    .RESET_B(net1005),
    .D(\u_top_module.u_filter.shift_reg[160] ),
    .Q_N(_1126_),
    .Q(\u_top_module.u_filter.shift_reg[161] ));
 sg13g2_dfrbp_1 _2450_ (.CLK(net916),
    .RESET_B(net1005),
    .D(\u_top_module.u_filter.shift_reg[161] ),
    .Q_N(_1127_),
    .Q(\u_top_module.u_filter.shift_reg[162] ));
 sg13g2_dfrbp_1 _2451_ (.CLK(net916),
    .RESET_B(net1007),
    .D(\u_top_module.u_filter.shift_reg[162] ),
    .Q_N(_1128_),
    .Q(\u_top_module.u_filter.shift_reg[163] ));
 sg13g2_dfrbp_1 _2452_ (.CLK(net918),
    .RESET_B(net1005),
    .D(\u_top_module.u_filter.shift_reg[163] ),
    .Q_N(_1129_),
    .Q(\u_top_module.u_filter.shift_reg[164] ));
 sg13g2_dfrbp_1 _2453_ (.CLK(net918),
    .RESET_B(net1009),
    .D(\u_top_module.u_filter.shift_reg[164] ),
    .Q_N(_1130_),
    .Q(\u_top_module.u_filter.shift_reg[165] ));
 sg13g2_dfrbp_1 _2454_ (.CLK(net918),
    .RESET_B(net1009),
    .D(\u_top_module.u_filter.shift_reg[165] ),
    .Q_N(_1131_),
    .Q(\u_top_module.u_filter.shift_reg[166] ));
 sg13g2_dfrbp_1 _2455_ (.CLK(net918),
    .RESET_B(net1009),
    .D(\u_top_module.u_filter.shift_reg[166] ),
    .Q_N(_1132_),
    .Q(\u_top_module.u_filter.shift_reg[167] ));
 sg13g2_dfrbp_1 _2456_ (.CLK(net916),
    .RESET_B(net1005),
    .D(\u_top_module.u_filter.shift_reg[167] ),
    .Q_N(_1133_),
    .Q(\u_top_module.u_filter.shift_reg[168] ));
 sg13g2_dfrbp_1 _2457_ (.CLK(net916),
    .RESET_B(net1005),
    .D(\u_top_module.u_filter.shift_reg[168] ),
    .Q_N(_1134_),
    .Q(\u_top_module.u_filter.shift_reg[169] ));
 sg13g2_dfrbp_1 _2458_ (.CLK(net916),
    .RESET_B(net1005),
    .D(\u_top_module.u_filter.shift_reg[169] ),
    .Q_N(_1135_),
    .Q(\u_top_module.u_filter.shift_reg[170] ));
 sg13g2_dfrbp_1 _2459_ (.CLK(net916),
    .RESET_B(net1005),
    .D(\u_top_module.u_filter.shift_reg[170] ),
    .Q_N(_1136_),
    .Q(\u_top_module.u_filter.shift_reg[171] ));
 sg13g2_dfrbp_1 _2460_ (.CLK(net907),
    .RESET_B(net997),
    .D(\u_top_module.u_filter.shift_reg[171] ),
    .Q_N(_1137_),
    .Q(\u_top_module.u_filter.shift_reg[172] ));
 sg13g2_dfrbp_1 _2461_ (.CLK(net906),
    .RESET_B(net997),
    .D(\u_top_module.u_filter.shift_reg[172] ),
    .Q_N(_1138_),
    .Q(\u_top_module.u_filter.shift_reg[173] ));
 sg13g2_dfrbp_1 _2462_ (.CLK(net906),
    .RESET_B(net993),
    .D(\u_top_module.u_filter.shift_reg[173] ),
    .Q_N(_1139_),
    .Q(\u_top_module.u_filter.shift_reg[174] ));
 sg13g2_dfrbp_1 _2463_ (.CLK(net905),
    .RESET_B(net993),
    .D(\u_top_module.u_filter.shift_reg[174] ),
    .Q_N(_1140_),
    .Q(\u_top_module.u_filter.shift_reg[175] ));
 sg13g2_dfrbp_1 _2464_ (.CLK(net905),
    .RESET_B(net988),
    .D(\u_top_module.u_filter.shift_reg[175] ),
    .Q_N(_1141_),
    .Q(\u_top_module.u_filter.shift_reg[176] ));
 sg13g2_dfrbp_1 _2465_ (.CLK(net898),
    .RESET_B(net987),
    .D(\u_top_module.u_filter.shift_reg[176] ),
    .Q_N(_1142_),
    .Q(\u_top_module.u_filter.shift_reg[177] ));
 sg13g2_dfrbp_1 _2466_ (.CLK(net897),
    .RESET_B(net988),
    .D(\u_top_module.u_filter.shift_reg[177] ),
    .Q_N(_1143_),
    .Q(\u_top_module.u_filter.shift_reg[178] ));
 sg13g2_dfrbp_1 _2467_ (.CLK(net897),
    .RESET_B(net987),
    .D(\u_top_module.u_filter.shift_reg[178] ),
    .Q_N(_1144_),
    .Q(\u_top_module.u_filter.shift_reg[179] ));
 sg13g2_dfrbp_1 _2468_ (.CLK(net899),
    .RESET_B(net986),
    .D(\u_top_module.u_filter.shift_reg[179] ),
    .Q_N(_1145_),
    .Q(\u_top_module.u_filter.shift_reg[180] ));
 sg13g2_dfrbp_1 _2469_ (.CLK(net899),
    .RESET_B(net986),
    .D(\u_top_module.u_filter.shift_reg[180] ),
    .Q_N(_1146_),
    .Q(\u_top_module.u_filter.shift_reg[181] ));
 sg13g2_dfrbp_1 _2470_ (.CLK(net899),
    .RESET_B(net986),
    .D(\u_top_module.u_filter.shift_reg[181] ),
    .Q_N(_1147_),
    .Q(\u_top_module.u_filter.shift_reg[182] ));
 sg13g2_dfrbp_1 _2471_ (.CLK(net899),
    .RESET_B(net991),
    .D(\u_top_module.u_filter.shift_reg[182] ),
    .Q_N(_1148_),
    .Q(\u_top_module.u_filter.shift_reg[183] ));
 sg13g2_dfrbp_1 _2472_ (.CLK(net900),
    .RESET_B(net986),
    .D(\u_top_module.u_filter.shift_reg[183] ),
    .Q_N(_1149_),
    .Q(\u_top_module.u_filter.shift_reg[184] ));
 sg13g2_dfrbp_1 _2473_ (.CLK(net900),
    .RESET_B(net989),
    .D(\u_top_module.u_filter.shift_reg[184] ),
    .Q_N(_1150_),
    .Q(\u_top_module.u_filter.shift_reg[185] ));
 sg13g2_dfrbp_1 _2474_ (.CLK(net901),
    .RESET_B(net990),
    .D(\u_top_module.u_filter.shift_reg[185] ),
    .Q_N(_1151_),
    .Q(\u_top_module.u_filter.shift_reg[186] ));
 sg13g2_dfrbp_1 _2475_ (.CLK(net901),
    .RESET_B(net990),
    .D(\u_top_module.u_filter.shift_reg[186] ),
    .Q_N(_1152_),
    .Q(\u_top_module.u_filter.shift_reg[187] ));
 sg13g2_dfrbp_1 _2476_ (.CLK(net901),
    .RESET_B(net990),
    .D(\u_top_module.u_filter.shift_reg[187] ),
    .Q_N(_1153_),
    .Q(\u_top_module.u_filter.shift_reg[188] ));
 sg13g2_dfrbp_1 _2477_ (.CLK(net911),
    .RESET_B(net1001),
    .D(\u_top_module.u_filter.shift_reg[188] ),
    .Q_N(_1154_),
    .Q(\u_top_module.u_filter.shift_reg[189] ));
 sg13g2_dfrbp_1 _2478_ (.CLK(net911),
    .RESET_B(net1001),
    .D(\u_top_module.u_filter.shift_reg[189] ),
    .Q_N(_1155_),
    .Q(\u_top_module.u_filter.shift_reg[190] ));
 sg13g2_dfrbp_1 _2479_ (.CLK(net911),
    .RESET_B(net1000),
    .D(\u_top_module.u_filter.shift_reg[190] ),
    .Q_N(_1156_),
    .Q(\u_top_module.u_filter.shift_reg[191] ));
 sg13g2_dfrbp_1 _2480_ (.CLK(net918),
    .RESET_B(net1001),
    .D(\u_top_module.u_filter.shift_reg[191] ),
    .Q_N(_1157_),
    .Q(\u_top_module.u_filter.shift_reg[192] ));
 sg13g2_dfrbp_1 _2481_ (.CLK(net927),
    .RESET_B(net1034),
    .D(\u_top_module.u_filter.shift_reg[192] ),
    .Q_N(_1158_),
    .Q(\u_top_module.u_filter.shift_reg[193] ));
 sg13g2_dfrbp_1 _2482_ (.CLK(net927),
    .RESET_B(net1036),
    .D(\u_top_module.u_filter.shift_reg[193] ),
    .Q_N(_1159_),
    .Q(\u_top_module.u_filter.shift_reg[194] ));
 sg13g2_dfrbp_1 _2483_ (.CLK(net922),
    .RESET_B(net1031),
    .D(\u_top_module.u_filter.shift_reg[194] ),
    .Q_N(_1160_),
    .Q(\u_top_module.u_filter.shift_reg[195] ));
 sg13g2_dfrbp_1 _2484_ (.CLK(net922),
    .RESET_B(net1031),
    .D(\u_top_module.u_filter.shift_reg[195] ),
    .Q_N(_1161_),
    .Q(\u_top_module.u_filter.shift_reg[196] ));
 sg13g2_dfrbp_1 _2485_ (.CLK(net929),
    .RESET_B(net1030),
    .D(\u_top_module.u_filter.shift_reg[196] ),
    .Q_N(_1162_),
    .Q(\u_top_module.u_filter.shift_reg[197] ));
 sg13g2_dfrbp_1 _2486_ (.CLK(net922),
    .RESET_B(net1030),
    .D(\u_top_module.u_filter.shift_reg[197] ),
    .Q_N(_1163_),
    .Q(\u_top_module.u_filter.shift_reg[198] ));
 sg13g2_dfrbp_1 _2487_ (.CLK(net929),
    .RESET_B(net1030),
    .D(\u_top_module.u_filter.shift_reg[198] ),
    .Q_N(_1164_),
    .Q(\u_top_module.u_filter.shift_reg[199] ));
 sg13g2_dfrbp_1 _2488_ (.CLK(net922),
    .RESET_B(net1030),
    .D(\u_top_module.u_filter.shift_reg[199] ),
    .Q_N(_1165_),
    .Q(\u_top_module.u_filter.shift_reg[200] ));
 sg13g2_dfrbp_1 _2489_ (.CLK(net933),
    .RESET_B(net1030),
    .D(\u_top_module.u_filter.shift_reg[200] ),
    .Q_N(_1166_),
    .Q(\u_top_module.u_filter.shift_reg[201] ));
 sg13g2_dfrbp_1 _2490_ (.CLK(net933),
    .RESET_B(net1031),
    .D(\u_top_module.u_filter.shift_reg[201] ),
    .Q_N(_1167_),
    .Q(\u_top_module.u_filter.shift_reg[202] ));
 sg13g2_dfrbp_1 _2491_ (.CLK(net933),
    .RESET_B(net1030),
    .D(\u_top_module.u_filter.shift_reg[202] ),
    .Q_N(_1168_),
    .Q(\u_top_module.u_filter.shift_reg[203] ));
 sg13g2_dfrbp_1 _2492_ (.CLK(net922),
    .RESET_B(net1031),
    .D(\u_top_module.u_filter.shift_reg[203] ),
    .Q_N(_1169_),
    .Q(\u_top_module.u_filter.shift_reg[204] ));
 sg13g2_dfrbp_1 _2493_ (.CLK(net922),
    .RESET_B(net1030),
    .D(\u_top_module.u_filter.shift_reg[204] ),
    .Q_N(_1170_),
    .Q(\u_top_module.u_filter.shift_reg[205] ));
 sg13g2_dfrbp_1 _2494_ (.CLK(net927),
    .RESET_B(net1030),
    .D(\u_top_module.u_filter.shift_reg[205] ),
    .Q_N(_1171_),
    .Q(\u_top_module.u_filter.shift_reg[206] ));
 sg13g2_dfrbp_1 _2495_ (.CLK(net927),
    .RESET_B(net1036),
    .D(\u_top_module.u_filter.shift_reg[206] ),
    .Q_N(_1172_),
    .Q(\u_top_module.u_filter.shift_reg[207] ));
 sg13g2_dfrbp_1 _2496_ (.CLK(net927),
    .RESET_B(net1036),
    .D(\u_top_module.u_filter.shift_reg[207] ),
    .Q_N(_1173_),
    .Q(\u_top_module.u_filter.shift_reg[208] ));
 sg13g2_dfrbp_1 _2497_ (.CLK(net935),
    .RESET_B(net1036),
    .D(\u_top_module.u_filter.shift_reg[208] ),
    .Q_N(_1174_),
    .Q(\u_top_module.u_filter.shift_reg[209] ));
 sg13g2_dfrbp_1 _2498_ (.CLK(net935),
    .RESET_B(net1036),
    .D(\u_top_module.u_filter.shift_reg[209] ),
    .Q_N(_1175_),
    .Q(\u_top_module.u_filter.shift_reg[210] ));
 sg13g2_dfrbp_1 _2499_ (.CLK(net935),
    .RESET_B(net1045),
    .D(\u_top_module.u_filter.shift_reg[210] ),
    .Q_N(_1176_),
    .Q(\u_top_module.u_filter.shift_reg[211] ));
 sg13g2_dfrbp_1 _2500_ (.CLK(net934),
    .RESET_B(net1043),
    .D(\u_top_module.u_filter.shift_reg[211] ),
    .Q_N(_1177_),
    .Q(\u_top_module.u_filter.shift_reg[212] ));
 sg13g2_dfrbp_1 _2501_ (.CLK(net935),
    .RESET_B(net1043),
    .D(\u_top_module.u_filter.shift_reg[212] ),
    .Q_N(_1178_),
    .Q(\u_top_module.u_filter.shift_reg[213] ));
 sg13g2_dfrbp_1 _2502_ (.CLK(net940),
    .RESET_B(net1043),
    .D(\u_top_module.u_filter.shift_reg[213] ),
    .Q_N(_1179_),
    .Q(\u_top_module.u_filter.shift_reg[214] ));
 sg13g2_dfrbp_1 _2503_ (.CLK(net940),
    .RESET_B(net1044),
    .D(\u_top_module.u_filter.shift_reg[214] ),
    .Q_N(_1180_),
    .Q(\u_top_module.u_filter.shift_reg[215] ));
 sg13g2_dfrbp_1 _2504_ (.CLK(net936),
    .RESET_B(net1045),
    .D(\u_top_module.u_filter.shift_reg[215] ),
    .Q_N(_1181_),
    .Q(\u_top_module.u_filter.shift_reg[216] ));
 sg13g2_dfrbp_1 _2505_ (.CLK(net936),
    .RESET_B(net1045),
    .D(\u_top_module.u_filter.shift_reg[216] ),
    .Q_N(_1182_),
    .Q(\u_top_module.u_filter.shift_reg[217] ));
 sg13g2_dfrbp_1 _2506_ (.CLK(net936),
    .RESET_B(net1045),
    .D(\u_top_module.u_filter.shift_reg[217] ),
    .Q_N(_1183_),
    .Q(\u_top_module.u_filter.shift_reg[218] ));
 sg13g2_dfrbp_1 _2507_ (.CLK(net936),
    .RESET_B(net1046),
    .D(\u_top_module.u_filter.shift_reg[218] ),
    .Q_N(_1184_),
    .Q(\u_top_module.u_filter.shift_reg[219] ));
 sg13g2_dfrbp_1 _2508_ (.CLK(net936),
    .RESET_B(net1046),
    .D(\u_top_module.u_filter.shift_reg[219] ),
    .Q_N(_1185_),
    .Q(\u_top_module.u_filter.shift_reg[220] ));
 sg13g2_dfrbp_1 _2509_ (.CLK(net937),
    .RESET_B(net1046),
    .D(\u_top_module.u_filter.shift_reg[220] ),
    .Q_N(_1186_),
    .Q(\u_top_module.u_filter.shift_reg[221] ));
 sg13g2_dfrbp_1 _2510_ (.CLK(net937),
    .RESET_B(net1046),
    .D(\u_top_module.u_filter.shift_reg[221] ),
    .Q_N(_1187_),
    .Q(\u_top_module.u_filter.shift_reg[222] ));
 sg13g2_dfrbp_1 _2511_ (.CLK(net938),
    .RESET_B(net1046),
    .D(\u_top_module.u_filter.shift_reg[222] ),
    .Q_N(_1188_),
    .Q(\u_top_module.u_filter.shift_reg[223] ));
 sg13g2_dfrbp_1 _2512_ (.CLK(net938),
    .RESET_B(net1048),
    .D(\u_top_module.u_filter.shift_reg[223] ),
    .Q_N(_1189_),
    .Q(\u_top_module.u_filter.shift_reg[224] ));
 sg13g2_dfrbp_1 _2513_ (.CLK(net938),
    .RESET_B(net1047),
    .D(\u_top_module.u_filter.shift_reg[224] ),
    .Q_N(_1190_),
    .Q(\u_top_module.u_filter.shift_reg[225] ));
 sg13g2_dfrbp_1 _2514_ (.CLK(net938),
    .RESET_B(net1047),
    .D(\u_top_module.u_filter.shift_reg[225] ),
    .Q_N(_1191_),
    .Q(\u_top_module.u_filter.shift_reg[226] ));
 sg13g2_dfrbp_1 _2515_ (.CLK(net938),
    .RESET_B(net1048),
    .D(\u_top_module.u_filter.shift_reg[226] ),
    .Q_N(_1192_),
    .Q(\u_top_module.u_filter.shift_reg[227] ));
 sg13g2_dfrbp_1 _2516_ (.CLK(net938),
    .RESET_B(net1047),
    .D(\u_top_module.u_filter.shift_reg[227] ),
    .Q_N(_1193_),
    .Q(\u_top_module.u_filter.shift_reg[228] ));
 sg13g2_dfrbp_1 _2517_ (.CLK(net938),
    .RESET_B(net1047),
    .D(\u_top_module.u_filter.shift_reg[228] ),
    .Q_N(_1194_),
    .Q(\u_top_module.u_filter.shift_reg[229] ));
 sg13g2_dfrbp_1 _2518_ (.CLK(net939),
    .RESET_B(net1048),
    .D(\u_top_module.u_filter.shift_reg[229] ),
    .Q_N(_1195_),
    .Q(\u_top_module.u_filter.shift_reg[230] ));
 sg13g2_dfrbp_1 _2519_ (.CLK(net939),
    .RESET_B(net1047),
    .D(\u_top_module.u_filter.shift_reg[230] ),
    .Q_N(_1196_),
    .Q(\u_top_module.u_filter.shift_reg[231] ));
 sg13g2_dfrbp_1 _2520_ (.CLK(net939),
    .RESET_B(net1047),
    .D(\u_top_module.u_filter.shift_reg[231] ),
    .Q_N(_1197_),
    .Q(\u_top_module.u_filter.shift_reg[232] ));
 sg13g2_dfrbp_1 _2521_ (.CLK(net938),
    .RESET_B(net1047),
    .D(\u_top_module.u_filter.shift_reg[232] ),
    .Q_N(_1198_),
    .Q(\u_top_module.u_filter.shift_reg[233] ));
 sg13g2_dfrbp_1 _2522_ (.CLK(net939),
    .RESET_B(net1047),
    .D(\u_top_module.u_filter.shift_reg[233] ),
    .Q_N(_1199_),
    .Q(\u_top_module.u_filter.shift_reg[234] ));
 sg13g2_dfrbp_1 _2523_ (.CLK(net939),
    .RESET_B(net1044),
    .D(\u_top_module.u_filter.shift_reg[234] ),
    .Q_N(_1200_),
    .Q(\u_top_module.u_filter.shift_reg[235] ));
 sg13g2_dfrbp_1 _2524_ (.CLK(net939),
    .RESET_B(net1043),
    .D(\u_top_module.u_filter.shift_reg[235] ),
    .Q_N(_1201_),
    .Q(\u_top_module.u_filter.shift_reg[236] ));
 sg13g2_dfrbp_1 _2525_ (.CLK(net934),
    .RESET_B(net1043),
    .D(\u_top_module.u_filter.shift_reg[236] ),
    .Q_N(_1202_),
    .Q(\u_top_module.u_filter.shift_reg[237] ));
 sg13g2_dfrbp_1 _2526_ (.CLK(net934),
    .RESET_B(net1044),
    .D(\u_top_module.u_filter.shift_reg[237] ),
    .Q_N(_1203_),
    .Q(\u_top_module.u_filter.shift_reg[238] ));
 sg13g2_dfrbp_1 _2527_ (.CLK(net934),
    .RESET_B(net1044),
    .D(\u_top_module.u_filter.shift_reg[238] ),
    .Q_N(_1204_),
    .Q(\u_top_module.u_filter.shift_reg[239] ));
 sg13g2_dfrbp_1 _2528_ (.CLK(net934),
    .RESET_B(net1043),
    .D(\u_top_module.u_filter.shift_reg[239] ),
    .Q_N(_1205_),
    .Q(\u_top_module.u_filter.shift_reg[240] ));
 sg13g2_dfrbp_1 _2529_ (.CLK(net934),
    .RESET_B(net1043),
    .D(\u_top_module.u_filter.shift_reg[240] ),
    .Q_N(_1206_),
    .Q(\u_top_module.u_filter.shift_reg[241] ));
 sg13g2_dfrbp_1 _2530_ (.CLK(net934),
    .RESET_B(net1043),
    .D(\u_top_module.u_filter.shift_reg[241] ),
    .Q_N(_1207_),
    .Q(\u_top_module.u_filter.shift_reg[242] ));
 sg13g2_dfrbp_1 _2531_ (.CLK(net934),
    .RESET_B(net1037),
    .D(\u_top_module.u_filter.shift_reg[242] ),
    .Q_N(_1208_),
    .Q(\u_top_module.u_filter.shift_reg[243] ));
 sg13g2_dfrbp_1 _2532_ (.CLK(net928),
    .RESET_B(net1037),
    .D(\u_top_module.u_filter.shift_reg[243] ),
    .Q_N(_1209_),
    .Q(\u_top_module.u_filter.shift_reg[244] ));
 sg13g2_dfrbp_1 _2533_ (.CLK(net926),
    .RESET_B(net1037),
    .D(\u_top_module.u_filter.shift_reg[244] ),
    .Q_N(_1210_),
    .Q(\u_top_module.u_filter.shift_reg[245] ));
 sg13g2_dfrbp_1 _2534_ (.CLK(net928),
    .RESET_B(net1035),
    .D(\u_top_module.u_filter.shift_reg[245] ),
    .Q_N(_1211_),
    .Q(\u_top_module.u_filter.shift_reg[246] ));
 sg13g2_dfrbp_1 _2535_ (.CLK(net927),
    .RESET_B(net1035),
    .D(\u_top_module.u_filter.shift_reg[246] ),
    .Q_N(_1212_),
    .Q(\u_top_module.u_filter.shift_reg[247] ));
 sg13g2_dfrbp_1 _2536_ (.CLK(net926),
    .RESET_B(net1035),
    .D(\u_top_module.u_filter.shift_reg[247] ),
    .Q_N(_1213_),
    .Q(\u_top_module.u_filter.shift_reg[248] ));
 sg13g2_dfrbp_1 _2537_ (.CLK(net926),
    .RESET_B(net1035),
    .D(\u_top_module.u_filter.shift_reg[248] ),
    .Q_N(_1214_),
    .Q(\u_top_module.u_filter.shift_reg[249] ));
 sg13g2_dfrbp_1 _2538_ (.CLK(net926),
    .RESET_B(net1035),
    .D(\u_top_module.u_filter.shift_reg[249] ),
    .Q_N(_1215_),
    .Q(\u_top_module.u_filter.shift_reg[250] ));
 sg13g2_dfrbp_1 _2539_ (.CLK(net926),
    .RESET_B(net1035),
    .D(\u_top_module.u_filter.shift_reg[250] ),
    .Q_N(_1216_),
    .Q(\u_top_module.u_filter.shift_reg[251] ));
 sg13g2_dfrbp_1 _2540_ (.CLK(net926),
    .RESET_B(net1035),
    .D(\u_top_module.u_filter.shift_reg[251] ),
    .Q_N(_1217_),
    .Q(\u_top_module.u_filter.shift_reg[252] ));
 sg13g2_dfrbp_1 _2541_ (.CLK(net926),
    .RESET_B(net1036),
    .D(\u_top_module.u_filter.shift_reg[252] ),
    .Q_N(_1218_),
    .Q(\u_top_module.u_filter.shift_reg[253] ));
 sg13g2_dfrbp_1 _2542_ (.CLK(net926),
    .RESET_B(net1035),
    .D(\u_top_module.u_filter.shift_reg[253] ),
    .Q_N(_0774_),
    .Q(\u_top_module.u_filter.shift_reg[254] ));
 sg13g2_dfrbp_1 _2543_ (.CLK(net980),
    .RESET_B(net1039),
    .D(_0196_),
    .Q_N(_0010_),
    .Q(\u_top_module.dec_clk ));
 sg13g2_dfrbp_1 _2544_ (.CLK(net981),
    .RESET_B(net1026),
    .D(_0002_),
    .Q_N(_1219_),
    .Q(\u_top_module.u_decimator.counter[0] ));
 sg13g2_dfrbp_1 _2545_ (.CLK(net978),
    .RESET_B(net1026),
    .D(_0003_),
    .Q_N(_1220_),
    .Q(\u_top_module.u_decimator.counter[1] ));
 sg13g2_dfrbp_1 _2546_ (.CLK(net978),
    .RESET_B(net1026),
    .D(_0004_),
    .Q_N(_0773_),
    .Q(\u_top_module.u_decimator.counter[2] ));
 sg13g2_tiehi _2085__28 (.L_HI(net28));
 sg13g2_tiehi _2086__29 (.L_HI(net29));
 sg13g2_tiehi _2087__30 (.L_HI(net30));
 sg13g2_tiehi _2088__31 (.L_HI(net31));
 sg13g2_tiehi _2089__32 (.L_HI(net32));
 sg13g2_tiehi _2090__33 (.L_HI(net33));
 sg13g2_tiehi _2091__34 (.L_HI(net34));
 sg13g2_tiehi _2092__35 (.L_HI(net35));
 sg13g2_tiehi _2093__36 (.L_HI(net36));
 sg13g2_tiehi _2094__37 (.L_HI(net37));
 sg13g2_tiehi _2095__38 (.L_HI(net38));
 sg13g2_tiehi _2096__39 (.L_HI(net39));
 sg13g2_tiehi _2097__40 (.L_HI(net40));
 sg13g2_tiehi _2098__41 (.L_HI(net41));
 sg13g2_tiehi _2099__42 (.L_HI(net42));
 sg13g2_tiehi _2100__43 (.L_HI(net43));
 sg13g2_tiehi _2101__44 (.L_HI(net44));
 sg13g2_tiehi _2102__45 (.L_HI(net45));
 sg13g2_tiehi _2103__46 (.L_HI(net46));
 sg13g2_tiehi _2104__47 (.L_HI(net47));
 sg13g2_tiehi _2105__48 (.L_HI(net48));
 sg13g2_tiehi _2108__49 (.L_HI(net49));
 sg13g2_tiehi _2107__50 (.L_HI(net50));
 sg13g2_tiehi _2286__51 (.L_HI(net51));
 sg13g2_tiehi _2285__52 (.L_HI(net52));
 sg13g2_tiehi _2284__53 (.L_HI(net53));
 sg13g2_tiehi _2283__54 (.L_HI(net54));
 sg13g2_tiehi _2282__55 (.L_HI(net55));
 sg13g2_tiehi _2281__56 (.L_HI(net56));
 sg13g2_tiehi _2280__57 (.L_HI(net57));
 sg13g2_tiehi _2279__58 (.L_HI(net58));
 sg13g2_tiehi _2278__59 (.L_HI(net59));
 sg13g2_tiehi _2277__60 (.L_HI(net60));
 sg13g2_tiehi _2276__61 (.L_HI(net61));
 sg13g2_tiehi _2275__62 (.L_HI(net62));
 sg13g2_tiehi _2274__63 (.L_HI(net63));
 sg13g2_tiehi _2273__64 (.L_HI(net64));
 sg13g2_tiehi _2272__65 (.L_HI(net65));
 sg13g2_tiehi _2271__66 (.L_HI(net66));
 sg13g2_tiehi _2270__67 (.L_HI(net67));
 sg13g2_tiehi _2269__68 (.L_HI(net68));
 sg13g2_tiehi _2268__69 (.L_HI(net69));
 sg13g2_tiehi _2267__70 (.L_HI(net70));
 sg13g2_tiehi _2266__71 (.L_HI(net71));
 sg13g2_tiehi _2265__72 (.L_HI(net72));
 sg13g2_tiehi _2264__73 (.L_HI(net73));
 sg13g2_tiehi _2263__74 (.L_HI(net74));
 sg13g2_tiehi _2262__75 (.L_HI(net75));
 sg13g2_tiehi _2261__76 (.L_HI(net76));
 sg13g2_tiehi _2260__77 (.L_HI(net77));
 sg13g2_tiehi _2259__78 (.L_HI(net78));
 sg13g2_tiehi _2258__79 (.L_HI(net79));
 sg13g2_tiehi _2257__80 (.L_HI(net80));
 sg13g2_tiehi _2256__81 (.L_HI(net81));
 sg13g2_tiehi _2255__82 (.L_HI(net82));
 sg13g2_tiehi _2254__83 (.L_HI(net83));
 sg13g2_tiehi _2253__84 (.L_HI(net84));
 sg13g2_tiehi _2252__85 (.L_HI(net85));
 sg13g2_tiehi _2251__86 (.L_HI(net86));
 sg13g2_tiehi _2250__87 (.L_HI(net87));
 sg13g2_tiehi _2249__88 (.L_HI(net88));
 sg13g2_tiehi _2248__89 (.L_HI(net89));
 sg13g2_tiehi _2247__90 (.L_HI(net90));
 sg13g2_tiehi _2246__91 (.L_HI(net91));
 sg13g2_tiehi _2245__92 (.L_HI(net92));
 sg13g2_tiehi _2243__93 (.L_HI(net93));
 sg13g2_tiehi _2241__94 (.L_HI(net94));
 sg13g2_tiehi _2240__95 (.L_HI(net95));
 sg13g2_tiehi _2239__96 (.L_HI(net96));
 sg13g2_tiehi _2238__97 (.L_HI(net97));
 sg13g2_tiehi _2237__98 (.L_HI(net98));
 sg13g2_tiehi _2235__99 (.L_HI(net99));
 sg13g2_tiehi _2233__100 (.L_HI(net100));
 sg13g2_tiehi _2231__101 (.L_HI(net101));
 sg13g2_tiehi _2229__102 (.L_HI(net102));
 sg13g2_tiehi _2227__103 (.L_HI(net103));
 sg13g2_tiehi _2225__104 (.L_HI(net104));
 sg13g2_tiehi _2223__105 (.L_HI(net105));
 sg13g2_tiehi _2222__106 (.L_HI(net106));
 sg13g2_tiehi _2106__107 (.L_HI(net107));
 sg13g2_tiehi _2224__108 (.L_HI(net108));
 sg13g2_tiehi _2226__109 (.L_HI(net109));
 sg13g2_tiehi _2228__110 (.L_HI(net110));
 sg13g2_tiehi _2230__111 (.L_HI(net111));
 sg13g2_tiehi _2232__112 (.L_HI(net112));
 sg13g2_tiehi _2234__113 (.L_HI(net113));
 sg13g2_tiehi _2236__114 (.L_HI(net114));
 sg13g2_tiehi _2242__115 (.L_HI(net115));
 sg13g2_tiehi _2287__116 (.L_HI(net116));
 sg13g2_antennanp ANTENNA_1 (.A(rst_n));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_5 (.L_LO(net5));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_6 (.L_LO(net6));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_7 (.L_LO(net7));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_8 (.L_LO(net8));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_9 (.L_LO(net9));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_10 (.L_LO(net10));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_11 (.L_LO(net11));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_12 (.L_LO(net12));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_13 (.L_LO(net13));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_14 (.L_LO(net14));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_15 (.L_LO(net15));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_16 (.L_LO(net16));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_17 (.L_LO(net17));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_18 (.L_LO(net18));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_19 (.L_LO(net19));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_20 (.L_LO(net20));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_21 (.L_LO(net21));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_22 (.L_LO(net22));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_23 (.L_LO(net23));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_24 (.L_LO(net24));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_25 (.L_LO(net25));
 sg13g2_tielo _2221__26 (.L_LO(net26));
 sg13g2_tiehi _2084__27 (.L_HI(net27));
 sg13g2_buf_1 _2660_ (.A(\u_top_module.out ),
    .X(uo_out[0]));
 sg13g2_buf_1 _2661_ (.A(net980),
    .X(uo_out[1]));
 sg13g2_buf_2 fanout792 (.A(_0656_),
    .X(net792));
 sg13g2_buf_4 fanout793 (.X(net793),
    .A(net796));
 sg13g2_buf_4 fanout794 (.X(net794),
    .A(net795));
 sg13g2_buf_4 fanout795 (.X(net795),
    .A(net796));
 sg13g2_buf_2 fanout796 (.A(_0700_),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_0692_));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(_0689_));
 sg13g2_buf_2 fanout799 (.A(_0689_),
    .X(net799));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(net802));
 sg13g2_buf_1 fanout801 (.A(net802),
    .X(net801));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(_0688_));
 sg13g2_buf_4 fanout803 (.X(net803),
    .A(_0688_));
 sg13g2_buf_2 fanout804 (.A(_0688_),
    .X(net804));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(net806));
 sg13g2_buf_4 fanout806 (.X(net806),
    .A(_0680_));
 sg13g2_buf_2 fanout807 (.A(_0680_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_0680_),
    .X(net808));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(net811));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(net811));
 sg13g2_buf_4 fanout811 (.X(net811),
    .A(_0685_));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(net816));
 sg13g2_buf_2 fanout813 (.A(net816),
    .X(net813));
 sg13g2_buf_4 fanout814 (.X(net814),
    .A(net816));
 sg13g2_buf_1 fanout815 (.A(net816),
    .X(net815));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(_0683_));
 sg13g2_buf_4 fanout817 (.X(net817),
    .A(net818));
 sg13g2_buf_4 fanout818 (.X(net818),
    .A(_0682_));
 sg13g2_buf_4 fanout819 (.X(net819),
    .A(_0675_));
 sg13g2_buf_2 fanout820 (.A(_0675_),
    .X(net820));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(net822));
 sg13g2_buf_2 fanout822 (.A(_0675_),
    .X(net822));
 sg13g2_buf_4 fanout823 (.X(net823),
    .A(net825));
 sg13g2_buf_2 fanout824 (.A(net825),
    .X(net824));
 sg13g2_buf_4 fanout825 (.X(net825),
    .A(_0673_));
 sg13g2_buf_4 fanout826 (.X(net826),
    .A(net828));
 sg13g2_buf_4 fanout827 (.X(net827),
    .A(_0673_));
 sg13g2_buf_1 fanout828 (.A(_0673_),
    .X(net828));
 sg13g2_buf_8 fanout829 (.A(_0672_),
    .X(net829));
 sg13g2_buf_4 fanout830 (.X(net830),
    .A(_0561_));
 sg13g2_buf_2 fanout831 (.A(_0561_),
    .X(net831));
 sg13g2_buf_4 fanout832 (.X(net832),
    .A(_0560_));
 sg13g2_buf_2 fanout833 (.A(_0560_),
    .X(net833));
 sg13g2_buf_4 fanout834 (.X(net834),
    .A(net838));
 sg13g2_buf_2 fanout835 (.A(net838),
    .X(net835));
 sg13g2_buf_4 fanout836 (.X(net836),
    .A(net838));
 sg13g2_buf_4 fanout837 (.X(net837),
    .A(net838));
 sg13g2_buf_2 fanout838 (.A(\u_top_module.filter_length[2] ),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(net842),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(net842),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(\u_top_module.filter_length[1] ),
    .X(net842));
 sg13g2_buf_4 fanout843 (.X(net843),
    .A(net846));
 sg13g2_buf_2 fanout844 (.A(net846),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(net846),
    .X(net845));
 sg13g2_buf_1 fanout846 (.A(\u_top_module.filter_length[1] ),
    .X(net846));
 sg13g2_buf_4 fanout847 (.X(net847),
    .A(net850));
 sg13g2_buf_2 fanout848 (.A(net850),
    .X(net848));
 sg13g2_buf_1 fanout849 (.A(net850),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(net855),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(net855),
    .X(net851));
 sg13g2_buf_1 fanout852 (.A(net855),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(net854),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(net855),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(\u_top_module.filter_length[1] ),
    .X(net855));
 sg13g2_buf_4 fanout856 (.X(net856),
    .A(net858));
 sg13g2_buf_4 fanout857 (.X(net857),
    .A(net858));
 sg13g2_buf_4 fanout858 (.X(net858),
    .A(net870));
 sg13g2_buf_4 fanout859 (.X(net859),
    .A(net862));
 sg13g2_buf_4 fanout860 (.X(net860),
    .A(net862));
 sg13g2_buf_2 fanout861 (.A(net862),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(net870),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(net865),
    .X(net863));
 sg13g2_buf_4 fanout864 (.X(net864),
    .A(net870));
 sg13g2_buf_1 fanout865 (.A(net870),
    .X(net865));
 sg13g2_buf_4 fanout866 (.X(net866),
    .A(net869));
 sg13g2_buf_2 fanout867 (.A(net869),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(net869),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(net870),
    .X(net869));
 sg13g2_buf_4 fanout870 (.X(net870),
    .A(\u_top_module.filter_length[0] ));
 sg13g2_buf_4 fanout871 (.X(net871),
    .A(_0571_));
 sg13g2_buf_4 fanout872 (.X(net872),
    .A(_0571_));
 sg13g2_buf_4 fanout873 (.X(net873),
    .A(_0570_));
 sg13g2_buf_4 fanout874 (.X(net874),
    .A(_0570_));
 sg13g2_buf_4 fanout875 (.X(net875),
    .A(_0581_));
 sg13g2_buf_4 fanout876 (.X(net876),
    .A(_0581_));
 sg13g2_buf_4 fanout877 (.X(net877),
    .A(_0576_));
 sg13g2_buf_4 fanout878 (.X(net878),
    .A(_0576_));
 sg13g2_buf_4 fanout879 (.X(net879),
    .A(_0574_));
 sg13g2_buf_4 fanout880 (.X(net880),
    .A(_0574_));
 sg13g2_buf_4 fanout881 (.X(net881),
    .A(_0573_));
 sg13g2_buf_4 fanout882 (.X(net882),
    .A(_0573_));
 sg13g2_buf_4 fanout883 (.X(net883),
    .A(_0671_));
 sg13g2_buf_4 fanout884 (.X(net884),
    .A(_0671_));
 sg13g2_buf_4 fanout885 (.X(net885),
    .A(net886));
 sg13g2_buf_4 fanout886 (.X(net886),
    .A(_0669_));
 sg13g2_buf_2 fanout887 (.A(net890),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(net890),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(net890),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(net892),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(net892),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(_0640_),
    .X(net892));
 sg13g2_buf_4 fanout893 (.X(net893),
    .A(_0580_));
 sg13g2_buf_4 fanout894 (.X(net894),
    .A(_0580_));
 sg13g2_buf_4 fanout895 (.X(net895),
    .A(net896));
 sg13g2_buf_4 fanout896 (.X(net896),
    .A(_0577_));
 sg13g2_buf_2 fanout897 (.A(net898),
    .X(net897));
 sg13g2_buf_1 fanout898 (.A(net899),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(net909),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(net909),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(net909),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(net905),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(net904),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(net905),
    .X(net904));
 sg13g2_buf_1 fanout905 (.A(net908),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(net907),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(net908),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(net909),
    .X(net908));
 sg13g2_buf_1 fanout909 (.A(net942),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(net911),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(net914),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(net914),
    .X(net912));
 sg13g2_buf_1 fanout913 (.A(net914),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(net942),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(net919),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(net919),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(net918),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(net919),
    .X(net918));
 sg13g2_buf_1 fanout919 (.A(net942),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(net922),
    .X(net920));
 sg13g2_buf_1 fanout921 (.A(net922),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(net929),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(net925),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(net925),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(net928),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(net927),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(net928),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(net929),
    .X(net928));
 sg13g2_buf_1 fanout929 (.A(net942),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(net932),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(net941),
    .X(net931));
 sg13g2_buf_1 fanout932 (.A(net941),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(net941),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(net935),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(net940),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(net940),
    .X(net936));
 sg13g2_buf_1 fanout937 (.A(net940),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(net939),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(net940),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(net941),
    .X(net940));
 sg13g2_buf_1 fanout941 (.A(net942),
    .X(net941));
 sg13g2_buf_4 fanout942 (.X(net942),
    .A(\u_top_module.dec_clk ));
 sg13g2_buf_4 fanout943 (.X(net943),
    .A(\u_top_module.capture_reg[7] ));
 sg13g2_buf_2 fanout944 (.A(\u_top_module.capture_reg[6] ),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(\u_top_module.capture_reg[5] ),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(\u_top_module.capture_reg[4] ),
    .X(net946));
 sg13g2_buf_4 fanout947 (.X(net947),
    .A(\u_top_module.capture_reg[3] ));
 sg13g2_buf_2 fanout948 (.A(\u_top_module.capture_reg[2] ),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(\u_top_module.capture_reg[1] ),
    .X(net949));
 sg13g2_buf_4 fanout950 (.X(net950),
    .A(\u_top_module.capture_reg[0] ));
 sg13g2_buf_2 fanout951 (.A(net952),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(net955),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(net955),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(net955),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(net983),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(net957),
    .X(net956));
 sg13g2_buf_1 fanout957 (.A(net958),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(net983),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(net961),
    .X(net959));
 sg13g2_buf_1 fanout960 (.A(net961),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(net962),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(net966),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(net966),
    .X(net963));
 sg13g2_buf_1 fanout964 (.A(net966),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(net966),
    .X(net965));
 sg13g2_buf_1 fanout966 (.A(net983),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(net970),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(net970),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(net970),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(net982),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(net982),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(net982),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(net977),
    .X(net973));
 sg13g2_buf_1 fanout974 (.A(net977),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(net977),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(net977),
    .X(net976));
 sg13g2_buf_1 fanout977 (.A(net982),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(net981),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(net980),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(net981),
    .X(net980));
 sg13g2_buf_1 fanout981 (.A(net982),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(net983),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(ui_in[0]),
    .X(net983));
 sg13g2_buf_4 fanout984 (.X(net984),
    .A(net985));
 sg13g2_buf_4 fanout985 (.X(net985),
    .A(net1051));
 sg13g2_buf_4 fanout986 (.X(net986),
    .A(net991));
 sg13g2_buf_4 fanout987 (.X(net987),
    .A(net988));
 sg13g2_buf_2 fanout988 (.A(net991),
    .X(net988));
 sg13g2_buf_4 fanout989 (.X(net989),
    .A(net991));
 sg13g2_buf_4 fanout990 (.X(net990),
    .A(net991));
 sg13g2_buf_2 fanout991 (.A(net999),
    .X(net991));
 sg13g2_buf_4 fanout992 (.X(net992),
    .A(net996));
 sg13g2_buf_2 fanout993 (.A(net996),
    .X(net993));
 sg13g2_buf_4 fanout994 (.X(net994),
    .A(net996));
 sg13g2_buf_2 fanout995 (.A(net996),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(net999),
    .X(net996));
 sg13g2_buf_4 fanout997 (.X(net997),
    .A(net999));
 sg13g2_buf_4 fanout998 (.X(net998),
    .A(net999));
 sg13g2_buf_2 fanout999 (.A(net1010),
    .X(net999));
 sg13g2_buf_4 fanout1000 (.X(net1000),
    .A(net1004));
 sg13g2_buf_4 fanout1001 (.X(net1001),
    .A(net1004));
 sg13g2_buf_4 fanout1002 (.X(net1002),
    .A(net1004));
 sg13g2_buf_4 fanout1003 (.X(net1003),
    .A(net1004));
 sg13g2_buf_2 fanout1004 (.A(net1010),
    .X(net1004));
 sg13g2_buf_4 fanout1005 (.X(net1005),
    .A(net1007));
 sg13g2_buf_4 fanout1006 (.X(net1006),
    .A(net1007));
 sg13g2_buf_2 fanout1007 (.A(net1010),
    .X(net1007));
 sg13g2_buf_4 fanout1008 (.X(net1008),
    .A(net1009));
 sg13g2_buf_4 fanout1009 (.X(net1009),
    .A(net1010));
 sg13g2_buf_2 fanout1010 (.A(net1051),
    .X(net1010));
 sg13g2_buf_4 fanout1011 (.X(net1011),
    .A(net1014));
 sg13g2_buf_2 fanout1012 (.A(net1014),
    .X(net1012));
 sg13g2_buf_4 fanout1013 (.X(net1013),
    .A(net1014));
 sg13g2_buf_2 fanout1014 (.A(net1016),
    .X(net1014));
 sg13g2_buf_4 fanout1015 (.X(net1015),
    .A(net1016));
 sg13g2_buf_2 fanout1016 (.A(net1028),
    .X(net1016));
 sg13g2_buf_4 fanout1017 (.X(net1017),
    .A(net1028));
 sg13g2_buf_2 fanout1018 (.A(net1028),
    .X(net1018));
 sg13g2_buf_4 fanout1019 (.X(net1019),
    .A(net1023));
 sg13g2_buf_4 fanout1020 (.X(net1020),
    .A(net1023));
 sg13g2_buf_4 fanout1021 (.X(net1021),
    .A(net1022));
 sg13g2_buf_4 fanout1022 (.X(net1022),
    .A(net1023));
 sg13g2_buf_4 fanout1023 (.X(net1023),
    .A(net1027));
 sg13g2_buf_4 fanout1024 (.X(net1024),
    .A(net1027));
 sg13g2_buf_2 fanout1025 (.A(net1027),
    .X(net1025));
 sg13g2_buf_4 fanout1026 (.X(net1026),
    .A(net1027));
 sg13g2_buf_2 fanout1027 (.A(net1028),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(net1050),
    .X(net1028));
 sg13g2_buf_4 fanout1029 (.X(net1029),
    .A(net1032));
 sg13g2_buf_4 fanout1030 (.X(net1030),
    .A(net1032));
 sg13g2_buf_2 fanout1031 (.A(net1032),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(net1050),
    .X(net1032));
 sg13g2_buf_4 fanout1033 (.X(net1033),
    .A(net1034));
 sg13g2_buf_4 fanout1034 (.X(net1034),
    .A(net1037));
 sg13g2_buf_4 fanout1035 (.X(net1035),
    .A(net1036));
 sg13g2_buf_4 fanout1036 (.X(net1036),
    .A(net1037));
 sg13g2_buf_4 fanout1037 (.X(net1037),
    .A(net1050));
 sg13g2_buf_4 fanout1038 (.X(net1038),
    .A(net1042));
 sg13g2_buf_4 fanout1039 (.X(net1039),
    .A(net1041));
 sg13g2_buf_4 fanout1040 (.X(net1040),
    .A(net1041));
 sg13g2_buf_2 fanout1041 (.A(net1042),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(net1049),
    .X(net1042));
 sg13g2_buf_4 fanout1043 (.X(net1043),
    .A(net1049));
 sg13g2_buf_2 fanout1044 (.A(net1045),
    .X(net1044));
 sg13g2_buf_4 fanout1045 (.X(net1045),
    .A(net1049));
 sg13g2_buf_4 fanout1046 (.X(net1046),
    .A(net1048));
 sg13g2_buf_4 fanout1047 (.X(net1047),
    .A(net1048));
 sg13g2_buf_2 fanout1048 (.A(net1049),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(net1050),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(net1051),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(rst_n),
    .X(net1051));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_tielo tt_um_pdm_pitch_filter_arghunter_4 (.L_LO(net4));
 sg13g2_antennanp ANTENNA_2 (.A(rst_n));
 sg13g2_antennanp ANTENNA_3 (.A(ui_in[0]));
 sg13g2_antennanp ANTENNA_4 (.A(ui_in[0]));
 sg13g2_antennanp ANTENNA_5 (.A(ui_in[0]));
 sg13g2_antennanp ANTENNA_6 (.A(ui_in[0]));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_fill_1 FILLER_2_266 ();
 sg13g2_fill_2 FILLER_2_293 ();
 sg13g2_decap_8 FILLER_2_321 ();
 sg13g2_fill_2 FILLER_2_328 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_4 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_261 ();
 sg13g2_decap_8 FILLER_4_268 ();
 sg13g2_decap_8 FILLER_4_275 ();
 sg13g2_decap_4 FILLER_4_282 ();
 sg13g2_decap_8 FILLER_4_312 ();
 sg13g2_fill_1 FILLER_4_319 ();
 sg13g2_fill_2 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_4 FILLER_5_245 ();
 sg13g2_fill_2 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_277 ();
 sg13g2_decap_4 FILLER_5_284 ();
 sg13g2_fill_1 FILLER_5_288 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_4 FILLER_5_340 ();
 sg13g2_fill_1 FILLER_5_344 ();
 sg13g2_fill_1 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_fill_2 FILLER_6_224 ();
 sg13g2_fill_1 FILLER_6_226 ();
 sg13g2_fill_1 FILLER_6_264 ();
 sg13g2_fill_2 FILLER_6_271 ();
 sg13g2_fill_1 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_285 ();
 sg13g2_decap_8 FILLER_6_292 ();
 sg13g2_fill_2 FILLER_6_324 ();
 sg13g2_decap_8 FILLER_6_358 ();
 sg13g2_decap_8 FILLER_6_365 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_4 FILLER_7_224 ();
 sg13g2_fill_2 FILLER_7_228 ();
 sg13g2_fill_1 FILLER_7_261 ();
 sg13g2_fill_2 FILLER_7_319 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_4 FILLER_8_210 ();
 sg13g2_fill_1 FILLER_8_214 ();
 sg13g2_decap_8 FILLER_8_246 ();
 sg13g2_decap_8 FILLER_8_253 ();
 sg13g2_fill_2 FILLER_8_260 ();
 sg13g2_fill_1 FILLER_8_262 ();
 sg13g2_decap_8 FILLER_8_272 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_fill_2 FILLER_8_317 ();
 sg13g2_fill_1 FILLER_8_319 ();
 sg13g2_fill_1 FILLER_8_345 ();
 sg13g2_decap_8 FILLER_8_376 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_decap_4 FILLER_9_188 ();
 sg13g2_fill_2 FILLER_9_192 ();
 sg13g2_decap_8 FILLER_9_197 ();
 sg13g2_decap_8 FILLER_9_204 ();
 sg13g2_decap_4 FILLER_9_211 ();
 sg13g2_fill_2 FILLER_9_241 ();
 sg13g2_fill_2 FILLER_9_247 ();
 sg13g2_fill_1 FILLER_9_249 ();
 sg13g2_fill_2 FILLER_9_262 ();
 sg13g2_decap_4 FILLER_9_269 ();
 sg13g2_fill_2 FILLER_9_278 ();
 sg13g2_decap_8 FILLER_9_288 ();
 sg13g2_decap_8 FILLER_9_295 ();
 sg13g2_decap_4 FILLER_9_302 ();
 sg13g2_fill_2 FILLER_9_311 ();
 sg13g2_fill_1 FILLER_9_313 ();
 sg13g2_decap_8 FILLER_9_318 ();
 sg13g2_decap_8 FILLER_9_325 ();
 sg13g2_fill_1 FILLER_9_332 ();
 sg13g2_decap_4 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_fill_2 FILLER_10_131 ();
 sg13g2_fill_1 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_138 ();
 sg13g2_decap_8 FILLER_10_145 ();
 sg13g2_decap_8 FILLER_10_152 ();
 sg13g2_decap_8 FILLER_10_159 ();
 sg13g2_decap_8 FILLER_10_166 ();
 sg13g2_decap_8 FILLER_10_206 ();
 sg13g2_decap_8 FILLER_10_213 ();
 sg13g2_decap_8 FILLER_10_220 ();
 sg13g2_fill_2 FILLER_10_227 ();
 sg13g2_fill_1 FILLER_10_233 ();
 sg13g2_fill_1 FILLER_10_264 ();
 sg13g2_decap_4 FILLER_10_299 ();
 sg13g2_fill_2 FILLER_10_342 ();
 sg13g2_fill_1 FILLER_10_344 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_4 FILLER_11_84 ();
 sg13g2_fill_2 FILLER_11_120 ();
 sg13g2_fill_1 FILLER_11_122 ();
 sg13g2_decap_8 FILLER_11_149 ();
 sg13g2_fill_2 FILLER_11_156 ();
 sg13g2_fill_2 FILLER_11_240 ();
 sg13g2_fill_1 FILLER_11_242 ();
 sg13g2_fill_1 FILLER_11_326 ();
 sg13g2_decap_4 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_4 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_135 ();
 sg13g2_fill_2 FILLER_12_188 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_fill_1 FILLER_12_322 ();
 sg13g2_decap_4 FILLER_12_328 ();
 sg13g2_fill_2 FILLER_12_337 ();
 sg13g2_fill_1 FILLER_12_339 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_4 FILLER_13_64 ();
 sg13g2_fill_2 FILLER_13_68 ();
 sg13g2_fill_1 FILLER_13_96 ();
 sg13g2_decap_4 FILLER_13_162 ();
 sg13g2_fill_1 FILLER_13_187 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_decap_4 FILLER_13_200 ();
 sg13g2_decap_8 FILLER_13_212 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_4 FILLER_13_252 ();
 sg13g2_decap_4 FILLER_13_268 ();
 sg13g2_fill_2 FILLER_13_272 ();
 sg13g2_decap_8 FILLER_13_279 ();
 sg13g2_decap_8 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_298 ();
 sg13g2_decap_8 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_312 ();
 sg13g2_fill_2 FILLER_13_319 ();
 sg13g2_fill_1 FILLER_13_321 ();
 sg13g2_fill_1 FILLER_13_327 ();
 sg13g2_fill_2 FILLER_13_333 ();
 sg13g2_fill_1 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_4 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_32 ();
 sg13g2_fill_2 FILLER_14_59 ();
 sg13g2_fill_2 FILLER_14_99 ();
 sg13g2_fill_1 FILLER_14_101 ();
 sg13g2_decap_4 FILLER_14_113 ();
 sg13g2_decap_4 FILLER_14_130 ();
 sg13g2_fill_2 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_139 ();
 sg13g2_fill_1 FILLER_14_146 ();
 sg13g2_decap_8 FILLER_14_155 ();
 sg13g2_decap_8 FILLER_14_162 ();
 sg13g2_decap_8 FILLER_14_169 ();
 sg13g2_decap_4 FILLER_14_176 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_decap_4 FILLER_14_213 ();
 sg13g2_fill_2 FILLER_14_243 ();
 sg13g2_fill_1 FILLER_14_245 ();
 sg13g2_decap_4 FILLER_14_277 ();
 sg13g2_decap_4 FILLER_14_286 ();
 sg13g2_fill_2 FILLER_14_290 ();
 sg13g2_decap_4 FILLER_14_301 ();
 sg13g2_fill_2 FILLER_14_305 ();
 sg13g2_fill_1 FILLER_14_333 ();
 sg13g2_decap_4 FILLER_14_352 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_fill_2 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_44 ();
 sg13g2_fill_1 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_102 ();
 sg13g2_decap_8 FILLER_15_109 ();
 sg13g2_decap_4 FILLER_15_116 ();
 sg13g2_fill_1 FILLER_15_120 ();
 sg13g2_decap_4 FILLER_15_147 ();
 sg13g2_fill_1 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_155 ();
 sg13g2_fill_2 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_172 ();
 sg13g2_decap_8 FILLER_15_179 ();
 sg13g2_decap_4 FILLER_15_186 ();
 sg13g2_fill_1 FILLER_15_190 ();
 sg13g2_fill_2 FILLER_15_195 ();
 sg13g2_fill_1 FILLER_15_197 ();
 sg13g2_decap_8 FILLER_15_212 ();
 sg13g2_decap_8 FILLER_15_219 ();
 sg13g2_fill_2 FILLER_15_226 ();
 sg13g2_fill_1 FILLER_15_228 ();
 sg13g2_fill_1 FILLER_15_255 ();
 sg13g2_decap_8 FILLER_15_328 ();
 sg13g2_fill_2 FILLER_15_335 ();
 sg13g2_decap_4 FILLER_15_340 ();
 sg13g2_fill_1 FILLER_15_344 ();
 sg13g2_fill_1 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_fill_1 FILLER_16_85 ();
 sg13g2_fill_2 FILLER_16_117 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_fill_1 FILLER_16_129 ();
 sg13g2_fill_2 FILLER_16_187 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_decap_4 FILLER_16_222 ();
 sg13g2_fill_1 FILLER_16_226 ();
 sg13g2_decap_4 FILLER_16_243 ();
 sg13g2_fill_2 FILLER_16_286 ();
 sg13g2_decap_4 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_4 FILLER_17_42 ();
 sg13g2_fill_2 FILLER_17_46 ();
 sg13g2_decap_4 FILLER_17_51 ();
 sg13g2_fill_2 FILLER_17_55 ();
 sg13g2_decap_4 FILLER_17_61 ();
 sg13g2_fill_2 FILLER_17_70 ();
 sg13g2_decap_4 FILLER_17_75 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_fill_2 FILLER_17_91 ();
 sg13g2_fill_1 FILLER_17_93 ();
 sg13g2_fill_2 FILLER_17_99 ();
 sg13g2_fill_1 FILLER_17_101 ();
 sg13g2_decap_8 FILLER_17_106 ();
 sg13g2_fill_1 FILLER_17_113 ();
 sg13g2_fill_2 FILLER_17_192 ();
 sg13g2_fill_1 FILLER_17_259 ();
 sg13g2_decap_4 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_30 ();
 sg13g2_decap_4 FILLER_18_57 ();
 sg13g2_fill_1 FILLER_18_61 ();
 sg13g2_fill_1 FILLER_18_67 ();
 sg13g2_fill_2 FILLER_18_97 ();
 sg13g2_fill_1 FILLER_18_99 ();
 sg13g2_decap_8 FILLER_18_104 ();
 sg13g2_fill_2 FILLER_18_116 ();
 sg13g2_fill_2 FILLER_18_123 ();
 sg13g2_fill_1 FILLER_18_125 ();
 sg13g2_fill_2 FILLER_18_138 ();
 sg13g2_fill_1 FILLER_18_140 ();
 sg13g2_fill_2 FILLER_18_184 ();
 sg13g2_fill_1 FILLER_18_191 ();
 sg13g2_decap_8 FILLER_18_218 ();
 sg13g2_fill_1 FILLER_18_225 ();
 sg13g2_decap_8 FILLER_18_257 ();
 sg13g2_decap_8 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_271 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_fill_2 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_4 FILLER_18_324 ();
 sg13g2_fill_2 FILLER_18_328 ();
 sg13g2_fill_2 FILLER_18_335 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_4 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_32 ();
 sg13g2_fill_2 FILLER_19_115 ();
 sg13g2_fill_2 FILLER_19_121 ();
 sg13g2_fill_1 FILLER_19_123 ();
 sg13g2_decap_4 FILLER_19_127 ();
 sg13g2_fill_1 FILLER_19_135 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_fill_1 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_159 ();
 sg13g2_fill_2 FILLER_19_165 ();
 sg13g2_decap_8 FILLER_19_171 ();
 sg13g2_decap_8 FILLER_19_178 ();
 sg13g2_decap_8 FILLER_19_185 ();
 sg13g2_fill_2 FILLER_19_192 ();
 sg13g2_fill_1 FILLER_19_194 ();
 sg13g2_decap_4 FILLER_19_198 ();
 sg13g2_fill_1 FILLER_19_202 ();
 sg13g2_decap_8 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_218 ();
 sg13g2_fill_1 FILLER_19_245 ();
 sg13g2_fill_2 FILLER_19_250 ();
 sg13g2_fill_1 FILLER_19_252 ();
 sg13g2_fill_1 FILLER_19_257 ();
 sg13g2_decap_8 FILLER_19_267 ();
 sg13g2_decap_8 FILLER_19_274 ();
 sg13g2_fill_1 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_4 FILLER_19_294 ();
 sg13g2_fill_2 FILLER_19_306 ();
 sg13g2_decap_4 FILLER_19_318 ();
 sg13g2_fill_1 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_fill_1 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_377 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_fill_2 FILLER_20_76 ();
 sg13g2_decap_4 FILLER_20_104 ();
 sg13g2_fill_1 FILLER_20_108 ();
 sg13g2_fill_1 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_146 ();
 sg13g2_decap_8 FILLER_20_153 ();
 sg13g2_decap_8 FILLER_20_160 ();
 sg13g2_decap_4 FILLER_20_167 ();
 sg13g2_fill_1 FILLER_20_171 ();
 sg13g2_fill_2 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_209 ();
 sg13g2_decap_8 FILLER_20_216 ();
 sg13g2_decap_8 FILLER_20_223 ();
 sg13g2_decap_8 FILLER_20_230 ();
 sg13g2_decap_8 FILLER_20_237 ();
 sg13g2_decap_4 FILLER_20_244 ();
 sg13g2_fill_2 FILLER_20_248 ();
 sg13g2_fill_1 FILLER_20_281 ();
 sg13g2_fill_2 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_341 ();
 sg13g2_fill_2 FILLER_20_348 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_4 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_65 ();
 sg13g2_decap_8 FILLER_21_72 ();
 sg13g2_decap_4 FILLER_21_87 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_2 FILLER_21_173 ();
 sg13g2_decap_4 FILLER_21_179 ();
 sg13g2_fill_1 FILLER_21_183 ();
 sg13g2_decap_8 FILLER_21_240 ();
 sg13g2_decap_8 FILLER_21_247 ();
 sg13g2_decap_4 FILLER_21_254 ();
 sg13g2_fill_1 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_4 FILLER_22_84 ();
 sg13g2_fill_1 FILLER_22_88 ();
 sg13g2_fill_2 FILLER_22_93 ();
 sg13g2_fill_1 FILLER_22_95 ();
 sg13g2_fill_1 FILLER_22_101 ();
 sg13g2_fill_1 FILLER_22_137 ();
 sg13g2_decap_8 FILLER_22_205 ();
 sg13g2_decap_4 FILLER_22_212 ();
 sg13g2_fill_1 FILLER_22_216 ();
 sg13g2_decap_8 FILLER_22_243 ();
 sg13g2_decap_8 FILLER_22_250 ();
 sg13g2_fill_2 FILLER_22_257 ();
 sg13g2_decap_4 FILLER_22_285 ();
 sg13g2_fill_2 FILLER_22_297 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_4 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_95 ();
 sg13g2_decap_8 FILLER_23_107 ();
 sg13g2_decap_4 FILLER_23_114 ();
 sg13g2_decap_8 FILLER_23_122 ();
 sg13g2_decap_4 FILLER_23_129 ();
 sg13g2_fill_1 FILLER_23_133 ();
 sg13g2_decap_4 FILLER_23_147 ();
 sg13g2_fill_2 FILLER_23_155 ();
 sg13g2_decap_4 FILLER_23_161 ();
 sg13g2_fill_1 FILLER_23_165 ();
 sg13g2_decap_8 FILLER_23_174 ();
 sg13g2_fill_2 FILLER_23_181 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_decap_4 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_264 ();
 sg13g2_decap_4 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_275 ();
 sg13g2_fill_1 FILLER_23_286 ();
 sg13g2_decap_8 FILLER_23_296 ();
 sg13g2_decap_4 FILLER_23_303 ();
 sg13g2_fill_2 FILLER_23_307 ();
 sg13g2_decap_8 FILLER_23_314 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_335 ();
 sg13g2_decap_8 FILLER_23_376 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_4 FILLER_24_77 ();
 sg13g2_fill_1 FILLER_24_81 ();
 sg13g2_fill_1 FILLER_24_108 ();
 sg13g2_fill_2 FILLER_24_135 ();
 sg13g2_fill_1 FILLER_24_163 ();
 sg13g2_fill_2 FILLER_24_169 ();
 sg13g2_fill_2 FILLER_24_200 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_decap_4 FILLER_24_211 ();
 sg13g2_fill_2 FILLER_24_215 ();
 sg13g2_decap_4 FILLER_24_269 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_299 ();
 sg13g2_decap_8 FILLER_24_323 ();
 sg13g2_decap_8 FILLER_24_330 ();
 sg13g2_decap_8 FILLER_24_337 ();
 sg13g2_fill_2 FILLER_24_344 ();
 sg13g2_decap_8 FILLER_24_356 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_4 FILLER_25_77 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_decap_4 FILLER_25_139 ();
 sg13g2_fill_2 FILLER_25_143 ();
 sg13g2_decap_8 FILLER_25_178 ();
 sg13g2_fill_1 FILLER_25_189 ();
 sg13g2_fill_1 FILLER_25_194 ();
 sg13g2_decap_8 FILLER_25_214 ();
 sg13g2_decap_8 FILLER_25_221 ();
 sg13g2_decap_8 FILLER_25_228 ();
 sg13g2_decap_8 FILLER_25_235 ();
 sg13g2_decap_4 FILLER_25_242 ();
 sg13g2_decap_4 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_319 ();
 sg13g2_decap_4 FILLER_25_326 ();
 sg13g2_fill_1 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_4 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_4 FILLER_25_370 ();
 sg13g2_fill_2 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_4 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_81 ();
 sg13g2_fill_1 FILLER_26_117 ();
 sg13g2_decap_8 FILLER_26_128 ();
 sg13g2_decap_4 FILLER_26_135 ();
 sg13g2_fill_1 FILLER_26_169 ();
 sg13g2_fill_1 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_180 ();
 sg13g2_decap_4 FILLER_26_187 ();
 sg13g2_decap_8 FILLER_26_225 ();
 sg13g2_decap_8 FILLER_26_232 ();
 sg13g2_decap_4 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_243 ();
 sg13g2_fill_1 FILLER_26_254 ();
 sg13g2_decap_8 FILLER_26_260 ();
 sg13g2_fill_1 FILLER_26_304 ();
 sg13g2_fill_2 FILLER_26_331 ();
 sg13g2_fill_1 FILLER_26_338 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_108 ();
 sg13g2_decap_8 FILLER_27_115 ();
 sg13g2_decap_8 FILLER_27_122 ();
 sg13g2_decap_8 FILLER_27_129 ();
 sg13g2_decap_8 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_143 ();
 sg13g2_decap_8 FILLER_27_153 ();
 sg13g2_decap_4 FILLER_27_160 ();
 sg13g2_fill_1 FILLER_27_164 ();
 sg13g2_fill_2 FILLER_27_191 ();
 sg13g2_fill_1 FILLER_27_193 ();
 sg13g2_fill_2 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_204 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_decap_4 FILLER_28_216 ();
 sg13g2_fill_1 FILLER_28_220 ();
 sg13g2_fill_1 FILLER_28_251 ();
 sg13g2_fill_2 FILLER_28_278 ();
 sg13g2_fill_1 FILLER_28_280 ();
 sg13g2_fill_2 FILLER_28_299 ();
 sg13g2_decap_8 FILLER_28_306 ();
 sg13g2_fill_2 FILLER_28_355 ();
 sg13g2_fill_1 FILLER_28_357 ();
 sg13g2_fill_2 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_4 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_95 ();
 sg13g2_decap_4 FILLER_29_157 ();
 sg13g2_fill_2 FILLER_29_169 ();
 sg13g2_fill_1 FILLER_29_171 ();
 sg13g2_decap_8 FILLER_29_181 ();
 sg13g2_decap_4 FILLER_29_188 ();
 sg13g2_fill_1 FILLER_29_192 ();
 sg13g2_fill_2 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_230 ();
 sg13g2_decap_8 FILLER_29_237 ();
 sg13g2_decap_8 FILLER_29_244 ();
 sg13g2_decap_8 FILLER_29_251 ();
 sg13g2_decap_8 FILLER_29_258 ();
 sg13g2_decap_8 FILLER_29_265 ();
 sg13g2_decap_8 FILLER_29_272 ();
 sg13g2_decap_8 FILLER_29_279 ();
 sg13g2_decap_4 FILLER_29_286 ();
 sg13g2_fill_1 FILLER_29_290 ();
 sg13g2_fill_2 FILLER_29_301 ();
 sg13g2_decap_4 FILLER_29_363 ();
 sg13g2_fill_2 FILLER_29_379 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_4 FILLER_30_84 ();
 sg13g2_fill_1 FILLER_30_88 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_2 FILLER_30_134 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_decap_8 FILLER_30_163 ();
 sg13g2_decap_4 FILLER_30_170 ();
 sg13g2_fill_2 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_fill_2 FILLER_30_215 ();
 sg13g2_decap_8 FILLER_30_243 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_fill_1 FILLER_30_252 ();
 sg13g2_fill_1 FILLER_30_279 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_fill_1 FILLER_30_328 ();
 sg13g2_decap_8 FILLER_30_338 ();
 sg13g2_decap_8 FILLER_30_345 ();
 sg13g2_decap_8 FILLER_30_352 ();
 sg13g2_decap_8 FILLER_30_359 ();
 sg13g2_fill_2 FILLER_30_366 ();
 sg13g2_fill_1 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_decap_8 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_4 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_fill_1 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_131 ();
 sg13g2_decap_4 FILLER_31_138 ();
 sg13g2_decap_4 FILLER_31_146 ();
 sg13g2_fill_1 FILLER_31_242 ();
 sg13g2_fill_2 FILLER_31_248 ();
 sg13g2_fill_2 FILLER_31_258 ();
 sg13g2_fill_2 FILLER_31_293 ();
 sg13g2_fill_2 FILLER_31_308 ();
 sg13g2_fill_1 FILLER_31_310 ();
 sg13g2_decap_8 FILLER_31_316 ();
 sg13g2_fill_2 FILLER_31_323 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_4 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_107 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_147 ();
 sg13g2_decap_4 FILLER_32_155 ();
 sg13g2_fill_2 FILLER_32_159 ();
 sg13g2_fill_1 FILLER_32_194 ();
 sg13g2_fill_2 FILLER_32_211 ();
 sg13g2_decap_4 FILLER_32_268 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_fill_2 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_32_384 ();
 sg13g2_decap_8 FILLER_32_391 ();
 sg13g2_decap_8 FILLER_32_398 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_fill_2 FILLER_33_77 ();
 sg13g2_decap_4 FILLER_33_105 ();
 sg13g2_fill_2 FILLER_33_135 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_decap_4 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_151 ();
 sg13g2_fill_2 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_208 ();
 sg13g2_decap_4 FILLER_33_215 ();
 sg13g2_fill_2 FILLER_33_222 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_257 ();
 sg13g2_decap_8 FILLER_33_262 ();
 sg13g2_decap_8 FILLER_33_269 ();
 sg13g2_decap_8 FILLER_33_276 ();
 sg13g2_decap_4 FILLER_33_283 ();
 sg13g2_fill_1 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_4 FILLER_33_308 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_fill_2 FILLER_34_63 ();
 sg13g2_fill_2 FILLER_34_116 ();
 sg13g2_fill_1 FILLER_34_118 ();
 sg13g2_fill_1 FILLER_34_145 ();
 sg13g2_decap_4 FILLER_34_156 ();
 sg13g2_fill_1 FILLER_34_160 ();
 sg13g2_decap_4 FILLER_34_165 ();
 sg13g2_fill_1 FILLER_34_169 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_4 FILLER_34_189 ();
 sg13g2_fill_1 FILLER_34_193 ();
 sg13g2_fill_1 FILLER_34_197 ();
 sg13g2_decap_4 FILLER_34_202 ();
 sg13g2_fill_2 FILLER_34_206 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_fill_2 FILLER_34_238 ();
 sg13g2_fill_1 FILLER_34_240 ();
 sg13g2_fill_2 FILLER_34_250 ();
 sg13g2_decap_4 FILLER_34_278 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_decap_8 FILLER_34_309 ();
 sg13g2_decap_8 FILLER_34_316 ();
 sg13g2_decap_4 FILLER_34_323 ();
 sg13g2_fill_1 FILLER_34_327 ();
 sg13g2_decap_8 FILLER_34_340 ();
 sg13g2_decap_8 FILLER_34_347 ();
 sg13g2_fill_2 FILLER_34_354 ();
 sg13g2_fill_1 FILLER_34_356 ();
 sg13g2_decap_8 FILLER_34_397 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_65 ();
 sg13g2_fill_2 FILLER_35_92 ();
 sg13g2_fill_1 FILLER_35_104 ();
 sg13g2_decap_8 FILLER_35_141 ();
 sg13g2_decap_8 FILLER_35_148 ();
 sg13g2_fill_1 FILLER_35_155 ();
 sg13g2_fill_2 FILLER_35_160 ();
 sg13g2_decap_4 FILLER_35_191 ();
 sg13g2_fill_1 FILLER_35_195 ();
 sg13g2_decap_8 FILLER_35_222 ();
 sg13g2_decap_8 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_236 ();
 sg13g2_decap_8 FILLER_35_289 ();
 sg13g2_decap_4 FILLER_35_296 ();
 sg13g2_fill_1 FILLER_35_324 ();
 sg13g2_decap_8 FILLER_35_351 ();
 sg13g2_decap_8 FILLER_35_358 ();
 sg13g2_decap_8 FILLER_35_374 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_89 ();
 sg13g2_fill_2 FILLER_36_113 ();
 sg13g2_fill_1 FILLER_36_115 ();
 sg13g2_fill_2 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_134 ();
 sg13g2_decap_4 FILLER_36_157 ();
 sg13g2_fill_1 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_218 ();
 sg13g2_fill_2 FILLER_36_251 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_fill_2 FILLER_36_304 ();
 sg13g2_fill_1 FILLER_36_306 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_decap_4 FILLER_36_350 ();
 sg13g2_fill_2 FILLER_36_354 ();
 sg13g2_decap_8 FILLER_36_376 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_4 FILLER_37_77 ();
 sg13g2_fill_1 FILLER_37_81 ();
 sg13g2_fill_1 FILLER_37_92 ();
 sg13g2_decap_8 FILLER_37_99 ();
 sg13g2_decap_8 FILLER_37_106 ();
 sg13g2_decap_4 FILLER_37_113 ();
 sg13g2_decap_4 FILLER_37_169 ();
 sg13g2_fill_2 FILLER_37_181 ();
 sg13g2_fill_2 FILLER_37_226 ();
 sg13g2_decap_4 FILLER_37_249 ();
 sg13g2_fill_2 FILLER_37_253 ();
 sg13g2_decap_8 FILLER_37_290 ();
 sg13g2_decap_8 FILLER_37_297 ();
 sg13g2_fill_2 FILLER_37_304 ();
 sg13g2_fill_2 FILLER_37_311 ();
 sg13g2_fill_1 FILLER_37_313 ();
 sg13g2_fill_2 FILLER_37_337 ();
 sg13g2_fill_1 FILLER_37_339 ();
 sg13g2_fill_2 FILLER_37_366 ();
 sg13g2_decap_8 FILLER_37_394 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_4 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_67 ();
 sg13g2_fill_2 FILLER_38_95 ();
 sg13g2_decap_4 FILLER_38_103 ();
 sg13g2_decap_8 FILLER_38_117 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_fill_2 FILLER_38_131 ();
 sg13g2_decap_8 FILLER_38_169 ();
 sg13g2_decap_8 FILLER_38_176 ();
 sg13g2_decap_8 FILLER_38_183 ();
 sg13g2_decap_4 FILLER_38_190 ();
 sg13g2_fill_1 FILLER_38_209 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_4 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_decap_4 FILLER_38_274 ();
 sg13g2_fill_2 FILLER_38_278 ();
 sg13g2_decap_4 FILLER_38_291 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_313 ();
 sg13g2_fill_2 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_329 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_decap_4 FILLER_38_340 ();
 sg13g2_fill_1 FILLER_38_344 ();
 sg13g2_decap_4 FILLER_38_405 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_fill_1 FILLER_39_77 ();
 sg13g2_fill_2 FILLER_39_104 ();
 sg13g2_decap_4 FILLER_39_132 ();
 sg13g2_decap_8 FILLER_39_172 ();
 sg13g2_fill_2 FILLER_39_179 ();
 sg13g2_fill_2 FILLER_39_185 ();
 sg13g2_decap_8 FILLER_39_191 ();
 sg13g2_fill_1 FILLER_39_198 ();
 sg13g2_decap_8 FILLER_39_204 ();
 sg13g2_fill_1 FILLER_39_237 ();
 sg13g2_decap_8 FILLER_39_264 ();
 sg13g2_fill_2 FILLER_39_271 ();
 sg13g2_decap_4 FILLER_39_306 ();
 sg13g2_decap_8 FILLER_39_314 ();
 sg13g2_decap_4 FILLER_39_321 ();
 sg13g2_decap_4 FILLER_39_339 ();
 sg13g2_fill_1 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_370 ();
 sg13g2_decap_4 FILLER_39_377 ();
 sg13g2_fill_2 FILLER_39_381 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_fill_1 FILLER_40_97 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_fill_2 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_155 ();
 sg13g2_decap_4 FILLER_40_162 ();
 sg13g2_fill_1 FILLER_40_166 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_fill_1 FILLER_40_217 ();
 sg13g2_fill_2 FILLER_40_244 ();
 sg13g2_fill_1 FILLER_40_246 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_4 FILLER_40_280 ();
 sg13g2_fill_1 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_318 ();
 sg13g2_decap_4 FILLER_40_325 ();
 sg13g2_fill_2 FILLER_40_329 ();
 sg13g2_fill_1 FILLER_40_342 ();
 sg13g2_decap_8 FILLER_40_358 ();
 sg13g2_decap_8 FILLER_40_365 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_decap_8 FILLER_40_387 ();
 sg13g2_decap_8 FILLER_40_394 ();
 sg13g2_decap_8 FILLER_40_401 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_fill_1 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_102 ();
 sg13g2_fill_2 FILLER_41_109 ();
 sg13g2_fill_1 FILLER_41_111 ();
 sg13g2_fill_1 FILLER_41_122 ();
 sg13g2_fill_2 FILLER_41_134 ();
 sg13g2_fill_1 FILLER_41_136 ();
 sg13g2_decap_4 FILLER_41_228 ();
 sg13g2_fill_1 FILLER_41_232 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_fill_1 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_279 ();
 sg13g2_decap_8 FILLER_41_286 ();
 sg13g2_decap_8 FILLER_41_293 ();
 sg13g2_decap_8 FILLER_41_300 ();
 sg13g2_fill_2 FILLER_41_307 ();
 sg13g2_decap_8 FILLER_41_314 ();
 sg13g2_decap_8 FILLER_41_321 ();
 sg13g2_fill_2 FILLER_41_328 ();
 sg13g2_fill_1 FILLER_41_330 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_fill_1 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_359 ();
 sg13g2_fill_2 FILLER_41_366 ();
 sg13g2_fill_1 FILLER_41_368 ();
 sg13g2_decap_4 FILLER_41_377 ();
 sg13g2_fill_2 FILLER_41_381 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_4 FILLER_42_63 ();
 sg13g2_fill_2 FILLER_42_67 ();
 sg13g2_decap_8 FILLER_42_73 ();
 sg13g2_fill_2 FILLER_42_80 ();
 sg13g2_fill_1 FILLER_42_82 ();
 sg13g2_decap_4 FILLER_42_145 ();
 sg13g2_fill_1 FILLER_42_149 ();
 sg13g2_decap_8 FILLER_42_156 ();
 sg13g2_decap_8 FILLER_42_163 ();
 sg13g2_fill_1 FILLER_42_196 ();
 sg13g2_fill_1 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_decap_8 FILLER_42_277 ();
 sg13g2_decap_8 FILLER_42_284 ();
 sg13g2_decap_4 FILLER_42_302 ();
 sg13g2_fill_1 FILLER_42_306 ();
 sg13g2_fill_1 FILLER_42_317 ();
 sg13g2_decap_8 FILLER_42_344 ();
 sg13g2_decap_8 FILLER_42_351 ();
 sg13g2_decap_8 FILLER_42_358 ();
 sg13g2_decap_4 FILLER_42_403 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_4 FILLER_43_56 ();
 sg13g2_fill_2 FILLER_43_60 ();
 sg13g2_decap_4 FILLER_43_88 ();
 sg13g2_fill_1 FILLER_43_92 ();
 sg13g2_decap_8 FILLER_43_106 ();
 sg13g2_decap_4 FILLER_43_113 ();
 sg13g2_fill_2 FILLER_43_117 ();
 sg13g2_decap_8 FILLER_43_171 ();
 sg13g2_decap_8 FILLER_43_186 ();
 sg13g2_decap_4 FILLER_43_193 ();
 sg13g2_fill_2 FILLER_43_222 ();
 sg13g2_fill_1 FILLER_43_224 ();
 sg13g2_fill_1 FILLER_43_254 ();
 sg13g2_fill_2 FILLER_43_281 ();
 sg13g2_decap_8 FILLER_43_340 ();
 sg13g2_fill_2 FILLER_43_347 ();
 sg13g2_fill_1 FILLER_43_349 ();
 sg13g2_decap_8 FILLER_43_381 ();
 sg13g2_decap_8 FILLER_43_388 ();
 sg13g2_decap_8 FILLER_43_395 ();
 sg13g2_decap_8 FILLER_43_402 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_99 ();
 sg13g2_decap_8 FILLER_44_106 ();
 sg13g2_fill_1 FILLER_44_113 ();
 sg13g2_decap_8 FILLER_44_122 ();
 sg13g2_decap_4 FILLER_44_129 ();
 sg13g2_decap_8 FILLER_44_179 ();
 sg13g2_decap_8 FILLER_44_186 ();
 sg13g2_decap_8 FILLER_44_193 ();
 sg13g2_decap_8 FILLER_44_200 ();
 sg13g2_decap_8 FILLER_44_207 ();
 sg13g2_decap_8 FILLER_44_214 ();
 sg13g2_decap_8 FILLER_44_221 ();
 sg13g2_fill_2 FILLER_44_228 ();
 sg13g2_fill_2 FILLER_44_242 ();
 sg13g2_fill_2 FILLER_44_282 ();
 sg13g2_fill_1 FILLER_44_370 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_4 FILLER_45_56 ();
 sg13g2_fill_2 FILLER_45_102 ();
 sg13g2_fill_1 FILLER_45_104 ();
 sg13g2_decap_8 FILLER_45_131 ();
 sg13g2_decap_4 FILLER_45_138 ();
 sg13g2_fill_1 FILLER_45_142 ();
 sg13g2_fill_2 FILLER_45_149 ();
 sg13g2_fill_1 FILLER_45_151 ();
 sg13g2_decap_8 FILLER_45_157 ();
 sg13g2_decap_8 FILLER_45_164 ();
 sg13g2_decap_8 FILLER_45_171 ();
 sg13g2_fill_2 FILLER_45_178 ();
 sg13g2_decap_8 FILLER_45_206 ();
 sg13g2_decap_8 FILLER_45_213 ();
 sg13g2_decap_8 FILLER_45_220 ();
 sg13g2_fill_1 FILLER_45_227 ();
 sg13g2_fill_2 FILLER_45_254 ();
 sg13g2_fill_1 FILLER_45_256 ();
 sg13g2_fill_2 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_401 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_93 ();
 sg13g2_fill_2 FILLER_46_110 ();
 sg13g2_decap_8 FILLER_46_143 ();
 sg13g2_decap_8 FILLER_46_150 ();
 sg13g2_decap_4 FILLER_46_157 ();
 sg13g2_fill_2 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_fill_1 FILLER_46_175 ();
 sg13g2_fill_2 FILLER_46_179 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_fill_1 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_229 ();
 sg13g2_decap_8 FILLER_46_236 ();
 sg13g2_decap_8 FILLER_46_243 ();
 sg13g2_decap_8 FILLER_46_250 ();
 sg13g2_decap_8 FILLER_46_257 ();
 sg13g2_decap_8 FILLER_46_264 ();
 sg13g2_decap_8 FILLER_46_271 ();
 sg13g2_decap_8 FILLER_46_278 ();
 sg13g2_fill_2 FILLER_46_285 ();
 sg13g2_decap_8 FILLER_46_297 ();
 sg13g2_decap_8 FILLER_46_325 ();
 sg13g2_decap_8 FILLER_46_332 ();
 sg13g2_decap_4 FILLER_46_339 ();
 sg13g2_fill_2 FILLER_46_343 ();
 sg13g2_fill_2 FILLER_46_363 ();
 sg13g2_fill_2 FILLER_46_372 ();
 sg13g2_fill_1 FILLER_46_374 ();
 sg13g2_decap_8 FILLER_46_401 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_4 FILLER_47_70 ();
 sg13g2_fill_2 FILLER_47_74 ();
 sg13g2_fill_2 FILLER_47_86 ();
 sg13g2_decap_4 FILLER_47_109 ();
 sg13g2_fill_2 FILLER_47_113 ();
 sg13g2_fill_2 FILLER_47_125 ();
 sg13g2_fill_1 FILLER_47_132 ();
 sg13g2_fill_2 FILLER_47_141 ();
 sg13g2_fill_2 FILLER_47_184 ();
 sg13g2_fill_1 FILLER_47_186 ();
 sg13g2_decap_8 FILLER_47_199 ();
 sg13g2_decap_4 FILLER_47_206 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_305 ();
 sg13g2_decap_8 FILLER_47_320 ();
 sg13g2_fill_2 FILLER_47_327 ();
 sg13g2_fill_1 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_335 ();
 sg13g2_decap_8 FILLER_47_342 ();
 sg13g2_decap_4 FILLER_47_349 ();
 sg13g2_fill_1 FILLER_47_353 ();
 sg13g2_fill_2 FILLER_47_380 ();
 sg13g2_fill_1 FILLER_47_382 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_fill_2 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_110 ();
 sg13g2_fill_1 FILLER_48_117 ();
 sg13g2_decap_4 FILLER_48_126 ();
 sg13g2_fill_1 FILLER_48_154 ();
 sg13g2_fill_1 FILLER_48_204 ();
 sg13g2_fill_2 FILLER_48_297 ();
 sg13g2_fill_1 FILLER_48_299 ();
 sg13g2_fill_2 FILLER_48_312 ();
 sg13g2_fill_1 FILLER_48_340 ();
 sg13g2_decap_4 FILLER_48_351 ();
 sg13g2_fill_2 FILLER_48_355 ();
 sg13g2_decap_8 FILLER_48_362 ();
 sg13g2_fill_1 FILLER_48_369 ();
 sg13g2_fill_2 FILLER_48_381 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_4 FILLER_49_56 ();
 sg13g2_fill_2 FILLER_49_97 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_fill_1 FILLER_49_147 ();
 sg13g2_fill_2 FILLER_49_164 ();
 sg13g2_fill_2 FILLER_49_195 ();
 sg13g2_fill_2 FILLER_49_202 ();
 sg13g2_fill_1 FILLER_49_228 ();
 sg13g2_fill_2 FILLER_49_233 ();
 sg13g2_fill_1 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_266 ();
 sg13g2_fill_2 FILLER_49_273 ();
 sg13g2_fill_2 FILLER_49_293 ();
 sg13g2_fill_1 FILLER_49_295 ();
 sg13g2_decap_8 FILLER_49_374 ();
 sg13g2_fill_2 FILLER_49_381 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_4 FILLER_50_56 ();
 sg13g2_fill_1 FILLER_50_60 ();
 sg13g2_fill_2 FILLER_50_97 ();
 sg13g2_fill_1 FILLER_50_99 ();
 sg13g2_decap_4 FILLER_50_108 ();
 sg13g2_decap_4 FILLER_50_117 ();
 sg13g2_fill_1 FILLER_50_121 ();
 sg13g2_decap_8 FILLER_50_132 ();
 sg13g2_decap_8 FILLER_50_139 ();
 sg13g2_decap_8 FILLER_50_146 ();
 sg13g2_fill_1 FILLER_50_153 ();
 sg13g2_decap_4 FILLER_50_162 ();
 sg13g2_fill_1 FILLER_50_166 ();
 sg13g2_decap_4 FILLER_50_170 ();
 sg13g2_fill_2 FILLER_50_200 ();
 sg13g2_decap_8 FILLER_50_218 ();
 sg13g2_decap_8 FILLER_50_225 ();
 sg13g2_decap_8 FILLER_50_232 ();
 sg13g2_decap_4 FILLER_50_239 ();
 sg13g2_fill_2 FILLER_50_327 ();
 sg13g2_fill_1 FILLER_50_329 ();
 sg13g2_decap_4 FILLER_50_364 ();
 sg13g2_fill_2 FILLER_50_381 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_4 FILLER_51_77 ();
 sg13g2_fill_2 FILLER_51_91 ();
 sg13g2_fill_1 FILLER_51_93 ();
 sg13g2_fill_2 FILLER_51_109 ();
 sg13g2_fill_2 FILLER_51_137 ();
 sg13g2_fill_2 FILLER_51_144 ();
 sg13g2_fill_1 FILLER_51_146 ();
 sg13g2_decap_4 FILLER_51_155 ();
 sg13g2_fill_2 FILLER_51_159 ();
 sg13g2_fill_1 FILLER_51_174 ();
 sg13g2_decap_4 FILLER_51_210 ();
 sg13g2_decap_8 FILLER_51_234 ();
 sg13g2_decap_4 FILLER_51_241 ();
 sg13g2_fill_2 FILLER_51_245 ();
 sg13g2_decap_8 FILLER_51_286 ();
 sg13g2_decap_8 FILLER_51_293 ();
 sg13g2_decap_8 FILLER_51_300 ();
 sg13g2_fill_2 FILLER_51_307 ();
 sg13g2_decap_4 FILLER_51_314 ();
 sg13g2_decap_8 FILLER_51_323 ();
 sg13g2_decap_8 FILLER_51_330 ();
 sg13g2_decap_4 FILLER_51_337 ();
 sg13g2_fill_2 FILLER_51_341 ();
 sg13g2_decap_8 FILLER_51_348 ();
 sg13g2_decap_8 FILLER_51_391 ();
 sg13g2_decap_8 FILLER_51_398 ();
 sg13g2_decap_4 FILLER_51_405 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_fill_2 FILLER_52_118 ();
 sg13g2_fill_1 FILLER_52_133 ();
 sg13g2_fill_2 FILLER_52_144 ();
 sg13g2_fill_2 FILLER_52_183 ();
 sg13g2_decap_4 FILLER_52_189 ();
 sg13g2_decap_8 FILLER_52_245 ();
 sg13g2_fill_2 FILLER_52_252 ();
 sg13g2_fill_1 FILLER_52_254 ();
 sg13g2_decap_4 FILLER_52_263 ();
 sg13g2_decap_8 FILLER_52_272 ();
 sg13g2_decap_8 FILLER_52_279 ();
 sg13g2_decap_8 FILLER_52_291 ();
 sg13g2_fill_2 FILLER_52_312 ();
 sg13g2_fill_1 FILLER_52_314 ();
 sg13g2_decap_4 FILLER_52_341 ();
 sg13g2_fill_1 FILLER_52_350 ();
 sg13g2_decap_8 FILLER_52_387 ();
 sg13g2_decap_8 FILLER_52_394 ();
 sg13g2_decap_8 FILLER_52_401 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_fill_1 FILLER_53_84 ();
 sg13g2_decap_4 FILLER_53_95 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_4 FILLER_53_119 ();
 sg13g2_fill_1 FILLER_53_123 ();
 sg13g2_decap_8 FILLER_53_178 ();
 sg13g2_decap_8 FILLER_53_185 ();
 sg13g2_decap_4 FILLER_53_192 ();
 sg13g2_fill_1 FILLER_53_196 ();
 sg13g2_fill_1 FILLER_53_221 ();
 sg13g2_fill_2 FILLER_53_226 ();
 sg13g2_decap_8 FILLER_53_248 ();
 sg13g2_fill_2 FILLER_53_255 ();
 sg13g2_decap_4 FILLER_53_265 ();
 sg13g2_fill_1 FILLER_53_295 ();
 sg13g2_fill_2 FILLER_53_348 ();
 sg13g2_fill_1 FILLER_53_350 ();
 sg13g2_fill_2 FILLER_53_368 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_fill_2 FILLER_54_70 ();
 sg13g2_fill_1 FILLER_54_72 ();
 sg13g2_fill_2 FILLER_54_115 ();
 sg13g2_decap_4 FILLER_54_143 ();
 sg13g2_fill_1 FILLER_54_147 ();
 sg13g2_fill_2 FILLER_54_156 ();
 sg13g2_fill_1 FILLER_54_158 ();
 sg13g2_decap_8 FILLER_54_167 ();
 sg13g2_decap_8 FILLER_54_174 ();
 sg13g2_fill_2 FILLER_54_181 ();
 sg13g2_fill_1 FILLER_54_183 ();
 sg13g2_decap_8 FILLER_54_193 ();
 sg13g2_decap_8 FILLER_54_200 ();
 sg13g2_decap_8 FILLER_54_207 ();
 sg13g2_decap_4 FILLER_54_214 ();
 sg13g2_fill_1 FILLER_54_218 ();
 sg13g2_decap_4 FILLER_54_222 ();
 sg13g2_fill_1 FILLER_54_226 ();
 sg13g2_decap_4 FILLER_54_321 ();
 sg13g2_fill_2 FILLER_54_325 ();
 sg13g2_decap_4 FILLER_54_331 ();
 sg13g2_fill_2 FILLER_54_335 ();
 sg13g2_decap_4 FILLER_54_340 ();
 sg13g2_fill_1 FILLER_54_344 ();
 sg13g2_fill_1 FILLER_54_368 ();
 sg13g2_decap_8 FILLER_54_374 ();
 sg13g2_fill_2 FILLER_54_381 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_fill_2 FILLER_55_70 ();
 sg13g2_decap_4 FILLER_55_98 ();
 sg13g2_decap_4 FILLER_55_128 ();
 sg13g2_fill_1 FILLER_55_132 ();
 sg13g2_decap_8 FILLER_55_149 ();
 sg13g2_decap_8 FILLER_55_162 ();
 sg13g2_decap_4 FILLER_55_169 ();
 sg13g2_decap_4 FILLER_55_208 ();
 sg13g2_decap_8 FILLER_55_222 ();
 sg13g2_decap_8 FILLER_55_229 ();
 sg13g2_fill_2 FILLER_55_297 ();
 sg13g2_fill_1 FILLER_55_309 ();
 sg13g2_decap_8 FILLER_55_314 ();
 sg13g2_decap_8 FILLER_55_321 ();
 sg13g2_decap_8 FILLER_55_328 ();
 sg13g2_decap_4 FILLER_55_335 ();
 sg13g2_fill_1 FILLER_55_339 ();
 sg13g2_fill_1 FILLER_55_351 ();
 sg13g2_fill_1 FILLER_55_361 ();
 sg13g2_fill_1 FILLER_55_372 ();
 sg13g2_decap_8 FILLER_55_399 ();
 sg13g2_fill_2 FILLER_55_406 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_fill_1 FILLER_56_77 ();
 sg13g2_fill_1 FILLER_56_104 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_fill_2 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_145 ();
 sg13g2_fill_2 FILLER_56_188 ();
 sg13g2_fill_2 FILLER_56_216 ();
 sg13g2_fill_1 FILLER_56_238 ();
 sg13g2_decap_8 FILLER_56_265 ();
 sg13g2_fill_1 FILLER_56_272 ();
 sg13g2_fill_1 FILLER_56_299 ();
 sg13g2_decap_8 FILLER_56_334 ();
 sg13g2_fill_2 FILLER_56_341 ();
 sg13g2_fill_1 FILLER_56_343 ();
 sg13g2_fill_1 FILLER_56_357 ();
 sg13g2_decap_8 FILLER_56_394 ();
 sg13g2_decap_8 FILLER_56_401 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_4 FILLER_57_70 ();
 sg13g2_fill_2 FILLER_57_100 ();
 sg13g2_fill_1 FILLER_57_128 ();
 sg13g2_fill_2 FILLER_57_189 ();
 sg13g2_fill_2 FILLER_57_217 ();
 sg13g2_decap_4 FILLER_57_237 ();
 sg13g2_fill_1 FILLER_57_241 ();
 sg13g2_decap_8 FILLER_57_256 ();
 sg13g2_decap_4 FILLER_57_263 ();
 sg13g2_decap_4 FILLER_57_353 ();
 sg13g2_decap_8 FILLER_57_387 ();
 sg13g2_decap_8 FILLER_57_394 ();
 sg13g2_decap_8 FILLER_57_401 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_4 FILLER_58_70 ();
 sg13g2_fill_2 FILLER_58_74 ();
 sg13g2_decap_4 FILLER_58_112 ();
 sg13g2_fill_2 FILLER_58_116 ();
 sg13g2_fill_2 FILLER_58_190 ();
 sg13g2_fill_1 FILLER_58_192 ();
 sg13g2_fill_2 FILLER_58_198 ();
 sg13g2_fill_2 FILLER_58_213 ();
 sg13g2_decap_8 FILLER_58_241 ();
 sg13g2_decap_4 FILLER_58_248 ();
 sg13g2_decap_8 FILLER_58_278 ();
 sg13g2_decap_8 FILLER_58_285 ();
 sg13g2_fill_1 FILLER_58_292 ();
 sg13g2_fill_2 FILLER_58_311 ();
 sg13g2_decap_8 FILLER_58_339 ();
 sg13g2_decap_8 FILLER_58_346 ();
 sg13g2_fill_2 FILLER_58_353 ();
 sg13g2_fill_1 FILLER_58_355 ();
 sg13g2_decap_8 FILLER_58_373 ();
 sg13g2_fill_2 FILLER_58_380 ();
 sg13g2_fill_1 FILLER_58_382 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_fill_2 FILLER_59_84 ();
 sg13g2_fill_1 FILLER_59_86 ();
 sg13g2_decap_8 FILLER_59_92 ();
 sg13g2_decap_8 FILLER_59_99 ();
 sg13g2_decap_8 FILLER_59_106 ();
 sg13g2_decap_8 FILLER_59_113 ();
 sg13g2_decap_8 FILLER_59_120 ();
 sg13g2_decap_8 FILLER_59_127 ();
 sg13g2_fill_2 FILLER_59_150 ();
 sg13g2_decap_8 FILLER_59_173 ();
 sg13g2_decap_8 FILLER_59_180 ();
 sg13g2_decap_8 FILLER_59_187 ();
 sg13g2_decap_8 FILLER_59_194 ();
 sg13g2_decap_4 FILLER_59_205 ();
 sg13g2_fill_1 FILLER_59_209 ();
 sg13g2_decap_4 FILLER_59_215 ();
 sg13g2_fill_2 FILLER_59_228 ();
 sg13g2_fill_1 FILLER_59_230 ();
 sg13g2_fill_1 FILLER_59_250 ();
 sg13g2_decap_8 FILLER_59_259 ();
 sg13g2_decap_8 FILLER_59_266 ();
 sg13g2_decap_8 FILLER_59_273 ();
 sg13g2_decap_8 FILLER_59_280 ();
 sg13g2_decap_8 FILLER_59_287 ();
 sg13g2_decap_4 FILLER_59_294 ();
 sg13g2_fill_2 FILLER_59_303 ();
 sg13g2_fill_1 FILLER_59_305 ();
 sg13g2_decap_8 FILLER_59_310 ();
 sg13g2_decap_8 FILLER_59_317 ();
 sg13g2_fill_1 FILLER_59_324 ();
 sg13g2_decap_8 FILLER_59_351 ();
 sg13g2_decap_8 FILLER_59_358 ();
 sg13g2_decap_8 FILLER_59_365 ();
 sg13g2_decap_8 FILLER_59_372 ();
 sg13g2_decap_4 FILLER_59_379 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_fill_1 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_95 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_fill_1 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_130 ();
 sg13g2_fill_1 FILLER_60_137 ();
 sg13g2_decap_8 FILLER_60_144 ();
 sg13g2_decap_8 FILLER_60_151 ();
 sg13g2_decap_8 FILLER_60_158 ();
 sg13g2_fill_1 FILLER_60_165 ();
 sg13g2_fill_2 FILLER_60_171 ();
 sg13g2_fill_1 FILLER_60_173 ();
 sg13g2_decap_4 FILLER_60_177 ();
 sg13g2_decap_4 FILLER_60_215 ();
 sg13g2_fill_1 FILLER_60_219 ();
 sg13g2_fill_1 FILLER_60_246 ();
 sg13g2_fill_2 FILLER_60_277 ();
 sg13g2_fill_1 FILLER_60_279 ();
 sg13g2_fill_2 FILLER_60_289 ();
 sg13g2_decap_8 FILLER_60_304 ();
 sg13g2_decap_8 FILLER_60_311 ();
 sg13g2_decap_8 FILLER_60_318 ();
 sg13g2_fill_2 FILLER_60_359 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_4 FILLER_61_77 ();
 sg13g2_fill_1 FILLER_61_117 ();
 sg13g2_decap_4 FILLER_61_220 ();
 sg13g2_fill_2 FILLER_61_300 ();
 sg13g2_decap_4 FILLER_61_320 ();
 sg13g2_fill_2 FILLER_61_324 ();
 sg13g2_fill_1 FILLER_61_334 ();
 sg13g2_fill_2 FILLER_61_380 ();
 sg13g2_fill_1 FILLER_61_382 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_4 FILLER_62_70 ();
 sg13g2_fill_1 FILLER_62_106 ();
 sg13g2_fill_2 FILLER_62_133 ();
 sg13g2_fill_1 FILLER_62_135 ();
 sg13g2_decap_8 FILLER_62_162 ();
 sg13g2_decap_8 FILLER_62_172 ();
 sg13g2_decap_8 FILLER_62_179 ();
 sg13g2_decap_8 FILLER_62_186 ();
 sg13g2_decap_8 FILLER_62_193 ();
 sg13g2_fill_2 FILLER_62_233 ();
 sg13g2_fill_1 FILLER_62_235 ();
 sg13g2_decap_8 FILLER_62_246 ();
 sg13g2_decap_4 FILLER_62_294 ();
 sg13g2_fill_1 FILLER_62_303 ();
 sg13g2_fill_2 FILLER_62_330 ();
 sg13g2_fill_1 FILLER_62_358 ();
 sg13g2_fill_2 FILLER_62_369 ();
 sg13g2_fill_1 FILLER_62_371 ();
 sg13g2_decap_8 FILLER_62_398 ();
 sg13g2_decap_4 FILLER_62_405 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_4 FILLER_63_70 ();
 sg13g2_fill_1 FILLER_63_100 ();
 sg13g2_fill_2 FILLER_63_117 ();
 sg13g2_fill_1 FILLER_63_165 ();
 sg13g2_fill_1 FILLER_63_170 ();
 sg13g2_fill_2 FILLER_63_205 ();
 sg13g2_fill_1 FILLER_63_212 ();
 sg13g2_decap_4 FILLER_63_222 ();
 sg13g2_decap_8 FILLER_63_262 ();
 sg13g2_decap_8 FILLER_63_269 ();
 sg13g2_decap_8 FILLER_63_276 ();
 sg13g2_decap_4 FILLER_63_283 ();
 sg13g2_fill_1 FILLER_63_287 ();
 sg13g2_fill_2 FILLER_63_327 ();
 sg13g2_fill_1 FILLER_63_352 ();
 sg13g2_fill_2 FILLER_63_370 ();
 sg13g2_fill_2 FILLER_63_381 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_fill_2 FILLER_64_105 ();
 sg13g2_fill_1 FILLER_64_107 ();
 sg13g2_decap_4 FILLER_64_113 ();
 sg13g2_fill_2 FILLER_64_117 ();
 sg13g2_decap_8 FILLER_64_134 ();
 sg13g2_fill_2 FILLER_64_141 ();
 sg13g2_fill_1 FILLER_64_169 ();
 sg13g2_fill_1 FILLER_64_173 ();
 sg13g2_fill_2 FILLER_64_181 ();
 sg13g2_fill_1 FILLER_64_183 ();
 sg13g2_decap_8 FILLER_64_203 ();
 sg13g2_decap_4 FILLER_64_210 ();
 sg13g2_fill_2 FILLER_64_214 ();
 sg13g2_decap_8 FILLER_64_230 ();
 sg13g2_decap_8 FILLER_64_237 ();
 sg13g2_decap_8 FILLER_64_244 ();
 sg13g2_decap_8 FILLER_64_251 ();
 sg13g2_decap_8 FILLER_64_258 ();
 sg13g2_decap_8 FILLER_64_265 ();
 sg13g2_decap_4 FILLER_64_324 ();
 sg13g2_fill_1 FILLER_64_333 ();
 sg13g2_fill_2 FILLER_64_347 ();
 sg13g2_fill_1 FILLER_64_349 ();
 sg13g2_fill_1 FILLER_64_357 ();
 sg13g2_decap_8 FILLER_64_384 ();
 sg13g2_decap_8 FILLER_64_391 ();
 sg13g2_decap_8 FILLER_64_398 ();
 sg13g2_decap_4 FILLER_64_405 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_fill_2 FILLER_65_70 ();
 sg13g2_fill_1 FILLER_65_72 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_4 FILLER_65_129 ();
 sg13g2_fill_2 FILLER_65_133 ();
 sg13g2_decap_4 FILLER_65_157 ();
 sg13g2_fill_2 FILLER_65_161 ();
 sg13g2_fill_1 FILLER_65_194 ();
 sg13g2_fill_1 FILLER_65_221 ();
 sg13g2_decap_8 FILLER_65_240 ();
 sg13g2_fill_2 FILLER_65_304 ();
 sg13g2_decap_8 FILLER_65_316 ();
 sg13g2_decap_8 FILLER_65_323 ();
 sg13g2_decap_8 FILLER_65_330 ();
 sg13g2_decap_4 FILLER_65_337 ();
 sg13g2_fill_2 FILLER_65_341 ();
 sg13g2_decap_4 FILLER_65_353 ();
 sg13g2_fill_2 FILLER_65_357 ();
 sg13g2_decap_8 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_399 ();
 sg13g2_fill_2 FILLER_65_406 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_4 FILLER_66_70 ();
 sg13g2_fill_1 FILLER_66_74 ();
 sg13g2_fill_2 FILLER_66_117 ();
 sg13g2_decap_8 FILLER_66_145 ();
 sg13g2_decap_8 FILLER_66_152 ();
 sg13g2_fill_2 FILLER_66_159 ();
 sg13g2_fill_2 FILLER_66_239 ();
 sg13g2_fill_2 FILLER_66_267 ();
 sg13g2_fill_1 FILLER_66_269 ();
 sg13g2_fill_1 FILLER_66_288 ();
 sg13g2_fill_2 FILLER_66_294 ();
 sg13g2_fill_1 FILLER_66_301 ();
 sg13g2_decap_8 FILLER_66_311 ();
 sg13g2_decap_4 FILLER_66_318 ();
 sg13g2_fill_2 FILLER_66_327 ();
 sg13g2_fill_1 FILLER_66_329 ();
 sg13g2_fill_1 FILLER_66_335 ();
 sg13g2_fill_2 FILLER_66_349 ();
 sg13g2_fill_1 FILLER_66_351 ();
 sg13g2_decap_8 FILLER_66_369 ();
 sg13g2_decap_8 FILLER_66_376 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_120 ();
 sg13g2_decap_8 FILLER_67_127 ();
 sg13g2_decap_4 FILLER_67_134 ();
 sg13g2_fill_1 FILLER_67_138 ();
 sg13g2_decap_8 FILLER_67_175 ();
 sg13g2_fill_2 FILLER_67_182 ();
 sg13g2_fill_1 FILLER_67_184 ();
 sg13g2_decap_8 FILLER_67_197 ();
 sg13g2_fill_2 FILLER_67_213 ();
 sg13g2_decap_8 FILLER_67_275 ();
 sg13g2_decap_4 FILLER_67_282 ();
 sg13g2_decap_4 FILLER_67_290 ();
 sg13g2_fill_1 FILLER_67_294 ();
 sg13g2_decap_4 FILLER_67_306 ();
 sg13g2_fill_2 FILLER_67_341 ();
 sg13g2_fill_1 FILLER_67_343 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_fill_2 FILLER_68_84 ();
 sg13g2_decap_4 FILLER_68_126 ();
 sg13g2_fill_2 FILLER_68_162 ();
 sg13g2_decap_8 FILLER_68_173 ();
 sg13g2_decap_8 FILLER_68_180 ();
 sg13g2_fill_2 FILLER_68_187 ();
 sg13g2_fill_1 FILLER_68_189 ();
 sg13g2_decap_8 FILLER_68_195 ();
 sg13g2_decap_8 FILLER_68_202 ();
 sg13g2_decap_8 FILLER_68_209 ();
 sg13g2_fill_1 FILLER_68_216 ();
 sg13g2_decap_8 FILLER_68_226 ();
 sg13g2_decap_8 FILLER_68_233 ();
 sg13g2_decap_8 FILLER_68_240 ();
 sg13g2_fill_2 FILLER_68_247 ();
 sg13g2_fill_1 FILLER_68_249 ();
 sg13g2_decap_4 FILLER_68_255 ();
 sg13g2_fill_2 FILLER_68_259 ();
 sg13g2_decap_4 FILLER_68_287 ();
 sg13g2_fill_1 FILLER_68_291 ();
 sg13g2_fill_2 FILLER_68_298 ();
 sg13g2_fill_1 FILLER_68_300 ();
 sg13g2_decap_4 FILLER_68_343 ();
 sg13g2_fill_1 FILLER_68_347 ();
 sg13g2_decap_4 FILLER_68_371 ();
 sg13g2_fill_2 FILLER_68_380 ();
 sg13g2_fill_1 FILLER_68_382 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_fill_2 FILLER_69_70 ();
 sg13g2_decap_4 FILLER_69_98 ();
 sg13g2_fill_2 FILLER_69_102 ();
 sg13g2_fill_2 FILLER_69_114 ();
 sg13g2_decap_8 FILLER_69_160 ();
 sg13g2_decap_4 FILLER_69_167 ();
 sg13g2_fill_2 FILLER_69_205 ();
 sg13g2_decap_8 FILLER_69_211 ();
 sg13g2_fill_2 FILLER_69_218 ();
 sg13g2_decap_8 FILLER_69_224 ();
 sg13g2_decap_8 FILLER_69_231 ();
 sg13g2_decap_8 FILLER_69_238 ();
 sg13g2_decap_4 FILLER_69_245 ();
 sg13g2_decap_8 FILLER_69_253 ();
 sg13g2_decap_4 FILLER_69_260 ();
 sg13g2_fill_1 FILLER_69_264 ();
 sg13g2_fill_1 FILLER_69_291 ();
 sg13g2_decap_8 FILLER_69_304 ();
 sg13g2_fill_2 FILLER_69_311 ();
 sg13g2_fill_2 FILLER_69_321 ();
 sg13g2_decap_8 FILLER_69_349 ();
 sg13g2_fill_2 FILLER_69_361 ();
 sg13g2_fill_1 FILLER_69_363 ();
 sg13g2_decap_8 FILLER_69_390 ();
 sg13g2_decap_8 FILLER_69_397 ();
 sg13g2_decap_4 FILLER_69_404 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_fill_2 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_94 ();
 sg13g2_decap_8 FILLER_70_101 ();
 sg13g2_decap_4 FILLER_70_108 ();
 sg13g2_fill_2 FILLER_70_120 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_fill_1 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_144 ();
 sg13g2_decap_8 FILLER_70_151 ();
 sg13g2_decap_4 FILLER_70_158 ();
 sg13g2_fill_2 FILLER_70_162 ();
 sg13g2_decap_8 FILLER_70_174 ();
 sg13g2_fill_2 FILLER_70_181 ();
 sg13g2_decap_8 FILLER_70_232 ();
 sg13g2_fill_2 FILLER_70_239 ();
 sg13g2_fill_1 FILLER_70_241 ();
 sg13g2_decap_8 FILLER_70_250 ();
 sg13g2_fill_2 FILLER_70_257 ();
 sg13g2_fill_1 FILLER_70_259 ();
 sg13g2_decap_8 FILLER_70_269 ();
 sg13g2_fill_2 FILLER_70_276 ();
 sg13g2_fill_1 FILLER_70_278 ();
 sg13g2_fill_1 FILLER_70_284 ();
 sg13g2_decap_8 FILLER_70_316 ();
 sg13g2_decap_8 FILLER_70_323 ();
 sg13g2_decap_8 FILLER_70_330 ();
 sg13g2_decap_8 FILLER_70_337 ();
 sg13g2_decap_8 FILLER_70_344 ();
 sg13g2_decap_8 FILLER_70_351 ();
 sg13g2_fill_1 FILLER_70_358 ();
 sg13g2_fill_2 FILLER_70_364 ();
 sg13g2_fill_2 FILLER_70_379 ();
 sg13g2_fill_1 FILLER_70_381 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_fill_2 FILLER_71_77 ();
 sg13g2_fill_1 FILLER_71_79 ();
 sg13g2_decap_8 FILLER_71_90 ();
 sg13g2_decap_8 FILLER_71_97 ();
 sg13g2_decap_8 FILLER_71_104 ();
 sg13g2_decap_4 FILLER_71_111 ();
 sg13g2_fill_1 FILLER_71_115 ();
 sg13g2_fill_2 FILLER_71_121 ();
 sg13g2_fill_1 FILLER_71_123 ();
 sg13g2_decap_8 FILLER_71_137 ();
 sg13g2_decap_8 FILLER_71_190 ();
 sg13g2_fill_1 FILLER_71_205 ();
 sg13g2_fill_2 FILLER_71_242 ();
 sg13g2_fill_2 FILLER_71_270 ();
 sg13g2_fill_2 FILLER_71_279 ();
 sg13g2_decap_8 FILLER_71_297 ();
 sg13g2_decap_4 FILLER_71_304 ();
 sg13g2_decap_4 FILLER_71_348 ();
 sg13g2_fill_1 FILLER_71_357 ();
 sg13g2_fill_2 FILLER_71_368 ();
 sg13g2_fill_1 FILLER_71_370 ();
 sg13g2_fill_1 FILLER_71_380 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_4 FILLER_72_63 ();
 sg13g2_fill_1 FILLER_72_67 ();
 sg13g2_decap_4 FILLER_72_130 ();
 sg13g2_fill_2 FILLER_72_134 ();
 sg13g2_fill_2 FILLER_72_162 ();
 sg13g2_fill_1 FILLER_72_164 ();
 sg13g2_decap_8 FILLER_72_191 ();
 sg13g2_decap_8 FILLER_72_198 ();
 sg13g2_decap_8 FILLER_72_205 ();
 sg13g2_decap_8 FILLER_72_212 ();
 sg13g2_fill_1 FILLER_72_297 ();
 sg13g2_fill_2 FILLER_72_323 ();
 sg13g2_fill_1 FILLER_72_325 ();
 sg13g2_fill_1 FILLER_72_357 ();
 sg13g2_fill_2 FILLER_72_378 ();
 sg13g2_fill_1 FILLER_72_380 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_fill_2 FILLER_73_56 ();
 sg13g2_fill_1 FILLER_73_58 ();
 sg13g2_fill_1 FILLER_73_142 ();
 sg13g2_decap_4 FILLER_73_221 ();
 sg13g2_fill_1 FILLER_73_225 ();
 sg13g2_fill_2 FILLER_73_283 ();
 sg13g2_fill_1 FILLER_73_285 ();
 sg13g2_fill_2 FILLER_73_348 ();
 sg13g2_fill_1 FILLER_73_350 ();
 sg13g2_fill_2 FILLER_73_356 ();
 sg13g2_fill_1 FILLER_73_358 ();
 sg13g2_fill_2 FILLER_73_364 ();
 sg13g2_fill_1 FILLER_73_366 ();
 sg13g2_fill_2 FILLER_73_406 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_4 FILLER_74_70 ();
 sg13g2_decap_4 FILLER_74_104 ();
 sg13g2_fill_2 FILLER_74_123 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_4 FILLER_74_168 ();
 sg13g2_fill_2 FILLER_74_172 ();
 sg13g2_decap_4 FILLER_74_184 ();
 sg13g2_fill_1 FILLER_74_188 ();
 sg13g2_decap_8 FILLER_74_199 ();
 sg13g2_fill_1 FILLER_74_206 ();
 sg13g2_decap_8 FILLER_74_223 ();
 sg13g2_decap_8 FILLER_74_230 ();
 sg13g2_decap_8 FILLER_74_237 ();
 sg13g2_decap_8 FILLER_74_244 ();
 sg13g2_decap_8 FILLER_74_251 ();
 sg13g2_decap_8 FILLER_74_258 ();
 sg13g2_fill_2 FILLER_74_265 ();
 sg13g2_decap_8 FILLER_74_271 ();
 sg13g2_decap_8 FILLER_74_278 ();
 sg13g2_fill_1 FILLER_74_285 ();
 sg13g2_decap_4 FILLER_74_291 ();
 sg13g2_fill_1 FILLER_74_295 ();
 sg13g2_fill_2 FILLER_74_316 ();
 sg13g2_decap_8 FILLER_74_396 ();
 sg13g2_decap_4 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_fill_1 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_88 ();
 sg13g2_decap_8 FILLER_75_95 ();
 sg13g2_decap_8 FILLER_75_102 ();
 sg13g2_decap_8 FILLER_75_109 ();
 sg13g2_decap_8 FILLER_75_116 ();
 sg13g2_decap_8 FILLER_75_123 ();
 sg13g2_decap_8 FILLER_75_150 ();
 sg13g2_fill_2 FILLER_75_157 ();
 sg13g2_decap_4 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_232 ();
 sg13g2_decap_4 FILLER_75_270 ();
 sg13g2_fill_1 FILLER_75_274 ();
 sg13g2_fill_2 FILLER_75_280 ();
 sg13g2_decap_8 FILLER_75_291 ();
 sg13g2_decap_4 FILLER_75_298 ();
 sg13g2_fill_2 FILLER_75_302 ();
 sg13g2_decap_8 FILLER_75_308 ();
 sg13g2_fill_1 FILLER_75_315 ();
 sg13g2_decap_8 FILLER_75_337 ();
 sg13g2_decap_8 FILLER_75_344 ();
 sg13g2_decap_4 FILLER_75_351 ();
 sg13g2_fill_1 FILLER_75_355 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_fill_1 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_88 ();
 sg13g2_decap_8 FILLER_76_95 ();
 sg13g2_fill_1 FILLER_76_102 ();
 sg13g2_fill_2 FILLER_76_113 ();
 sg13g2_fill_1 FILLER_76_115 ();
 sg13g2_decap_4 FILLER_76_126 ();
 sg13g2_fill_2 FILLER_76_166 ();
 sg13g2_fill_1 FILLER_76_168 ();
 sg13g2_fill_2 FILLER_76_177 ();
 sg13g2_decap_8 FILLER_76_215 ();
 sg13g2_decap_4 FILLER_76_222 ();
 sg13g2_fill_1 FILLER_76_226 ();
 sg13g2_decap_8 FILLER_76_335 ();
 sg13g2_fill_2 FILLER_76_342 ();
 sg13g2_fill_2 FILLER_76_378 ();
 sg13g2_fill_1 FILLER_76_380 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_fill_2 FILLER_77_70 ();
 sg13g2_decap_4 FILLER_77_98 ();
 sg13g2_decap_4 FILLER_77_138 ();
 sg13g2_fill_1 FILLER_77_142 ();
 sg13g2_fill_1 FILLER_77_195 ();
 sg13g2_fill_1 FILLER_77_232 ();
 sg13g2_decap_4 FILLER_77_327 ();
 sg13g2_decap_4 FILLER_77_357 ();
 sg13g2_fill_1 FILLER_77_361 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_fill_2 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_4 FILLER_78_63 ();
 sg13g2_fill_1 FILLER_78_67 ();
 sg13g2_fill_2 FILLER_78_94 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_fill_2 FILLER_78_133 ();
 sg13g2_fill_1 FILLER_78_161 ();
 sg13g2_fill_2 FILLER_78_205 ();
 sg13g2_decap_8 FILLER_78_233 ();
 sg13g2_decap_8 FILLER_78_240 ();
 sg13g2_fill_1 FILLER_78_299 ();
 sg13g2_decap_4 FILLER_78_404 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_fill_2 FILLER_79_63 ();
 sg13g2_fill_2 FILLER_79_153 ();
 sg13g2_decap_4 FILLER_79_163 ();
 sg13g2_fill_1 FILLER_79_167 ();
 sg13g2_decap_8 FILLER_79_223 ();
 sg13g2_decap_8 FILLER_79_230 ();
 sg13g2_decap_8 FILLER_79_237 ();
 sg13g2_decap_8 FILLER_79_244 ();
 sg13g2_decap_4 FILLER_79_251 ();
 sg13g2_fill_2 FILLER_79_259 ();
 sg13g2_fill_1 FILLER_79_261 ();
 sg13g2_fill_2 FILLER_79_314 ();
 sg13g2_fill_1 FILLER_79_342 ();
 sg13g2_decap_8 FILLER_79_351 ();
 sg13g2_decap_8 FILLER_79_358 ();
 sg13g2_decap_8 FILLER_79_391 ();
 sg13g2_decap_8 FILLER_79_398 ();
 sg13g2_decap_4 FILLER_79_405 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_fill_2 FILLER_80_68 ();
 sg13g2_fill_1 FILLER_80_70 ();
 sg13g2_fill_1 FILLER_80_93 ();
 sg13g2_fill_2 FILLER_80_104 ();
 sg13g2_fill_2 FILLER_80_118 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_4 FILLER_80_180 ();
 sg13g2_decap_4 FILLER_80_188 ();
 sg13g2_decap_4 FILLER_80_196 ();
 sg13g2_decap_4 FILLER_80_204 ();
 sg13g2_decap_4 FILLER_80_212 ();
 sg13g2_decap_4 FILLER_80_220 ();
 sg13g2_decap_8 FILLER_80_228 ();
 sg13g2_decap_8 FILLER_80_235 ();
 sg13g2_decap_8 FILLER_80_242 ();
 sg13g2_decap_8 FILLER_80_249 ();
 sg13g2_decap_8 FILLER_80_256 ();
 sg13g2_decap_8 FILLER_80_263 ();
 sg13g2_decap_8 FILLER_80_270 ();
 sg13g2_decap_8 FILLER_80_277 ();
 sg13g2_decap_8 FILLER_80_284 ();
 sg13g2_decap_8 FILLER_80_291 ();
 sg13g2_decap_8 FILLER_80_298 ();
 sg13g2_decap_8 FILLER_80_305 ();
 sg13g2_decap_8 FILLER_80_312 ();
 sg13g2_decap_8 FILLER_80_319 ();
 sg13g2_decap_8 FILLER_80_326 ();
 sg13g2_decap_8 FILLER_80_333 ();
 sg13g2_decap_4 FILLER_80_340 ();
 sg13g2_decap_4 FILLER_80_348 ();
 sg13g2_decap_4 FILLER_80_356 ();
 sg13g2_decap_8 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_371 ();
 sg13g2_fill_2 FILLER_80_378 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
 assign uo_out[2] = net20;
 assign uo_out[3] = net21;
 assign uo_out[4] = net22;
 assign uo_out[5] = net23;
 assign uo_out[6] = net24;
 assign uo_out[7] = net25;
endmodule

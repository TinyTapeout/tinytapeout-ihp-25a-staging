module tt_um_spi_pwm_djuara (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire clknet_0_clk;
 wire \addr_reg_clk[0] ;
 wire \addr_reg_clk[1] ;
 wire \addr_reg_clk[2] ;
 wire \addr_reg_sampled[0] ;
 wire \addr_reg_sampled[1] ;
 wire \addr_reg_sampled[2] ;
 wire \cycles_freq[0] ;
 wire \cycles_freq[10] ;
 wire \cycles_freq[11] ;
 wire \cycles_freq[12] ;
 wire \cycles_freq[13] ;
 wire \cycles_freq[14] ;
 wire \cycles_freq[15] ;
 wire \cycles_freq[1] ;
 wire \cycles_freq[2] ;
 wire \cycles_freq[3] ;
 wire \cycles_freq[4] ;
 wire \cycles_freq[5] ;
 wire \cycles_freq[6] ;
 wire \cycles_freq[7] ;
 wire \cycles_freq[8] ;
 wire \cycles_freq[9] ;
 wire \cycles_high[0] ;
 wire \cycles_high[10] ;
 wire \cycles_high[11] ;
 wire \cycles_high[12] ;
 wire \cycles_high[13] ;
 wire \cycles_high[14] ;
 wire \cycles_high[15] ;
 wire \cycles_high[1] ;
 wire \cycles_high[2] ;
 wire \cycles_high[3] ;
 wire \cycles_high[4] ;
 wire \cycles_high[5] ;
 wire \cycles_high[6] ;
 wire \cycles_high[7] ;
 wire \cycles_high[8] ;
 wire \cycles_high[9] ;
 wire \data_wr_z1[0] ;
 wire \data_wr_z1[1] ;
 wire \data_wr_z1[2] ;
 wire \data_wr_z1[3] ;
 wire \data_wr_z1[4] ;
 wire \data_wr_z1[5] ;
 wire \data_wr_z1[6] ;
 wire \data_wr_z1[7] ;
 wire \dev_regs[0][0] ;
 wire \dev_regs[0][1] ;
 wire \dev_regs[0][2] ;
 wire \dev_regs[0][3] ;
 wire \dev_regs[0][4] ;
 wire \dev_regs[0][5] ;
 wire \dev_regs[0][6] ;
 wire \dev_regs[0][7] ;
 wire \dev_regs[1][0] ;
 wire \dev_regs[1][1] ;
 wire \dev_regs[1][2] ;
 wire \dev_regs[1][3] ;
 wire \dev_regs[1][4] ;
 wire \dev_regs[1][5] ;
 wire \dev_regs[1][6] ;
 wire \dev_regs[1][7] ;
 wire miso_clk;
 wire miso_sampled;
 wire pwm;
 wire \pwm_inst.counter[0] ;
 wire \pwm_inst.counter[10] ;
 wire \pwm_inst.counter[11] ;
 wire \pwm_inst.counter[12] ;
 wire \pwm_inst.counter[13] ;
 wire \pwm_inst.counter[14] ;
 wire \pwm_inst.counter[15] ;
 wire \pwm_inst.counter[1] ;
 wire \pwm_inst.counter[2] ;
 wire \pwm_inst.counter[3] ;
 wire \pwm_inst.counter[4] ;
 wire \pwm_inst.counter[5] ;
 wire \pwm_inst.counter[6] ;
 wire \pwm_inst.counter[7] ;
 wire \pwm_inst.counter[8] ;
 wire \pwm_inst.counter[9] ;
 wire \spi_own_clock_ins.data_rd[0] ;
 wire \spi_own_clock_ins.data_rd[1] ;
 wire \spi_own_clock_ins.data_rd[2] ;
 wire \spi_own_clock_ins.data_rd[3] ;
 wire \spi_own_clock_ins.data_rd[4] ;
 wire \spi_own_clock_ins.data_rd[5] ;
 wire \spi_own_clock_ins.data_rd[6] ;
 wire \spi_own_clock_ins.data_rd[7] ;
 wire \spi_own_clock_ins.data_rd_z1[0] ;
 wire \spi_own_clock_ins.data_rd_z1[1] ;
 wire \spi_own_clock_ins.data_rd_z1[2] ;
 wire \spi_own_clock_ins.data_rd_z1[3] ;
 wire \spi_own_clock_ins.data_rd_z1[4] ;
 wire \spi_own_clock_ins.data_rd_z1[5] ;
 wire \spi_own_clock_ins.data_rd_z1[6] ;
 wire \spi_own_clock_ins.data_rd_z1[7] ;
 wire \spi_own_clock_ins.index[0] ;
 wire \spi_own_clock_ins.index[1] ;
 wire \spi_own_clock_ins.index[2] ;
 wire \spi_own_clock_ins.index[3] ;
 wire \spi_own_clock_ins.spi_data_reg[0] ;
 wire \spi_own_clock_ins.spi_data_reg[1] ;
 wire \spi_own_clock_ins.spi_data_reg[2] ;
 wire \spi_own_clock_ins.spi_data_reg[3] ;
 wire \spi_own_clock_ins.spi_data_reg[4] ;
 wire \spi_own_clock_ins.spi_data_reg[5] ;
 wire \spi_own_clock_ins.spi_data_reg[6] ;
 wire \spi_own_clock_ins.spi_data_reg[7] ;
 wire \spi_own_clock_ins.spi_state[0] ;
 wire \spi_own_clock_ins.spi_state[1] ;
 wire \spi_own_clock_ins.spi_state[2] ;
 wire \spi_own_clock_ins.spi_state[3] ;
 wire \spi_sampled_ins.cs ;
 wire \spi_sampled_ins.cs_z1 ;
 wire \spi_sampled_ins.index[0] ;
 wire \spi_sampled_ins.index[1] ;
 wire \spi_sampled_ins.index[2] ;
 wire \spi_sampled_ins.index[3] ;
 wire \spi_sampled_ins.mosi ;
 wire \spi_sampled_ins.mosi_z1 ;
 wire \spi_sampled_ins.neg_edge_det.signal ;
 wire \spi_sampled_ins.neg_edge_det.signal_z1 ;
 wire \spi_sampled_ins.sclk_z1 ;
 wire \spi_sampled_ins.spi_data_reg[0] ;
 wire \spi_sampled_ins.spi_data_reg[1] ;
 wire \spi_sampled_ins.spi_data_reg[2] ;
 wire \spi_sampled_ins.spi_data_reg[3] ;
 wire \spi_sampled_ins.spi_data_reg[4] ;
 wire \spi_sampled_ins.spi_data_reg[5] ;
 wire \spi_sampled_ins.spi_data_reg[6] ;
 wire \spi_sampled_ins.spi_data_reg[7] ;
 wire \spi_sampled_ins.spi_state[0] ;
 wire \spi_sampled_ins.spi_state[1] ;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;

 sg13g2_inv_1 _0842_ (.Y(_0213_),
    .A(net115));
 sg13g2_inv_1 _0843_ (.Y(_0214_),
    .A(net164));
 sg13g2_inv_2 _0844_ (.Y(_0215_),
    .A(net170));
 sg13g2_inv_1 _0845_ (.Y(_0082_),
    .A(net285));
 sg13g2_inv_2 _0846_ (.Y(_0216_),
    .A(\addr_reg_clk[1] ));
 sg13g2_inv_1 _0847_ (.Y(_0217_),
    .A(\addr_reg_clk[0] ));
 sg13g2_inv_1 _0848_ (.Y(_0218_),
    .A(\spi_own_clock_ins.index[2] ));
 sg13g2_inv_1 _0849_ (.Y(_0219_),
    .A(\spi_own_clock_ins.index[1] ));
 sg13g2_inv_1 _0850_ (.Y(_0220_),
    .A(\spi_sampled_ins.spi_data_reg[7] ));
 sg13g2_inv_1 _0851_ (.Y(_0221_),
    .A(\spi_own_clock_ins.spi_state[1] ));
 sg13g2_inv_1 _0852_ (.Y(_0222_),
    .A(\spi_own_clock_ins.spi_state[3] ));
 sg13g2_inv_1 _0853_ (.Y(_0223_),
    .A(_0020_));
 sg13g2_inv_1 _0854_ (.Y(_0224_),
    .A(_0021_));
 sg13g2_inv_1 _0855_ (.Y(_0225_),
    .A(\cycles_freq[15] ));
 sg13g2_inv_1 _0856_ (.Y(_0226_),
    .A(\cycles_freq[14] ));
 sg13g2_inv_1 _0857_ (.Y(_0227_),
    .A(net161));
 sg13g2_inv_1 _0858_ (.Y(_0228_),
    .A(net130));
 sg13g2_inv_1 _0859_ (.Y(_0229_),
    .A(\cycles_freq[12] ));
 sg13g2_inv_2 _0860_ (.Y(_0230_),
    .A(net63));
 sg13g2_inv_2 _0861_ (.Y(_0231_),
    .A(net169));
 sg13g2_inv_2 _0862_ (.Y(_0232_),
    .A(net159));
 sg13g2_inv_2 _0863_ (.Y(_0233_),
    .A(net163));
 sg13g2_inv_2 _0864_ (.Y(_0234_),
    .A(net155));
 sg13g2_inv_1 _0865_ (.Y(_0235_),
    .A(\pwm_inst.counter[6] ));
 sg13g2_inv_1 _0866_ (.Y(_0236_),
    .A(\cycles_freq[5] ));
 sg13g2_inv_2 _0867_ (.Y(_0237_),
    .A(net153));
 sg13g2_inv_1 _0868_ (.Y(_0238_),
    .A(\cycles_freq[4] ));
 sg13g2_inv_1 _0869_ (.Y(_0239_),
    .A(net165));
 sg13g2_inv_1 _0870_ (.Y(_0240_),
    .A(net128));
 sg13g2_inv_1 _0871_ (.Y(_0241_),
    .A(\cycles_high[13] ));
 sg13g2_inv_1 _0872_ (.Y(_0242_),
    .A(\cycles_high[12] ));
 sg13g2_inv_1 _0873_ (.Y(_0243_),
    .A(\cycles_high[10] ));
 sg13g2_inv_1 _0874_ (.Y(_0244_),
    .A(net113));
 sg13g2_inv_1 _0875_ (.Y(_0245_),
    .A(\dev_regs[0][1] ));
 sg13g2_inv_1 _0876_ (.Y(_0246_),
    .A(\dev_regs[0][2] ));
 sg13g2_inv_1 _0877_ (.Y(_0247_),
    .A(\dev_regs[0][4] ));
 sg13g2_inv_1 _0878_ (.Y(_0248_),
    .A(\dev_regs[0][7] ));
 sg13g2_inv_1 _0879_ (.Y(_0069_),
    .A(net293));
 sg13g2_nor2b_1 _0880_ (.A(\spi_sampled_ins.spi_state[1] ),
    .B_N(\spi_sampled_ins.spi_state[0] ),
    .Y(_0249_));
 sg13g2_nand2b_2 _0881_ (.Y(_0250_),
    .B(\spi_sampled_ins.spi_state[0] ),
    .A_N(\spi_sampled_ins.spi_state[1] ));
 sg13g2_nor2b_2 _0882_ (.A(\spi_sampled_ins.spi_state[0] ),
    .B_N(\spi_sampled_ins.spi_state[1] ),
    .Y(_0251_));
 sg13g2_nor2_1 _0883_ (.A(_0249_),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_nand2b_1 _0884_ (.Y(_0253_),
    .B(\spi_sampled_ins.neg_edge_det.signal ),
    .A_N(\spi_sampled_ins.neg_edge_det.signal_z1 ));
 sg13g2_nand2_2 _0885_ (.Y(_0254_),
    .A(_0214_),
    .B(_0215_));
 sg13g2_nor3_2 _0886_ (.A(\spi_sampled_ins.index[2] ),
    .B(\spi_sampled_ins.index[1] ),
    .C(\spi_sampled_ins.index[0] ),
    .Y(_0255_));
 sg13g2_and2_1 _0887_ (.A(\spi_sampled_ins.index[3] ),
    .B(_0255_),
    .X(_0256_));
 sg13g2_nand2b_1 _0888_ (.Y(_0257_),
    .B(_0256_),
    .A_N(_0253_));
 sg13g2_and2_1 _0889_ (.A(_0252_),
    .B(_0257_),
    .X(_0258_));
 sg13g2_nand2_1 _0890_ (.Y(_0259_),
    .A(\spi_sampled_ins.index[1] ),
    .B(\spi_sampled_ins.index[0] ));
 sg13g2_nor2_1 _0891_ (.A(_0027_),
    .B(_0259_),
    .Y(_0260_));
 sg13g2_or2_1 _0892_ (.X(_0261_),
    .B(_0259_),
    .A(_0027_));
 sg13g2_nor2b_2 _0893_ (.A(net38),
    .B_N(net81),
    .Y(_0262_));
 sg13g2_nand2b_2 _0894_ (.Y(_0263_),
    .B(net81),
    .A_N(net38));
 sg13g2_o21ai_1 _0895_ (.B1(_0028_),
    .Y(_0264_),
    .A1(_0261_),
    .A2(_0263_));
 sg13g2_or2_1 _0896_ (.X(_0265_),
    .B(\spi_sampled_ins.spi_state[0] ),
    .A(\spi_sampled_ins.spi_state[1] ));
 sg13g2_nor2b_1 _0897_ (.A(\spi_sampled_ins.index[3] ),
    .B_N(_0255_),
    .Y(_0266_));
 sg13g2_nor2_1 _0898_ (.A(\spi_sampled_ins.spi_state[1] ),
    .B(_0266_),
    .Y(_0267_));
 sg13g2_nor2_1 _0899_ (.A(\spi_sampled_ins.spi_state[0] ),
    .B(_0256_),
    .Y(_0268_));
 sg13g2_nor2_1 _0900_ (.A(_0267_),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_a21oi_2 _0901_ (.B1(_0269_),
    .Y(_0270_),
    .A2(_0265_),
    .A1(_0253_));
 sg13g2_a22oi_1 _0902_ (.Y(_0271_),
    .B1(_0260_),
    .B2(_0251_),
    .A2(_0255_),
    .A1(_0249_));
 sg13g2_nand2b_1 _0903_ (.Y(_0272_),
    .B(_0028_),
    .A_N(_0271_));
 sg13g2_nor2_1 _0904_ (.A(_0250_),
    .B(_0255_),
    .Y(_0273_));
 sg13g2_a21oi_1 _0905_ (.A1(_0251_),
    .A2(_0261_),
    .Y(_0274_),
    .B1(_0273_));
 sg13g2_o21ai_1 _0906_ (.B1(_0272_),
    .Y(_0275_),
    .A1(_0028_),
    .A2(_0274_));
 sg13g2_a21oi_1 _0907_ (.A1(_0258_),
    .A2(_0264_),
    .Y(_0276_),
    .B1(_0275_));
 sg13g2_nor2_1 _0908_ (.A(net101),
    .B(_0270_),
    .Y(_0277_));
 sg13g2_a21oi_1 _0909_ (.A1(_0270_),
    .A2(_0276_),
    .Y(_0212_),
    .B1(_0277_));
 sg13g2_xor2_1 _0910_ (.B(_0254_),
    .A(_0027_),
    .X(_0278_));
 sg13g2_xnor2_1 _0911_ (.Y(_0279_),
    .A(_0027_),
    .B(_0259_));
 sg13g2_o21ai_1 _0912_ (.B1(_0252_),
    .Y(_0280_),
    .A1(_0220_),
    .A2(_0257_));
 sg13g2_nor2_2 _0913_ (.A(net101),
    .B(_0263_),
    .Y(_0281_));
 sg13g2_nor2b_1 _0914_ (.A(_0280_),
    .B_N(_0281_),
    .Y(_0282_));
 sg13g2_o21ai_1 _0915_ (.B1(_0279_),
    .Y(_0283_),
    .A1(_0251_),
    .A2(_0282_));
 sg13g2_o21ai_1 _0916_ (.B1(_0283_),
    .Y(_0284_),
    .A1(_0250_),
    .A2(_0278_));
 sg13g2_o21ai_1 _0917_ (.B1(_0270_),
    .Y(_0285_),
    .A1(_0280_),
    .A2(_0281_));
 sg13g2_a22oi_1 _0918_ (.Y(_0211_),
    .B1(_0285_),
    .B2(_0213_),
    .A2(_0284_),
    .A1(_0270_));
 sg13g2_nand2_1 _0919_ (.Y(_0286_),
    .A(\spi_sampled_ins.index[0] ),
    .B(_0281_));
 sg13g2_xnor2_1 _0920_ (.Y(_0287_),
    .A(\spi_sampled_ins.index[1] ),
    .B(_0286_));
 sg13g2_nand2_1 _0921_ (.Y(_0288_),
    .A(_0254_),
    .B(_0259_));
 sg13g2_nand2_1 _0922_ (.Y(_0289_),
    .A(_0251_),
    .B(_0288_));
 sg13g2_o21ai_1 _0923_ (.B1(_0289_),
    .Y(_0290_),
    .A1(_0250_),
    .A2(_0288_));
 sg13g2_nor2b_1 _0924_ (.A(_0290_),
    .B_N(_0270_),
    .Y(_0291_));
 sg13g2_o21ai_1 _0925_ (.B1(_0291_),
    .Y(_0292_),
    .A1(_0280_),
    .A2(_0287_));
 sg13g2_o21ai_1 _0926_ (.B1(_0292_),
    .Y(_0210_),
    .A1(_0214_),
    .A2(_0270_));
 sg13g2_a21oi_1 _0927_ (.A1(\spi_sampled_ins.index[0] ),
    .A2(_0281_),
    .Y(_0293_),
    .B1(_0256_));
 sg13g2_nand2b_1 _0928_ (.Y(_0294_),
    .B(_0258_),
    .A_N(_0293_));
 sg13g2_o21ai_1 _0929_ (.B1(_0294_),
    .Y(_0295_),
    .A1(_0215_),
    .A2(_0252_));
 sg13g2_nand2b_1 _0930_ (.Y(_0296_),
    .B(_0258_),
    .A_N(_0281_));
 sg13g2_nand2_1 _0931_ (.Y(_0297_),
    .A(_0270_),
    .B(_0296_));
 sg13g2_a22oi_1 _0932_ (.Y(_0209_),
    .B1(_0297_),
    .B2(_0215_),
    .A2(_0295_),
    .A1(_0270_));
 sg13g2_nor2_1 _0933_ (.A(\spi_sampled_ins.spi_state[1] ),
    .B(_0253_),
    .Y(_0298_));
 sg13g2_o21ai_1 _0934_ (.B1(_0298_),
    .Y(_0299_),
    .A1(_0250_),
    .A2(_0266_));
 sg13g2_nor2_1 _0935_ (.A(_0268_),
    .B(_0299_),
    .Y(_0300_));
 sg13g2_nand3_1 _0936_ (.B(_0250_),
    .C(_0300_),
    .A(net55),
    .Y(_0301_));
 sg13g2_nand2b_1 _0937_ (.Y(_0208_),
    .B(_0301_),
    .A_N(\spi_sampled_ins.spi_state[1] ));
 sg13g2_nor2_1 _0938_ (.A(net125),
    .B(_0220_),
    .Y(_0302_));
 sg13g2_a22oi_1 _0939_ (.Y(_0303_),
    .B1(_0300_),
    .B2(_0302_),
    .A2(_0299_),
    .A1(net125));
 sg13g2_inv_1 _0940_ (.Y(_0207_),
    .A(net126));
 sg13g2_nand2b_1 _0941_ (.Y(_0304_),
    .B(\spi_own_clock_ins.data_rd_z1[7] ),
    .A_N(net283));
 sg13g2_nor3_2 _0942_ (.A(\addr_reg_clk[1] ),
    .B(\addr_reg_clk[0] ),
    .C(_0223_),
    .Y(_0305_));
 sg13g2_nor2_1 _0943_ (.A(_0216_),
    .B(_0020_),
    .Y(_0306_));
 sg13g2_nor3_1 _0944_ (.A(_0216_),
    .B(\addr_reg_clk[0] ),
    .C(_0020_),
    .Y(_0307_));
 sg13g2_inv_1 _0945_ (.Y(_0308_),
    .A(_0307_));
 sg13g2_nor3_2 _0946_ (.A(\addr_reg_clk[1] ),
    .B(_0217_),
    .C(_0223_),
    .Y(_0309_));
 sg13g2_nor3_1 _0947_ (.A(\addr_reg_clk[1] ),
    .B(_0217_),
    .C(_0020_),
    .Y(_0310_));
 sg13g2_nand3_1 _0948_ (.B(\addr_reg_clk[1] ),
    .C(\addr_reg_clk[0] ),
    .A(\addr_reg_clk[2] ),
    .Y(_0311_));
 sg13g2_nor3_1 _0949_ (.A(\addr_reg_clk[2] ),
    .B(_0216_),
    .C(_0217_),
    .Y(_0312_));
 sg13g2_nor3_1 _0950_ (.A(_0216_),
    .B(\addr_reg_clk[0] ),
    .C(_0223_),
    .Y(_0313_));
 sg13g2_inv_1 _0951_ (.Y(_0314_),
    .A(net263));
 sg13g2_nand2_1 _0952_ (.Y(_0315_),
    .A(\cycles_high[7] ),
    .B(net263));
 sg13g2_nor3_1 _0953_ (.A(\addr_reg_clk[1] ),
    .B(\addr_reg_clk[0] ),
    .C(_0020_),
    .Y(_0316_));
 sg13g2_a22oi_1 _0954_ (.Y(_0317_),
    .B1(net264),
    .B2(\cycles_high[15] ),
    .A2(net267),
    .A1(uio_oe[7]));
 sg13g2_a22oi_1 _0955_ (.Y(_0318_),
    .B1(net274),
    .B2(\cycles_freq[7] ),
    .A2(net265),
    .A1(\cycles_freq[15] ));
 sg13g2_nand4_1 _0956_ (.B(_0315_),
    .C(_0317_),
    .A(net276),
    .Y(_0319_),
    .D(_0318_));
 sg13g2_a221oi_1 _0957_ (.B2(\dev_regs[1][7] ),
    .C1(_0319_),
    .B1(_0309_),
    .A1(\dev_regs[0][7] ),
    .Y(_0320_),
    .A2(net268));
 sg13g2_o21ai_1 _0958_ (.B1(net284),
    .Y(_0321_),
    .A1(net15),
    .A2(_0311_));
 sg13g2_o21ai_1 _0959_ (.B1(_0304_),
    .Y(_0206_),
    .A1(_0320_),
    .A2(_0321_));
 sg13g2_nand2b_1 _0960_ (.Y(_0322_),
    .B(\spi_own_clock_ins.data_rd_z1[6] ),
    .A_N(net281));
 sg13g2_nand2_1 _0961_ (.Y(_0323_),
    .A(\cycles_freq[14] ),
    .B(net265));
 sg13g2_a22oi_1 _0962_ (.Y(_0324_),
    .B1(net263),
    .B2(\cycles_high[6] ),
    .A2(net264),
    .A1(\cycles_high[14] ));
 sg13g2_a22oi_1 _0963_ (.Y(_0325_),
    .B1(net274),
    .B2(\cycles_freq[6] ),
    .A2(net266),
    .A1(\dev_regs[1][6] ));
 sg13g2_nand2_1 _0964_ (.Y(_0326_),
    .A(net276),
    .B(_0323_));
 sg13g2_a22oi_1 _0965_ (.Y(_0327_),
    .B1(net267),
    .B2(uio_oe[6]),
    .A2(net268),
    .A1(\dev_regs[0][6] ));
 sg13g2_nand3_1 _0966_ (.B(_0325_),
    .C(_0327_),
    .A(_0324_),
    .Y(_0328_));
 sg13g2_nor2_1 _0967_ (.A(_0326_),
    .B(_0328_),
    .Y(_0329_));
 sg13g2_o21ai_1 _0968_ (.B1(net284),
    .Y(_0330_),
    .A1(net14),
    .A2(_0311_));
 sg13g2_o21ai_1 _0969_ (.B1(_0322_),
    .Y(_0205_),
    .A1(_0329_),
    .A2(_0330_));
 sg13g2_nand2b_1 _0970_ (.Y(_0331_),
    .B(\spi_own_clock_ins.data_rd_z1[5] ),
    .A_N(net281));
 sg13g2_a22oi_1 _0971_ (.Y(_0332_),
    .B1(net267),
    .B2(uio_oe[5]),
    .A2(net268),
    .A1(\dev_regs[0][5] ));
 sg13g2_a22oi_1 _0972_ (.Y(_0333_),
    .B1(net264),
    .B2(\cycles_high[13] ),
    .A2(net266),
    .A1(\dev_regs[1][5] ));
 sg13g2_nand2_1 _0973_ (.Y(_0334_),
    .A(_0332_),
    .B(_0333_));
 sg13g2_nand2_1 _0974_ (.Y(_0335_),
    .A(\cycles_high[5] ),
    .B(net263));
 sg13g2_a22oi_1 _0975_ (.Y(_0336_),
    .B1(net274),
    .B2(\cycles_freq[5] ),
    .A2(net265),
    .A1(\cycles_freq[13] ));
 sg13g2_nand3_1 _0976_ (.B(_0335_),
    .C(_0336_),
    .A(net276),
    .Y(_0337_));
 sg13g2_nor2_1 _0977_ (.A(_0334_),
    .B(_0337_),
    .Y(_0338_));
 sg13g2_o21ai_1 _0978_ (.B1(net283),
    .Y(_0339_),
    .A1(net13),
    .A2(net275));
 sg13g2_o21ai_1 _0979_ (.B1(_0331_),
    .Y(_0204_),
    .A1(_0338_),
    .A2(_0339_));
 sg13g2_nand2b_1 _0980_ (.Y(_0340_),
    .B(\spi_own_clock_ins.data_rd_z1[4] ),
    .A_N(net283));
 sg13g2_a22oi_1 _0981_ (.Y(_0341_),
    .B1(net264),
    .B2(\cycles_high[12] ),
    .A2(net265),
    .A1(\cycles_freq[12] ));
 sg13g2_nand2_1 _0982_ (.Y(_0342_),
    .A(uio_oe[4]),
    .B(net267));
 sg13g2_a22oi_1 _0983_ (.Y(_0343_),
    .B1(net263),
    .B2(\cycles_high[4] ),
    .A2(net266),
    .A1(\dev_regs[1][4] ));
 sg13g2_a22oi_1 _0984_ (.Y(_0344_),
    .B1(net274),
    .B2(\cycles_freq[4] ),
    .A2(net268),
    .A1(\dev_regs[0][4] ));
 sg13g2_nand2_1 _0985_ (.Y(_0345_),
    .A(_0343_),
    .B(_0344_));
 sg13g2_nand3_1 _0986_ (.B(_0341_),
    .C(_0342_),
    .A(net276),
    .Y(_0346_));
 sg13g2_nor2_1 _0987_ (.A(_0345_),
    .B(_0346_),
    .Y(_0347_));
 sg13g2_o21ai_1 _0988_ (.B1(net283),
    .Y(_0348_),
    .A1(net12),
    .A2(net275));
 sg13g2_o21ai_1 _0989_ (.B1(_0340_),
    .Y(_0203_),
    .A1(_0347_),
    .A2(_0348_));
 sg13g2_nand2b_1 _0990_ (.Y(_0349_),
    .B(\spi_own_clock_ins.data_rd_z1[3] ),
    .A_N(net281));
 sg13g2_a22oi_1 _0991_ (.Y(_0350_),
    .B1(net265),
    .B2(\cycles_freq[11] ),
    .A2(net266),
    .A1(\dev_regs[1][3] ));
 sg13g2_a22oi_1 _0992_ (.Y(_0351_),
    .B1(_0313_),
    .B2(\cycles_high[3] ),
    .A2(_0312_),
    .A1(\cycles_high[11] ));
 sg13g2_nand2_1 _0993_ (.Y(_0352_),
    .A(_0350_),
    .B(_0351_));
 sg13g2_nand2_1 _0994_ (.Y(_0353_),
    .A(\cycles_freq[3] ),
    .B(_0316_));
 sg13g2_a22oi_1 _0995_ (.Y(_0354_),
    .B1(net267),
    .B2(uio_oe[3]),
    .A2(_0305_),
    .A1(\dev_regs[0][3] ));
 sg13g2_nand3_1 _0996_ (.B(_0353_),
    .C(_0354_),
    .A(net275),
    .Y(_0355_));
 sg13g2_nor2_1 _0997_ (.A(_0352_),
    .B(_0355_),
    .Y(_0356_));
 sg13g2_o21ai_1 _0998_ (.B1(net283),
    .Y(_0357_),
    .A1(net11),
    .A2(net275));
 sg13g2_o21ai_1 _0999_ (.B1(_0349_),
    .Y(_0202_),
    .A1(_0356_),
    .A2(_0357_));
 sg13g2_nand2b_1 _1000_ (.Y(_0358_),
    .B(\spi_own_clock_ins.data_rd_z1[2] ),
    .A_N(net284));
 sg13g2_nand2_1 _1001_ (.Y(_0359_),
    .A(\cycles_freq[10] ),
    .B(_0310_));
 sg13g2_a22oi_1 _1002_ (.Y(_0360_),
    .B1(net266),
    .B2(\dev_regs[1][2] ),
    .A2(_0305_),
    .A1(\dev_regs[0][2] ));
 sg13g2_a22oi_1 _1003_ (.Y(_0361_),
    .B1(net263),
    .B2(\cycles_high[2] ),
    .A2(net264),
    .A1(\cycles_high[10] ));
 sg13g2_nand4_1 _1004_ (.B(_0359_),
    .C(_0360_),
    .A(net276),
    .Y(_0362_),
    .D(_0361_));
 sg13g2_a221oi_1 _1005_ (.B2(\cycles_freq[2] ),
    .C1(_0362_),
    .B1(net274),
    .A1(uio_oe[2]),
    .Y(_0363_),
    .A2(net267));
 sg13g2_o21ai_1 _1006_ (.B1(net283),
    .Y(_0364_),
    .A1(net10),
    .A2(net275));
 sg13g2_o21ai_1 _1007_ (.B1(_0358_),
    .Y(_0201_),
    .A1(_0363_),
    .A2(_0364_));
 sg13g2_nand2b_1 _1008_ (.Y(_0365_),
    .B(\spi_own_clock_ins.data_rd_z1[1] ),
    .A_N(net284));
 sg13g2_nand2_1 _1009_ (.Y(_0366_),
    .A(\cycles_freq[9] ),
    .B(net265));
 sg13g2_a22oi_1 _1010_ (.Y(_0367_),
    .B1(net264),
    .B2(\cycles_high[9] ),
    .A2(net268),
    .A1(\dev_regs[0][1] ));
 sg13g2_a22oi_1 _1011_ (.Y(_0368_),
    .B1(net274),
    .B2(\cycles_freq[1] ),
    .A2(net267),
    .A1(uio_oe[1]));
 sg13g2_nand4_1 _1012_ (.B(_0366_),
    .C(_0367_),
    .A(net276),
    .Y(_0369_),
    .D(_0368_));
 sg13g2_a221oi_1 _1013_ (.B2(\cycles_high[1] ),
    .C1(_0369_),
    .B1(net263),
    .A1(\dev_regs[1][1] ),
    .Y(_0370_),
    .A2(net266));
 sg13g2_o21ai_1 _1014_ (.B1(net283),
    .Y(_0371_),
    .A1(net9),
    .A2(net275));
 sg13g2_o21ai_1 _1015_ (.B1(_0365_),
    .Y(_0200_),
    .A1(_0370_),
    .A2(_0371_));
 sg13g2_nand2b_1 _1016_ (.Y(_0372_),
    .B(\spi_own_clock_ins.data_rd_z1[0] ),
    .A_N(net284));
 sg13g2_nand2_1 _1017_ (.Y(_0373_),
    .A(\cycles_freq[8] ),
    .B(net265));
 sg13g2_a22oi_1 _1018_ (.Y(_0374_),
    .B1(net263),
    .B2(\cycles_high[0] ),
    .A2(net264),
    .A1(\cycles_high[8] ));
 sg13g2_a22oi_1 _1019_ (.Y(_0375_),
    .B1(net274),
    .B2(\cycles_freq[0] ),
    .A2(net267),
    .A1(uio_oe[0]));
 sg13g2_nand4_1 _1020_ (.B(_0373_),
    .C(_0374_),
    .A(net276),
    .Y(_0376_),
    .D(_0375_));
 sg13g2_a221oi_1 _1021_ (.B2(\dev_regs[1][0] ),
    .C1(_0376_),
    .B1(net266),
    .A1(\dev_regs[0][0] ),
    .Y(_0377_),
    .A2(net268));
 sg13g2_o21ai_1 _1022_ (.B1(net283),
    .Y(_0378_),
    .A1(net8),
    .A2(net275));
 sg13g2_o21ai_1 _1023_ (.B1(_0372_),
    .Y(_0199_),
    .A1(_0377_),
    .A2(_0378_));
 sg13g2_or2_1 _1024_ (.X(_0379_),
    .B(_0265_),
    .A(_0257_));
 sg13g2_mux2_1 _1025_ (.A0(net76),
    .A1(\addr_reg_sampled[2] ),
    .S(_0379_),
    .X(_0198_));
 sg13g2_mux2_1 _1026_ (.A0(net74),
    .A1(\addr_reg_sampled[1] ),
    .S(_0379_),
    .X(_0197_));
 sg13g2_mux2_1 _1027_ (.A0(net71),
    .A1(\addr_reg_sampled[0] ),
    .S(_0379_),
    .X(_0196_));
 sg13g2_mux2_1 _1028_ (.A0(\spi_own_clock_ins.data_rd[7] ),
    .A1(\spi_own_clock_ins.data_rd_z1[7] ),
    .S(net282),
    .X(_0195_));
 sg13g2_mux2_1 _1029_ (.A0(\spi_own_clock_ins.data_rd[6] ),
    .A1(\spi_own_clock_ins.data_rd_z1[6] ),
    .S(net281),
    .X(_0194_));
 sg13g2_mux2_1 _1030_ (.A0(\spi_own_clock_ins.data_rd[5] ),
    .A1(\spi_own_clock_ins.data_rd_z1[5] ),
    .S(net281),
    .X(_0193_));
 sg13g2_mux2_1 _1031_ (.A0(\spi_own_clock_ins.data_rd[4] ),
    .A1(\spi_own_clock_ins.data_rd_z1[4] ),
    .S(net281),
    .X(_0192_));
 sg13g2_mux2_1 _1032_ (.A0(\spi_own_clock_ins.data_rd[3] ),
    .A1(\spi_own_clock_ins.data_rd_z1[3] ),
    .S(net281),
    .X(_0191_));
 sg13g2_mux2_1 _1033_ (.A0(\spi_own_clock_ins.data_rd[2] ),
    .A1(\spi_own_clock_ins.data_rd_z1[2] ),
    .S(net281),
    .X(_0190_));
 sg13g2_mux2_1 _1034_ (.A0(\spi_own_clock_ins.data_rd[1] ),
    .A1(\spi_own_clock_ins.data_rd_z1[1] ),
    .S(net284),
    .X(_0189_));
 sg13g2_mux2_1 _1035_ (.A0(\spi_own_clock_ins.data_rd[0] ),
    .A1(\spi_own_clock_ins.data_rd_z1[0] ),
    .S(net284),
    .X(_0188_));
 sg13g2_nor2_1 _1036_ (.A(\spi_own_clock_ins.index[1] ),
    .B(\spi_own_clock_ins.index[0] ),
    .Y(_0380_));
 sg13g2_nor3_1 _1037_ (.A(\spi_own_clock_ins.index[2] ),
    .B(\spi_own_clock_ins.index[1] ),
    .C(\spi_own_clock_ins.index[0] ),
    .Y(_0381_));
 sg13g2_nand2_2 _1038_ (.Y(_0382_),
    .A(_0218_),
    .B(_0380_));
 sg13g2_and2_2 _1039_ (.A(\spi_own_clock_ins.index[3] ),
    .B(_0381_),
    .X(_0383_));
 sg13g2_nand2_1 _1040_ (.Y(_0384_),
    .A(\spi_own_clock_ins.index[3] ),
    .B(_0381_));
 sg13g2_nand2_2 _1041_ (.Y(_0385_),
    .A(\spi_own_clock_ins.spi_state[0] ),
    .B(_0383_));
 sg13g2_mux2_1 _1042_ (.A0(\spi_own_clock_ins.spi_data_reg[2] ),
    .A1(\addr_reg_clk[2] ),
    .S(_0385_),
    .X(_0186_));
 sg13g2_nor2_1 _1043_ (.A(\spi_own_clock_ins.spi_data_reg[1] ),
    .B(_0385_),
    .Y(_0386_));
 sg13g2_a21oi_1 _1044_ (.A1(_0216_),
    .A2(_0385_),
    .Y(_0185_),
    .B1(_0386_));
 sg13g2_nor2_1 _1045_ (.A(\spi_own_clock_ins.spi_data_reg[0] ),
    .B(_0385_),
    .Y(_0387_));
 sg13g2_a21oi_1 _1046_ (.A1(_0217_),
    .A2(_0385_),
    .Y(_0184_),
    .B1(_0387_));
 sg13g2_nor4_1 _1047_ (.A(net282),
    .B(\spi_own_clock_ins.spi_state[1] ),
    .C(\spi_own_clock_ins.spi_state[3] ),
    .D(\spi_own_clock_ins.spi_state[0] ),
    .Y(_0388_));
 sg13g2_nand2_2 _1048_ (.Y(_0389_),
    .A(\spi_own_clock_ins.spi_state[3] ),
    .B(_0383_));
 sg13g2_nand2b_1 _1049_ (.Y(_0390_),
    .B(_0389_),
    .A_N(_0388_));
 sg13g2_nor3_1 _1050_ (.A(\spi_own_clock_ins.index[3] ),
    .B(_0023_),
    .C(_0382_),
    .Y(_0391_));
 sg13g2_nor2_1 _1051_ (.A(_0390_),
    .B(_0391_),
    .Y(_0392_));
 sg13g2_inv_1 _1052_ (.Y(_0393_),
    .A(_0392_));
 sg13g2_a21oi_1 _1053_ (.A1(_0026_),
    .A2(_0382_),
    .Y(_0394_),
    .B1(_0221_));
 sg13g2_o21ai_1 _1054_ (.B1(_0394_),
    .Y(_0395_),
    .A1(_0026_),
    .A2(_0382_));
 sg13g2_o21ai_1 _1055_ (.B1(_0022_),
    .Y(_0396_),
    .A1(\spi_own_clock_ins.spi_state[1] ),
    .A2(\spi_own_clock_ins.spi_state[3] ));
 sg13g2_a21oi_1 _1056_ (.A1(_0384_),
    .A2(_0396_),
    .Y(_0397_),
    .B1(\spi_own_clock_ins.spi_state[3] ));
 sg13g2_nand2_1 _1057_ (.Y(_0398_),
    .A(\spi_own_clock_ins.index[1] ),
    .B(net280));
 sg13g2_nor2_1 _1058_ (.A(_0025_),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_xor2_1 _1059_ (.B(_0399_),
    .A(_0026_),
    .X(_0400_));
 sg13g2_o21ai_1 _1060_ (.B1(_0395_),
    .Y(_0401_),
    .A1(_0397_),
    .A2(_0400_));
 sg13g2_a22oi_1 _1061_ (.Y(_0402_),
    .B1(_0392_),
    .B2(_0401_),
    .A2(_0390_),
    .A1(\spi_own_clock_ins.index[3] ));
 sg13g2_inv_1 _1062_ (.Y(_0183_),
    .A(_0402_));
 sg13g2_nand3_1 _1063_ (.B(_0222_),
    .C(_0022_),
    .A(_0221_),
    .Y(_0403_));
 sg13g2_nand2_1 _1064_ (.Y(_0404_),
    .A(net282),
    .B(_0383_));
 sg13g2_xor2_1 _1065_ (.B(_0380_),
    .A(_0025_),
    .X(_0405_));
 sg13g2_o21ai_1 _1066_ (.B1(_0404_),
    .Y(_0406_),
    .A1(_0221_),
    .A2(_0405_));
 sg13g2_nor2_1 _1067_ (.A(_0384_),
    .B(_0403_),
    .Y(_0407_));
 sg13g2_nand3b_1 _1068_ (.B(_0222_),
    .C(_0403_),
    .Y(_0408_),
    .A_N(net282));
 sg13g2_nand2_1 _1069_ (.Y(_0409_),
    .A(_0025_),
    .B(_0398_));
 sg13g2_nand3b_1 _1070_ (.B(_0408_),
    .C(_0409_),
    .Y(_0410_),
    .A_N(_0399_));
 sg13g2_o21ai_1 _1071_ (.B1(_0392_),
    .Y(_0411_),
    .A1(_0407_),
    .A2(_0410_));
 sg13g2_a21oi_1 _1072_ (.A1(_0403_),
    .A2(_0406_),
    .Y(_0412_),
    .B1(_0411_));
 sg13g2_a21oi_1 _1073_ (.A1(_0218_),
    .A2(_0393_),
    .Y(_0182_),
    .B1(_0412_));
 sg13g2_xor2_1 _1074_ (.B(net280),
    .A(\spi_own_clock_ins.index[1] ),
    .X(_0413_));
 sg13g2_o21ai_1 _1075_ (.B1(_0404_),
    .Y(_0414_),
    .A1(_0221_),
    .A2(_0413_));
 sg13g2_a221oi_1 _1076_ (.B2(_0403_),
    .C1(_0393_),
    .B1(_0414_),
    .A1(_0408_),
    .Y(_0415_),
    .A2(_0413_));
 sg13g2_a21oi_1 _1077_ (.A1(_0219_),
    .A2(_0393_),
    .Y(_0181_),
    .B1(_0415_));
 sg13g2_nor4_1 _1078_ (.A(net282),
    .B(\spi_own_clock_ins.spi_state[1] ),
    .C(\spi_own_clock_ins.spi_state[3] ),
    .D(_0022_),
    .Y(_0416_));
 sg13g2_nor3_1 _1079_ (.A(net280),
    .B(_0393_),
    .C(_0416_),
    .Y(_0417_));
 sg13g2_a21o_1 _1080_ (.A2(_0393_),
    .A1(net280),
    .B1(_0417_),
    .X(_0180_));
 sg13g2_a21oi_1 _1081_ (.A1(\spi_own_clock_ins.spi_state[0] ),
    .A2(_0384_),
    .Y(_0048_),
    .B1(_0391_));
 sg13g2_nor2_1 _1082_ (.A(net59),
    .B(_0263_),
    .Y(_0418_));
 sg13g2_a21oi_1 _1083_ (.A1(_0220_),
    .A2(_0263_),
    .Y(_0116_),
    .B1(net60));
 sg13g2_mux2_1 _1084_ (.A0(net59),
    .A1(net85),
    .S(_0262_),
    .X(_0115_));
 sg13g2_mux2_1 _1085_ (.A0(net85),
    .A1(net79),
    .S(_0262_),
    .X(_0114_));
 sg13g2_mux2_1 _1086_ (.A0(net79),
    .A1(\spi_sampled_ins.spi_data_reg[3] ),
    .S(_0262_),
    .X(_0113_));
 sg13g2_mux2_1 _1087_ (.A0(net76),
    .A1(net89),
    .S(_0263_),
    .X(_0112_));
 sg13g2_mux2_1 _1088_ (.A0(net76),
    .A1(net74),
    .S(_0262_),
    .X(_0111_));
 sg13g2_mux2_1 _1089_ (.A0(net74),
    .A1(net71),
    .S(_0262_),
    .X(_0110_));
 sg13g2_mux2_1 _1090_ (.A0(\spi_sampled_ins.spi_data_reg[0] ),
    .A1(net67),
    .S(_0262_),
    .X(_0109_));
 sg13g2_o21ai_1 _1091_ (.B1(\spi_own_clock_ins.spi_state[1] ),
    .Y(_0419_),
    .A1(\spi_own_clock_ins.index[3] ),
    .A2(_0382_));
 sg13g2_nand2_1 _1092_ (.Y(_0001_),
    .A(_0404_),
    .B(_0419_));
 sg13g2_o21ai_1 _1093_ (.B1(_0222_),
    .Y(_0003_),
    .A1(\spi_own_clock_ins.spi_data_reg[7] ),
    .A2(_0385_));
 sg13g2_nand3_1 _1094_ (.B(\spi_own_clock_ins.spi_state[0] ),
    .C(_0383_),
    .A(\spi_own_clock_ins.spi_data_reg[7] ),
    .Y(_0420_));
 sg13g2_o21ai_1 _1095_ (.B1(_0420_),
    .Y(_0002_),
    .A1(_0022_),
    .A2(_0383_));
 sg13g2_nand2_1 _1096_ (.Y(_0421_),
    .A(net1),
    .B(net7));
 sg13g2_nor2_1 _1097_ (.A(net268),
    .B(_0389_),
    .Y(_0422_));
 sg13g2_nand2_1 _1098_ (.Y(_0423_),
    .A(_0309_),
    .B(net251));
 sg13g2_nor2b_1 _1099_ (.A(\addr_reg_sampled[1] ),
    .B_N(\addr_reg_sampled[0] ),
    .Y(_0424_));
 sg13g2_nor2b_1 _1100_ (.A(\addr_reg_sampled[2] ),
    .B_N(_0424_),
    .Y(_0425_));
 sg13g2_nor2_1 _1101_ (.A(\addr_reg_sampled[1] ),
    .B(\addr_reg_sampled[0] ),
    .Y(_0426_));
 sg13g2_and2_1 _1102_ (.A(_0251_),
    .B(_0256_),
    .X(_0427_));
 sg13g2_o21ai_1 _1103_ (.B1(net257),
    .Y(_0428_),
    .A1(net268),
    .A2(_0389_));
 sg13g2_a21oi_2 _1104_ (.B1(_0428_),
    .Y(_0429_),
    .A2(_0426_),
    .A1(_0021_));
 sg13g2_a22oi_1 _1105_ (.Y(_0430_),
    .B1(net262),
    .B2(_0429_),
    .A2(net254),
    .A1(net266));
 sg13g2_nand2b_1 _1106_ (.Y(_0431_),
    .B(net257),
    .A_N(net55));
 sg13g2_nand3_1 _1107_ (.B(_0429_),
    .C(_0431_),
    .A(_0425_),
    .Y(_0432_));
 sg13g2_o21ai_1 _1108_ (.B1(_0432_),
    .Y(_0433_),
    .A1(net151),
    .A2(_0423_));
 sg13g2_a21oi_1 _1109_ (.A1(_0421_),
    .A2(net250),
    .Y(_0000_),
    .B1(_0433_));
 sg13g2_nand2b_1 _1110_ (.Y(_0434_),
    .B(\pwm_inst.counter[2] ),
    .A_N(\cycles_high[2] ));
 sg13g2_nand2b_1 _1111_ (.Y(_0435_),
    .B(\pwm_inst.counter[3] ),
    .A_N(\cycles_high[3] ));
 sg13g2_nand2_1 _1112_ (.Y(_0436_),
    .A(_0434_),
    .B(_0435_));
 sg13g2_nand2b_1 _1113_ (.Y(_0437_),
    .B(\cycles_high[3] ),
    .A_N(\pwm_inst.counter[3] ));
 sg13g2_nand2b_1 _1114_ (.Y(_0438_),
    .B(\pwm_inst.counter[1] ),
    .A_N(\cycles_high[1] ));
 sg13g2_nor2b_1 _1115_ (.A(net278),
    .B_N(\cycles_high[1] ),
    .Y(_0439_));
 sg13g2_nor2b_1 _1116_ (.A(\pwm_inst.counter[0] ),
    .B_N(\cycles_high[0] ),
    .Y(_0440_));
 sg13g2_o21ai_1 _1117_ (.B1(_0438_),
    .Y(_0441_),
    .A1(_0439_),
    .A2(_0440_));
 sg13g2_nand2b_1 _1118_ (.Y(_0442_),
    .B(\cycles_high[2] ),
    .A_N(\pwm_inst.counter[2] ));
 sg13g2_and4_1 _1119_ (.A(_0434_),
    .B(_0435_),
    .C(_0437_),
    .D(_0442_),
    .X(_0443_));
 sg13g2_a22oi_1 _1120_ (.Y(_0444_),
    .B1(_0441_),
    .B2(_0443_),
    .A2(_0437_),
    .A1(_0436_));
 sg13g2_nor2_1 _1121_ (.A(_0237_),
    .B(\cycles_high[4] ),
    .Y(_0445_));
 sg13g2_nand2_1 _1122_ (.Y(_0446_),
    .A(_0237_),
    .B(\cycles_high[4] ));
 sg13g2_nand2b_1 _1123_ (.Y(_0447_),
    .B(\cycles_high[5] ),
    .A_N(\pwm_inst.counter[5] ));
 sg13g2_nand3b_1 _1124_ (.B(_0446_),
    .C(_0447_),
    .Y(_0448_),
    .A_N(_0445_));
 sg13g2_nor2b_1 _1125_ (.A(\cycles_high[5] ),
    .B_N(net277),
    .Y(_0449_));
 sg13g2_a21oi_1 _1126_ (.A1(_0445_),
    .A2(_0447_),
    .Y(_0450_),
    .B1(_0449_));
 sg13g2_o21ai_1 _1127_ (.B1(_0450_),
    .Y(_0451_),
    .A1(_0444_),
    .A2(_0448_));
 sg13g2_nor2_1 _1128_ (.A(_0235_),
    .B(\cycles_high[6] ),
    .Y(_0452_));
 sg13g2_nand2_1 _1129_ (.Y(_0453_),
    .A(_0234_),
    .B(\cycles_high[7] ));
 sg13g2_o21ai_1 _1130_ (.B1(_0453_),
    .Y(_0454_),
    .A1(\pwm_inst.counter[6] ),
    .A2(_0244_));
 sg13g2_nor2_1 _1131_ (.A(_0452_),
    .B(_0454_),
    .Y(_0455_));
 sg13g2_nor2_1 _1132_ (.A(_0234_),
    .B(\cycles_high[7] ),
    .Y(_0456_));
 sg13g2_a221oi_1 _1133_ (.B2(_0451_),
    .C1(_0456_),
    .B1(_0455_),
    .A1(_0452_),
    .Y(_0457_),
    .A2(_0453_));
 sg13g2_nor2_1 _1134_ (.A(_0233_),
    .B(\cycles_high[8] ),
    .Y(_0458_));
 sg13g2_nand2_1 _1135_ (.Y(_0459_),
    .A(_0232_),
    .B(\cycles_high[9] ));
 sg13g2_a22oi_1 _1136_ (.Y(_0460_),
    .B1(\cycles_high[8] ),
    .B2(_0233_),
    .A2(\cycles_high[9] ),
    .A1(_0232_));
 sg13g2_nand2b_1 _1137_ (.Y(_0461_),
    .B(_0460_),
    .A_N(_0458_));
 sg13g2_nor2_1 _1138_ (.A(_0232_),
    .B(\cycles_high[9] ),
    .Y(_0462_));
 sg13g2_a21oi_1 _1139_ (.A1(_0458_),
    .A2(_0459_),
    .Y(_0463_),
    .B1(_0462_));
 sg13g2_o21ai_1 _1140_ (.B1(_0463_),
    .Y(_0464_),
    .A1(_0457_),
    .A2(_0461_));
 sg13g2_nor2_1 _1141_ (.A(_0230_),
    .B(\cycles_high[11] ),
    .Y(_0465_));
 sg13g2_nor2_1 _1142_ (.A(_0231_),
    .B(\cycles_high[10] ),
    .Y(_0466_));
 sg13g2_nand2_1 _1143_ (.Y(_0467_),
    .A(_0230_),
    .B(\cycles_high[11] ));
 sg13g2_o21ai_1 _1144_ (.B1(_0467_),
    .Y(_0468_),
    .A1(\pwm_inst.counter[10] ),
    .A2(_0243_));
 sg13g2_nor3_1 _1145_ (.A(_0465_),
    .B(_0466_),
    .C(_0468_),
    .Y(_0469_));
 sg13g2_a221oi_1 _1146_ (.B2(_0464_),
    .C1(_0465_),
    .B1(_0469_),
    .A1(_0466_),
    .Y(_0470_),
    .A2(_0467_));
 sg13g2_nand2b_1 _1147_ (.Y(_0471_),
    .B(\pwm_inst.counter[15] ),
    .A_N(\cycles_high[15] ));
 sg13g2_o21ai_1 _1148_ (.B1(_0471_),
    .Y(_0472_),
    .A1(_0227_),
    .A2(\cycles_high[14] ));
 sg13g2_nand2b_1 _1149_ (.Y(_0473_),
    .B(\cycles_high[15] ),
    .A_N(\pwm_inst.counter[15] ));
 sg13g2_a21oi_1 _1150_ (.A1(_0227_),
    .A2(\cycles_high[14] ),
    .Y(_0474_),
    .B1(_0472_));
 sg13g2_and2_1 _1151_ (.A(_0473_),
    .B(_0474_),
    .X(_0475_));
 sg13g2_a22oi_1 _1152_ (.Y(_0476_),
    .B1(_0242_),
    .B2(\pwm_inst.counter[12] ),
    .A2(_0241_),
    .A1(\pwm_inst.counter[13] ));
 sg13g2_nand2b_1 _1153_ (.Y(_0477_),
    .B(\cycles_high[12] ),
    .A_N(\pwm_inst.counter[12] ));
 sg13g2_nand2_1 _1154_ (.Y(_0478_),
    .A(_0228_),
    .B(\cycles_high[13] ));
 sg13g2_nand4_1 _1155_ (.B(_0476_),
    .C(_0477_),
    .A(_0475_),
    .Y(_0479_),
    .D(_0478_));
 sg13g2_nor2b_1 _1156_ (.A(_0476_),
    .B_N(_0478_),
    .Y(_0480_));
 sg13g2_a22oi_1 _1157_ (.Y(_0481_),
    .B1(_0475_),
    .B2(_0480_),
    .A2(_0473_),
    .A1(_0472_));
 sg13g2_o21ai_1 _1158_ (.B1(_0481_),
    .Y(_0482_),
    .A1(_0470_),
    .A2(_0479_));
 sg13g2_nand2b_1 _1159_ (.Y(_0483_),
    .B(\pwm_inst.counter[10] ),
    .A_N(\cycles_freq[10] ));
 sg13g2_o21ai_1 _1160_ (.B1(_0483_),
    .Y(_0484_),
    .A1(\cycles_freq[11] ),
    .A2(_0230_));
 sg13g2_nand2_1 _1161_ (.Y(_0485_),
    .A(\cycles_freq[11] ),
    .B(_0230_));
 sg13g2_a22oi_1 _1162_ (.Y(_0486_),
    .B1(\cycles_freq[9] ),
    .B2(_0232_),
    .A2(_0231_),
    .A1(\cycles_freq[10] ));
 sg13g2_nand2_1 _1163_ (.Y(_0487_),
    .A(_0485_),
    .B(_0486_));
 sg13g2_nand2b_1 _1164_ (.Y(_0488_),
    .B(\pwm_inst.counter[8] ),
    .A_N(\cycles_freq[8] ));
 sg13g2_o21ai_1 _1165_ (.B1(_0488_),
    .Y(_0489_),
    .A1(\cycles_freq[9] ),
    .A2(_0232_));
 sg13g2_nand2b_1 _1166_ (.Y(_0490_),
    .B(net278),
    .A_N(\cycles_freq[1] ));
 sg13g2_nor2b_1 _1167_ (.A(\pwm_inst.counter[0] ),
    .B_N(\cycles_freq[0] ),
    .Y(_0491_));
 sg13g2_nor2b_1 _1168_ (.A(net278),
    .B_N(\cycles_freq[1] ),
    .Y(_0492_));
 sg13g2_a221oi_1 _1169_ (.B2(_0491_),
    .C1(_0492_),
    .B1(_0490_),
    .A1(\cycles_freq[2] ),
    .Y(_0493_),
    .A2(_0240_));
 sg13g2_nand2b_1 _1170_ (.Y(_0494_),
    .B(\pwm_inst.counter[2] ),
    .A_N(\cycles_freq[2] ));
 sg13g2_o21ai_1 _1171_ (.B1(_0494_),
    .Y(_0495_),
    .A1(\cycles_freq[3] ),
    .A2(_0239_));
 sg13g2_a22oi_1 _1172_ (.Y(_0496_),
    .B1(\cycles_freq[3] ),
    .B2(_0239_),
    .A2(\cycles_freq[4] ),
    .A1(_0237_));
 sg13g2_o21ai_1 _1173_ (.B1(_0496_),
    .Y(_0497_),
    .A1(_0493_),
    .A2(_0495_));
 sg13g2_a22oi_1 _1174_ (.Y(_0498_),
    .B1(\pwm_inst.counter[4] ),
    .B2(_0238_),
    .A2(net277),
    .A1(_0236_));
 sg13g2_nor2_1 _1175_ (.A(_0236_),
    .B(net277),
    .Y(_0499_));
 sg13g2_a221oi_1 _1176_ (.B2(_0498_),
    .C1(_0499_),
    .B1(_0497_),
    .A1(\cycles_freq[6] ),
    .Y(_0500_),
    .A2(_0235_));
 sg13g2_nand2b_1 _1177_ (.Y(_0501_),
    .B(\pwm_inst.counter[6] ),
    .A_N(\cycles_freq[6] ));
 sg13g2_o21ai_1 _1178_ (.B1(_0501_),
    .Y(_0502_),
    .A1(\cycles_freq[7] ),
    .A2(_0234_));
 sg13g2_nor2_1 _1179_ (.A(_0500_),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_a22oi_1 _1180_ (.Y(_0504_),
    .B1(\cycles_freq[7] ),
    .B2(_0234_),
    .A2(\cycles_freq[8] ),
    .A1(_0233_));
 sg13g2_a22oi_1 _1181_ (.Y(_0505_),
    .B1(_0226_),
    .B2(\pwm_inst.counter[14] ),
    .A2(_0225_),
    .A1(\pwm_inst.counter[15] ));
 sg13g2_nor2_1 _1182_ (.A(\pwm_inst.counter[15] ),
    .B(_0225_),
    .Y(_0506_));
 sg13g2_nor2b_1 _1183_ (.A(_0506_),
    .B_N(_0505_),
    .Y(_0507_));
 sg13g2_o21ai_1 _1184_ (.B1(_0507_),
    .Y(_0508_),
    .A1(_0226_),
    .A2(\pwm_inst.counter[14] ));
 sg13g2_nand2_1 _1185_ (.Y(_0509_),
    .A(\pwm_inst.counter[12] ),
    .B(_0229_));
 sg13g2_o21ai_1 _1186_ (.B1(_0509_),
    .Y(_0510_),
    .A1(\cycles_freq[13] ),
    .A2(_0228_));
 sg13g2_nand2_1 _1187_ (.Y(_0511_),
    .A(\cycles_freq[13] ),
    .B(_0228_));
 sg13g2_o21ai_1 _1188_ (.B1(_0511_),
    .Y(_0512_),
    .A1(\pwm_inst.counter[12] ),
    .A2(_0229_));
 sg13g2_nor2_1 _1189_ (.A(_0484_),
    .B(_0487_),
    .Y(_0513_));
 sg13g2_nand3b_1 _1190_ (.B(_0504_),
    .C(_0513_),
    .Y(_0514_),
    .A_N(_0489_));
 sg13g2_a22oi_1 _1191_ (.Y(_0515_),
    .B1(_0489_),
    .B2(_0513_),
    .A2(_0485_),
    .A1(_0484_));
 sg13g2_o21ai_1 _1192_ (.B1(_0515_),
    .Y(_0516_),
    .A1(_0503_),
    .A2(_0514_));
 sg13g2_nor3_1 _1193_ (.A(_0508_),
    .B(_0510_),
    .C(_0512_),
    .Y(_0517_));
 sg13g2_nand3b_1 _1194_ (.B(_0510_),
    .C(_0511_),
    .Y(_0518_),
    .A_N(_0508_));
 sg13g2_o21ai_1 _1195_ (.B1(_0518_),
    .Y(_0519_),
    .A1(_0505_),
    .A2(_0506_));
 sg13g2_a21o_2 _1196_ (.A2(_0517_),
    .A1(_0516_),
    .B1(_0519_),
    .X(_0520_));
 sg13g2_nor2_1 _1197_ (.A(net6),
    .B(\dev_regs[1][0] ),
    .Y(_0521_));
 sg13g2_or2_1 _1198_ (.X(_0522_),
    .B(net117),
    .A(net6));
 sg13g2_nand2b_1 _1199_ (.Y(_0523_),
    .B(_0522_),
    .A_N(net149));
 sg13g2_a21oi_1 _1200_ (.A1(net240),
    .A2(_0520_),
    .Y(_0004_),
    .B1(_0523_));
 sg13g2_nand2_1 _1201_ (.Y(_0524_),
    .A(net278),
    .B(\pwm_inst.counter[0] ));
 sg13g2_o21ai_1 _1202_ (.B1(_0522_),
    .Y(_0525_),
    .A1(net278),
    .A2(net149));
 sg13g2_a221oi_1 _1203_ (.B2(net249),
    .C1(_0525_),
    .B1(net240),
    .A1(net278),
    .Y(_0011_),
    .A2(net149));
 sg13g2_nand3_1 _1204_ (.B(net278),
    .C(net149),
    .A(net128),
    .Y(_0526_));
 sg13g2_nand2_1 _1205_ (.Y(_0527_),
    .A(net272),
    .B(_0526_));
 sg13g2_a221oi_1 _1206_ (.B2(_0240_),
    .C1(_0527_),
    .B1(_0524_),
    .A1(net240),
    .Y(_0012_),
    .A2(net249));
 sg13g2_nand4_1 _1207_ (.B(net128),
    .C(net278),
    .A(net165),
    .Y(_0528_),
    .D(\pwm_inst.counter[0] ));
 sg13g2_a21oi_1 _1208_ (.A1(_0239_),
    .A2(_0526_),
    .Y(_0529_),
    .B1(_0521_));
 sg13g2_nand2_1 _1209_ (.Y(_0530_),
    .A(_0528_),
    .B(net166));
 sg13g2_a21oi_1 _1210_ (.A1(_0482_),
    .A2(net249),
    .Y(_0013_),
    .B1(net167));
 sg13g2_nor2_2 _1211_ (.A(_0237_),
    .B(_0528_),
    .Y(_0531_));
 sg13g2_a21oi_1 _1212_ (.A1(_0237_),
    .A2(_0528_),
    .Y(_0532_),
    .B1(net273));
 sg13g2_nand2b_1 _1213_ (.Y(_0533_),
    .B(net154),
    .A_N(_0531_));
 sg13g2_a21oi_1 _1214_ (.A1(_0482_),
    .A2(_0520_),
    .Y(_0014_),
    .B1(_0533_));
 sg13g2_o21ai_1 _1215_ (.B1(net272),
    .Y(_0534_),
    .A1(net277),
    .A2(_0531_));
 sg13g2_a221oi_1 _1216_ (.B2(net277),
    .C1(_0534_),
    .B1(_0531_),
    .A1(net240),
    .Y(_0015_),
    .A2(net249));
 sg13g2_nand3_1 _1217_ (.B(net277),
    .C(_0531_),
    .A(net168),
    .Y(_0535_));
 sg13g2_a21o_1 _1218_ (.A2(_0531_),
    .A1(net277),
    .B1(net168),
    .X(_0536_));
 sg13g2_nand3_1 _1219_ (.B(_0535_),
    .C(_0536_),
    .A(net272),
    .Y(_0537_));
 sg13g2_a21oi_1 _1220_ (.A1(net239),
    .A2(net248),
    .Y(_0016_),
    .B1(_0537_));
 sg13g2_nand4_1 _1221_ (.B(net172),
    .C(net277),
    .A(net155),
    .Y(_0538_),
    .D(_0531_));
 sg13g2_a21oi_1 _1222_ (.A1(_0234_),
    .A2(_0535_),
    .Y(_0539_),
    .B1(net273));
 sg13g2_nand2_1 _1223_ (.Y(_0540_),
    .A(_0538_),
    .B(net156));
 sg13g2_a21oi_1 _1224_ (.A1(net239),
    .A2(net248),
    .Y(_0017_),
    .B1(_0540_));
 sg13g2_a21oi_1 _1225_ (.A1(_0233_),
    .A2(_0538_),
    .Y(_0541_),
    .B1(net273));
 sg13g2_o21ai_1 _1226_ (.B1(_0541_),
    .Y(_0542_),
    .A1(_0233_),
    .A2(_0538_));
 sg13g2_a21oi_1 _1227_ (.A1(net239),
    .A2(net248),
    .Y(_0018_),
    .B1(_0542_));
 sg13g2_or3_2 _1228_ (.A(_0232_),
    .B(_0233_),
    .C(_0538_),
    .X(_0543_));
 sg13g2_o21ai_1 _1229_ (.B1(_0232_),
    .Y(_0544_),
    .A1(_0233_),
    .A2(_0538_));
 sg13g2_nand3_1 _1230_ (.B(_0543_),
    .C(net160),
    .A(net272),
    .Y(_0545_));
 sg13g2_a21oi_1 _1231_ (.A1(net240),
    .A2(net249),
    .Y(_0019_),
    .B1(_0545_));
 sg13g2_nor2_1 _1232_ (.A(_0231_),
    .B(_0543_),
    .Y(_0546_));
 sg13g2_a21oi_1 _1233_ (.A1(_0231_),
    .A2(_0543_),
    .Y(_0547_),
    .B1(net273));
 sg13g2_nand2b_1 _1234_ (.Y(_0548_),
    .B(_0547_),
    .A_N(_0546_));
 sg13g2_a21oi_1 _1235_ (.A1(net240),
    .A2(net249),
    .Y(_0005_),
    .B1(_0548_));
 sg13g2_nor3_2 _1236_ (.A(_0230_),
    .B(_0231_),
    .C(_0543_),
    .Y(_0549_));
 sg13g2_o21ai_1 _1237_ (.B1(net272),
    .Y(_0550_),
    .A1(net63),
    .A2(_0546_));
 sg13g2_a221oi_1 _1238_ (.B2(net63),
    .C1(_0550_),
    .B1(_0546_),
    .A1(net239),
    .Y(_0006_),
    .A2(net248));
 sg13g2_nand2_1 _1239_ (.Y(_0551_),
    .A(\pwm_inst.counter[12] ),
    .B(_0549_));
 sg13g2_o21ai_1 _1240_ (.B1(net272),
    .Y(_0552_),
    .A1(net143),
    .A2(_0549_));
 sg13g2_a221oi_1 _1241_ (.B2(net143),
    .C1(_0552_),
    .B1(_0549_),
    .A1(net239),
    .Y(_0007_),
    .A2(net248));
 sg13g2_nand3_1 _1242_ (.B(\pwm_inst.counter[12] ),
    .C(_0549_),
    .A(net130),
    .Y(_0553_));
 sg13g2_nand2_1 _1243_ (.Y(_0554_),
    .A(net272),
    .B(_0553_));
 sg13g2_a221oi_1 _1244_ (.B2(_0228_),
    .C1(_0554_),
    .B1(_0551_),
    .A1(net239),
    .Y(_0008_),
    .A2(net248));
 sg13g2_nor2_1 _1245_ (.A(_0227_),
    .B(_0553_),
    .Y(_0555_));
 sg13g2_a21oi_1 _1246_ (.A1(_0227_),
    .A2(_0553_),
    .Y(_0556_),
    .B1(net273));
 sg13g2_nand2b_1 _1247_ (.Y(_0557_),
    .B(net162),
    .A_N(_0555_));
 sg13g2_a21oi_1 _1248_ (.A1(net239),
    .A2(net248),
    .Y(_0009_),
    .B1(_0557_));
 sg13g2_o21ai_1 _1249_ (.B1(net272),
    .Y(_0558_),
    .A1(net111),
    .A2(_0555_));
 sg13g2_a221oi_1 _1250_ (.B2(net111),
    .C1(_0558_),
    .B1(_0555_),
    .A1(net239),
    .Y(_0010_),
    .A2(net248));
 sg13g2_mux4_1 _1251_ (.S0(net280),
    .A0(\spi_own_clock_ins.data_rd[0] ),
    .A1(\spi_own_clock_ins.data_rd[1] ),
    .A2(\spi_own_clock_ins.data_rd[2] ),
    .A3(\spi_own_clock_ins.data_rd[3] ),
    .S1(\spi_own_clock_ins.index[1] ),
    .X(_0559_));
 sg13g2_nor2_1 _1252_ (.A(\spi_own_clock_ins.index[2] ),
    .B(_0559_),
    .Y(_0560_));
 sg13g2_mux2_1 _1253_ (.A0(\spi_own_clock_ins.data_rd[4] ),
    .A1(\spi_own_clock_ins.data_rd[5] ),
    .S(net280),
    .X(_0561_));
 sg13g2_nor2b_1 _1254_ (.A(\spi_own_clock_ins.data_rd[7] ),
    .B_N(net280),
    .Y(_0562_));
 sg13g2_o21ai_1 _1255_ (.B1(\spi_own_clock_ins.index[1] ),
    .Y(_0563_),
    .A1(\spi_own_clock_ins.data_rd[6] ),
    .A2(net280));
 sg13g2_o21ai_1 _1256_ (.B1(\spi_own_clock_ins.index[2] ),
    .Y(_0564_),
    .A1(_0562_),
    .A2(_0563_));
 sg13g2_a21oi_1 _1257_ (.A1(_0219_),
    .A2(_0561_),
    .Y(_0565_),
    .B1(_0564_));
 sg13g2_nor3_1 _1258_ (.A(_0023_),
    .B(_0560_),
    .C(_0565_),
    .Y(miso_clk));
 sg13g2_nand2_1 _1259_ (.Y(_0566_),
    .A(\addr_reg_sampled[1] ),
    .B(\addr_reg_sampled[0] ));
 sg13g2_nor2_1 _1260_ (.A(\addr_reg_sampled[2] ),
    .B(_0566_),
    .Y(_0567_));
 sg13g2_nor3_2 _1261_ (.A(\addr_reg_sampled[1] ),
    .B(\addr_reg_sampled[0] ),
    .C(_0021_),
    .Y(_0568_));
 sg13g2_and2_1 _1262_ (.A(\cycles_freq[6] ),
    .B(_0568_),
    .X(_0569_));
 sg13g2_nor2b_1 _1263_ (.A(\addr_reg_sampled[0] ),
    .B_N(\addr_reg_sampled[1] ),
    .Y(_0570_));
 sg13g2_and2_1 _1264_ (.A(_0224_),
    .B(_0570_),
    .X(_0571_));
 sg13g2_a221oi_1 _1265_ (.B2(uio_oe[6]),
    .C1(_0569_),
    .B1(net260),
    .A1(\cycles_high[14] ),
    .Y(_0572_),
    .A2(net261));
 sg13g2_and2_1 _1266_ (.A(_0224_),
    .B(_0424_),
    .X(_0573_));
 sg13g2_nor2_1 _1267_ (.A(\addr_reg_sampled[2] ),
    .B(_0426_),
    .Y(_0574_));
 sg13g2_a21oi_1 _1268_ (.A1(_0224_),
    .A2(_0566_),
    .Y(_0575_),
    .B1(_0574_));
 sg13g2_a21oi_1 _1269_ (.A1(\cycles_freq[14] ),
    .A2(net259),
    .Y(_0576_),
    .B1(net256));
 sg13g2_nor2b_1 _1270_ (.A(\addr_reg_sampled[2] ),
    .B_N(_0570_),
    .Y(_0577_));
 sg13g2_inv_1 _1271_ (.Y(_0578_),
    .A(_0577_));
 sg13g2_a22oi_1 _1272_ (.Y(_0579_),
    .B1(net258),
    .B2(\cycles_high[6] ),
    .A2(net262),
    .A1(\dev_regs[1][6] ));
 sg13g2_nand3_1 _1273_ (.B(_0576_),
    .C(_0579_),
    .A(_0572_),
    .Y(_0580_));
 sg13g2_and3_1 _1274_ (.X(_0581_),
    .A(\addr_reg_sampled[2] ),
    .B(\addr_reg_sampled[1] ),
    .C(\addr_reg_sampled[0] ));
 sg13g2_a21oi_1 _1275_ (.A1(_0032_),
    .A2(net256),
    .Y(_0582_),
    .B1(net271));
 sg13g2_a221oi_1 _1276_ (.B2(_0580_),
    .C1(\spi_sampled_ins.index[0] ),
    .B1(_0582_),
    .A1(net14),
    .Y(_0583_),
    .A2(net269));
 sg13g2_and2_1 _1277_ (.A(\cycles_freq[15] ),
    .B(net259),
    .X(_0584_));
 sg13g2_a221oi_1 _1278_ (.B2(uio_oe[7]),
    .C1(_0584_),
    .B1(net260),
    .A1(\cycles_high[15] ),
    .Y(_0585_),
    .A2(net261));
 sg13g2_a21oi_1 _1279_ (.A1(\dev_regs[1][7] ),
    .A2(net262),
    .Y(_0586_),
    .B1(net256));
 sg13g2_a22oi_1 _1280_ (.Y(_0587_),
    .B1(net258),
    .B2(\cycles_high[7] ),
    .A2(_0568_),
    .A1(\cycles_freq[7] ));
 sg13g2_nand3_1 _1281_ (.B(_0586_),
    .C(_0587_),
    .A(_0585_),
    .Y(_0588_));
 sg13g2_a21oi_1 _1282_ (.A1(_0248_),
    .A2(_0575_),
    .Y(_0589_),
    .B1(net269));
 sg13g2_a221oi_1 _1283_ (.B2(_0589_),
    .C1(_0215_),
    .B1(_0588_),
    .A1(net15),
    .Y(_0590_),
    .A2(net269));
 sg13g2_o21ai_1 _1284_ (.B1(\spi_sampled_ins.index[1] ),
    .Y(_0591_),
    .A1(_0583_),
    .A2(_0590_));
 sg13g2_nand2_1 _1285_ (.Y(_0592_),
    .A(uio_oe[5]),
    .B(net260));
 sg13g2_a22oi_1 _1286_ (.Y(_0593_),
    .B1(_0568_),
    .B2(\cycles_freq[5] ),
    .A2(net261),
    .A1(\cycles_high[13] ));
 sg13g2_a22oi_1 _1287_ (.Y(_0594_),
    .B1(net258),
    .B2(\cycles_high[5] ),
    .A2(net262),
    .A1(\dev_regs[1][5] ));
 sg13g2_a21oi_1 _1288_ (.A1(\cycles_freq[13] ),
    .A2(net259),
    .Y(_0595_),
    .B1(net256));
 sg13g2_nand4_1 _1289_ (.B(_0593_),
    .C(_0594_),
    .A(_0592_),
    .Y(_0596_),
    .D(_0595_));
 sg13g2_a21oi_1 _1290_ (.A1(_0031_),
    .A2(net255),
    .Y(_0597_),
    .B1(net271));
 sg13g2_nand2b_1 _1291_ (.Y(_0598_),
    .B(\spi_sampled_ins.index[0] ),
    .A_N(\spi_sampled_ins.index[1] ));
 sg13g2_a221oi_1 _1292_ (.B2(_0597_),
    .C1(_0598_),
    .B1(_0596_),
    .A1(net13),
    .Y(_0599_),
    .A2(net269));
 sg13g2_and2_1 _1293_ (.A(\cycles_freq[4] ),
    .B(_0568_),
    .X(_0600_));
 sg13g2_a221oi_1 _1294_ (.B2(\cycles_high[4] ),
    .C1(_0600_),
    .B1(net258),
    .A1(uio_oe[4]),
    .Y(_0601_),
    .A2(net260));
 sg13g2_a21oi_1 _1295_ (.A1(\cycles_freq[12] ),
    .A2(net259),
    .Y(_0602_),
    .B1(net256));
 sg13g2_a22oi_1 _1296_ (.Y(_0603_),
    .B1(net261),
    .B2(\cycles_high[12] ),
    .A2(net262),
    .A1(\dev_regs[1][4] ));
 sg13g2_nand3_1 _1297_ (.B(_0602_),
    .C(_0603_),
    .A(_0601_),
    .Y(_0604_));
 sg13g2_a21oi_1 _1298_ (.A1(_0247_),
    .A2(net255),
    .Y(_0605_),
    .B1(net271));
 sg13g2_a221oi_1 _1299_ (.B2(_0605_),
    .C1(_0254_),
    .B1(_0604_),
    .A1(net12),
    .Y(_0606_),
    .A2(net270));
 sg13g2_nor2_1 _1300_ (.A(_0599_),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_a21oi_1 _1301_ (.A1(_0591_),
    .A2(_0607_),
    .Y(_0608_),
    .B1(_0213_));
 sg13g2_a22oi_1 _1302_ (.Y(_0609_),
    .B1(net260),
    .B2(uio_oe[3]),
    .A2(_0567_),
    .A1(\cycles_high[11] ));
 sg13g2_a221oi_1 _1303_ (.B2(\cycles_freq[11] ),
    .C1(net255),
    .B1(_0573_),
    .A1(\dev_regs[1][3] ),
    .Y(_0610_),
    .A2(net262));
 sg13g2_a22oi_1 _1304_ (.Y(_0611_),
    .B1(net258),
    .B2(\cycles_high[3] ),
    .A2(_0568_),
    .A1(\cycles_freq[3] ));
 sg13g2_nand3_1 _1305_ (.B(_0610_),
    .C(_0611_),
    .A(_0609_),
    .Y(_0612_));
 sg13g2_a21oi_1 _1306_ (.A1(_0030_),
    .A2(net255),
    .Y(_0613_),
    .B1(net269));
 sg13g2_a221oi_1 _1307_ (.B2(_0613_),
    .C1(_0215_),
    .B1(_0612_),
    .A1(net11),
    .Y(_0614_),
    .A2(net270));
 sg13g2_a221oi_1 _1308_ (.B2(\cycles_freq[10] ),
    .C1(net255),
    .B1(net259),
    .A1(\cycles_freq[2] ),
    .Y(_0615_),
    .A2(_0568_));
 sg13g2_a22oi_1 _1309_ (.Y(_0616_),
    .B1(_0571_),
    .B2(uio_oe[2]),
    .A2(_0425_),
    .A1(\dev_regs[1][2] ));
 sg13g2_a22oi_1 _1310_ (.Y(_0617_),
    .B1(net258),
    .B2(\cycles_high[2] ),
    .A2(net261),
    .A1(\cycles_high[10] ));
 sg13g2_nand3_1 _1311_ (.B(_0616_),
    .C(_0617_),
    .A(_0615_),
    .Y(_0618_));
 sg13g2_a21oi_1 _1312_ (.A1(_0246_),
    .A2(net255),
    .Y(_0619_),
    .B1(net269));
 sg13g2_a221oi_1 _1313_ (.B2(_0619_),
    .C1(\spi_sampled_ins.index[0] ),
    .B1(_0618_),
    .A1(net10),
    .Y(_0620_),
    .A2(net270));
 sg13g2_o21ai_1 _1314_ (.B1(\spi_sampled_ins.index[1] ),
    .Y(_0621_),
    .A1(_0614_),
    .A2(_0620_));
 sg13g2_and2_1 _1315_ (.A(\cycles_freq[0] ),
    .B(_0568_),
    .X(_0622_));
 sg13g2_a22oi_1 _1316_ (.Y(_0623_),
    .B1(net259),
    .B2(\cycles_freq[8] ),
    .A2(net262),
    .A1(\dev_regs[1][0] ));
 sg13g2_a21oi_1 _1317_ (.A1(uio_oe[0]),
    .A2(net260),
    .Y(_0624_),
    .B1(net256));
 sg13g2_a221oi_1 _1318_ (.B2(\cycles_high[0] ),
    .C1(_0622_),
    .B1(net258),
    .A1(\cycles_high[8] ),
    .Y(_0625_),
    .A2(net261));
 sg13g2_nand3_1 _1319_ (.B(_0624_),
    .C(_0625_),
    .A(_0623_),
    .Y(_0626_));
 sg13g2_a21oi_1 _1320_ (.A1(_0029_),
    .A2(net255),
    .Y(_0627_),
    .B1(net269));
 sg13g2_a221oi_1 _1321_ (.B2(_0627_),
    .C1(_0254_),
    .B1(_0626_),
    .A1(net8),
    .Y(_0628_),
    .A2(net270));
 sg13g2_nand2_1 _1322_ (.Y(_0629_),
    .A(uio_oe[1]),
    .B(net260));
 sg13g2_a22oi_1 _1323_ (.Y(_0630_),
    .B1(net259),
    .B2(\cycles_freq[9] ),
    .A2(net261),
    .A1(\cycles_high[9] ));
 sg13g2_a22oi_1 _1324_ (.Y(_0631_),
    .B1(net258),
    .B2(\cycles_high[1] ),
    .A2(net262),
    .A1(\dev_regs[1][1] ));
 sg13g2_a21oi_1 _1325_ (.A1(\cycles_freq[1] ),
    .A2(_0568_),
    .Y(_0632_),
    .B1(net256));
 sg13g2_nand4_1 _1326_ (.B(_0630_),
    .C(_0631_),
    .A(_0629_),
    .Y(_0633_),
    .D(_0632_));
 sg13g2_a21oi_1 _1327_ (.A1(_0245_),
    .A2(net255),
    .Y(_0634_),
    .B1(net271));
 sg13g2_a221oi_1 _1328_ (.B2(_0634_),
    .C1(_0598_),
    .B1(_0633_),
    .A1(net9),
    .Y(_0635_),
    .A2(net269));
 sg13g2_nor2_1 _1329_ (.A(_0628_),
    .B(_0635_),
    .Y(_0636_));
 sg13g2_a21oi_1 _1330_ (.A1(_0621_),
    .A2(_0636_),
    .Y(_0637_),
    .B1(\spi_sampled_ins.index[2] ));
 sg13g2_nor3_1 _1331_ (.A(_0250_),
    .B(_0608_),
    .C(_0637_),
    .Y(miso_sampled));
 sg13g2_nor3_1 _1332_ (.A(_0306_),
    .B(_0309_),
    .C(net273),
    .Y(_0638_));
 sg13g2_nor2b_2 _1333_ (.A(_0638_),
    .B_N(net251),
    .Y(_0639_));
 sg13g2_inv_1 _1334_ (.Y(_0640_),
    .A(_0639_));
 sg13g2_nand2_2 _1335_ (.Y(_0641_),
    .A(net311),
    .B(_0639_));
 sg13g2_mux2_1 _1336_ (.A0(\spi_own_clock_ins.spi_data_reg[0] ),
    .A1(net98),
    .S(_0641_),
    .X(_0101_));
 sg13g2_mux2_1 _1337_ (.A0(\spi_own_clock_ins.spi_data_reg[1] ),
    .A1(net109),
    .S(_0641_),
    .X(_0102_));
 sg13g2_mux2_1 _1338_ (.A0(\spi_own_clock_ins.spi_data_reg[2] ),
    .A1(net95),
    .S(_0641_),
    .X(_0103_));
 sg13g2_mux2_1 _1339_ (.A0(\spi_own_clock_ins.spi_data_reg[3] ),
    .A1(net104),
    .S(_0641_),
    .X(_0104_));
 sg13g2_mux2_1 _1340_ (.A0(\spi_own_clock_ins.spi_data_reg[4] ),
    .A1(net118),
    .S(_0641_),
    .X(_0105_));
 sg13g2_mux2_1 _1341_ (.A0(\spi_own_clock_ins.spi_data_reg[5] ),
    .A1(net110),
    .S(_0641_),
    .X(_0106_));
 sg13g2_mux2_1 _1342_ (.A0(\spi_own_clock_ins.spi_data_reg[6] ),
    .A1(net114),
    .S(_0641_),
    .X(_0107_));
 sg13g2_mux2_1 _1343_ (.A0(\spi_own_clock_ins.spi_data_reg[7] ),
    .A1(net151),
    .S(_0641_),
    .X(_0108_));
 sg13g2_nand2_1 _1344_ (.Y(_0642_),
    .A(\data_wr_z1[0] ),
    .B(net252));
 sg13g2_nand2_1 _1345_ (.Y(_0643_),
    .A(\spi_sampled_ins.spi_data_reg[0] ),
    .B(net257));
 sg13g2_o21ai_1 _1346_ (.B1(_0642_),
    .Y(_0644_),
    .A1(net253),
    .A2(_0643_));
 sg13g2_inv_2 _1347_ (.Y(_0645_),
    .A(_0644_));
 sg13g2_nand2_1 _1348_ (.Y(_0646_),
    .A(net117),
    .B(net250));
 sg13g2_o21ai_1 _1349_ (.B1(_0646_),
    .Y(_0125_),
    .A1(net250),
    .A2(_0645_));
 sg13g2_nand2_1 _1350_ (.Y(_0647_),
    .A(\data_wr_z1[1] ),
    .B(net252));
 sg13g2_nand2_1 _1351_ (.Y(_0648_),
    .A(\spi_sampled_ins.spi_data_reg[1] ),
    .B(net257));
 sg13g2_o21ai_1 _1352_ (.B1(_0647_),
    .Y(_0649_),
    .A1(net253),
    .A2(_0648_));
 sg13g2_inv_2 _1353_ (.Y(_0650_),
    .A(_0649_));
 sg13g2_nand2_1 _1354_ (.Y(_0651_),
    .A(net70),
    .B(net250));
 sg13g2_o21ai_1 _1355_ (.B1(_0651_),
    .Y(_0126_),
    .A1(net250),
    .A2(_0650_));
 sg13g2_nand2_1 _1356_ (.Y(_0652_),
    .A(\data_wr_z1[2] ),
    .B(net251));
 sg13g2_nand2_1 _1357_ (.Y(_0653_),
    .A(\spi_sampled_ins.spi_data_reg[2] ),
    .B(net257));
 sg13g2_o21ai_1 _1358_ (.B1(_0652_),
    .Y(_0654_),
    .A1(net251),
    .A2(_0653_));
 sg13g2_mux2_1 _1359_ (.A0(_0654_),
    .A1(net103),
    .S(_0430_),
    .X(_0127_));
 sg13g2_nand2_1 _1360_ (.Y(_0655_),
    .A(\data_wr_z1[3] ),
    .B(net252));
 sg13g2_nand2_1 _1361_ (.Y(_0656_),
    .A(\spi_sampled_ins.spi_data_reg[3] ),
    .B(net257));
 sg13g2_o21ai_1 _1362_ (.B1(_0655_),
    .Y(_0657_),
    .A1(net252),
    .A2(_0656_));
 sg13g2_mux2_1 _1363_ (.A0(_0657_),
    .A1(net90),
    .S(_0430_),
    .X(_0128_));
 sg13g2_nand2_1 _1364_ (.Y(_0658_),
    .A(\data_wr_z1[4] ),
    .B(net253));
 sg13g2_nand2_1 _1365_ (.Y(_0659_),
    .A(\spi_sampled_ins.spi_data_reg[4] ),
    .B(_0427_));
 sg13g2_o21ai_1 _1366_ (.B1(_0658_),
    .Y(_0660_),
    .A1(net252),
    .A2(_0659_));
 sg13g2_mux2_1 _1367_ (.A0(_0660_),
    .A1(net97),
    .S(net250),
    .X(_0129_));
 sg13g2_nand2_1 _1368_ (.Y(_0661_),
    .A(\data_wr_z1[5] ),
    .B(net253));
 sg13g2_nand2_1 _1369_ (.Y(_0662_),
    .A(\spi_sampled_ins.spi_data_reg[5] ),
    .B(net257));
 sg13g2_o21ai_1 _1370_ (.B1(_0661_),
    .Y(_0663_),
    .A1(net252),
    .A2(_0662_));
 sg13g2_mux2_1 _1371_ (.A0(_0663_),
    .A1(net96),
    .S(net250),
    .X(_0130_));
 sg13g2_nand2_1 _1372_ (.Y(_0664_),
    .A(\data_wr_z1[6] ),
    .B(net252));
 sg13g2_nand2_1 _1373_ (.Y(_0665_),
    .A(\spi_sampled_ins.spi_data_reg[6] ),
    .B(net257));
 sg13g2_o21ai_1 _1374_ (.B1(_0664_),
    .Y(_0666_),
    .A1(net252),
    .A2(_0665_));
 sg13g2_mux2_1 _1375_ (.A0(_0666_),
    .A1(net100),
    .S(net250),
    .X(_0131_));
 sg13g2_a22oi_1 _1376_ (.Y(_0667_),
    .B1(_0639_),
    .B2(_0314_),
    .A2(_0578_),
    .A1(_0429_));
 sg13g2_nor2_1 _1377_ (.A(_0429_),
    .B(_0639_),
    .Y(_0668_));
 sg13g2_a21oi_1 _1378_ (.A1(\addr_reg_sampled[2] ),
    .A2(\addr_reg_sampled[1] ),
    .Y(_0669_),
    .B1(net273));
 sg13g2_nand2b_1 _1379_ (.Y(_0670_),
    .B(_0669_),
    .A_N(_0425_));
 sg13g2_a21o_1 _1380_ (.A2(_0670_),
    .A1(_0429_),
    .B1(_0639_),
    .X(_0671_));
 sg13g2_nand2_1 _1381_ (.Y(_0672_),
    .A(_0667_),
    .B(_0671_));
 sg13g2_nand2_1 _1382_ (.Y(_0673_),
    .A(net84),
    .B(net247));
 sg13g2_o21ai_1 _1383_ (.B1(_0673_),
    .Y(_0132_),
    .A1(_0645_),
    .A2(net246));
 sg13g2_nand2_1 _1384_ (.Y(_0674_),
    .A(net107),
    .B(net247));
 sg13g2_o21ai_1 _1385_ (.B1(_0674_),
    .Y(_0133_),
    .A1(_0650_),
    .A2(net247));
 sg13g2_nand2_1 _1386_ (.Y(_0675_),
    .A(net52),
    .B(net247));
 sg13g2_o21ai_1 _1387_ (.B1(_0675_),
    .Y(_0134_),
    .A1(_0654_),
    .A2(net247));
 sg13g2_mux2_1 _1388_ (.A0(_0657_),
    .A1(net139),
    .S(net247),
    .X(_0135_));
 sg13g2_nand2_1 _1389_ (.Y(_0676_),
    .A(net44),
    .B(net246));
 sg13g2_o21ai_1 _1390_ (.B1(_0676_),
    .Y(_0136_),
    .A1(_0660_),
    .A2(net246));
 sg13g2_mux2_1 _1391_ (.A0(_0663_),
    .A1(net136),
    .S(net246),
    .X(_0137_));
 sg13g2_nor2_1 _1392_ (.A(_0666_),
    .B(net246),
    .Y(_0677_));
 sg13g2_a21oi_1 _1393_ (.A1(_0244_),
    .A2(net246),
    .Y(_0138_),
    .B1(_0677_));
 sg13g2_nor2_1 _1394_ (.A(net251),
    .B(_0431_),
    .Y(_0678_));
 sg13g2_a21oi_2 _1395_ (.B1(_0678_),
    .Y(_0679_),
    .A2(net254),
    .A1(\data_wr_z1[7] ));
 sg13g2_a21o_1 _1396_ (.A2(net254),
    .A1(\data_wr_z1[7] ),
    .B1(_0678_),
    .X(_0680_));
 sg13g2_nand2_1 _1397_ (.Y(_0681_),
    .A(net105),
    .B(net246));
 sg13g2_o21ai_1 _1398_ (.B1(_0681_),
    .Y(_0139_),
    .A1(net246),
    .A2(_0679_));
 sg13g2_nand2_1 _1399_ (.Y(_0682_),
    .A(net273),
    .B(net261));
 sg13g2_a21oi_1 _1400_ (.A1(_0429_),
    .A2(_0682_),
    .Y(_0683_),
    .B1(_0667_));
 sg13g2_o21ai_1 _1401_ (.B1(_0683_),
    .Y(_0684_),
    .A1(net264),
    .A2(_0640_));
 sg13g2_mux2_1 _1402_ (.A0(_0644_),
    .A1(net148),
    .S(_0684_),
    .X(_0140_));
 sg13g2_mux2_1 _1403_ (.A0(_0650_),
    .A1(net66),
    .S(_0684_),
    .X(_0141_));
 sg13g2_mux2_1 _1404_ (.A0(_0654_),
    .A1(net135),
    .S(_0684_),
    .X(_0142_));
 sg13g2_mux2_1 _1405_ (.A0(_0657_),
    .A1(net147),
    .S(_0684_),
    .X(_0143_));
 sg13g2_mux2_1 _1406_ (.A0(_0660_),
    .A1(net140),
    .S(_0684_),
    .X(_0144_));
 sg13g2_mux2_1 _1407_ (.A0(_0663_),
    .A1(net124),
    .S(_0684_),
    .X(_0145_));
 sg13g2_mux2_1 _1408_ (.A0(_0666_),
    .A1(net132),
    .S(_0684_),
    .X(_0146_));
 sg13g2_mux2_1 _1409_ (.A0(_0679_),
    .A1(net62),
    .S(_0684_),
    .X(_0147_));
 sg13g2_or2_1 _1410_ (.X(_0685_),
    .B(_0428_),
    .A(_0426_));
 sg13g2_nand2b_1 _1411_ (.Y(_0686_),
    .B(_0639_),
    .A_N(net274));
 sg13g2_nand3_1 _1412_ (.B(_0685_),
    .C(_0686_),
    .A(_0671_),
    .Y(_0687_));
 sg13g2_nand2_1 _1413_ (.Y(_0688_),
    .A(net78),
    .B(net245));
 sg13g2_o21ai_1 _1414_ (.B1(_0688_),
    .Y(_0148_),
    .A1(_0645_),
    .A2(net245));
 sg13g2_nand2_1 _1415_ (.Y(_0689_),
    .A(net99),
    .B(net245));
 sg13g2_o21ai_1 _1416_ (.B1(_0689_),
    .Y(_0149_),
    .A1(_0650_),
    .A2(net244));
 sg13g2_mux2_1 _1417_ (.A0(_0654_),
    .A1(net142),
    .S(net245),
    .X(_0150_));
 sg13g2_mux2_1 _1418_ (.A0(_0657_),
    .A1(net146),
    .S(net245),
    .X(_0151_));
 sg13g2_nand2_1 _1419_ (.Y(_0690_),
    .A(net46),
    .B(net244));
 sg13g2_o21ai_1 _1420_ (.B1(_0690_),
    .Y(_0152_),
    .A1(_0660_),
    .A2(net244));
 sg13g2_mux2_1 _1421_ (.A0(_0663_),
    .A1(net108),
    .S(net244),
    .X(_0153_));
 sg13g2_nand2_1 _1422_ (.Y(_0691_),
    .A(net45),
    .B(net244));
 sg13g2_o21ai_1 _1423_ (.B1(_0691_),
    .Y(_0154_),
    .A1(_0666_),
    .A2(net244));
 sg13g2_nand2_1 _1424_ (.Y(_0692_),
    .A(net93),
    .B(net244));
 sg13g2_o21ai_1 _1425_ (.B1(_0692_),
    .Y(_0155_),
    .A1(_0679_),
    .A2(net244));
 sg13g2_nand2b_1 _1426_ (.Y(_0693_),
    .B(_0639_),
    .A_N(net265));
 sg13g2_nand2b_1 _1427_ (.Y(_0694_),
    .B(_0429_),
    .A_N(net259));
 sg13g2_nand3_1 _1428_ (.B(_0693_),
    .C(_0694_),
    .A(_0671_),
    .Y(_0695_));
 sg13g2_mux2_1 _1429_ (.A0(_0645_),
    .A1(net65),
    .S(net243),
    .X(_0156_));
 sg13g2_nand2_1 _1430_ (.Y(_0696_),
    .A(net47),
    .B(net242));
 sg13g2_o21ai_1 _1431_ (.B1(_0696_),
    .Y(_0157_),
    .A1(_0649_),
    .A2(net242));
 sg13g2_mux2_1 _1432_ (.A0(_0654_),
    .A1(net138),
    .S(net243),
    .X(_0158_));
 sg13g2_mux2_1 _1433_ (.A0(_0657_),
    .A1(net152),
    .S(net243),
    .X(_0159_));
 sg13g2_mux2_1 _1434_ (.A0(_0660_),
    .A1(net133),
    .S(net242),
    .X(_0160_));
 sg13g2_mux2_1 _1435_ (.A0(_0663_),
    .A1(net134),
    .S(net242),
    .X(_0161_));
 sg13g2_nand2_1 _1436_ (.Y(_0697_),
    .A(net51),
    .B(net242));
 sg13g2_o21ai_1 _1437_ (.B1(_0697_),
    .Y(_0162_),
    .A1(_0666_),
    .A2(net242));
 sg13g2_nand2_1 _1438_ (.Y(_0698_),
    .A(net48),
    .B(net242));
 sg13g2_o21ai_1 _1439_ (.B1(_0698_),
    .Y(_0163_),
    .A1(_0680_),
    .A2(net242));
 sg13g2_o21ai_1 _1440_ (.B1(_0671_),
    .Y(_0699_),
    .A1(net251),
    .A2(net260));
 sg13g2_a21oi_2 _1441_ (.B1(_0699_),
    .Y(_0700_),
    .A2(_0639_),
    .A1(_0308_));
 sg13g2_mux2_1 _1442_ (.A0(net120),
    .A1(_0644_),
    .S(_0700_),
    .X(_0164_));
 sg13g2_mux2_1 _1443_ (.A0(net123),
    .A1(_0649_),
    .S(_0700_),
    .X(_0165_));
 sg13g2_mux2_1 _1444_ (.A0(net137),
    .A1(_0654_),
    .S(_0700_),
    .X(_0166_));
 sg13g2_mux2_1 _1445_ (.A0(net145),
    .A1(_0657_),
    .S(_0700_),
    .X(_0167_));
 sg13g2_mux2_1 _1446_ (.A0(net127),
    .A1(_0660_),
    .S(_0700_),
    .X(_0168_));
 sg13g2_mux2_1 _1447_ (.A0(net121),
    .A1(_0663_),
    .S(_0700_),
    .X(_0169_));
 sg13g2_mux2_1 _1448_ (.A0(net141),
    .A1(_0666_),
    .S(_0700_),
    .X(_0170_));
 sg13g2_mux2_1 _1449_ (.A0(net119),
    .A1(_0680_),
    .S(_0700_),
    .X(_0171_));
 sg13g2_nor2b_1 _1450_ (.A(net289),
    .B_N(net310),
    .Y(_0049_));
 sg13g2_nand2_1 _1451_ (.Y(_0701_),
    .A(net275),
    .B(net251));
 sg13g2_o21ai_1 _1452_ (.B1(_0701_),
    .Y(_0702_),
    .A1(net251),
    .A2(net271));
 sg13g2_nor2_2 _1453_ (.A(_0668_),
    .B(_0702_),
    .Y(_0703_));
 sg13g2_nor2_1 _1454_ (.A(net83),
    .B(_0703_),
    .Y(_0704_));
 sg13g2_a21oi_1 _1455_ (.A1(_0645_),
    .A2(_0703_),
    .Y(_0172_),
    .B1(_0704_));
 sg13g2_nor2_1 _1456_ (.A(net86),
    .B(_0703_),
    .Y(_0705_));
 sg13g2_a21oi_1 _1457_ (.A1(_0650_),
    .A2(net241),
    .Y(_0173_),
    .B1(_0705_));
 sg13g2_mux2_1 _1458_ (.A0(net73),
    .A1(_0654_),
    .S(net241),
    .X(_0174_));
 sg13g2_mux2_1 _1459_ (.A0(net69),
    .A1(_0657_),
    .S(net241),
    .X(_0175_));
 sg13g2_mux2_1 _1460_ (.A0(net82),
    .A1(_0660_),
    .S(net241),
    .X(_0176_));
 sg13g2_mux2_1 _1461_ (.A0(net92),
    .A1(_0663_),
    .S(net241),
    .X(_0177_));
 sg13g2_mux2_1 _1462_ (.A0(net91),
    .A1(_0666_),
    .S(net241),
    .X(_0178_));
 sg13g2_nor2_1 _1463_ (.A(net87),
    .B(net241),
    .Y(_0706_));
 sg13g2_a21oi_1 _1464_ (.A1(_0679_),
    .A2(net241),
    .Y(_0179_),
    .B1(_0706_));
 sg13g2_nand2_1 _1465_ (.Y(_0707_),
    .A(net57),
    .B(net249));
 sg13g2_a21oi_1 _1466_ (.A1(net240),
    .A2(_0707_),
    .Y(_0187_),
    .B1(_0521_));
 sg13g2_nor2b_1 _1467_ (.A(net279),
    .B_N(net314),
    .Y(_0084_));
 sg13g2_inv_1 _1468_ (.Y(_0080_),
    .A(net285));
 sg13g2_inv_1 _1469_ (.Y(_0078_),
    .A(net285));
 sg13g2_inv_1 _1470_ (.Y(_0076_),
    .A(net285));
 sg13g2_inv_1 _1471_ (.Y(_0074_),
    .A(net285));
 sg13g2_inv_1 _1472_ (.Y(_0072_),
    .A(net285));
 sg13g2_inv_1 _1473_ (.Y(_0070_),
    .A(net285));
 sg13g2_inv_1 _1474_ (.Y(_0068_),
    .A(net288));
 sg13g2_buf_1 _1475_ (.A(net50),
    .X(_0117_));
 sg13g2_buf_1 _1476_ (.A(net40),
    .X(_0118_));
 sg13g2_buf_1 _1477_ (.A(net41),
    .X(_0119_));
 sg13g2_buf_1 _1478_ (.A(net43),
    .X(_0120_));
 sg13g2_buf_1 _1479_ (.A(net42),
    .X(_0121_));
 sg13g2_buf_1 _1480_ (.A(net53),
    .X(_0122_));
 sg13g2_buf_1 _1481_ (.A(net54),
    .X(_0123_));
 sg13g2_buf_1 _1482_ (.A(net39),
    .X(_0124_));
 sg13g2_nor2b_1 _1483_ (.A(net287),
    .B_N(net308),
    .Y(_0050_));
 sg13g2_nor2b_1 _1484_ (.A(net287),
    .B_N(net308),
    .Y(_0051_));
 sg13g2_nor2b_1 _1485_ (.A(net287),
    .B_N(net308),
    .Y(_0052_));
 sg13g2_nor2b_1 _1486_ (.A(net287),
    .B_N(net308),
    .Y(_0053_));
 sg13g2_nor2b_1 _1487_ (.A(net287),
    .B_N(net308),
    .Y(_0054_));
 sg13g2_nor2b_1 _1488_ (.A(net289),
    .B_N(net308),
    .Y(_0055_));
 sg13g2_nor2b_1 _1489_ (.A(net289),
    .B_N(net308),
    .Y(_0056_));
 sg13g2_nor2b_1 _1490_ (.A(net286),
    .B_N(net311),
    .Y(_0057_));
 sg13g2_nor2b_1 _1491_ (.A(net286),
    .B_N(net311),
    .Y(_0058_));
 sg13g2_nor2b_1 _1492_ (.A(net285),
    .B_N(net311),
    .Y(_0059_));
 sg13g2_nor2b_1 _1493_ (.A(net289),
    .B_N(net309),
    .Y(_0060_));
 sg13g2_nor2b_1 _1494_ (.A(net289),
    .B_N(net310),
    .Y(_0061_));
 sg13g2_nor2b_1 _1495_ (.A(net288),
    .B_N(net309),
    .Y(_0062_));
 sg13g2_nor2b_1 _1496_ (.A(net288),
    .B_N(net309),
    .Y(_0063_));
 sg13g2_nor2b_1 _1497_ (.A(net287),
    .B_N(net309),
    .Y(_0064_));
 sg13g2_nor2b_1 _1498_ (.A(net287),
    .B_N(net309),
    .Y(_0065_));
 sg13g2_nor2b_1 _1499_ (.A(net287),
    .B_N(net308),
    .Y(_0066_));
 sg13g2_nor2b_1 _1500_ (.A(net288),
    .B_N(net309),
    .Y(_0067_));
 sg13g2_inv_1 _1501_ (.Y(_0071_),
    .A(net290));
 sg13g2_inv_1 _1502_ (.Y(_0073_),
    .A(net290));
 sg13g2_inv_1 _1503_ (.Y(_0075_),
    .A(net290));
 sg13g2_inv_1 _1504_ (.Y(_0077_),
    .A(net290));
 sg13g2_inv_1 _1505_ (.Y(_0079_),
    .A(net290));
 sg13g2_inv_1 _1506_ (.Y(_0081_),
    .A(net290));
 sg13g2_inv_1 _1507_ (.Y(_0083_),
    .A(net290));
 sg13g2_nor2b_1 _1508_ (.A(net279),
    .B_N(net314),
    .Y(_0085_));
 sg13g2_nor2b_1 _1509_ (.A(net279),
    .B_N(net312),
    .Y(_0086_));
 sg13g2_nor2b_1 _1510_ (.A(net288),
    .B_N(net314),
    .Y(_0087_));
 sg13g2_nor2b_1 _1511_ (.A(net288),
    .B_N(net314),
    .Y(_0088_));
 sg13g2_nor2b_1 _1512_ (.A(net288),
    .B_N(net309),
    .Y(_0089_));
 sg13g2_nor2b_1 _1513_ (.A(net288),
    .B_N(net309),
    .Y(_0090_));
 sg13g2_nor2b_1 _1514_ (.A(net286),
    .B_N(net311),
    .Y(_0091_));
 sg13g2_nor2b_1 _1515_ (.A(net286),
    .B_N(net311),
    .Y(_0092_));
 sg13g2_nor2b_1 _1516_ (.A(net286),
    .B_N(net311),
    .Y(_0093_));
 sg13g2_nor2b_1 _1517_ (.A(net286),
    .B_N(net312),
    .Y(_0094_));
 sg13g2_nor2b_1 _1518_ (.A(net122),
    .B_N(net315),
    .Y(_0095_));
 sg13g2_nor2b_1 _1519_ (.A(net279),
    .B_N(net314),
    .Y(_0096_));
 sg13g2_nor2b_1 _1520_ (.A(net279),
    .B_N(net314),
    .Y(_0097_));
 sg13g2_nor2b_1 _1521_ (.A(net279),
    .B_N(net312),
    .Y(_0098_));
 sg13g2_nor2b_1 _1522_ (.A(net279),
    .B_N(net313),
    .Y(_0099_));
 sg13g2_nor2b_1 _1523_ (.A(net279),
    .B_N(net314),
    .Y(_0100_));
 sg13g2_dfrbp_1 _1524_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net28),
    .D(_0101_),
    .Q_N(_0804_),
    .Q(\data_wr_z1[0] ));
 sg13g2_dfrbp_1 _1525_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net27),
    .D(_0102_),
    .Q_N(_0803_),
    .Q(\data_wr_z1[1] ));
 sg13g2_dfrbp_1 _1526_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net26),
    .D(_0103_),
    .Q_N(_0802_),
    .Q(\data_wr_z1[2] ));
 sg13g2_dfrbp_1 _1527_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net25),
    .D(_0104_),
    .Q_N(_0801_),
    .Q(\data_wr_z1[3] ));
 sg13g2_dfrbp_1 _1528_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net24),
    .D(_0105_),
    .Q_N(_0800_),
    .Q(\data_wr_z1[4] ));
 sg13g2_dfrbp_1 _1529_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net23),
    .D(_0106_),
    .Q_N(_0799_),
    .Q(\data_wr_z1[5] ));
 sg13g2_dfrbp_1 _1530_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net22),
    .D(_0107_),
    .Q_N(_0798_),
    .Q(\data_wr_z1[6] ));
 sg13g2_dfrbp_1 _1531_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net21),
    .D(_0108_),
    .Q_N(_0797_),
    .Q(\data_wr_z1[7] ));
 sg13g2_dfrbp_1 _1532_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net171),
    .D(net68),
    .Q_N(_0796_),
    .Q(\spi_sampled_ins.spi_data_reg[0] ));
 sg13g2_dfrbp_1 _1533_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net171),
    .D(_0110_),
    .Q_N(_0795_),
    .Q(\spi_sampled_ins.spi_data_reg[1] ));
 sg13g2_dfrbp_1 _1534_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net171),
    .D(_0111_),
    .Q_N(_0794_),
    .Q(\spi_sampled_ins.spi_data_reg[2] ));
 sg13g2_dfrbp_1 _1535_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net171),
    .D(_0112_),
    .Q_N(_0793_),
    .Q(\spi_sampled_ins.spi_data_reg[3] ));
 sg13g2_dfrbp_1 _1536_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net171),
    .D(net80),
    .Q_N(_0792_),
    .Q(\spi_sampled_ins.spi_data_reg[4] ));
 sg13g2_dfrbp_1 _1537_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net171),
    .D(_0114_),
    .Q_N(_0791_),
    .Q(\spi_sampled_ins.spi_data_reg[5] ));
 sg13g2_dfrbp_1 _1538_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net171),
    .D(_0115_),
    .Q_N(_0790_),
    .Q(\spi_sampled_ins.spi_data_reg[6] ));
 sg13g2_dfrbp_1 _1539_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net171),
    .D(net61),
    .Q_N(_0024_),
    .Q(\spi_sampled_ins.spi_data_reg[7] ));
 sg13g2_dfrbp_1 _1540_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net312),
    .D(_0117_),
    .Q_N(_0029_),
    .Q(\dev_regs[0][0] ));
 sg13g2_dfrbp_1 _1541_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net305),
    .D(_0118_),
    .Q_N(\dev_regs[0][1] ),
    .Q(_0033_));
 sg13g2_dfrbp_1 _1542_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net313),
    .D(_0119_),
    .Q_N(\dev_regs[0][2] ),
    .Q(_0034_));
 sg13g2_dfrbp_1 _1543_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net312),
    .D(_0120_),
    .Q_N(_0030_),
    .Q(\dev_regs[0][3] ));
 sg13g2_dfrbp_1 _1544_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net305),
    .D(_0121_),
    .Q_N(\dev_regs[0][4] ),
    .Q(_0035_));
 sg13g2_dfrbp_1 _1545_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net313),
    .D(_0122_),
    .Q_N(_0031_),
    .Q(\dev_regs[0][5] ));
 sg13g2_dfrbp_1 _1546_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net313),
    .D(_0123_),
    .Q_N(_0032_),
    .Q(\dev_regs[0][6] ));
 sg13g2_dfrbp_1 _1547_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net312),
    .D(_0124_),
    .Q_N(\dev_regs[0][7] ),
    .Q(_0036_));
 sg13g2_dfrbp_1 _1548_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net304),
    .D(_0125_),
    .Q_N(_0789_),
    .Q(\dev_regs[1][0] ));
 sg13g2_dfrbp_1 _1549_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net304),
    .D(_0126_),
    .Q_N(_0788_),
    .Q(\dev_regs[1][1] ));
 sg13g2_dfrbp_1 _1550_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net305),
    .D(_0127_),
    .Q_N(_0787_),
    .Q(\dev_regs[1][2] ));
 sg13g2_dfrbp_1 _1551_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net312),
    .D(_0128_),
    .Q_N(_0786_),
    .Q(\dev_regs[1][3] ));
 sg13g2_dfrbp_1 _1552_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net304),
    .D(_0129_),
    .Q_N(_0785_),
    .Q(\dev_regs[1][4] ));
 sg13g2_dfrbp_1 _1553_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net301),
    .D(_0130_),
    .Q_N(_0784_),
    .Q(\dev_regs[1][5] ));
 sg13g2_dfrbp_1 _1554_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net301),
    .D(_0131_),
    .Q_N(_0783_),
    .Q(\dev_regs[1][6] ));
 sg13g2_dfrbp_1 _1555_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net297),
    .D(_0132_),
    .Q_N(_0782_),
    .Q(\cycles_high[0] ));
 sg13g2_dfrbp_1 _1556_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net297),
    .D(_0133_),
    .Q_N(_0781_),
    .Q(\cycles_high[1] ));
 sg13g2_dfrbp_1 _1557_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net299),
    .D(_0134_),
    .Q_N(\cycles_high[2] ),
    .Q(_0037_));
 sg13g2_dfrbp_1 _1558_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net298),
    .D(_0135_),
    .Q_N(_0780_),
    .Q(\cycles_high[3] ));
 sg13g2_dfrbp_1 _1559_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net301),
    .D(_0136_),
    .Q_N(\cycles_high[4] ),
    .Q(_0038_));
 sg13g2_dfrbp_1 _1560_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net297),
    .D(_0137_),
    .Q_N(_0779_),
    .Q(\cycles_high[5] ));
 sg13g2_dfrbp_1 _1561_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net296),
    .D(_0138_),
    .Q_N(_0778_),
    .Q(\cycles_high[6] ));
 sg13g2_dfrbp_1 _1562_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net301),
    .D(net106),
    .Q_N(_0777_),
    .Q(\cycles_high[7] ));
 sg13g2_dfrbp_1 _1563_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net301),
    .D(_0140_),
    .Q_N(_0776_),
    .Q(\cycles_high[8] ));
 sg13g2_dfrbp_1 _1564_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net297),
    .D(_0141_),
    .Q_N(\cycles_high[9] ),
    .Q(_0039_));
 sg13g2_dfrbp_1 _1565_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net299),
    .D(_0142_),
    .Q_N(_0775_),
    .Q(\cycles_high[10] ));
 sg13g2_dfrbp_1 _1566_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net299),
    .D(_0143_),
    .Q_N(_0774_),
    .Q(\cycles_high[11] ));
 sg13g2_dfrbp_1 _1567_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net300),
    .D(_0144_),
    .Q_N(_0773_),
    .Q(\cycles_high[12] ));
 sg13g2_dfrbp_1 _1568_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net300),
    .D(_0145_),
    .Q_N(_0772_),
    .Q(\cycles_high[13] ));
 sg13g2_dfrbp_1 _1569_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net300),
    .D(_0146_),
    .Q_N(_0771_),
    .Q(\cycles_high[14] ));
 sg13g2_dfrbp_1 _1570_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net300),
    .D(_0147_),
    .Q_N(\cycles_high[15] ),
    .Q(_0040_));
 sg13g2_dfrbp_1 _1571_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net297),
    .D(_0148_),
    .Q_N(_0770_),
    .Q(\cycles_freq[0] ));
 sg13g2_dfrbp_1 _1572_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net297),
    .D(_0149_),
    .Q_N(_0769_),
    .Q(\cycles_freq[1] ));
 sg13g2_dfrbp_1 _1573_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net298),
    .D(_0150_),
    .Q_N(_0768_),
    .Q(\cycles_freq[2] ));
 sg13g2_dfrbp_1 _1574_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net298),
    .D(_0151_),
    .Q_N(_0767_),
    .Q(\cycles_freq[3] ));
 sg13g2_dfrbp_1 _1575_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net300),
    .D(_0152_),
    .Q_N(\cycles_freq[4] ),
    .Q(_0041_));
 sg13g2_dfrbp_1 _1576_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net296),
    .D(_0153_),
    .Q_N(_0766_),
    .Q(\cycles_freq[5] ));
 sg13g2_dfrbp_1 _1577_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net300),
    .D(_0154_),
    .Q_N(\cycles_freq[6] ),
    .Q(_0042_));
 sg13g2_dfrbp_1 _1578_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net301),
    .D(net94),
    .Q_N(_0765_),
    .Q(\cycles_freq[7] ));
 sg13g2_dfrbp_1 _1579_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net303),
    .D(_0156_),
    .Q_N(\cycles_freq[8] ),
    .Q(_0043_));
 sg13g2_dfrbp_1 _1580_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net302),
    .D(_0157_),
    .Q_N(\cycles_freq[9] ),
    .Q(_0044_));
 sg13g2_dfrbp_1 _1581_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net297),
    .D(_0158_),
    .Q_N(_0764_),
    .Q(\cycles_freq[10] ));
 sg13g2_dfrbp_1 _1582_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net297),
    .D(_0159_),
    .Q_N(_0763_),
    .Q(\cycles_freq[11] ));
 sg13g2_dfrbp_1 _1583_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net302),
    .D(_0160_),
    .Q_N(_0762_),
    .Q(\cycles_freq[12] ));
 sg13g2_dfrbp_1 _1584_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net300),
    .D(_0161_),
    .Q_N(_0761_),
    .Q(\cycles_freq[13] ));
 sg13g2_dfrbp_1 _1585_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net300),
    .D(_0162_),
    .Q_N(\cycles_freq[14] ),
    .Q(_0045_));
 sg13g2_dfrbp_1 _1586_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net302),
    .D(net49),
    .Q_N(\cycles_freq[15] ),
    .Q(_0046_));
 sg13g2_dfrbp_1 _1587_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net303),
    .D(_0164_),
    .Q_N(_0760_),
    .Q(uio_oe[0]));
 sg13g2_dfrbp_1 _1588_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net303),
    .D(_0165_),
    .Q_N(_0759_),
    .Q(uio_oe[1]));
 sg13g2_dfrbp_1 _1589_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net313),
    .D(_0166_),
    .Q_N(_0758_),
    .Q(uio_oe[2]));
 sg13g2_dfrbp_1 _1590_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net304),
    .D(_0167_),
    .Q_N(_0757_),
    .Q(uio_oe[3]));
 sg13g2_dfrbp_1 _1591_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net302),
    .D(_0168_),
    .Q_N(_0756_),
    .Q(uio_oe[4]));
 sg13g2_dfrbp_1 _1592_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net302),
    .D(_0169_),
    .Q_N(_0755_),
    .Q(uio_oe[5]));
 sg13g2_dfrbp_1 _1593_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net302),
    .D(_0170_),
    .Q_N(_0754_),
    .Q(uio_oe[6]));
 sg13g2_dfrbp_1 _1594_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net302),
    .D(_0171_),
    .Q_N(_0753_),
    .Q(uio_oe[7]));
 sg13g2_dfrbp_1 _1595_ (.CLK(net294),
    .RESET_B(_0049_),
    .D(_0048_),
    .Q_N(\spi_own_clock_ins.spi_state[0] ),
    .Q(_0047_));
 sg13g2_dfrbp_1 _1596_ (.CLK(net292),
    .RESET_B(_0050_),
    .D(_0001_),
    .Q_N(_0023_),
    .Q(\spi_own_clock_ins.spi_state[1] ));
 sg13g2_dfrbp_1 _1597_ (.CLK(net292),
    .RESET_B(_0051_),
    .D(_0002_),
    .Q_N(_0022_),
    .Q(\spi_own_clock_ins.spi_state[2] ));
 sg13g2_dfrbp_1 _1598_ (.CLK(net292),
    .RESET_B(_0052_),
    .D(_0003_),
    .Q_N(_0752_),
    .Q(\spi_own_clock_ins.spi_state[3] ));
 sg13g2_dfrbp_1 _1599_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net304),
    .D(_0172_),
    .Q_N(_0751_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _1600_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net304),
    .D(_0173_),
    .Q_N(_0750_),
    .Q(uio_out[1]));
 sg13g2_dfrbp_1 _1601_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net305),
    .D(_0174_),
    .Q_N(_0749_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _1602_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net304),
    .D(_0175_),
    .Q_N(_0748_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _1603_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net304),
    .D(_0176_),
    .Q_N(_0747_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _1604_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net302),
    .D(_0177_),
    .Q_N(_0746_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _1605_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net303),
    .D(_0178_),
    .Q_N(_0745_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _1606_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net303),
    .D(net88),
    .Q_N(_0744_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _1607_ (.CLK(net292),
    .RESET_B(_0053_),
    .D(_0180_),
    .Q_N(_0743_),
    .Q(\spi_own_clock_ins.index[0] ));
 sg13g2_dfrbp_1 _1608_ (.CLK(net292),
    .RESET_B(_0054_),
    .D(_0181_),
    .Q_N(_0742_),
    .Q(\spi_own_clock_ins.index[1] ));
 sg13g2_dfrbp_1 _1609_ (.CLK(net294),
    .RESET_B(_0055_),
    .D(_0182_),
    .Q_N(_0025_),
    .Q(\spi_own_clock_ins.index[2] ));
 sg13g2_dfrbp_1 _1610_ (.CLK(net294),
    .RESET_B(_0056_),
    .D(_0183_),
    .Q_N(_0026_),
    .Q(\spi_own_clock_ins.index[3] ));
 sg13g2_dfrbp_1 _1611_ (.CLK(net291),
    .RESET_B(_0057_),
    .D(_0184_),
    .Q_N(_0741_),
    .Q(\addr_reg_clk[0] ));
 sg13g2_dfrbp_1 _1612_ (.CLK(net291),
    .RESET_B(_0058_),
    .D(_0185_),
    .Q_N(_0740_),
    .Q(\addr_reg_clk[1] ));
 sg13g2_dfrbp_1 _1613_ (.CLK(net291),
    .RESET_B(_0059_),
    .D(_0186_),
    .Q_N(_0020_),
    .Q(\addr_reg_clk[2] ));
 sg13g2_dfrbp_1 _1614_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net298),
    .D(net58),
    .Q_N(_0739_),
    .Q(pwm));
 sg13g2_dfrbp_1 _1615_ (.CLK(net294),
    .RESET_B(_0060_),
    .D(_0188_),
    .Q_N(_0738_),
    .Q(\spi_own_clock_ins.data_rd[0] ));
 sg13g2_dfrbp_1 _1616_ (.CLK(net294),
    .RESET_B(_0061_),
    .D(_0189_),
    .Q_N(_0737_),
    .Q(\spi_own_clock_ins.data_rd[1] ));
 sg13g2_dfrbp_1 _1617_ (.CLK(net293),
    .RESET_B(_0062_),
    .D(_0190_),
    .Q_N(_0736_),
    .Q(\spi_own_clock_ins.data_rd[2] ));
 sg13g2_dfrbp_1 _1618_ (.CLK(net293),
    .RESET_B(_0063_),
    .D(_0191_),
    .Q_N(_0735_),
    .Q(\spi_own_clock_ins.data_rd[3] ));
 sg13g2_dfrbp_1 _1619_ (.CLK(net292),
    .RESET_B(_0064_),
    .D(_0192_),
    .Q_N(_0734_),
    .Q(\spi_own_clock_ins.data_rd[4] ));
 sg13g2_dfrbp_1 _1620_ (.CLK(net292),
    .RESET_B(_0065_),
    .D(_0193_),
    .Q_N(_0733_),
    .Q(\spi_own_clock_ins.data_rd[5] ));
 sg13g2_dfrbp_1 _1621_ (.CLK(net292),
    .RESET_B(_0066_),
    .D(_0194_),
    .Q_N(_0732_),
    .Q(\spi_own_clock_ins.data_rd[6] ));
 sg13g2_dfrbp_1 _1622_ (.CLK(net293),
    .RESET_B(_0067_),
    .D(_0195_),
    .Q_N(_0731_),
    .Q(\spi_own_clock_ins.data_rd[7] ));
 sg13g2_dfrbp_1 _1623_ (.CLK(_0069_),
    .RESET_B(_0068_),
    .D(net2),
    .Q_N(_0730_),
    .Q(\spi_own_clock_ins.spi_data_reg[0] ));
 sg13g2_dfrbp_1 _1624_ (.CLK(_0071_),
    .RESET_B(_0070_),
    .D(\spi_own_clock_ins.spi_data_reg[0] ),
    .Q_N(_0729_),
    .Q(\spi_own_clock_ins.spi_data_reg[1] ));
 sg13g2_dfrbp_1 _1625_ (.CLK(_0073_),
    .RESET_B(_0072_),
    .D(\spi_own_clock_ins.spi_data_reg[1] ),
    .Q_N(_0728_),
    .Q(\spi_own_clock_ins.spi_data_reg[2] ));
 sg13g2_dfrbp_1 _1626_ (.CLK(_0075_),
    .RESET_B(_0074_),
    .D(\spi_own_clock_ins.spi_data_reg[2] ),
    .Q_N(_0727_),
    .Q(\spi_own_clock_ins.spi_data_reg[3] ));
 sg13g2_dfrbp_1 _1627_ (.CLK(_0077_),
    .RESET_B(_0076_),
    .D(\spi_own_clock_ins.spi_data_reg[3] ),
    .Q_N(_0726_),
    .Q(\spi_own_clock_ins.spi_data_reg[4] ));
 sg13g2_dfrbp_1 _1628_ (.CLK(_0079_),
    .RESET_B(_0078_),
    .D(\spi_own_clock_ins.spi_data_reg[4] ),
    .Q_N(_0725_),
    .Q(\spi_own_clock_ins.spi_data_reg[5] ));
 sg13g2_dfrbp_1 _1629_ (.CLK(_0081_),
    .RESET_B(_0080_),
    .D(\spi_own_clock_ins.spi_data_reg[5] ),
    .Q_N(_0724_),
    .Q(\spi_own_clock_ins.spi_data_reg[6] ));
 sg13g2_dfrbp_1 _1630_ (.CLK(_0083_),
    .RESET_B(_0082_),
    .D(\spi_own_clock_ins.spi_data_reg[6] ),
    .Q_N(_0805_),
    .Q(\spi_own_clock_ins.spi_data_reg[7] ));
 sg13g2_dfrbp_1 _1631_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net314),
    .D(net38),
    .Q_N(_0806_),
    .Q(\spi_sampled_ins.neg_edge_det.signal_z1 ));
 sg13g2_dfrbp_1 _1632_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net312),
    .D(_0000_),
    .Q_N(_0723_),
    .Q(\dev_regs[1][7] ));
 sg13g2_dfrbp_1 _1633_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(_0084_),
    .D(net72),
    .Q_N(_0722_),
    .Q(\addr_reg_sampled[0] ));
 sg13g2_dfrbp_1 _1634_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(_0085_),
    .D(net75),
    .Q_N(_0721_),
    .Q(\addr_reg_sampled[1] ));
 sg13g2_dfrbp_1 _1635_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(_0086_),
    .D(net77),
    .Q_N(_0021_),
    .Q(\addr_reg_sampled[2] ));
 sg13g2_dfrbp_1 _1636_ (.CLK(net293),
    .RESET_B(_0087_),
    .D(_0199_),
    .Q_N(_0720_),
    .Q(\spi_own_clock_ins.data_rd_z1[0] ));
 sg13g2_dfrbp_1 _1637_ (.CLK(net293),
    .RESET_B(_0088_),
    .D(_0200_),
    .Q_N(_0719_),
    .Q(\spi_own_clock_ins.data_rd_z1[1] ));
 sg13g2_dfrbp_1 _1638_ (.CLK(net293),
    .RESET_B(_0089_),
    .D(_0201_),
    .Q_N(_0718_),
    .Q(\spi_own_clock_ins.data_rd_z1[2] ));
 sg13g2_dfrbp_1 _1639_ (.CLK(net293),
    .RESET_B(_0090_),
    .D(_0202_),
    .Q_N(_0717_),
    .Q(\spi_own_clock_ins.data_rd_z1[3] ));
 sg13g2_dfrbp_1 _1640_ (.CLK(net291),
    .RESET_B(_0091_),
    .D(_0203_),
    .Q_N(_0716_),
    .Q(\spi_own_clock_ins.data_rd_z1[4] ));
 sg13g2_dfrbp_1 _1641_ (.CLK(net291),
    .RESET_B(_0092_),
    .D(_0204_),
    .Q_N(_0715_),
    .Q(\spi_own_clock_ins.data_rd_z1[5] ));
 sg13g2_dfrbp_1 _1642_ (.CLK(net291),
    .RESET_B(_0093_),
    .D(_0205_),
    .Q_N(_0714_),
    .Q(\spi_own_clock_ins.data_rd_z1[6] ));
 sg13g2_dfrbp_1 _1643_ (.CLK(net290),
    .RESET_B(_0094_),
    .D(_0206_),
    .Q_N(_0713_),
    .Q(\spi_own_clock_ins.data_rd_z1[7] ));
 sg13g2_dfrbp_1 _1644_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(_0095_),
    .D(_0207_),
    .Q_N(_0712_),
    .Q(\spi_sampled_ins.spi_state[0] ));
 sg13g2_dfrbp_1 _1645_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(_0096_),
    .D(net56),
    .Q_N(_0711_),
    .Q(\spi_sampled_ins.spi_state[1] ));
 sg13g2_dfrbp_1 _1646_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(_0097_),
    .D(_0209_),
    .Q_N(_0710_),
    .Q(\spi_sampled_ins.index[0] ));
 sg13g2_dfrbp_1 _1647_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(_0098_),
    .D(_0210_),
    .Q_N(_0709_),
    .Q(\spi_sampled_ins.index[1] ));
 sg13g2_dfrbp_1 _1648_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(_0099_),
    .D(net116),
    .Q_N(_0027_),
    .Q(\spi_sampled_ins.index[2] ));
 sg13g2_dfrbp_1 _1649_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(_0100_),
    .D(net102),
    .Q_N(_0028_),
    .Q(\spi_sampled_ins.index[3] ));
 sg13g2_dfrbp_1 _1650_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net29),
    .D(net3),
    .Q_N(_0807_),
    .Q(\spi_sampled_ins.sclk_z1 ));
 sg13g2_dfrbp_1 _1651_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net30),
    .D(net35),
    .Q_N(_0808_),
    .Q(\spi_sampled_ins.neg_edge_det.signal ));
 sg13g2_dfrbp_1 _1652_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net31),
    .D(net4),
    .Q_N(_0809_),
    .Q(\spi_sampled_ins.mosi_z1 ));
 sg13g2_dfrbp_1 _1653_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net32),
    .D(net36),
    .Q_N(_0810_),
    .Q(\spi_sampled_ins.mosi ));
 sg13g2_dfrbp_1 _1654_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net33),
    .D(net5),
    .Q_N(_0811_),
    .Q(\spi_sampled_ins.cs_z1 ));
 sg13g2_dfrbp_1 _1655_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net34),
    .D(net37),
    .Q_N(_0812_),
    .Q(\spi_sampled_ins.cs ));
 sg13g2_dfrbp_1 _1656_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net298),
    .D(_0004_),
    .Q_N(_0813_),
    .Q(\pwm_inst.counter[0] ));
 sg13g2_dfrbp_1 _1657_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net298),
    .D(net150),
    .Q_N(_0814_),
    .Q(\pwm_inst.counter[1] ));
 sg13g2_dfrbp_1 _1658_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net298),
    .D(net129),
    .Q_N(_0815_),
    .Q(\pwm_inst.counter[2] ));
 sg13g2_dfrbp_1 _1659_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net298),
    .D(_0013_),
    .Q_N(_0816_),
    .Q(\pwm_inst.counter[3] ));
 sg13g2_dfrbp_1 _1660_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net295),
    .D(_0014_),
    .Q_N(_0817_),
    .Q(\pwm_inst.counter[4] ));
 sg13g2_dfrbp_1 _1661_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net295),
    .D(net158),
    .Q_N(_0818_),
    .Q(\pwm_inst.counter[5] ));
 sg13g2_dfrbp_1 _1662_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net295),
    .D(_0016_),
    .Q_N(_0819_),
    .Q(\pwm_inst.counter[6] ));
 sg13g2_dfrbp_1 _1663_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net295),
    .D(_0017_),
    .Q_N(_0820_),
    .Q(\pwm_inst.counter[7] ));
 sg13g2_dfrbp_1 _1664_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net295),
    .D(_0018_),
    .Q_N(_0821_),
    .Q(\pwm_inst.counter[8] ));
 sg13g2_dfrbp_1 _1665_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net295),
    .D(_0019_),
    .Q_N(_0822_),
    .Q(\pwm_inst.counter[9] ));
 sg13g2_dfrbp_1 _1666_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net295),
    .D(_0005_),
    .Q_N(_0823_),
    .Q(\pwm_inst.counter[10] ));
 sg13g2_dfrbp_1 _1667_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net296),
    .D(net64),
    .Q_N(_0824_),
    .Q(\pwm_inst.counter[11] ));
 sg13g2_dfrbp_1 _1668_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net295),
    .D(net144),
    .Q_N(_0825_),
    .Q(\pwm_inst.counter[12] ));
 sg13g2_dfrbp_1 _1669_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net296),
    .D(net131),
    .Q_N(_0826_),
    .Q(\pwm_inst.counter[13] ));
 sg13g2_dfrbp_1 _1670_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net296),
    .D(_0009_),
    .Q_N(_0827_),
    .Q(\pwm_inst.counter[14] ));
 sg13g2_dfrbp_1 _1671_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net296),
    .D(net112),
    .Q_N(_0708_),
    .Q(\pwm_inst.counter[15] ));
 sg13g2_tiehi _1530__22 (.L_HI(net22));
 sg13g2_tiehi _1529__23 (.L_HI(net23));
 sg13g2_tiehi _1528__24 (.L_HI(net24));
 sg13g2_tiehi _1527__25 (.L_HI(net25));
 sg13g2_tiehi _1526__26 (.L_HI(net26));
 sg13g2_tiehi _1525__27 (.L_HI(net27));
 sg13g2_tiehi _1524__28 (.L_HI(net28));
 sg13g2_tiehi _1650__29 (.L_HI(net29));
 sg13g2_tiehi _1651__30 (.L_HI(net30));
 sg13g2_tiehi _1652__31 (.L_HI(net31));
 sg13g2_tiehi _1653__32 (.L_HI(net32));
 sg13g2_tiehi _1654__33 (.L_HI(net33));
 sg13g2_tiehi _1655__34 (.L_HI(net34));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_spi_pwm_djuara_17 (.L_LO(net17));
 sg13g2_tielo tt_um_spi_pwm_djuara_18 (.L_LO(net18));
 sg13g2_tielo tt_um_spi_pwm_djuara_19 (.L_LO(net19));
 sg13g2_tielo tt_um_spi_pwm_djuara_20 (.L_LO(net20));
 sg13g2_tiehi _1531__21 (.L_HI(net21));
 sg13g2_buf_2 _1691_ (.A(miso_clk),
    .X(uo_out[0]));
 sg13g2_buf_1 _1692_ (.A(miso_sampled),
    .X(uo_out[1]));
 sg13g2_buf_2 _1693_ (.A(pwm),
    .X(uo_out[2]));
 sg13g2_buf_2 fanout239 (.A(net240),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_0482_),
    .X(net240));
 sg13g2_buf_4 fanout241 (.X(net241),
    .A(_0703_));
 sg13g2_buf_2 fanout242 (.A(net243),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_0695_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_0687_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_0687_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_0672_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_0672_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(net249),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_0520_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_0430_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(net254),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(net253),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(net254),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_0422_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(net256),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_0575_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_0427_),
    .X(net257));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(_0577_));
 sg13g2_buf_2 fanout259 (.A(_0573_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_0571_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_0567_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_0425_),
    .X(net262));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(_0313_));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(_0312_));
 sg13g2_buf_2 fanout265 (.A(_0310_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_0309_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_0307_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_0305_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(net271),
    .X(net269));
 sg13g2_buf_1 fanout270 (.A(net271),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_0581_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_0522_),
    .X(net272));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(_0521_));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(_0316_));
 sg13g2_buf_2 fanout275 (.A(net276),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_0311_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(net157),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(\pwm_inst.counter[1] ),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net122),
    .X(net279));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(\spi_own_clock_ins.index[0] ));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(\spi_own_clock_ins.spi_state[2] ));
 sg13g2_buf_2 fanout282 (.A(\spi_own_clock_ins.spi_state[2] ),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(net284),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(\spi_own_clock_ins.spi_state[2] ),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(ui_in[2]),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(ui_in[2]),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(net289),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(ui_in[2]),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(ui_in[0]),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(ui_in[0]),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(net294),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(net294),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(ui_in[0]),
    .X(net294));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(net296));
 sg13g2_buf_4 fanout296 (.X(net296),
    .A(net307));
 sg13g2_buf_4 fanout297 (.X(net297),
    .A(net299));
 sg13g2_buf_4 fanout298 (.X(net298),
    .A(net307));
 sg13g2_buf_2 fanout299 (.A(net307),
    .X(net299));
 sg13g2_buf_4 fanout300 (.X(net300),
    .A(net301));
 sg13g2_buf_4 fanout301 (.X(net301),
    .A(net306));
 sg13g2_buf_4 fanout302 (.X(net302),
    .A(net306));
 sg13g2_buf_4 fanout303 (.X(net303),
    .A(net306));
 sg13g2_buf_4 fanout304 (.X(net304),
    .A(net306));
 sg13g2_buf_2 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(net307),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(rst_n),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(net310),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(net310),
    .X(net309));
 sg13g2_buf_1 fanout310 (.A(net311),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(rst_n),
    .X(net311));
 sg13g2_buf_4 fanout312 (.X(net312),
    .A(net315));
 sg13g2_buf_2 fanout313 (.A(net315),
    .X(net313));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(net315));
 sg13g2_buf_2 fanout315 (.A(rst_n),
    .X(net315));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[0]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[3]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[4]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[6]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[7]),
    .X(net15));
 sg13g2_tielo tt_um_spi_pwm_djuara_16 (.L_LO(net16));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\spi_sampled_ins.sclk_z1 ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold2 (.A(\spi_sampled_ins.mosi_z1 ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold3 (.A(\spi_sampled_ins.cs_z1 ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold4 (.A(\spi_sampled_ins.neg_edge_det.signal ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0036_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0033_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0034_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0035_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold9 (.A(\dev_regs[0][3] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0038_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0042_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0041_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0044_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0046_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0163_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold16 (.A(\dev_regs[0][0] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0045_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0037_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold19 (.A(\dev_regs[0][5] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold20 (.A(\dev_regs[0][6] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0024_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0208_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold23 (.A(pwm),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0187_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold25 (.A(\spi_sampled_ins.spi_data_reg[6] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0418_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0116_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0040_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold29 (.A(\pwm_inst.counter[11] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0006_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0043_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0039_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold33 (.A(\spi_sampled_ins.mosi ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0109_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold35 (.A(uio_out[3]),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold36 (.A(\dev_regs[1][1] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold37 (.A(\spi_sampled_ins.spi_data_reg[0] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0196_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold39 (.A(uio_out[2]),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold40 (.A(\spi_sampled_ins.spi_data_reg[1] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0197_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold42 (.A(\spi_sampled_ins.spi_data_reg[2] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0198_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold44 (.A(\cycles_freq[0] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold45 (.A(\spi_sampled_ins.spi_data_reg[4] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0113_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold47 (.A(\spi_sampled_ins.neg_edge_det.signal_z1 ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold48 (.A(uio_out[4]),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold49 (.A(uio_out[0]),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold50 (.A(\cycles_high[0] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold51 (.A(\spi_sampled_ins.spi_data_reg[5] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold52 (.A(uio_out[1]),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold53 (.A(uio_out[7]),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0179_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold55 (.A(\spi_sampled_ins.spi_data_reg[3] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold56 (.A(\dev_regs[1][3] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold57 (.A(uio_out[6]),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold58 (.A(uio_out[5]),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold59 (.A(\cycles_freq[7] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0155_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold61 (.A(\data_wr_z1[2] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold62 (.A(\dev_regs[1][5] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold63 (.A(\dev_regs[1][4] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold64 (.A(\data_wr_z1[0] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold65 (.A(\cycles_freq[1] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold66 (.A(\dev_regs[1][6] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold67 (.A(\spi_sampled_ins.index[3] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0212_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold69 (.A(\dev_regs[1][2] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold70 (.A(\data_wr_z1[3] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cycles_high[7] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0139_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold73 (.A(\cycles_high[1] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold74 (.A(\cycles_freq[5] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold75 (.A(\data_wr_z1[1] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold76 (.A(\data_wr_z1[5] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold77 (.A(\pwm_inst.counter[15] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0010_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold79 (.A(\cycles_high[6] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold80 (.A(\data_wr_z1[6] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold81 (.A(\spi_sampled_ins.index[2] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0211_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold83 (.A(\dev_regs[1][0] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold84 (.A(\data_wr_z1[4] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold85 (.A(uio_oe[7]),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold86 (.A(uio_oe[0]),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold87 (.A(uio_oe[5]),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold88 (.A(\spi_sampled_ins.cs ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold89 (.A(uio_oe[1]),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cycles_high[13] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold91 (.A(\spi_sampled_ins.spi_state[0] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0303_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold93 (.A(uio_oe[4]),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold94 (.A(\pwm_inst.counter[2] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0012_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold96 (.A(\pwm_inst.counter[13] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0008_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold98 (.A(\cycles_high[14] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold99 (.A(\cycles_freq[12] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold100 (.A(\cycles_freq[13] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold101 (.A(\cycles_high[10] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cycles_high[5] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold103 (.A(uio_oe[2]),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cycles_freq[10] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold105 (.A(\cycles_high[3] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cycles_high[12] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold107 (.A(uio_oe[6]),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cycles_freq[2] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold109 (.A(\pwm_inst.counter[12] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0007_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold111 (.A(uio_oe[3]),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold112 (.A(\cycles_freq[3] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold113 (.A(\cycles_high[11] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold114 (.A(\cycles_high[8] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold115 (.A(\pwm_inst.counter[0] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0011_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold117 (.A(\data_wr_z1[7] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cycles_freq[11] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold119 (.A(\pwm_inst.counter[4] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0532_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold121 (.A(\pwm_inst.counter[7] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0539_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold123 (.A(\pwm_inst.counter[5] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0015_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold125 (.A(\pwm_inst.counter[9] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0544_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold127 (.A(\pwm_inst.counter[14] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0556_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold129 (.A(\pwm_inst.counter[8] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold130 (.A(\spi_sampled_ins.index[1] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold131 (.A(\pwm_inst.counter[3] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0529_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0530_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold134 (.A(\pwm_inst.counter[6] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold135 (.A(\pwm_inst.counter[10] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold136 (.A(\spi_sampled_ins.index[0] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0812_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold138 (.A(\pwm_inst.counter[6] ),
    .X(net172));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_fill_2 FILLER_9_42 ();
 sg13g2_fill_1 FILLER_9_44 ();
 sg13g2_fill_1 FILLER_9_75 ();
 sg13g2_decap_8 FILLER_9_81 ();
 sg13g2_decap_8 FILLER_9_88 ();
 sg13g2_decap_8 FILLER_9_99 ();
 sg13g2_decap_8 FILLER_9_106 ();
 sg13g2_decap_8 FILLER_9_113 ();
 sg13g2_decap_8 FILLER_9_120 ();
 sg13g2_decap_8 FILLER_9_127 ();
 sg13g2_fill_2 FILLER_9_134 ();
 sg13g2_decap_4 FILLER_9_140 ();
 sg13g2_fill_2 FILLER_9_144 ();
 sg13g2_decap_8 FILLER_9_150 ();
 sg13g2_decap_8 FILLER_9_157 ();
 sg13g2_decap_8 FILLER_9_164 ();
 sg13g2_decap_8 FILLER_9_171 ();
 sg13g2_decap_8 FILLER_9_178 ();
 sg13g2_decap_8 FILLER_9_185 ();
 sg13g2_decap_8 FILLER_9_192 ();
 sg13g2_decap_8 FILLER_9_199 ();
 sg13g2_decap_8 FILLER_9_206 ();
 sg13g2_decap_8 FILLER_9_213 ();
 sg13g2_decap_8 FILLER_9_220 ();
 sg13g2_decap_8 FILLER_9_227 ();
 sg13g2_decap_8 FILLER_9_234 ();
 sg13g2_decap_8 FILLER_9_241 ();
 sg13g2_decap_8 FILLER_9_248 ();
 sg13g2_decap_8 FILLER_9_255 ();
 sg13g2_decap_8 FILLER_9_262 ();
 sg13g2_decap_8 FILLER_9_269 ();
 sg13g2_decap_8 FILLER_9_276 ();
 sg13g2_decap_8 FILLER_9_283 ();
 sg13g2_decap_8 FILLER_9_290 ();
 sg13g2_decap_8 FILLER_9_297 ();
 sg13g2_decap_8 FILLER_9_304 ();
 sg13g2_decap_8 FILLER_9_311 ();
 sg13g2_decap_8 FILLER_9_318 ();
 sg13g2_decap_8 FILLER_9_325 ();
 sg13g2_decap_8 FILLER_9_332 ();
 sg13g2_decap_8 FILLER_9_339 ();
 sg13g2_decap_8 FILLER_9_346 ();
 sg13g2_decap_8 FILLER_9_353 ();
 sg13g2_decap_8 FILLER_9_360 ();
 sg13g2_decap_8 FILLER_9_367 ();
 sg13g2_decap_8 FILLER_9_374 ();
 sg13g2_decap_8 FILLER_9_381 ();
 sg13g2_decap_8 FILLER_9_388 ();
 sg13g2_decap_8 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_4 FILLER_10_28 ();
 sg13g2_fill_1 FILLER_10_32 ();
 sg13g2_fill_1 FILLER_10_38 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_4 FILLER_10_56 ();
 sg13g2_decap_4 FILLER_10_86 ();
 sg13g2_fill_1 FILLER_10_100 ();
 sg13g2_decap_4 FILLER_10_116 ();
 sg13g2_fill_2 FILLER_10_134 ();
 sg13g2_fill_1 FILLER_10_136 ();
 sg13g2_decap_8 FILLER_10_173 ();
 sg13g2_decap_8 FILLER_10_180 ();
 sg13g2_decap_8 FILLER_10_187 ();
 sg13g2_decap_8 FILLER_10_194 ();
 sg13g2_decap_8 FILLER_10_201 ();
 sg13g2_decap_8 FILLER_10_208 ();
 sg13g2_decap_8 FILLER_10_215 ();
 sg13g2_decap_8 FILLER_10_222 ();
 sg13g2_decap_8 FILLER_10_229 ();
 sg13g2_decap_8 FILLER_10_236 ();
 sg13g2_decap_8 FILLER_10_243 ();
 sg13g2_decap_8 FILLER_10_250 ();
 sg13g2_decap_8 FILLER_10_257 ();
 sg13g2_decap_8 FILLER_10_264 ();
 sg13g2_decap_8 FILLER_10_271 ();
 sg13g2_decap_8 FILLER_10_278 ();
 sg13g2_decap_8 FILLER_10_285 ();
 sg13g2_decap_8 FILLER_10_292 ();
 sg13g2_decap_8 FILLER_10_299 ();
 sg13g2_decap_8 FILLER_10_306 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_decap_8 FILLER_10_327 ();
 sg13g2_decap_8 FILLER_10_334 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_decap_8 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_362 ();
 sg13g2_decap_8 FILLER_10_369 ();
 sg13g2_decap_8 FILLER_10_376 ();
 sg13g2_decap_8 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_fill_1 FILLER_11_21 ();
 sg13g2_fill_2 FILLER_11_58 ();
 sg13g2_fill_1 FILLER_11_60 ();
 sg13g2_fill_1 FILLER_11_141 ();
 sg13g2_fill_2 FILLER_11_156 ();
 sg13g2_decap_8 FILLER_11_170 ();
 sg13g2_decap_8 FILLER_11_177 ();
 sg13g2_decap_8 FILLER_11_184 ();
 sg13g2_decap_8 FILLER_11_191 ();
 sg13g2_decap_8 FILLER_11_198 ();
 sg13g2_decap_8 FILLER_11_205 ();
 sg13g2_decap_8 FILLER_11_212 ();
 sg13g2_decap_8 FILLER_11_219 ();
 sg13g2_decap_8 FILLER_11_226 ();
 sg13g2_decap_8 FILLER_11_233 ();
 sg13g2_decap_8 FILLER_11_240 ();
 sg13g2_decap_8 FILLER_11_247 ();
 sg13g2_decap_4 FILLER_11_254 ();
 sg13g2_decap_8 FILLER_11_284 ();
 sg13g2_decap_8 FILLER_11_291 ();
 sg13g2_decap_8 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_9 ();
 sg13g2_fill_2 FILLER_12_18 ();
 sg13g2_fill_1 FILLER_12_20 ();
 sg13g2_fill_1 FILLER_12_34 ();
 sg13g2_fill_2 FILLER_12_45 ();
 sg13g2_fill_1 FILLER_12_47 ();
 sg13g2_fill_1 FILLER_12_68 ();
 sg13g2_fill_1 FILLER_12_78 ();
 sg13g2_fill_1 FILLER_12_104 ();
 sg13g2_decap_8 FILLER_12_181 ();
 sg13g2_decap_8 FILLER_12_188 ();
 sg13g2_decap_8 FILLER_12_195 ();
 sg13g2_decap_8 FILLER_12_202 ();
 sg13g2_decap_8 FILLER_12_209 ();
 sg13g2_decap_8 FILLER_12_216 ();
 sg13g2_decap_8 FILLER_12_223 ();
 sg13g2_fill_2 FILLER_12_230 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_fill_2 FILLER_12_242 ();
 sg13g2_fill_2 FILLER_12_247 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_fill_2 FILLER_12_266 ();
 sg13g2_decap_4 FILLER_12_284 ();
 sg13g2_fill_2 FILLER_12_288 ();
 sg13g2_decap_8 FILLER_12_300 ();
 sg13g2_fill_2 FILLER_12_307 ();
 sg13g2_fill_1 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_323 ();
 sg13g2_decap_8 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_337 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_decap_8 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_fill_1 FILLER_13_26 ();
 sg13g2_fill_2 FILLER_13_36 ();
 sg13g2_fill_1 FILLER_13_57 ();
 sg13g2_fill_2 FILLER_13_84 ();
 sg13g2_fill_1 FILLER_13_86 ();
 sg13g2_fill_2 FILLER_13_101 ();
 sg13g2_fill_1 FILLER_13_103 ();
 sg13g2_fill_1 FILLER_13_109 ();
 sg13g2_fill_1 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_180 ();
 sg13g2_decap_8 FILLER_13_187 ();
 sg13g2_decap_8 FILLER_13_327 ();
 sg13g2_decap_8 FILLER_13_334 ();
 sg13g2_decap_8 FILLER_13_341 ();
 sg13g2_decap_8 FILLER_13_348 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_decap_8 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_45 ();
 sg13g2_fill_2 FILLER_14_107 ();
 sg13g2_decap_8 FILLER_14_180 ();
 sg13g2_decap_8 FILLER_14_187 ();
 sg13g2_fill_2 FILLER_14_194 ();
 sg13g2_fill_2 FILLER_14_229 ();
 sg13g2_fill_1 FILLER_14_231 ();
 sg13g2_fill_2 FILLER_14_235 ();
 sg13g2_fill_1 FILLER_14_237 ();
 sg13g2_decap_8 FILLER_14_241 ();
 sg13g2_fill_2 FILLER_14_248 ();
 sg13g2_decap_8 FILLER_14_253 ();
 sg13g2_decap_8 FILLER_14_260 ();
 sg13g2_fill_2 FILLER_14_267 ();
 sg13g2_decap_8 FILLER_14_272 ();
 sg13g2_decap_8 FILLER_14_279 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_decap_4 FILLER_14_316 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_358 ();
 sg13g2_fill_2 FILLER_14_365 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_fill_1 FILLER_15_26 ();
 sg13g2_fill_1 FILLER_15_32 ();
 sg13g2_fill_2 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_44 ();
 sg13g2_fill_2 FILLER_15_125 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_fill_1 FILLER_15_201 ();
 sg13g2_fill_2 FILLER_15_228 ();
 sg13g2_decap_8 FILLER_15_256 ();
 sg13g2_fill_2 FILLER_15_263 ();
 sg13g2_fill_1 FILLER_15_265 ();
 sg13g2_decap_8 FILLER_15_310 ();
 sg13g2_decap_8 FILLER_15_317 ();
 sg13g2_fill_1 FILLER_15_324 ();
 sg13g2_fill_2 FILLER_15_343 ();
 sg13g2_fill_1 FILLER_15_345 ();
 sg13g2_fill_1 FILLER_15_364 ();
 sg13g2_decap_4 FILLER_15_383 ();
 sg13g2_fill_1 FILLER_15_387 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_fill_1 FILLER_16_47 ();
 sg13g2_fill_2 FILLER_16_63 ();
 sg13g2_fill_1 FILLER_16_65 ();
 sg13g2_fill_2 FILLER_16_94 ();
 sg13g2_fill_1 FILLER_16_96 ();
 sg13g2_fill_1 FILLER_16_106 ();
 sg13g2_fill_1 FILLER_16_123 ();
 sg13g2_fill_2 FILLER_16_143 ();
 sg13g2_decap_8 FILLER_16_155 ();
 sg13g2_fill_2 FILLER_16_162 ();
 sg13g2_fill_1 FILLER_16_164 ();
 sg13g2_decap_8 FILLER_16_219 ();
 sg13g2_decap_4 FILLER_16_241 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_fill_1 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_342 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_fill_2 FILLER_16_366 ();
 sg13g2_fill_1 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_4 FILLER_16_388 ();
 sg13g2_fill_2 FILLER_16_392 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_11 ();
 sg13g2_fill_1 FILLER_17_34 ();
 sg13g2_fill_1 FILLER_17_40 ();
 sg13g2_fill_2 FILLER_17_60 ();
 sg13g2_fill_1 FILLER_17_62 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_fill_1 FILLER_17_84 ();
 sg13g2_fill_2 FILLER_17_100 ();
 sg13g2_fill_2 FILLER_17_106 ();
 sg13g2_fill_1 FILLER_17_108 ();
 sg13g2_decap_4 FILLER_17_113 ();
 sg13g2_fill_1 FILLER_17_117 ();
 sg13g2_fill_2 FILLER_17_151 ();
 sg13g2_fill_1 FILLER_17_202 ();
 sg13g2_fill_2 FILLER_17_220 ();
 sg13g2_fill_2 FILLER_17_248 ();
 sg13g2_decap_8 FILLER_17_253 ();
 sg13g2_decap_4 FILLER_17_260 ();
 sg13g2_fill_2 FILLER_17_264 ();
 sg13g2_fill_2 FILLER_17_305 ();
 sg13g2_fill_1 FILLER_17_323 ();
 sg13g2_fill_2 FILLER_17_339 ();
 sg13g2_fill_1 FILLER_17_386 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_1 FILLER_18_26 ();
 sg13g2_fill_1 FILLER_18_35 ();
 sg13g2_fill_1 FILLER_18_79 ();
 sg13g2_fill_2 FILLER_18_97 ();
 sg13g2_fill_2 FILLER_18_185 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_1 FILLER_18_219 ();
 sg13g2_decap_4 FILLER_18_234 ();
 sg13g2_fill_2 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_279 ();
 sg13g2_fill_2 FILLER_18_294 ();
 sg13g2_fill_1 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_338 ();
 sg13g2_fill_2 FILLER_18_350 ();
 sg13g2_fill_1 FILLER_18_352 ();
 sg13g2_decap_4 FILLER_18_362 ();
 sg13g2_fill_1 FILLER_18_366 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_46 ();
 sg13g2_fill_1 FILLER_19_48 ();
 sg13g2_fill_1 FILLER_19_58 ();
 sg13g2_fill_1 FILLER_19_63 ();
 sg13g2_fill_2 FILLER_19_69 ();
 sg13g2_fill_1 FILLER_19_71 ();
 sg13g2_fill_1 FILLER_19_80 ();
 sg13g2_fill_2 FILLER_19_102 ();
 sg13g2_fill_2 FILLER_19_119 ();
 sg13g2_fill_1 FILLER_19_126 ();
 sg13g2_fill_2 FILLER_19_140 ();
 sg13g2_fill_1 FILLER_19_142 ();
 sg13g2_fill_1 FILLER_19_180 ();
 sg13g2_decap_8 FILLER_19_199 ();
 sg13g2_decap_4 FILLER_19_206 ();
 sg13g2_fill_1 FILLER_19_210 ();
 sg13g2_fill_1 FILLER_19_217 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_decap_4 FILLER_19_250 ();
 sg13g2_fill_1 FILLER_19_254 ();
 sg13g2_decap_4 FILLER_19_260 ();
 sg13g2_fill_2 FILLER_19_307 ();
 sg13g2_fill_2 FILLER_19_319 ();
 sg13g2_fill_1 FILLER_19_321 ();
 sg13g2_decap_8 FILLER_19_327 ();
 sg13g2_decap_4 FILLER_19_334 ();
 sg13g2_fill_1 FILLER_19_338 ();
 sg13g2_decap_4 FILLER_19_365 ();
 sg13g2_fill_1 FILLER_19_369 ();
 sg13g2_decap_4 FILLER_19_375 ();
 sg13g2_decap_4 FILLER_19_384 ();
 sg13g2_fill_1 FILLER_19_388 ();
 sg13g2_decap_4 FILLER_19_392 ();
 sg13g2_fill_1 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_fill_2 FILLER_20_36 ();
 sg13g2_fill_1 FILLER_20_85 ();
 sg13g2_fill_1 FILLER_20_93 ();
 sg13g2_fill_2 FILLER_20_151 ();
 sg13g2_decap_8 FILLER_20_205 ();
 sg13g2_decap_8 FILLER_20_212 ();
 sg13g2_fill_2 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_decap_4 FILLER_20_232 ();
 sg13g2_fill_1 FILLER_20_241 ();
 sg13g2_fill_1 FILLER_20_283 ();
 sg13g2_fill_1 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_345 ();
 sg13g2_fill_2 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_fill_2 FILLER_20_376 ();
 sg13g2_fill_1 FILLER_20_378 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_11 ();
 sg13g2_fill_2 FILLER_21_17 ();
 sg13g2_decap_4 FILLER_21_46 ();
 sg13g2_fill_2 FILLER_21_50 ();
 sg13g2_fill_2 FILLER_21_109 ();
 sg13g2_fill_1 FILLER_21_111 ();
 sg13g2_fill_2 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_151 ();
 sg13g2_decap_8 FILLER_21_183 ();
 sg13g2_fill_2 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_251 ();
 sg13g2_decap_8 FILLER_21_258 ();
 sg13g2_fill_2 FILLER_21_265 ();
 sg13g2_decap_4 FILLER_21_293 ();
 sg13g2_decap_8 FILLER_21_302 ();
 sg13g2_decap_4 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_313 ();
 sg13g2_fill_2 FILLER_21_319 ();
 sg13g2_fill_1 FILLER_21_321 ();
 sg13g2_decap_8 FILLER_21_327 ();
 sg13g2_decap_4 FILLER_21_334 ();
 sg13g2_decap_8 FILLER_21_374 ();
 sg13g2_fill_1 FILLER_21_381 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_fill_2 FILLER_22_26 ();
 sg13g2_decap_4 FILLER_22_48 ();
 sg13g2_fill_1 FILLER_22_52 ();
 sg13g2_fill_1 FILLER_22_79 ();
 sg13g2_fill_1 FILLER_22_85 ();
 sg13g2_fill_2 FILLER_22_89 ();
 sg13g2_fill_1 FILLER_22_91 ();
 sg13g2_fill_2 FILLER_22_144 ();
 sg13g2_fill_1 FILLER_22_146 ();
 sg13g2_fill_2 FILLER_22_157 ();
 sg13g2_decap_4 FILLER_22_185 ();
 sg13g2_fill_1 FILLER_22_206 ();
 sg13g2_decap_8 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_224 ();
 sg13g2_fill_1 FILLER_22_226 ();
 sg13g2_decap_8 FILLER_22_232 ();
 sg13g2_decap_4 FILLER_22_239 ();
 sg13g2_decap_8 FILLER_22_248 ();
 sg13g2_decap_4 FILLER_22_255 ();
 sg13g2_decap_4 FILLER_22_264 ();
 sg13g2_fill_1 FILLER_22_268 ();
 sg13g2_decap_8 FILLER_22_274 ();
 sg13g2_decap_8 FILLER_22_281 ();
 sg13g2_decap_4 FILLER_22_288 ();
 sg13g2_fill_1 FILLER_22_302 ();
 sg13g2_decap_8 FILLER_22_339 ();
 sg13g2_decap_4 FILLER_22_346 ();
 sg13g2_fill_1 FILLER_22_350 ();
 sg13g2_decap_4 FILLER_22_387 ();
 sg13g2_fill_1 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_34 ();
 sg13g2_fill_1 FILLER_23_36 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_4 FILLER_23_49 ();
 sg13g2_decap_4 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_67 ();
 sg13g2_fill_1 FILLER_23_77 ();
 sg13g2_decap_4 FILLER_23_82 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_fill_2 FILLER_23_101 ();
 sg13g2_fill_1 FILLER_23_103 ();
 sg13g2_decap_4 FILLER_23_155 ();
 sg13g2_fill_2 FILLER_23_188 ();
 sg13g2_fill_1 FILLER_23_190 ();
 sg13g2_fill_2 FILLER_23_236 ();
 sg13g2_decap_4 FILLER_23_316 ();
 sg13g2_fill_1 FILLER_23_320 ();
 sg13g2_decap_4 FILLER_23_326 ();
 sg13g2_decap_4 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_363 ();
 sg13g2_fill_2 FILLER_23_380 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_decap_4 FILLER_24_43 ();
 sg13g2_fill_1 FILLER_24_47 ();
 sg13g2_decap_4 FILLER_24_74 ();
 sg13g2_fill_2 FILLER_24_96 ();
 sg13g2_fill_2 FILLER_24_109 ();
 sg13g2_fill_2 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_fill_1 FILLER_24_127 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_fill_2 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_182 ();
 sg13g2_fill_1 FILLER_24_184 ();
 sg13g2_decap_8 FILLER_24_257 ();
 sg13g2_decap_8 FILLER_24_264 ();
 sg13g2_decap_4 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_fill_2 FILLER_24_287 ();
 sg13g2_decap_4 FILLER_24_299 ();
 sg13g2_fill_1 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_314 ();
 sg13g2_fill_2 FILLER_24_331 ();
 sg13g2_fill_1 FILLER_24_333 ();
 sg13g2_decap_8 FILLER_24_365 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_51 ();
 sg13g2_fill_1 FILLER_25_53 ();
 sg13g2_fill_2 FILLER_25_59 ();
 sg13g2_fill_1 FILLER_25_78 ();
 sg13g2_decap_4 FILLER_25_102 ();
 sg13g2_decap_4 FILLER_25_120 ();
 sg13g2_fill_1 FILLER_25_124 ();
 sg13g2_fill_1 FILLER_25_145 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_192 ();
 sg13g2_fill_1 FILLER_25_198 ();
 sg13g2_fill_2 FILLER_25_207 ();
 sg13g2_fill_1 FILLER_25_209 ();
 sg13g2_fill_1 FILLER_25_283 ();
 sg13g2_decap_8 FILLER_25_325 ();
 sg13g2_fill_2 FILLER_25_377 ();
 sg13g2_fill_1 FILLER_26_44 ();
 sg13g2_fill_1 FILLER_26_80 ();
 sg13g2_decap_4 FILLER_26_106 ();
 sg13g2_decap_8 FILLER_26_116 ();
 sg13g2_fill_2 FILLER_26_123 ();
 sg13g2_fill_1 FILLER_26_125 ();
 sg13g2_decap_8 FILLER_26_156 ();
 sg13g2_decap_8 FILLER_26_163 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_fill_2 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_fill_1 FILLER_26_223 ();
 sg13g2_fill_2 FILLER_26_227 ();
 sg13g2_fill_1 FILLER_26_253 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_fill_2 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_331 ();
 sg13g2_fill_2 FILLER_26_337 ();
 sg13g2_fill_2 FILLER_26_366 ();
 sg13g2_fill_1 FILLER_26_372 ();
 sg13g2_fill_1 FILLER_26_400 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_58 ();
 sg13g2_fill_2 FILLER_27_78 ();
 sg13g2_fill_2 FILLER_27_96 ();
 sg13g2_fill_1 FILLER_27_98 ();
 sg13g2_decap_4 FILLER_27_109 ();
 sg13g2_decap_8 FILLER_27_123 ();
 sg13g2_fill_2 FILLER_27_130 ();
 sg13g2_decap_4 FILLER_27_164 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_fill_2 FILLER_27_191 ();
 sg13g2_fill_1 FILLER_27_193 ();
 sg13g2_decap_4 FILLER_27_213 ();
 sg13g2_fill_2 FILLER_27_217 ();
 sg13g2_fill_2 FILLER_27_224 ();
 sg13g2_fill_1 FILLER_27_249 ();
 sg13g2_fill_2 FILLER_27_285 ();
 sg13g2_fill_1 FILLER_27_287 ();
 sg13g2_decap_4 FILLER_27_298 ();
 sg13g2_fill_2 FILLER_27_380 ();
 sg13g2_fill_1 FILLER_27_382 ();
 sg13g2_decap_4 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_132 ();
 sg13g2_fill_2 FILLER_28_139 ();
 sg13g2_decap_4 FILLER_28_156 ();
 sg13g2_fill_2 FILLER_28_160 ();
 sg13g2_decap_8 FILLER_28_188 ();
 sg13g2_fill_1 FILLER_28_195 ();
 sg13g2_fill_1 FILLER_28_225 ();
 sg13g2_fill_1 FILLER_28_239 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_fill_2 FILLER_28_269 ();
 sg13g2_decap_8 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_283 ();
 sg13g2_fill_1 FILLER_28_285 ();
 sg13g2_fill_1 FILLER_28_295 ();
 sg13g2_fill_1 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_315 ();
 sg13g2_fill_2 FILLER_28_326 ();
 sg13g2_fill_2 FILLER_28_338 ();
 sg13g2_fill_2 FILLER_28_345 ();
 sg13g2_fill_1 FILLER_28_365 ();
 sg13g2_fill_2 FILLER_28_381 ();
 sg13g2_fill_2 FILLER_29_51 ();
 sg13g2_fill_1 FILLER_29_75 ();
 sg13g2_fill_1 FILLER_29_87 ();
 sg13g2_fill_2 FILLER_29_98 ();
 sg13g2_fill_2 FILLER_29_120 ();
 sg13g2_fill_1 FILLER_29_122 ();
 sg13g2_fill_2 FILLER_29_151 ();
 sg13g2_fill_2 FILLER_29_165 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_4 FILLER_29_210 ();
 sg13g2_fill_2 FILLER_29_214 ();
 sg13g2_decap_8 FILLER_29_225 ();
 sg13g2_decap_8 FILLER_29_232 ();
 sg13g2_decap_4 FILLER_29_239 ();
 sg13g2_fill_2 FILLER_29_243 ();
 sg13g2_decap_8 FILLER_29_270 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_47 ();
 sg13g2_fill_1 FILLER_30_49 ();
 sg13g2_fill_1 FILLER_30_115 ();
 sg13g2_fill_2 FILLER_30_134 ();
 sg13g2_decap_4 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_162 ();
 sg13g2_decap_4 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_178 ();
 sg13g2_fill_1 FILLER_30_187 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_fill_2 FILLER_30_214 ();
 sg13g2_fill_1 FILLER_30_216 ();
 sg13g2_decap_4 FILLER_30_236 ();
 sg13g2_decap_4 FILLER_30_253 ();
 sg13g2_fill_1 FILLER_30_257 ();
 sg13g2_fill_2 FILLER_30_316 ();
 sg13g2_fill_2 FILLER_30_361 ();
 sg13g2_fill_2 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_58 ();
 sg13g2_fill_2 FILLER_31_82 ();
 sg13g2_fill_1 FILLER_31_112 ();
 sg13g2_fill_2 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_145 ();
 sg13g2_fill_2 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_214 ();
 sg13g2_fill_2 FILLER_31_219 ();
 sg13g2_decap_8 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_240 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_decap_8 FILLER_31_260 ();
 sg13g2_fill_2 FILLER_31_267 ();
 sg13g2_fill_1 FILLER_31_269 ();
 sg13g2_fill_2 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_290 ();
 sg13g2_fill_1 FILLER_31_292 ();
 sg13g2_fill_2 FILLER_31_307 ();
 sg13g2_fill_1 FILLER_31_309 ();
 sg13g2_fill_1 FILLER_31_327 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_4 ();
 sg13g2_fill_2 FILLER_32_37 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_112 ();
 sg13g2_decap_4 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_144 ();
 sg13g2_decap_4 FILLER_32_149 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_decap_8 FILLER_32_158 ();
 sg13g2_fill_2 FILLER_32_165 ();
 sg13g2_decap_4 FILLER_32_176 ();
 sg13g2_fill_2 FILLER_32_180 ();
 sg13g2_decap_4 FILLER_32_186 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_decap_4 FILLER_32_228 ();
 sg13g2_fill_1 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_375 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_4 FILLER_33_150 ();
 sg13g2_fill_1 FILLER_33_185 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_73 ();
 sg13g2_fill_2 FILLER_34_110 ();
 sg13g2_fill_1 FILLER_34_131 ();
 sg13g2_fill_2 FILLER_34_163 ();
 sg13g2_fill_2 FILLER_34_191 ();
 sg13g2_fill_1 FILLER_34_193 ();
 sg13g2_fill_2 FILLER_34_233 ();
 sg13g2_fill_1 FILLER_34_235 ();
 sg13g2_fill_2 FILLER_34_285 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_293 ();
 sg13g2_fill_2 FILLER_34_299 ();
 sg13g2_fill_1 FILLER_34_327 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_fill_2 FILLER_35_59 ();
 sg13g2_fill_2 FILLER_35_146 ();
 sg13g2_fill_2 FILLER_35_157 ();
 sg13g2_fill_1 FILLER_35_169 ();
 sg13g2_fill_1 FILLER_35_205 ();
 sg13g2_fill_1 FILLER_35_286 ();
 sg13g2_fill_2 FILLER_35_302 ();
 sg13g2_fill_1 FILLER_35_314 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_fill_2 FILLER_36_36 ();
 sg13g2_fill_2 FILLER_36_57 ();
 sg13g2_fill_1 FILLER_36_75 ();
 sg13g2_decap_4 FILLER_36_214 ();
 sg13g2_fill_2 FILLER_36_218 ();
 sg13g2_fill_2 FILLER_36_262 ();
 sg13g2_fill_2 FILLER_36_277 ();
 sg13g2_fill_1 FILLER_36_279 ();
 sg13g2_fill_2 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_297 ();
 sg13g2_fill_2 FILLER_36_309 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_fill_2 FILLER_36_331 ();
 sg13g2_fill_1 FILLER_36_346 ();
 sg13g2_fill_2 FILLER_36_373 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_53 ();
 sg13g2_fill_1 FILLER_37_65 ();
 sg13g2_fill_2 FILLER_37_111 ();
 sg13g2_fill_1 FILLER_37_113 ();
 sg13g2_fill_1 FILLER_37_186 ();
 sg13g2_fill_2 FILLER_37_226 ();
 sg13g2_fill_1 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_286 ();
 sg13g2_fill_2 FILLER_37_297 ();
 sg13g2_fill_1 FILLER_37_304 ();
 sg13g2_fill_2 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_46 ();
 sg13g2_fill_1 FILLER_38_129 ();
 sg13g2_fill_2 FILLER_38_201 ();
 sg13g2_fill_2 FILLER_38_220 ();
 sg13g2_fill_1 FILLER_38_222 ();
 sg13g2_fill_2 FILLER_38_270 ();
 sg13g2_fill_1 FILLER_38_298 ();
 sg13g2_fill_1 FILLER_38_309 ();
 sg13g2_fill_2 FILLER_38_356 ();
 sg13g2_fill_2 FILLER_38_389 ();
 assign uo_out[3] = net16;
 assign uo_out[4] = net17;
 assign uo_out[5] = net18;
 assign uo_out[6] = net19;
 assign uo_out[7] = net20;
endmodule

module tt_um_wokwi_group_8 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire \proj_10.net10 ;
 wire \proj_10.net16 ;
 wire \proj_10.net17 ;
 wire \proj_10.net18 ;
 wire \proj_10.net19 ;
 wire \proj_10.net9 ;
 wire \proj_11.net4 ;
 wire \proj_11.net5 ;
 wire \proj_12.net10 ;
 wire \proj_12.net16 ;
 wire \proj_12.net17 ;
 wire \proj_12.net18 ;
 wire \proj_12.net9 ;
 wire \proj_13.net7 ;
 wire \proj_13.net8 ;
 wire \proj_13.net9 ;
 wire \proj_14.net13 ;
 wire \proj_14.net14 ;
 wire \proj_14.net15 ;
 wire \proj_14.net16 ;
 wire \proj_14.net17 ;
 wire \proj_14.net18 ;
 wire \proj_14.net19 ;
 wire \proj_14.net20 ;
 wire \proj_14.net21 ;
 wire \proj_14.net22 ;
 wire \proj_14.net23 ;
 wire \proj_14.net24 ;
 wire \proj_14.net25 ;
 wire \proj_14.net26 ;
 wire \proj_14.net27 ;
 wire \proj_14.net28 ;
 wire \proj_14.net29 ;
 wire \proj_14.net3 ;
 wire \proj_14.net30 ;
 wire \proj_14.net31 ;
 wire \proj_14.net32 ;
 wire \proj_14.net4 ;
 wire \proj_14.net5 ;
 wire \proj_14.net6 ;
 wire \proj_14.net7 ;
 wire \proj__0.net12 ;
 wire \proj__0.net13 ;
 wire \proj__0.net14 ;
 wire \proj__0.net15 ;
 wire \proj__0.net16 ;
 wire \proj__0.net17 ;
 wire \proj__0.net18 ;
 wire \proj__0.net19 ;
 wire \proj__0.net20 ;
 wire \proj__0.net21 ;
 wire \proj__0.net22 ;
 wire \proj__0.net23 ;
 wire \proj__0.net24 ;
 wire \proj__0.net4 ;
 wire \proj__0.net5 ;
 wire \proj__0.net6 ;
 wire \proj__1.net8 ;
 wire \proj__1.net9 ;
 wire \proj__2.net10 ;
 wire \proj__2.net11 ;
 wire \proj__2.net12 ;
 wire \proj__2.net5 ;
 wire \proj__2.net6 ;
 wire \proj__2.net7 ;
 wire \proj__2.net8 ;
 wire \proj__2.net9 ;
 wire \proj__3.net10 ;
 wire \proj__3.net11 ;
 wire \proj__3.net12 ;
 wire \proj__3.net9 ;
 wire \proj__5.net10 ;
 wire \proj__5.net8 ;
 wire \proj__5.net9 ;
 wire \proj__6.net10 ;
 wire \proj__6.net11 ;
 wire \proj__6.net7 ;
 wire \proj__6.net8 ;
 wire \proj__6.net9 ;
 wire \proj__7.net10 ;
 wire \proj__7.net11 ;
 wire \proj__7.net12 ;
 wire \proj__7.net13 ;
 wire \proj__7.net14 ;
 wire \proj__7.net9 ;
 wire \proj__8.net14 ;
 wire \proj__8.net15 ;
 wire \proj__8.net16 ;
 wire \proj__8.net17 ;
 wire \proj__8.net18 ;
 wire \proj__8.net19 ;
 wire \proj__8.net2 ;
 wire \proj__8.net20 ;
 wire \proj__8.net21 ;
 wire \proj__8.net22 ;
 wire \proj__8.net23 ;
 wire \proj__8.net24 ;
 wire \proj__8.net25 ;
 wire \proj__8.net26 ;
 wire \proj__8.net27 ;
 wire \proj__8.net28 ;
 wire \proj__8.net29 ;
 wire \proj__8.net3 ;
 wire \proj__8.net30 ;
 wire \proj__8.net31 ;
 wire \proj__8.net32 ;
 wire \proj__8.net33 ;
 wire \proj__8.net34 ;
 wire \proj__8.net35 ;
 wire \proj__8.net36 ;
 wire \proj__8.net37 ;
 wire \proj__8.net38 ;
 wire \proj__8.net39 ;
 wire \proj__8.net4 ;
 wire \proj__8.net40 ;
 wire \proj__8.net41 ;
 wire \proj__8.net42 ;
 wire \proj__8.net43 ;
 wire \proj__8.net44 ;
 wire \proj__8.net45 ;
 wire \proj__8.net46 ;
 wire \proj__8.net47 ;
 wire \proj__8.net48 ;
 wire \proj__8.net49 ;
 wire \proj__8.net5 ;
 wire \proj__8.net50 ;
 wire \proj__8.net51 ;
 wire \proj__8.net52 ;
 wire \proj__8.net53 ;
 wire \proj__8.net54 ;
 wire \proj__8.net55 ;
 wire \proj__8.net56 ;
 wire \proj__8.net57 ;
 wire \proj__8.net58 ;
 wire \proj__8.net59 ;
 wire \proj__8.net6 ;
 wire \proj__8.net60 ;
 wire \proj__8.net61 ;
 wire \proj__8.net62 ;
 wire \proj__8.net63 ;
 wire \proj__8.net64 ;
 wire \proj__8.net65 ;
 wire \proj__8.net66 ;
 wire \proj__8.net67 ;
 wire \proj__8.net68 ;
 wire \proj__8.net69 ;
 wire \proj__8.net7 ;
 wire \proj__8.net8 ;
 wire \proj__9.net10 ;
 wire \proj__9.net11 ;
 wire \proj__9.net12 ;
 wire \proj__9.net9 ;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire \proj__2.flop1/_0_ ;
 wire \proj__2.flop1/_1_ ;
 wire net28;
 wire net29;
 wire \proj__2.flop1/notq ;
 wire \proj__2.flop2/_0_ ;
 wire \proj__2.flop2/_1_ ;
 wire net30;
 wire net31;
 wire \proj__2.flop2/notq ;
 wire \proj__2.flop3/_0_ ;
 wire \proj__2.flop3/_1_ ;
 wire net32;
 wire net33;
 wire \proj__2.flop3/notq ;
 wire \proj__2.flop4/_0_ ;
 wire \proj__2.flop4/_1_ ;
 wire net34;
 wire net35;
 wire \proj__2.flop4/notq ;
 wire \proj__2.flop5/_0_ ;
 wire \proj__2.flop5/_1_ ;
 wire net36;
 wire net37;
 wire \proj__2.flop5/notq ;
 wire \proj__2.flop6/_0_ ;
 wire \proj__2.flop6/_1_ ;
 wire net38;
 wire net39;
 wire \proj__2.flop6/notq ;
 wire \proj__2.flop7/_0_ ;
 wire \proj__2.flop7/_1_ ;
 wire net40;
 wire net41;
 wire \proj__2.flop7/notq ;
 wire \proj__2.flop8/_0_ ;
 wire \proj__2.flop8/_1_ ;
 wire net42;
 wire net58;
 wire \proj__2.flop8/notq ;
 wire net64;
 wire net65;
 wire net66;
 wire clknet_0_clk;
 wire \proj__8.flop4/q ;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;

 sg13g2_inv_1 _071_ (.Y(_048_),
    .A(net6));
 sg13g2_inv_1 _072_ (.Y(_049_),
    .A(\proj__0.net5 ));
 sg13g2_inv_1 _073_ (.Y(_050_),
    .A(\proj__0.net6 ));
 sg13g2_nand2_2 _074_ (.Y(_051_),
    .A(net10),
    .B(net9));
 sg13g2_nor3_2 _075_ (.A(net7),
    .B(net8),
    .C(_051_),
    .Y(_052_));
 sg13g2_nand2_2 _076_ (.Y(_053_),
    .A(net7),
    .B(net8));
 sg13g2_nor3_2 _077_ (.A(net10),
    .B(net9),
    .C(_053_),
    .Y(_054_));
 sg13g2_nand2b_2 _078_ (.Y(_055_),
    .B(net7),
    .A_N(net8));
 sg13g2_nor2b_1 _079_ (.A(_055_),
    .B_N(_051_),
    .Y(_056_));
 sg13g2_nand2b_2 _080_ (.Y(_057_),
    .B(net8),
    .A_N(net7));
 sg13g2_nor2_2 _081_ (.A(_051_),
    .B(_057_),
    .Y(_058_));
 sg13g2_nor4_1 _082_ (.A(_052_),
    .B(_054_),
    .C(_056_),
    .D(_058_),
    .Y(_059_));
 sg13g2_nor3_2 _083_ (.A(net10),
    .B(net9),
    .C(_057_),
    .Y(_060_));
 sg13g2_nand2b_2 _084_ (.Y(_061_),
    .B(net10),
    .A_N(net9));
 sg13g2_nor2_1 _085_ (.A(_057_),
    .B(_061_),
    .Y(_062_));
 sg13g2_a22oi_1 _086_ (.Y(_063_),
    .B1(_062_),
    .B2(\proj_10.net10 ),
    .A2(_060_),
    .A1(\proj__2.net12 ));
 sg13g2_o21ai_1 _087_ (.B1(_063_),
    .Y(uo_out[7]),
    .A1(_048_),
    .A2(_059_));
 sg13g2_nor2_2 _088_ (.A(_055_),
    .B(_061_),
    .Y(_064_));
 sg13g2_nor2_2 _089_ (.A(_051_),
    .B(_055_),
    .Y(_065_));
 sg13g2_nand2b_2 _090_ (.Y(_066_),
    .B(net9),
    .A_N(net10));
 sg13g2_nor2_2 _091_ (.A(_057_),
    .B(_066_),
    .Y(_067_));
 sg13g2_nor3_2 _092_ (.A(net7),
    .B(net8),
    .C(_061_),
    .Y(_068_));
 sg13g2_a22oi_1 _093_ (.Y(_069_),
    .B1(_068_),
    .B2(\proj__8.net2 ),
    .A2(_054_),
    .A1(\proj__3.net9 ));
 sg13g2_nor2_2 _094_ (.A(_053_),
    .B(_066_),
    .Y(_070_));
 sg13g2_nor4_2 _095_ (.A(net7),
    .B(net8),
    .C(net10),
    .Y(_000_),
    .D(net9));
 sg13g2_and2_1 _096_ (.A(\proj__0.net4 ),
    .B(_000_),
    .X(_001_));
 sg13g2_nor2_1 _097_ (.A(_053_),
    .B(_061_),
    .Y(_002_));
 sg13g2_a22oi_1 _098_ (.Y(_003_),
    .B1(_064_),
    .B2(\proj__9.net9 ),
    .A2(_062_),
    .A1(\proj_10.net9 ));
 sg13g2_a22oi_1 _099_ (.Y(_004_),
    .B1(_065_),
    .B2(\proj_13.net7 ),
    .A2(_060_),
    .A1(\proj__2.net5 ));
 sg13g2_a22oi_1 _100_ (.Y(_005_),
    .B1(_002_),
    .B2(\proj_11.net4 ),
    .A2(_070_),
    .A1(\proj__7.net9 ));
 sg13g2_a22oi_1 _101_ (.Y(_006_),
    .B1(_067_),
    .B2(\proj__6.net7 ),
    .A2(_058_),
    .A1(\proj_14.net3 ));
 sg13g2_a21oi_1 _102_ (.A1(\proj_12.net9 ),
    .A2(_052_),
    .Y(_007_),
    .B1(_001_));
 sg13g2_and4_1 _103_ (.A(_069_),
    .B(_005_),
    .C(_006_),
    .D(_007_),
    .X(_008_));
 sg13g2_nand3_1 _104_ (.B(_004_),
    .C(_008_),
    .A(_003_),
    .Y(uo_out[0]));
 sg13g2_nor3_2 _105_ (.A(net7),
    .B(net8),
    .C(_066_),
    .Y(_009_));
 sg13g2_a21oi_1 _106_ (.A1(\proj__2.net6 ),
    .A2(_060_),
    .Y(_010_),
    .B1(_001_));
 sg13g2_a22oi_1 _107_ (.Y(_011_),
    .B1(_068_),
    .B2(\proj__8.net3 ),
    .A2(_067_),
    .A1(\proj__6.net8 ));
 sg13g2_a22oi_1 _108_ (.Y(_012_),
    .B1(_002_),
    .B2(\proj_11.net5 ),
    .A2(_064_),
    .A1(net52));
 sg13g2_a22oi_1 _109_ (.Y(_013_),
    .B1(_070_),
    .B2(\proj__7.net10 ),
    .A2(_058_),
    .A1(\proj_14.net4 ));
 sg13g2_a22oi_1 _110_ (.Y(_014_),
    .B1(_065_),
    .B2(\proj_13.net8 ),
    .A2(_052_),
    .A1(\proj_12.net10 ));
 sg13g2_and4_1 _111_ (.A(_010_),
    .B(_012_),
    .C(_013_),
    .D(_014_),
    .X(_015_));
 sg13g2_a22oi_1 _112_ (.Y(_016_),
    .B1(_009_),
    .B2(net6),
    .A2(_054_),
    .A1(\proj__3.net10 ));
 sg13g2_nand3_1 _113_ (.B(_015_),
    .C(_016_),
    .A(_011_),
    .Y(uo_out[1]));
 sg13g2_nor3_2 _114_ (.A(net10),
    .B(net9),
    .C(_055_),
    .Y(_017_));
 sg13g2_a22oi_1 _115_ (.Y(_018_),
    .B1(_017_),
    .B2(\proj__1.net8 ),
    .A2(_060_),
    .A1(\proj__2.net7 ));
 sg13g2_a22oi_1 _116_ (.Y(_019_),
    .B1(_065_),
    .B2(\proj_13.net9 ),
    .A2(_058_),
    .A1(\proj_14.net5 ));
 sg13g2_a21oi_1 _117_ (.A1(\proj__7.net11 ),
    .A2(_070_),
    .Y(_020_),
    .B1(_001_));
 sg13g2_a22oi_1 _118_ (.Y(_021_),
    .B1(_009_),
    .B2(net52),
    .A2(_054_),
    .A1(\proj__3.net11 ));
 sg13g2_a22oi_1 _119_ (.Y(_022_),
    .B1(_068_),
    .B2(\proj__8.net4 ),
    .A2(_064_),
    .A1(\proj__9.net10 ));
 sg13g2_and3_1 _120_ (.X(_023_),
    .A(_020_),
    .B(_021_),
    .C(_022_));
 sg13g2_nand3_1 _121_ (.B(_019_),
    .C(_023_),
    .A(_018_),
    .Y(uo_out[2]));
 sg13g2_and2_1 _122_ (.A(\proj__8.net5 ),
    .B(_068_),
    .X(_024_));
 sg13g2_a221oi_1 _123_ (.B2(\proj__7.net12 ),
    .C1(_024_),
    .B1(_070_),
    .A1(\proj__2.net8 ),
    .Y(_025_),
    .A2(_060_));
 sg13g2_a21oi_1 _124_ (.A1(\proj_14.net3 ),
    .A2(_058_),
    .Y(_026_),
    .B1(_000_));
 sg13g2_o21ai_1 _125_ (.B1(net49),
    .Y(_027_),
    .A1(_052_),
    .A2(_064_));
 sg13g2_a22oi_1 _126_ (.Y(_028_),
    .B1(_017_),
    .B2(\proj__1.net9 ),
    .A2(_054_),
    .A1(\proj__3.net12 ));
 sg13g2_nor2_2 _127_ (.A(_055_),
    .B(_066_),
    .Y(_029_));
 sg13g2_a22oi_1 _128_ (.Y(_030_),
    .B1(_029_),
    .B2(\proj__5.net8 ),
    .A2(_067_),
    .A1(\proj__6.net9 ));
 sg13g2_and4_1 _129_ (.A(_026_),
    .B(_027_),
    .C(_028_),
    .D(_030_),
    .X(_031_));
 sg13g2_a22oi_1 _130_ (.Y(uo_out[3]),
    .B1(_025_),
    .B2(_031_),
    .A2(_000_),
    .A1(_049_));
 sg13g2_or3_1 _131_ (.A(_052_),
    .B(_054_),
    .C(_017_),
    .X(_032_));
 sg13g2_a22oi_1 _132_ (.Y(_033_),
    .B1(_009_),
    .B2(net50),
    .A2(_064_),
    .A1(\proj__9.net11 ));
 sg13g2_a22oi_1 _133_ (.Y(_034_),
    .B1(_029_),
    .B2(\proj__5.net9 ),
    .A2(_068_),
    .A1(\proj__8.net6 ));
 sg13g2_a21oi_1 _134_ (.A1(\proj_14.net6 ),
    .A2(_058_),
    .Y(_035_),
    .B1(_001_));
 sg13g2_a22oi_1 _135_ (.Y(_036_),
    .B1(_070_),
    .B2(\proj__7.net13 ),
    .A2(_060_),
    .A1(\proj__2.net9 ));
 sg13g2_nand4_1 _136_ (.B(_034_),
    .C(_035_),
    .A(_033_),
    .Y(_037_),
    .D(_036_));
 sg13g2_a21o_1 _137_ (.A2(_032_),
    .A1(net48),
    .B1(_037_),
    .X(uo_out[4]));
 sg13g2_o21ai_1 _138_ (.B1(net4),
    .Y(_038_),
    .A1(_064_),
    .A2(_032_));
 sg13g2_a22oi_1 _139_ (.Y(_039_),
    .B1(_067_),
    .B2(\proj__6.net10 ),
    .A2(_060_),
    .A1(\proj__2.net10 ));
 sg13g2_nand2_1 _140_ (.Y(_040_),
    .A(\proj__7.net14 ),
    .B(_070_));
 sg13g2_a22oi_1 _141_ (.Y(_041_),
    .B1(_009_),
    .B2(net49),
    .A2(_068_),
    .A1(\proj__8.net7 ));
 sg13g2_and4_1 _142_ (.A(_026_),
    .B(_039_),
    .C(_040_),
    .D(_041_),
    .X(_042_));
 sg13g2_a22oi_1 _143_ (.Y(uo_out[5]),
    .B1(_038_),
    .B2(_042_),
    .A2(_000_),
    .A1(_050_));
 sg13g2_nand2_1 _144_ (.Y(_043_),
    .A(net5),
    .B(_032_));
 sg13g2_a22oi_1 _145_ (.Y(_044_),
    .B1(_067_),
    .B2(\proj__6.net11 ),
    .A2(_064_),
    .A1(\proj__9.net12 ));
 sg13g2_and2_1 _146_ (.A(\proj__5.net10 ),
    .B(_029_),
    .X(_045_));
 sg13g2_a22oi_1 _147_ (.Y(_046_),
    .B1(_068_),
    .B2(\proj__8.net8 ),
    .A2(_060_),
    .A1(\proj__2.net11 ));
 sg13g2_a221oi_1 _148_ (.B2(net48),
    .C1(_045_),
    .B1(_009_),
    .A1(\proj_14.net7 ),
    .Y(_047_),
    .A2(_058_));
 sg13g2_nand4_1 _149_ (.B(_044_),
    .C(_046_),
    .A(_043_),
    .Y(uo_out[6]),
    .D(_047_));
 sg13g2_tielo tt_um_wokwi_group_8_12 (.L_LO(net12));
 sg13g2_tielo tt_um_wokwi_group_8_13 (.L_LO(net13));
 sg13g2_tielo tt_um_wokwi_group_8_14 (.L_LO(net14));
 sg13g2_tielo tt_um_wokwi_group_8_15 (.L_LO(net15));
 sg13g2_tielo tt_um_wokwi_group_8_16 (.L_LO(net16));
 sg13g2_tielo tt_um_wokwi_group_8_17 (.L_LO(net17));
 sg13g2_tielo tt_um_wokwi_group_8_18 (.L_LO(net18));
 sg13g2_tielo tt_um_wokwi_group_8_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wokwi_group_8_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wokwi_group_8_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wokwi_group_8_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wokwi_group_8_23 (.L_LO(net23));
 sg13g2_tielo tt_um_wokwi_group_8_24 (.L_LO(net24));
 sg13g2_tielo tt_um_wokwi_group_8_25 (.L_LO(net25));
 sg13g2_tielo tt_um_wokwi_group_8_26 (.L_LO(net26));
 sg13g2_tielo \proj__2.flop1/dffsr_27  (.L_LO(net27));
 sg13g2_and2_1 \proj_10.and1/_0_  (.A(\proj_10.net16 ),
    .B(net53),
    .X(\proj_10.net9 ));
 sg13g2_and2_1 \proj_10.and2/_0_  (.A(net4),
    .B(net3),
    .X(\proj_10.net16 ));
 sg13g2_or2_1 \proj_10.or1/_0_  (.X(\proj_10.net17 ),
    .B(net5),
    .A(net6));
 sg13g2_or2_1 \proj_10.or3/_0_  (.X(\proj_10.net18 ),
    .B(net51),
    .A(net49));
 sg13g2_or2_1 \proj_10.or5/_0_  (.X(\proj_10.net19 ),
    .B(\proj_10.net18 ),
    .A(\proj_10.net17 ));
 sg13g2_or2_1 \proj_10.or6/_0_  (.X(\proj_10.net10 ),
    .B(net56),
    .A(\proj_10.net19 ));
 sg13g2_and2_1 \proj_11.and1/_0_  (.A(net53),
    .B(net56),
    .X(\proj_11.net4 ));
 sg13g2_inv_1 \proj_11.not1/_0_  (.Y(\proj_11.net5 ),
    .A(net51));
 sg13g2_and2_1 \proj_12.and1/_0_  (.A(net53),
    .B(net56),
    .X(\proj_12.net17 ));
 sg13g2_and2_1 \proj_12.and2/_0_  (.A(\proj_12.net16 ),
    .B(net50),
    .X(\proj_12.net18 ));
 sg13g2_or2_1 \proj_12.or1/_0_  (.X(\proj_12.net10 ),
    .B(\proj_12.net18 ),
    .A(\proj_12.net17 ));
 sg13g2_xor2_1 \proj_12.xor1/_0_  (.B(net56),
    .A(net52),
    .X(\proj_12.net16 ));
 sg13g2_xor2_1 \proj_12.xor2/_0_  (.B(\proj_12.net16 ),
    .A(net51),
    .X(\proj_12.net9 ));
 sg13g2_and2_1 \proj_13.and1/_0_  (.A(net53),
    .B(net56),
    .X(\proj_13.net7 ));
 sg13g2_or2_1 \proj_13.or1/_0_  (.X(\proj_13.net9 ),
    .B(net51),
    .A(net2));
 sg13g2_xor2_1 \proj_13.xor1/_0_  (.B(net48),
    .A(net4),
    .X(\proj_13.net8 ));
 sg13g2_and2_1 \proj_14.and1/_0_  (.A(\proj_14.net14 ),
    .B(\proj_14.net20 ),
    .X(\proj_14.net21 ));
 sg13g2_and2_1 \proj_14.and10/_0_  (.A(\proj_14.net15 ),
    .B(\proj_14.net19 ),
    .X(\proj_14.net30 ));
 sg13g2_and2_1 \proj_14.and11/_0_  (.A(\proj_14.net17 ),
    .B(\proj_14.net30 ),
    .X(\proj_14.net31 ));
 sg13g2_and2_1 \proj_14.and2/_0_  (.A(\proj_14.net19 ),
    .B(\proj_14.net15 ),
    .X(\proj_14.net22 ));
 sg13g2_and2_1 \proj_14.and3/_0_  (.A(\proj_14.net22 ),
    .B(\proj_14.net18 ),
    .X(\proj_14.net23 ));
 sg13g2_and2_1 \proj_14.and4/_0_  (.A(\proj_14.net20 ),
    .B(\proj_14.net24 ),
    .X(\proj_14.net25 ));
 sg13g2_and2_1 \proj_14.and5/_0_  (.A(\proj_14.net14 ),
    .B(\proj_14.net18 ),
    .X(\proj_14.net24 ));
 sg13g2_and2_1 \proj_14.and6/_0_  (.A(\proj_14.net20 ),
    .B(\proj_14.net26 ),
    .X(\proj_14.net27 ));
 sg13g2_and2_1 \proj_14.and7/_0_  (.A(\proj_14.net15 ),
    .B(\proj_14.net18 ),
    .X(\proj_14.net26 ));
 sg13g2_and2_1 \proj_14.and8/_0_  (.A(\proj_14.net14 ),
    .B(\proj_14.net18 ),
    .X(\proj_14.net28 ));
 sg13g2_and2_1 \proj_14.and9/_0_  (.A(\proj_14.net19 ),
    .B(\proj_14.net28 ),
    .X(\proj_14.net29 ));
 sg13g2_dfrbp_1 \proj_14.flop1/_1_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net58),
    .D(net73),
    .Q_N(\proj_14.net15 ),
    .Q(\proj_14.net14 ));
 sg13g2_tiehi \proj_14.flop2/_1__44  (.L_HI(net59));
 sg13g2_dfrbp_1 \proj_14.flop2/_1_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net59),
    .D(net70),
    .Q_N(\proj_14.net18 ),
    .Q(\proj_14.net17 ));
 sg13g2_tiehi \proj_14.flop3/_1__45  (.L_HI(net60));
 sg13g2_dfrbp_1 \proj_14.flop3/_1_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net60),
    .D(net68),
    .Q_N(\proj_14.net19 ),
    .Q(\proj_14.net20 ));
 sg13g2_tiehi \proj__0.flop1/_1__46  (.L_HI(net61));
 sg13g2_or2_1 \proj_14.or1/_0_  (.X(\proj_14.net4 ),
    .B(\proj_14.net27 ),
    .A(\proj_14.net25 ));
 sg13g2_or2_1 \proj_14.or2/_0_  (.X(\proj_14.net3 ),
    .B(\proj_14.net23 ),
    .A(\proj_14.net4 ));
 sg13g2_or2_1 \proj_14.or3/_0_  (.X(\proj_14.net5 ),
    .B(\proj_14.net4 ),
    .A(\proj_14.net29 ));
 sg13g2_or2_1 \proj_14.or4/_0_  (.X(\proj_14.net32 ),
    .B(\proj_14.net23 ),
    .A(\proj_14.net4 ));
 sg13g2_or2_1 \proj_14.or5/_0_  (.X(\proj_14.net7 ),
    .B(\proj_14.net29 ),
    .A(\proj_14.net31 ));
 sg13g2_or2_1 \proj_14.or6/_0_  (.X(\proj_14.net6 ),
    .B(\proj_14.net32 ),
    .A(\proj_14.net7 ));
 sg13g2_xor2_1 \proj_14.xor1/_0_  (.B(net72),
    .A(\proj_14.net20 ),
    .X(\proj_14.net13 ));
 sg13g2_xor2_1 \proj_14.xor2/_0_  (.B(net69),
    .A(\proj_14.net21 ),
    .X(\proj_14.net16 ));
 sg13g2_and2_1 \proj__0.and1/_0_  (.A(\proj__0.net12 ),
    .B(net57),
    .X(\proj__0.net13 ));
 sg13g2_and2_1 \proj__0.and2/_0_  (.A(net52),
    .B(\proj__0.net12 ),
    .X(\proj__0.net14 ));
 sg13g2_and2_1 \proj__0.and3/_0_  (.A(\proj__0.net17 ),
    .B(\proj__0.net16 ),
    .X(\proj__0.net20 ));
 sg13g2_and2_1 \proj__0.and4/_0_  (.A(\proj__0.net15 ),
    .B(\proj__0.net18 ),
    .X(\proj__0.net21 ));
 sg13g2_and2_1 \proj__0.and5/_0_  (.A(\proj__0.net16 ),
    .B(\proj__0.net18 ),
    .X(\proj__0.net23 ));
 sg13g2_dfrbp_1 \proj__0.flop1/_1_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net61),
    .D(net67),
    .Q_N(\proj__0.net15 ),
    .Q(\proj__0.net16 ));
 sg13g2_tiehi \proj__0.flop2/_1__47  (.L_HI(net62));
 sg13g2_dfrbp_1 \proj__0.flop2/_1_  (.CLK(\proj__0.net15 ),
    .RESET_B(net62),
    .D(\proj__0.net17 ),
    .Q_N(\proj__0.net17 ),
    .Q(\proj__0.net18 ));
 sg13g2_tiehi \proj__8.flop1/_1__48  (.L_HI(net63));
 sg13g2_mux2_1 \proj__0.mux1/_0_  (.A0(\proj__0.net24 ),
    .A1(\proj__0.net14 ),
    .S(\proj__0.net12 ),
    .X(\proj__0.net6 ));
 sg13g2_mux2_1 \proj__0.mux2/_0_  (.A0(\proj__0.net22 ),
    .A1(\proj__0.net13 ),
    .S(\proj__0.net12 ),
    .X(\proj__0.net5 ));
 sg13g2_mux2_1 \proj__0.mux3/_0_  (.A0(\proj__0.net19 ),
    .A1(\proj__0.net12 ),
    .S(\proj__0.net12 ),
    .X(\proj__0.net4 ));
 sg13g2_or2_1 \proj__0.or1/_0_  (.X(\proj__0.net19 ),
    .B(\proj__0.net16 ),
    .A(\proj__0.net18 ));
 sg13g2_or2_2 \proj__0.or4/_0_  (.X(\proj__0.net12 ),
    .B(net57),
    .A(net52));
 sg13g2_xor2_1 \proj__0.xor4/_0_  (.B(\proj__0.net20 ),
    .A(\proj__0.net21 ),
    .X(\proj__0.net22 ));
 sg13g2_xor2_1 \proj__0.xor5/_0_  (.B(\proj__0.net21 ),
    .A(\proj__0.net23 ),
    .X(\proj__0.net24 ));
 sg13g2_inv_1 \proj__1.not3/_0_  (.Y(\proj__1.net8 ),
    .A(net50));
 sg13g2_inv_1 \proj__1.not4/_0_  (.Y(\proj__1.net9 ),
    .A(net49));
 sg13g2_inv_1 \proj__2.flop1/_4_  (.Y(\proj__2.flop1/_0_ ),
    .A(net1));
 sg13g2_inv_1 \proj__2.flop1/_5_  (.Y(\proj__2.flop1/_1_ ),
    .A(net53));
 sg13g2_tielo \proj__2.flop1/dffsr_28  (.L_LO(net28));
 sg13g2_tielo \proj__2.flop2/dffsr_29  (.L_LO(net29));
 sg13g2_sdfbbp_1 \proj__2.flop1/dffsr  (.Q(\proj__2.net5 ),
    .Q_N(\proj__2.flop1/notq ),
    .RESET_B(\proj__2.flop1/_0_ ),
    .SET_B(\proj__2.flop1/_1_ ),
    .D(net57),
    .SCE(net28),
    .SCD(net27),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_inv_1 \proj__2.flop2/_4_  (.Y(\proj__2.flop2/_0_ ),
    .A(net1));
 sg13g2_inv_1 \proj__2.flop2/_5_  (.Y(\proj__2.flop2/_1_ ),
    .A(net54));
 sg13g2_tielo \proj__2.flop2/dffsr_30  (.L_LO(net30));
 sg13g2_tielo \proj__2.flop3/dffsr_31  (.L_LO(net31));
 sg13g2_sdfbbp_1 \proj__2.flop2/dffsr  (.Q(\proj__2.net6 ),
    .Q_N(\proj__2.flop2/notq ),
    .RESET_B(\proj__2.flop2/_0_ ),
    .SET_B(\proj__2.flop2/_1_ ),
    .D(net75),
    .SCE(net30),
    .SCD(net29),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_inv_1 \proj__2.flop3/_4_  (.Y(\proj__2.flop3/_0_ ),
    .A(net1));
 sg13g2_inv_1 \proj__2.flop3/_5_  (.Y(\proj__2.flop3/_1_ ),
    .A(net54));
 sg13g2_tielo \proj__2.flop3/dffsr_32  (.L_LO(net32));
 sg13g2_tielo \proj__2.flop4/dffsr_33  (.L_LO(net33));
 sg13g2_sdfbbp_1 \proj__2.flop3/dffsr  (.Q(\proj__2.net7 ),
    .Q_N(\proj__2.flop3/notq ),
    .RESET_B(\proj__2.flop3/_0_ ),
    .SET_B(\proj__2.flop3/_1_ ),
    .D(net80),
    .SCE(net32),
    .SCD(net31),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_inv_1 \proj__2.flop4/_4_  (.Y(\proj__2.flop4/_0_ ),
    .A(net1));
 sg13g2_inv_1 \proj__2.flop4/_5_  (.Y(\proj__2.flop4/_1_ ),
    .A(net54));
 sg13g2_tielo \proj__2.flop4/dffsr_34  (.L_LO(net34));
 sg13g2_tielo \proj__2.flop5/dffsr_35  (.L_LO(net35));
 sg13g2_sdfbbp_1 \proj__2.flop4/dffsr  (.Q(\proj__2.net8 ),
    .Q_N(\proj__2.flop4/notq ),
    .RESET_B(\proj__2.flop4/_0_ ),
    .SET_B(\proj__2.flop4/_1_ ),
    .D(net78),
    .SCE(net34),
    .SCD(net33),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_inv_1 \proj__2.flop5/_4_  (.Y(\proj__2.flop5/_0_ ),
    .A(net1));
 sg13g2_inv_1 \proj__2.flop5/_5_  (.Y(\proj__2.flop5/_1_ ),
    .A(net54));
 sg13g2_tielo \proj__2.flop5/dffsr_36  (.L_LO(net36));
 sg13g2_tielo \proj__2.flop6/dffsr_37  (.L_LO(net37));
 sg13g2_sdfbbp_1 \proj__2.flop5/dffsr  (.Q(\proj__2.net9 ),
    .Q_N(\proj__2.flop5/notq ),
    .RESET_B(\proj__2.flop5/_0_ ),
    .SET_B(\proj__2.flop5/_1_ ),
    .D(net79),
    .SCE(net36),
    .SCD(net35),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_inv_1 \proj__2.flop6/_4_  (.Y(\proj__2.flop6/_0_ ),
    .A(net1));
 sg13g2_inv_1 \proj__2.flop6/_5_  (.Y(\proj__2.flop6/_1_ ),
    .A(net54));
 sg13g2_tielo \proj__2.flop6/dffsr_38  (.L_LO(net38));
 sg13g2_tielo \proj__2.flop7/dffsr_39  (.L_LO(net39));
 sg13g2_sdfbbp_1 \proj__2.flop6/dffsr  (.Q(\proj__2.net10 ),
    .Q_N(\proj__2.flop6/notq ),
    .RESET_B(\proj__2.flop6/_0_ ),
    .SET_B(\proj__2.flop6/_1_ ),
    .D(net76),
    .SCE(net38),
    .SCD(net37),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_inv_1 \proj__2.flop7/_4_  (.Y(\proj__2.flop7/_0_ ),
    .A(net1));
 sg13g2_inv_1 \proj__2.flop7/_5_  (.Y(\proj__2.flop7/_1_ ),
    .A(net53));
 sg13g2_tielo \proj__2.flop7/dffsr_40  (.L_LO(net40));
 sg13g2_tielo \proj__2.flop8/dffsr_41  (.L_LO(net41));
 sg13g2_sdfbbp_1 \proj__2.flop7/dffsr  (.Q(\proj__2.net11 ),
    .Q_N(\proj__2.flop7/notq ),
    .RESET_B(\proj__2.flop7/_0_ ),
    .SET_B(\proj__2.flop7/_1_ ),
    .D(net74),
    .SCE(net40),
    .SCD(net39),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_inv_1 \proj__2.flop8/_4_  (.Y(\proj__2.flop8/_0_ ),
    .A(net1));
 sg13g2_inv_1 \proj__2.flop8/_5_  (.Y(\proj__2.flop8/_1_ ),
    .A(net53));
 sg13g2_tielo \proj__2.flop8/dffsr_42  (.L_LO(net42));
 sg13g2_tiehi \proj_14.flop1/_1__43  (.L_HI(net58));
 sg13g2_sdfbbp_1 \proj__2.flop8/dffsr  (.Q(\proj__2.net12 ),
    .Q_N(\proj__2.flop8/notq ),
    .RESET_B(\proj__2.flop8/_0_ ),
    .SET_B(\proj__2.flop8/_1_ ),
    .D(net77),
    .SCE(net42),
    .SCD(net41),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_inv_1 \proj__3.not1/_0_  (.Y(\proj__3.net9 ),
    .A(net57));
 sg13g2_inv_1 \proj__3.not2/_0_  (.Y(\proj__3.net10 ),
    .A(net52));
 sg13g2_inv_1 \proj__3.not3/_0_  (.Y(\proj__3.net11 ),
    .A(net50));
 sg13g2_inv_1 \proj__3.not4/_0_  (.Y(\proj__3.net12 ),
    .A(net49));
 sg13g2_and2_1 \proj__5.and1/_0_  (.A(net52),
    .B(net57),
    .X(\proj__5.net10 ));
 sg13g2_or2_1 \proj__5.or1/_0_  (.X(\proj__5.net9 ),
    .B(net48),
    .A(net4));
 sg13g2_xor2_1 \proj__5.xor1/_0_  (.B(net50),
    .A(net49),
    .X(\proj__5.net8 ));
 sg13g2_and2_1 \proj__6.and1/_0_  (.A(net50),
    .B(net52),
    .X(\proj__6.net8 ));
 sg13g2_and2_1 \proj__6.and2/_0_  (.A(net6),
    .B(net48),
    .X(\proj__6.net11 ));
 sg13g2_inv_1 \proj__6.not1/_0_  (.Y(\proj__6.net7 ),
    .A(net56));
 sg13g2_inv_1 \proj__6.not2/_0_  (.Y(\proj__6.net9 ),
    .A(net49));
 sg13g2_xor2_1 \proj__6.xor1/_0_  (.B(net48),
    .A(net6),
    .X(\proj__6.net10 ));
 sg13g2_inv_1 \proj__7.not1/_0_  (.Y(\proj__7.net12 ),
    .A(net5));
 sg13g2_inv_1 \proj__7.not2/_0_  (.Y(\proj__7.net10 ),
    .A(net50));
 sg13g2_inv_1 \proj__7.not3/_0_  (.Y(\proj__7.net11 ),
    .A(net49));
 sg13g2_inv_1 \proj__7.not4/_0_  (.Y(\proj__7.net13 ),
    .A(net48));
 sg13g2_or2_1 \proj__7.or1/_0_  (.X(\proj__7.net14 ),
    .B(net4),
    .A(net6));
 sg13g2_xor2_1 \proj__7.xor1/_0_  (.B(net56),
    .A(net55),
    .X(\proj__7.net9 ));
 sg13g2_and2_1 \proj__8.and1/_0_  (.A(\proj__8.net22 ),
    .B(net44),
    .X(\proj__8.net25 ));
 sg13g2_and2_1 \proj__8.and10/_0_  (.A(\proj__8.net23 ),
    .B(net43),
    .X(\proj__8.net39 ));
 sg13g2_and2_1 \proj__8.and11/_0_  (.A(\proj__8.net19 ),
    .B(\proj__8.net22 ),
    .X(\proj__8.net40 ));
 sg13g2_and2_1 \proj__8.and12/_0_  (.A(net45),
    .B(net43),
    .X(\proj__8.net41 ));
 sg13g2_and2_1 \proj__8.and13/_0_  (.A(\proj__8.net21 ),
    .B(\proj__8.net22 ),
    .X(\proj__8.net42 ));
 sg13g2_and2_1 \proj__8.and14/_0_  (.A(\proj__8.net44 ),
    .B(\proj__8.net43 ),
    .X(\proj__8.net34 ));
 sg13g2_and2_1 \proj__8.and15/_0_  (.A(\proj__8.net14 ),
    .B(net43),
    .X(\proj__8.net43 ));
 sg13g2_and2_1 \proj__8.and16/_0_  (.A(net47),
    .B(net46),
    .X(\proj__8.net44 ));
 sg13g2_and2_1 \proj__8.and17/_0_  (.A(\proj__8.net46 ),
    .B(\proj__8.net45 ),
    .X(\proj__8.net47 ));
 sg13g2_and2_1 \proj__8.and18/_0_  (.A(net45),
    .B(net44),
    .X(\proj__8.net45 ));
 sg13g2_and2_1 \proj__8.and19/_0_  (.A(\proj__8.net21 ),
    .B(\proj__8.net17 ),
    .X(\proj__8.net46 ));
 sg13g2_and2_1 \proj__8.and2/_0_  (.A(\proj__8.net26 ),
    .B(\proj__8.net25 ),
    .X(\proj__8.net27 ));
 sg13g2_and2_1 \proj__8.and20/_0_  (.A(\proj__8.net49 ),
    .B(\proj__8.net48 ),
    .X(\proj__8.net50 ));
 sg13g2_and2_1 \proj__8.and21/_0_  (.A(\proj__8.net23 ),
    .B(\proj__8.net20 ),
    .X(\proj__8.net48 ));
 sg13g2_and2_1 \proj__8.and22/_0_  (.A(\proj__8.net21 ),
    .B(\proj__8.net22 ),
    .X(\proj__8.net49 ));
 sg13g2_and2_1 \proj__8.and23/_0_  (.A(\proj__8.net21 ),
    .B(\proj__8.net51 ),
    .X(\proj__8.net52 ));
 sg13g2_and2_1 \proj__8.and24/_0_  (.A(\proj__8.net23 ),
    .B(net44),
    .X(\proj__8.net51 ));
 sg13g2_and2_1 \proj__8.and25/_0_  (.A(\proj__8.net55 ),
    .B(\proj__8.net54 ),
    .X(\proj__8.net56 ));
 sg13g2_and2_1 \proj__8.and26/_0_  (.A(\proj__8.net23 ),
    .B(net43),
    .X(\proj__8.net54 ));
 sg13g2_and2_1 \proj__8.and27/_0_  (.A(net47),
    .B(\proj__8.net22 ),
    .X(\proj__8.net55 ));
 sg13g2_and2_1 \proj__8.and28/_0_  (.A(\proj__8.net58 ),
    .B(\proj__8.net57 ),
    .X(\proj__8.net59 ));
 sg13g2_and2_1 \proj__8.and29/_0_  (.A(net45),
    .B(net43),
    .X(\proj__8.net57 ));
 sg13g2_and2_1 \proj__8.and3/_0_  (.A(net45),
    .B(net43),
    .X(\proj__8.net28 ));
 sg13g2_and2_1 \proj__8.and30/_0_  (.A(net47),
    .B(net46),
    .X(\proj__8.net58 ));
 sg13g2_and2_1 \proj__8.and31/_0_  (.A(net46),
    .B(\proj__8.net60 ),
    .X(\proj__8.net61 ));
 sg13g2_and2_1 \proj__8.and32/_0_  (.A(\proj__8.net23 ),
    .B(net43),
    .X(\proj__8.net60 ));
 sg13g2_and2_1 \proj__8.and33/_0_  (.A(\proj__8.net22 ),
    .B(\proj__8.net64 ),
    .X(\proj__8.net65 ));
 sg13g2_and2_1 \proj__8.and34/_0_  (.A(\proj__8.net23 ),
    .B(net43),
    .X(\proj__8.net64 ));
 sg13g2_and2_1 \proj__8.and35/_0_  (.A(\proj__8.net67 ),
    .B(\proj__8.net66 ),
    .X(\proj__8.net68 ));
 sg13g2_and2_1 \proj__8.and36/_0_  (.A(net45),
    .B(net44),
    .X(\proj__8.net66 ));
 sg13g2_and2_1 \proj__8.and37/_0_  (.A(net47),
    .B(net46),
    .X(\proj__8.net67 ));
 sg13g2_and2_1 \proj__8.and4/_0_  (.A(\proj__8.net29 ),
    .B(\proj__8.net28 ),
    .X(\proj__8.net30 ));
 sg13g2_and2_1 \proj__8.and5/_0_  (.A(\proj__8.net23 ),
    .B(net44),
    .X(\proj__8.net31 ));
 sg13g2_and2_1 \proj__8.and6/_0_  (.A(\proj__8.net21 ),
    .B(net46),
    .X(\proj__8.net32 ));
 sg13g2_and2_1 \proj__8.and7/_0_  (.A(\proj__8.net32 ),
    .B(\proj__8.net31 ),
    .X(\proj__8.net33 ));
 sg13g2_and2_1 \proj__8.and8/_0_  (.A(\proj__8.net40 ),
    .B(\proj__8.net39 ),
    .X(\proj__8.net37 ));
 sg13g2_and2_1 \proj__8.and9/_0_  (.A(\proj__8.net42 ),
    .B(\proj__8.net41 ),
    .X(\proj__8.net38 ));
 sg13g2_dfrbp_1 \proj__8.flop1/_1_  (.CLK(\proj__8.net15 ),
    .RESET_B(net63),
    .D(net45),
    .Q_N(\proj__8.net14 ),
    .Q(\proj__8.net16 ));
 sg13g2_tiehi \proj__8.flop2/_1__49  (.L_HI(net64));
 sg13g2_dfrbp_1 \proj__8.flop2/_1_  (.CLK(\proj__8.net18 ),
    .RESET_B(net64),
    .D(net46),
    .Q_N(\proj__8.net17 ),
    .Q(\proj__8.net15 ));
 sg13g2_tiehi \proj__8.flop3/_1__50  (.L_HI(net65));
 sg13g2_dfrbp_1 \proj__8.flop3/_1_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net65),
    .D(net47),
    .Q_N(\proj__8.net19 ),
    .Q(\proj__8.net18 ));
 sg13g2_tiehi \proj__8.flop4/_1__51  (.L_HI(net66));
 sg13g2_dfrbp_1 \proj__8.flop4/_1_  (.CLK(\proj__8.net16 ),
    .RESET_B(net66),
    .D(\proj__8.net20 ),
    .Q_N(\proj__8.net20 ),
    .Q(\proj__8.flop4/q ));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_inv_1 \proj__8.not1/_0_  (.Y(\proj__8.net21 ),
    .A(net47));
 sg13g2_inv_1 \proj__8.not10/_0_  (.Y(\proj__8.net8 ),
    .A(\proj__8.net69 ));
 sg13g2_inv_2 \proj__8.not2/_0_  (.Y(\proj__8.net22 ),
    .A(net46));
 sg13g2_inv_2 \proj__8.not3/_0_  (.Y(\proj__8.net23 ),
    .A(net45));
 sg13g2_inv_1 \proj__8.not4/_0_  (.Y(\proj__8.net24 ),
    .A(\proj__8.net20 ));
 sg13g2_inv_1 \proj__8.not5/_0_  (.Y(\proj__8.net2 ),
    .A(\proj__8.net27 ));
 sg13g2_inv_1 \proj__8.not6/_0_  (.Y(\proj__8.net3 ),
    .A(\proj__8.net30 ));
 sg13g2_inv_1 \proj__8.not7/_0_  (.Y(\proj__8.net4 ),
    .A(\proj__8.net33 ));
 sg13g2_inv_1 \proj__8.not8/_0_  (.Y(\proj__8.net5 ),
    .A(\proj__8.net36 ));
 sg13g2_inv_1 \proj__8.not9/_0_  (.Y(\proj__8.net7 ),
    .A(\proj__8.net63 ));
 sg13g2_or2_1 \proj__8.or1/_0_  (.X(\proj__8.net36 ),
    .B(\proj__8.net34 ),
    .A(\proj__8.net35 ));
 sg13g2_or2_1 \proj__8.or2/_0_  (.X(\proj__8.net35 ),
    .B(\proj__8.net37 ),
    .A(\proj__8.net38 ));
 sg13g2_or2_1 \proj__8.or3/_0_  (.X(\proj__8.net53 ),
    .B(\proj__8.net47 ),
    .A(\proj__8.net50 ));
 sg13g2_or2_1 \proj__8.or4/_0_  (.X(\proj__8.net6 ),
    .B(\proj__8.net53 ),
    .A(\proj__8.net52 ));
 sg13g2_or2_1 \proj__8.or5/_0_  (.X(\proj__8.net62 ),
    .B(\proj__8.net56 ),
    .A(\proj__8.net59 ));
 sg13g2_or2_1 \proj__8.or6/_0_  (.X(\proj__8.net63 ),
    .B(\proj__8.net62 ),
    .A(\proj__8.net61 ));
 sg13g2_or2_1 \proj__8.or7/_0_  (.X(\proj__8.net69 ),
    .B(\proj__8.net65 ),
    .A(\proj__8.net68 ));
 sg13g2_xor2_1 \proj__8.xor2/_0_  (.B(net45),
    .A(net47),
    .X(\proj__8.net26 ));
 sg13g2_xor2_1 \proj__8.xor3/_0_  (.B(net46),
    .A(net47),
    .X(\proj__8.net29 ));
 sg13g2_and2_1 \proj__9.and1/_0_  (.A(net53),
    .B(net56),
    .X(\proj__9.net9 ));
 sg13g2_inv_1 \proj__9.not1/_0_  (.Y(\proj__9.net10 ),
    .A(net50));
 sg13g2_inv_1 \proj__9.not2/_0_  (.Y(\proj__9.net12 ),
    .A(net5));
 sg13g2_inv_1 \proj__9.not4/_0_  (.Y(\proj__9.net11 ),
    .A(net48));
 sg13g2_buf_2 fanout43 (.A(net44),
    .X(net43));
 sg13g2_buf_1 fanout44 (.A(\proj__8.net24 ),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(\proj__8.net14 ),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(\proj__8.net17 ),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(net71),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(net3),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(net2),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(ui_in[2]),
    .X(net50));
 sg13g2_buf_1 fanout51 (.A(ui_in[2]),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(net55),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(net55),
    .X(net53));
 sg13g2_buf_1 fanout54 (.A(net55),
    .X(net54));
 sg13g2_buf_1 fanout55 (.A(ui_in[1]),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(net57),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(ui_in[0]),
    .X(net57));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_buf_4 input7 (.X(net7),
    .A(uio_in[0]));
 sg13g2_buf_4 input8 (.X(net8),
    .A(uio_in[1]));
 sg13g2_buf_4 input9 (.X(net9),
    .A(uio_in[2]));
 sg13g2_buf_2 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_tielo tt_um_wokwi_group_8_11 (.L_LO(net11));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\proj__0.net15 ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold2 (.A(\proj_14.net19 ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold3 (.A(\proj_14.net17 ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold4 (.A(\proj_14.net16 ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold5 (.A(\proj__8.net19 ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold6 (.A(\proj_14.net14 ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold7 (.A(\proj_14.net13 ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold8 (.A(\proj__2.net10 ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold9 (.A(\proj__2.net5 ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold10 (.A(\proj__2.net9 ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold11 (.A(\proj__2.net11 ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold12 (.A(\proj__2.net7 ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold13 (.A(\proj__2.net8 ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold14 (.A(\proj__2.net6 ),
    .X(net80));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_4 FILLER_23_252 ();
 sg13g2_decap_4 FILLER_23_260 ();
 sg13g2_fill_2 FILLER_23_264 ();
 sg13g2_decap_8 FILLER_23_271 ();
 sg13g2_decap_8 FILLER_23_278 ();
 sg13g2_decap_8 FILLER_23_285 ();
 sg13g2_decap_8 FILLER_23_292 ();
 sg13g2_decap_8 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_306 ();
 sg13g2_decap_8 FILLER_23_313 ();
 sg13g2_decap_8 FILLER_23_320 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_decap_8 FILLER_23_334 ();
 sg13g2_decap_8 FILLER_23_341 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_decap_8 FILLER_23_355 ();
 sg13g2_decap_8 FILLER_23_362 ();
 sg13g2_decap_8 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_376 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_4 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_199 ();
 sg13g2_fill_1 FILLER_24_206 ();
 sg13g2_fill_2 FILLER_24_233 ();
 sg13g2_fill_1 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_272 ();
 sg13g2_decap_4 FILLER_24_290 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_310 ();
 sg13g2_decap_8 FILLER_24_317 ();
 sg13g2_decap_8 FILLER_24_324 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_4 FILLER_25_179 ();
 sg13g2_fill_2 FILLER_25_183 ();
 sg13g2_decap_8 FILLER_25_211 ();
 sg13g2_fill_2 FILLER_25_222 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_decap_4 FILLER_25_277 ();
 sg13g2_decap_8 FILLER_25_307 ();
 sg13g2_decap_8 FILLER_25_314 ();
 sg13g2_decap_8 FILLER_25_321 ();
 sg13g2_decap_8 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_decap_8 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_349 ();
 sg13g2_decap_8 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_fill_2 FILLER_26_154 ();
 sg13g2_decap_4 FILLER_26_160 ();
 sg13g2_decap_4 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_199 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_fill_2 FILLER_26_217 ();
 sg13g2_fill_2 FILLER_26_226 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_decap_8 FILLER_26_246 ();
 sg13g2_fill_2 FILLER_26_253 ();
 sg13g2_decap_8 FILLER_26_285 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_309 ();
 sg13g2_decap_4 FILLER_26_316 ();
 sg13g2_decap_8 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_330 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_decap_8 FILLER_26_344 ();
 sg13g2_decap_4 FILLER_26_351 ();
 sg13g2_fill_1 FILLER_26_355 ();
 sg13g2_decap_8 FILLER_26_359 ();
 sg13g2_decap_8 FILLER_26_366 ();
 sg13g2_decap_8 FILLER_26_373 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_4 FILLER_27_140 ();
 sg13g2_fill_1 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_fill_2 FILLER_27_195 ();
 sg13g2_fill_1 FILLER_27_197 ();
 sg13g2_decap_4 FILLER_27_206 ();
 sg13g2_fill_1 FILLER_27_210 ();
 sg13g2_decap_4 FILLER_27_286 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_297 ();
 sg13g2_decap_8 FILLER_27_375 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_4 FILLER_28_154 ();
 sg13g2_fill_2 FILLER_28_193 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_4 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_243 ();
 sg13g2_decap_8 FILLER_28_250 ();
 sg13g2_decap_4 FILLER_28_257 ();
 sg13g2_fill_1 FILLER_28_261 ();
 sg13g2_fill_2 FILLER_28_266 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_291 ();
 sg13g2_decap_4 FILLER_28_311 ();
 sg13g2_decap_4 FILLER_28_325 ();
 sg13g2_fill_1 FILLER_28_329 ();
 sg13g2_fill_2 FILLER_28_335 ();
 sg13g2_fill_1 FILLER_28_337 ();
 sg13g2_fill_2 FILLER_28_359 ();
 sg13g2_decap_8 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_28_383 ();
 sg13g2_decap_8 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_fill_2 FILLER_29_161 ();
 sg13g2_fill_1 FILLER_29_163 ();
 sg13g2_decap_8 FILLER_29_183 ();
 sg13g2_decap_8 FILLER_29_190 ();
 sg13g2_fill_2 FILLER_29_197 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_fill_2 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_215 ();
 sg13g2_fill_1 FILLER_29_226 ();
 sg13g2_decap_8 FILLER_29_230 ();
 sg13g2_fill_2 FILLER_29_237 ();
 sg13g2_fill_1 FILLER_29_245 ();
 sg13g2_fill_2 FILLER_29_255 ();
 sg13g2_decap_8 FILLER_29_278 ();
 sg13g2_decap_8 FILLER_29_285 ();
 sg13g2_fill_1 FILLER_29_292 ();
 sg13g2_fill_2 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_313 ();
 sg13g2_decap_8 FILLER_29_328 ();
 sg13g2_decap_4 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_fill_2 FILLER_30_161 ();
 sg13g2_fill_2 FILLER_30_188 ();
 sg13g2_decap_8 FILLER_30_218 ();
 sg13g2_fill_2 FILLER_30_225 ();
 sg13g2_fill_1 FILLER_30_227 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_fill_2 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_268 ();
 sg13g2_fill_1 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_318 ();
 sg13g2_fill_2 FILLER_30_326 ();
 sg13g2_fill_1 FILLER_30_328 ();
 sg13g2_decap_8 FILLER_30_383 ();
 sg13g2_decap_8 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_4 FILLER_31_168 ();
 sg13g2_fill_2 FILLER_31_172 ();
 sg13g2_decap_8 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_191 ();
 sg13g2_fill_1 FILLER_31_193 ();
 sg13g2_decap_4 FILLER_31_197 ();
 sg13g2_fill_2 FILLER_31_201 ();
 sg13g2_fill_2 FILLER_31_208 ();
 sg13g2_fill_1 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_fill_2 FILLER_31_231 ();
 sg13g2_fill_1 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_251 ();
 sg13g2_fill_1 FILLER_31_262 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_decap_8 FILLER_31_278 ();
 sg13g2_decap_4 FILLER_31_285 ();
 sg13g2_fill_2 FILLER_31_315 ();
 sg13g2_decap_4 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_339 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_4 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_144 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_4 FILLER_32_182 ();
 sg13g2_fill_1 FILLER_32_186 ();
 sg13g2_decap_8 FILLER_32_197 ();
 sg13g2_decap_8 FILLER_32_204 ();
 sg13g2_fill_1 FILLER_32_211 ();
 sg13g2_decap_8 FILLER_32_222 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_decap_8 FILLER_32_325 ();
 sg13g2_decap_8 FILLER_32_332 ();
 sg13g2_fill_2 FILLER_32_339 ();
 sg13g2_fill_2 FILLER_32_345 ();
 sg13g2_fill_2 FILLER_32_355 ();
 sg13g2_fill_1 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_373 ();
 sg13g2_decap_8 FILLER_32_380 ();
 sg13g2_decap_8 FILLER_32_387 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_4 FILLER_33_147 ();
 sg13g2_decap_4 FILLER_33_186 ();
 sg13g2_decap_4 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_234 ();
 sg13g2_fill_2 FILLER_33_241 ();
 sg13g2_fill_1 FILLER_33_243 ();
 sg13g2_decap_4 FILLER_33_258 ();
 sg13g2_fill_1 FILLER_33_262 ();
 sg13g2_fill_2 FILLER_33_280 ();
 sg13g2_decap_4 FILLER_33_289 ();
 sg13g2_fill_1 FILLER_33_293 ();
 sg13g2_decap_8 FILLER_33_305 ();
 sg13g2_decap_4 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_316 ();
 sg13g2_decap_8 FILLER_33_325 ();
 sg13g2_fill_2 FILLER_33_332 ();
 sg13g2_fill_1 FILLER_33_334 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_fill_2 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_160 ();
 sg13g2_decap_8 FILLER_34_167 ();
 sg13g2_decap_8 FILLER_34_174 ();
 sg13g2_decap_4 FILLER_34_181 ();
 sg13g2_decap_8 FILLER_34_195 ();
 sg13g2_decap_8 FILLER_34_202 ();
 sg13g2_fill_1 FILLER_34_209 ();
 sg13g2_fill_2 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_251 ();
 sg13g2_fill_1 FILLER_34_258 ();
 sg13g2_decap_4 FILLER_34_264 ();
 sg13g2_fill_2 FILLER_34_268 ();
 sg13g2_fill_1 FILLER_34_287 ();
 sg13g2_decap_4 FILLER_34_306 ();
 sg13g2_decap_4 FILLER_34_334 ();
 sg13g2_fill_2 FILLER_34_338 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_fill_2 FILLER_35_238 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_fill_2 FILLER_35_266 ();
 sg13g2_fill_2 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_289 ();
 sg13g2_decap_8 FILLER_35_300 ();
 sg13g2_fill_2 FILLER_35_307 ();
 sg13g2_fill_1 FILLER_35_309 ();
 sg13g2_decap_4 FILLER_35_313 ();
 sg13g2_decap_4 FILLER_35_333 ();
 sg13g2_fill_1 FILLER_35_337 ();
 sg13g2_decap_8 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_380 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_fill_1 FILLER_36_231 ();
 sg13g2_decap_4 FILLER_36_264 ();
 sg13g2_decap_4 FILLER_36_283 ();
 sg13g2_fill_2 FILLER_36_287 ();
 sg13g2_fill_1 FILLER_36_299 ();
 sg13g2_decap_4 FILLER_36_306 ();
 sg13g2_fill_2 FILLER_36_310 ();
 sg13g2_decap_8 FILLER_36_323 ();
 sg13g2_fill_2 FILLER_36_330 ();
 sg13g2_fill_1 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_238 ();
 sg13g2_fill_2 FILLER_37_247 ();
 sg13g2_fill_1 FILLER_37_249 ();
 sg13g2_fill_2 FILLER_37_288 ();
 sg13g2_fill_1 FILLER_37_290 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_fill_2 FILLER_37_336 ();
 sg13g2_fill_1 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_4 FILLER_38_266 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_decap_4 FILLER_38_324 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_decap_4 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_decap_8 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_362 ();
 sg13g2_decap_8 FILLER_38_369 ();
 sg13g2_decap_8 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 assign uio_oe[0] = net11;
 assign uio_oe[1] = net12;
 assign uio_oe[2] = net13;
 assign uio_oe[3] = net14;
 assign uio_oe[4] = net15;
 assign uio_oe[5] = net16;
 assign uio_oe[6] = net17;
 assign uio_oe[7] = net18;
 assign uio_out[0] = net19;
 assign uio_out[1] = net20;
 assign uio_out[2] = net21;
 assign uio_out[3] = net22;
 assign uio_out[4] = net23;
 assign uio_out[5] = net24;
 assign uio_out[6] = net25;
 assign uio_out[7] = net26;
endmodule

module tt_um_rebeccargb_colorbars (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire clknet_0_clk;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;

 sg13g2_inv_2 _0767_ (.Y(_0053_),
    .A(\counter[3] ));
 sg13g2_inv_1 _0768_ (.Y(_0054_),
    .A(\hvsync_gen.vpos[7] ));
 sg13g2_inv_1 _0769_ (.Y(_0055_),
    .A(net59));
 sg13g2_inv_1 _0770_ (.Y(_0056_),
    .A(net165));
 sg13g2_inv_1 _0771_ (.Y(_0057_),
    .A(net166));
 sg13g2_inv_1 _0772_ (.Y(_0058_),
    .A(\hvsync_gen.vpos[2] ));
 sg13g2_inv_1 _0773_ (.Y(_0059_),
    .A(\hvsync_gen.vpos[1] ));
 sg13g2_inv_2 _0774_ (.Y(_0060_),
    .A(net185));
 sg13g2_inv_1 _0775_ (.Y(_0061_),
    .A(\hvsync_gen.hpos[9] ));
 sg13g2_inv_2 _0776_ (.Y(_0062_),
    .A(net168));
 sg13g2_inv_2 _0777_ (.Y(_0063_),
    .A(net178));
 sg13g2_inv_1 _0778_ (.Y(_0064_),
    .A(_0009_));
 sg13g2_inv_2 _0779_ (.Y(_0065_),
    .A(net68));
 sg13g2_inv_1 _0780_ (.Y(_0066_),
    .A(_0012_));
 sg13g2_inv_1 _0781_ (.Y(_0067_),
    .A(_0021_));
 sg13g2_inv_2 _0782_ (.Y(_0068_),
    .A(_0013_));
 sg13g2_inv_1 _0783_ (.Y(_0069_),
    .A(_0019_));
 sg13g2_nor2_1 _0784_ (.A(net166),
    .B(\hvsync_gen.vpos[3] ),
    .Y(_0070_));
 sg13g2_xor2_1 _0785_ (.B(\hvsync_gen.vpos[3] ),
    .A(\hvsync_gen.vpos[4] ),
    .X(_0071_));
 sg13g2_inv_1 _0786_ (.Y(_0072_),
    .A(_0071_));
 sg13g2_xnor2_1 _0787_ (.Y(_0073_),
    .A(_0003_),
    .B(_0070_));
 sg13g2_inv_1 _0788_ (.Y(_0074_),
    .A(_0073_));
 sg13g2_nor3_1 _0789_ (.A(net165),
    .B(\hvsync_gen.vpos[4] ),
    .C(\hvsync_gen.vpos[3] ),
    .Y(_0075_));
 sg13g2_or3_2 _0790_ (.A(net165),
    .B(net166),
    .C(net167),
    .X(_0076_));
 sg13g2_xnor2_1 _0791_ (.Y(_0077_),
    .A(net164),
    .B(_0076_));
 sg13g2_and2_1 _0792_ (.A(\hvsync_gen.vpos[7] ),
    .B(net164),
    .X(_0078_));
 sg13g2_nand2_2 _0793_ (.Y(_0079_),
    .A(\hvsync_gen.vpos[7] ),
    .B(net164));
 sg13g2_nor2_1 _0794_ (.A(_0075_),
    .B(_0079_),
    .Y(_0080_));
 sg13g2_nand2_1 _0795_ (.Y(_0081_),
    .A(_0076_),
    .B(_0078_));
 sg13g2_a21o_1 _0796_ (.A2(_0076_),
    .A1(net164),
    .B1(\hvsync_gen.vpos[7] ),
    .X(_0082_));
 sg13g2_nand2_1 _0797_ (.Y(_0083_),
    .A(_0081_),
    .B(_0082_));
 sg13g2_or2_1 _0798_ (.X(_0084_),
    .B(_0014_),
    .A(\hvsync_gen.vpos[8] ));
 sg13g2_a21oi_2 _0799_ (.B1(_0084_),
    .Y(_0085_),
    .A2(_0078_),
    .A1(_0076_));
 sg13g2_a21o_1 _0800_ (.A2(_0078_),
    .A1(_0076_),
    .B1(_0084_),
    .X(_0086_));
 sg13g2_nor2_1 _0801_ (.A(net162),
    .B(_0086_),
    .Y(_0087_));
 sg13g2_nand2b_2 _0802_ (.Y(_0088_),
    .B(_0085_),
    .A_N(\hvsync_gen.vpos[9] ));
 sg13g2_nand2_1 _0803_ (.Y(_0089_),
    .A(net162),
    .B(_0086_));
 sg13g2_nor3_1 _0804_ (.A(_0055_),
    .B(_0075_),
    .C(_0079_),
    .Y(_0090_));
 sg13g2_a21o_1 _0805_ (.A2(_0085_),
    .A1(net162),
    .B1(_0090_),
    .X(_0091_));
 sg13g2_a221oi_1 _0806_ (.B2(net162),
    .C1(_0090_),
    .B1(_0085_),
    .A1(_0081_),
    .Y(_0092_),
    .A2(_0082_));
 sg13g2_nor2_1 _0807_ (.A(_0089_),
    .B(_0092_),
    .Y(_0093_));
 sg13g2_o21ai_1 _0808_ (.B1(_0088_),
    .Y(_0094_),
    .A1(_0089_),
    .A2(_0092_));
 sg13g2_xor2_1 _0809_ (.B(_0094_),
    .A(_0083_),
    .X(_0095_));
 sg13g2_nand2_1 _0810_ (.Y(_0096_),
    .A(_0077_),
    .B(_0095_));
 sg13g2_nand4_1 _0811_ (.B(\hvsync_gen.vpos[8] ),
    .C(_0080_),
    .A(net162),
    .Y(_0097_),
    .D(_0083_));
 sg13g2_a21o_1 _0812_ (.A2(_0087_),
    .A1(_0083_),
    .B1(_0091_),
    .X(_0098_));
 sg13g2_nand2_1 _0813_ (.Y(_0099_),
    .A(_0097_),
    .B(_0098_));
 sg13g2_a21oi_1 _0814_ (.A1(_0077_),
    .A2(_0095_),
    .Y(_0100_),
    .B1(_0099_));
 sg13g2_o21ai_1 _0815_ (.B1(_0089_),
    .Y(_0101_),
    .A1(_0088_),
    .A2(_0092_));
 sg13g2_nor2b_1 _0816_ (.A(_0093_),
    .B_N(_0101_),
    .Y(_0102_));
 sg13g2_o21ai_1 _0817_ (.B1(_0077_),
    .Y(_0103_),
    .A1(_0100_),
    .A2(_0102_));
 sg13g2_or3_1 _0818_ (.A(_0077_),
    .B(_0100_),
    .C(_0102_),
    .X(_0104_));
 sg13g2_nand2_1 _0819_ (.Y(_0105_),
    .A(_0103_),
    .B(_0104_));
 sg13g2_nand3_1 _0820_ (.B(_0103_),
    .C(_0104_),
    .A(_0074_),
    .Y(_0106_));
 sg13g2_xor2_1 _0821_ (.B(_0103_),
    .A(_0095_),
    .X(_0107_));
 sg13g2_and2_1 _0822_ (.A(_0106_),
    .B(_0107_),
    .X(_0108_));
 sg13g2_a22oi_1 _0823_ (.Y(_0109_),
    .B1(_0102_),
    .B2(_0096_),
    .A2(_0098_),
    .A1(_0097_));
 sg13g2_o21ai_1 _0824_ (.B1(_0088_),
    .Y(_0110_),
    .A1(_0100_),
    .A2(_0109_));
 sg13g2_a21oi_2 _0825_ (.B1(_0110_),
    .Y(_0111_),
    .A2(_0107_),
    .A1(_0106_));
 sg13g2_a21oi_1 _0826_ (.A1(_0106_),
    .A2(_0110_),
    .Y(_0112_),
    .B1(_0107_));
 sg13g2_xnor2_1 _0827_ (.Y(_0113_),
    .A(_0074_),
    .B(_0111_));
 sg13g2_xnor2_1 _0828_ (.Y(_0114_),
    .A(_0073_),
    .B(_0111_));
 sg13g2_o21ai_1 _0829_ (.B1(_0105_),
    .Y(_0115_),
    .A1(_0073_),
    .A2(_0111_));
 sg13g2_nand2b_1 _0830_ (.Y(_0116_),
    .B(_0110_),
    .A_N(_0106_));
 sg13g2_and2_1 _0831_ (.A(_0115_),
    .B(_0116_),
    .X(_0117_));
 sg13g2_a22oi_1 _0832_ (.Y(_0118_),
    .B1(_0115_),
    .B2(_0116_),
    .A2(_0113_),
    .A1(_0071_));
 sg13g2_o21ai_1 _0833_ (.B1(_0088_),
    .Y(_0119_),
    .A1(_0108_),
    .A2(_0112_));
 sg13g2_o21ai_1 _0834_ (.B1(_0071_),
    .Y(_0120_),
    .A1(_0118_),
    .A2(_0119_));
 sg13g2_or3_1 _0835_ (.A(_0071_),
    .B(_0118_),
    .C(_0119_),
    .X(_0121_));
 sg13g2_and2_1 _0836_ (.A(_0120_),
    .B(_0121_),
    .X(_0122_));
 sg13g2_and3_1 _0837_ (.X(_0123_),
    .A(net167),
    .B(_0120_),
    .C(_0121_));
 sg13g2_xnor2_1 _0838_ (.Y(_0124_),
    .A(_0113_),
    .B(_0120_));
 sg13g2_o21ai_1 _0839_ (.B1(_0119_),
    .Y(_0125_),
    .A1(_0072_),
    .A2(_0114_));
 sg13g2_a21o_1 _0840_ (.A2(_0125_),
    .A1(_0117_),
    .B1(_0118_),
    .X(_0126_));
 sg13g2_and2_1 _0841_ (.A(_0088_),
    .B(_0126_),
    .X(_0127_));
 sg13g2_o21ai_1 _0842_ (.B1(_0127_),
    .Y(net157),
    .A1(_0123_),
    .A2(_0124_));
 sg13g2_inv_1 _0843_ (.Y(_0128_),
    .A(uio_out[7]));
 sg13g2_xor2_1 _0844_ (.B(uio_out[7]),
    .A(_0004_),
    .X(_0129_));
 sg13g2_xnor2_1 _0845_ (.Y(_0130_),
    .A(_0004_),
    .B(net157));
 sg13g2_a21o_1 _0846_ (.A2(net157),
    .A1(net167),
    .B1(_0122_),
    .X(_0131_));
 sg13g2_nand2b_1 _0847_ (.Y(_0132_),
    .B(_0123_),
    .A_N(_0127_));
 sg13g2_and2_1 _0848_ (.A(_0131_),
    .B(_0132_),
    .X(_0133_));
 sg13g2_a22oi_1 _0849_ (.Y(_0134_),
    .B1(_0131_),
    .B2(_0132_),
    .A2(_0130_),
    .A1(_0058_));
 sg13g2_nand4_1 _0850_ (.B(_0114_),
    .C(_0120_),
    .A(net167),
    .Y(_0135_),
    .D(_0121_));
 sg13g2_and2_1 _0851_ (.A(_0088_),
    .B(_0135_),
    .X(_0136_));
 sg13g2_o21ai_1 _0852_ (.B1(_0136_),
    .Y(_0137_),
    .A1(_0123_),
    .A2(_0126_));
 sg13g2_nor2_2 _0853_ (.A(_0134_),
    .B(_0137_),
    .Y(_0138_));
 sg13g2_inv_4 _0854_ (.A(_0138_),
    .Y(uio_out[6]));
 sg13g2_o21ai_1 _0855_ (.B1(_0005_),
    .Y(_0139_),
    .A1(_0134_),
    .A2(_0137_));
 sg13g2_xnor2_1 _0856_ (.Y(_0140_),
    .A(_0130_),
    .B(_0139_));
 sg13g2_o21ai_1 _0857_ (.B1(_0058_),
    .Y(_0141_),
    .A1(_0134_),
    .A2(_0137_));
 sg13g2_or3_1 _0858_ (.A(_0058_),
    .B(_0134_),
    .C(_0137_),
    .X(_0142_));
 sg13g2_and3_1 _0859_ (.X(_0143_),
    .A(_0059_),
    .B(_0141_),
    .C(_0142_));
 sg13g2_nor2_1 _0860_ (.A(_0140_),
    .B(_0143_),
    .Y(_0144_));
 sg13g2_o21ai_1 _0861_ (.B1(_0137_),
    .Y(_0145_),
    .A1(\hvsync_gen.vpos[2] ),
    .A2(_0129_));
 sg13g2_a21o_1 _0862_ (.A2(_0145_),
    .A1(_0133_),
    .B1(_0134_),
    .X(_0146_));
 sg13g2_and2_1 _0863_ (.A(_0088_),
    .B(_0146_),
    .X(_0147_));
 sg13g2_nor2b_2 _0864_ (.A(_0144_),
    .B_N(_0147_),
    .Y(_0148_));
 sg13g2_inv_1 _0865_ (.Y(net151),
    .A(_0148_));
 sg13g2_nand2b_1 _0866_ (.Y(_0149_),
    .B(\hvsync_gen.vpos[0] ),
    .A_N(_0006_));
 sg13g2_nor2b_1 _0867_ (.A(\hvsync_gen.vpos[0] ),
    .B_N(_0006_),
    .Y(_0150_));
 sg13g2_a221oi_1 _0868_ (.B2(_0149_),
    .C1(_0150_),
    .B1(net151),
    .A1(_0141_),
    .Y(_0151_),
    .A2(_0142_));
 sg13g2_nand3_1 _0869_ (.B(_0141_),
    .C(_0142_),
    .A(_0006_),
    .Y(_0152_));
 sg13g2_a22oi_1 _0870_ (.Y(_0153_),
    .B1(net151),
    .B2(_0152_),
    .A2(_0146_),
    .A1(_0140_));
 sg13g2_a21oi_1 _0871_ (.A1(_0140_),
    .A2(_0143_),
    .Y(_0154_),
    .B1(_0146_));
 sg13g2_or2_1 _0872_ (.X(_0155_),
    .B(_0154_),
    .A(_0087_));
 sg13g2_nor3_1 _0873_ (.A(_0151_),
    .B(_0153_),
    .C(_0155_),
    .Y(_0156_));
 sg13g2_inv_1 _0874_ (.Y(net147),
    .A(net149));
 sg13g2_xor2_1 _0875_ (.B(net177),
    .A(\counter[4] ),
    .X(_0157_));
 sg13g2_inv_1 _0876_ (.Y(_0158_),
    .A(_0157_));
 sg13g2_xnor2_1 _0877_ (.Y(_0159_),
    .A(\counter[2] ),
    .B(\hvsync_gen.hpos[2] ));
 sg13g2_nor2_1 _0878_ (.A(net159),
    .B(\hvsync_gen.hpos[1] ),
    .Y(_0160_));
 sg13g2_and2_1 _0879_ (.A(\hvsync_gen.hpos[0] ),
    .B(\counter[0] ),
    .X(_0161_));
 sg13g2_a22oi_1 _0880_ (.Y(_0162_),
    .B1(\hvsync_gen.hpos[1] ),
    .B2(net159),
    .A2(\counter[0] ),
    .A1(net181));
 sg13g2_xnor2_1 _0881_ (.Y(_0163_),
    .A(\counter[1] ),
    .B(\hvsync_gen.hpos[1] ));
 sg13g2_or2_1 _0882_ (.X(_0164_),
    .B(_0162_),
    .A(_0160_));
 sg13g2_nor2_1 _0883_ (.A(_0159_),
    .B(_0164_),
    .Y(_0165_));
 sg13g2_or3_1 _0884_ (.A(_0159_),
    .B(_0160_),
    .C(_0162_),
    .X(_0166_));
 sg13g2_a21oi_1 _0885_ (.A1(\counter[2] ),
    .A2(\hvsync_gen.hpos[2] ),
    .Y(_0167_),
    .B1(_0165_));
 sg13g2_a22oi_1 _0886_ (.Y(_0168_),
    .B1(net179),
    .B2(\counter[2] ),
    .A2(net178),
    .A1(\counter[3] ));
 sg13g2_a22oi_1 _0887_ (.Y(_0169_),
    .B1(_0166_),
    .B2(_0168_),
    .A2(_0063_),
    .A1(_0053_));
 sg13g2_a221oi_1 _0888_ (.B2(_0168_),
    .C1(_0158_),
    .B1(_0166_),
    .A1(_0053_),
    .Y(_0170_),
    .A2(_0063_));
 sg13g2_xnor2_1 _0889_ (.Y(_0171_),
    .A(_0157_),
    .B(_0169_));
 sg13g2_nor2_1 _0890_ (.A(net186),
    .B(net175),
    .Y(_0172_));
 sg13g2_a21oi_1 _0891_ (.A1(net186),
    .A2(_0171_),
    .Y(_0173_),
    .B1(_0172_));
 sg13g2_inv_2 _0892_ (.Y(_0174_),
    .A(_0173_));
 sg13g2_or2_1 _0893_ (.X(_0175_),
    .B(net172),
    .A(net185));
 sg13g2_nand2_1 _0894_ (.Y(_0176_),
    .A(\counter[6] ),
    .B(net172));
 sg13g2_xor2_1 _0895_ (.B(net172),
    .A(\counter[6] ),
    .X(_0177_));
 sg13g2_xnor2_1 _0896_ (.Y(_0178_),
    .A(\counter[6] ),
    .B(net172));
 sg13g2_nor2_1 _0897_ (.A(\counter[5] ),
    .B(net174),
    .Y(_0179_));
 sg13g2_or2_1 _0898_ (.X(_0180_),
    .B(net174),
    .A(\counter[5] ));
 sg13g2_a22oi_1 _0899_ (.Y(_0181_),
    .B1(\counter[4] ),
    .B2(net177),
    .A2(net174),
    .A1(\counter[5] ));
 sg13g2_inv_1 _0900_ (.Y(_0182_),
    .A(_0181_));
 sg13g2_a21oi_1 _0901_ (.A1(\counter[4] ),
    .A2(net177),
    .Y(_0183_),
    .B1(_0170_));
 sg13g2_or2_1 _0902_ (.X(_0184_),
    .B(_0181_),
    .A(_0179_));
 sg13g2_o21ai_1 _0903_ (.B1(_0180_),
    .Y(_0185_),
    .A1(_0170_),
    .A2(_0182_));
 sg13g2_xnor2_1 _0904_ (.Y(_0186_),
    .A(_0178_),
    .B(_0185_));
 sg13g2_nand2_1 _0905_ (.Y(_0187_),
    .A(net185),
    .B(_0186_));
 sg13g2_and2_1 _0906_ (.A(_0175_),
    .B(_0187_),
    .X(_0188_));
 sg13g2_inv_1 _0907_ (.Y(_0189_),
    .A(_0188_));
 sg13g2_nor2_1 _0908_ (.A(net185),
    .B(net168),
    .Y(_0190_));
 sg13g2_nand2_1 _0909_ (.Y(_0191_),
    .A(\counter[8] ),
    .B(net168));
 sg13g2_xor2_1 _0910_ (.B(net168),
    .A(\counter[8] ),
    .X(_0192_));
 sg13g2_nor2_1 _0911_ (.A(\counter[7] ),
    .B(net170),
    .Y(_0193_));
 sg13g2_xor2_1 _0912_ (.B(net170),
    .A(\counter[7] ),
    .X(_0194_));
 sg13g2_nand2_1 _0913_ (.Y(_0195_),
    .A(_0177_),
    .B(_0194_));
 sg13g2_xor2_1 _0914_ (.B(net174),
    .A(\counter[5] ),
    .X(_0196_));
 sg13g2_nand4_1 _0915_ (.B(_0177_),
    .C(_0194_),
    .A(_0157_),
    .Y(_0197_),
    .D(_0196_));
 sg13g2_a221oi_1 _0916_ (.B2(_0168_),
    .C1(_0197_),
    .B1(_0166_),
    .A1(_0053_),
    .Y(_0198_),
    .A2(_0063_));
 sg13g2_a22oi_1 _0917_ (.Y(_0199_),
    .B1(\counter[6] ),
    .B2(net172),
    .A2(net170),
    .A1(\counter[7] ));
 sg13g2_or2_1 _0918_ (.X(_0200_),
    .B(_0199_),
    .A(_0193_));
 sg13g2_o21ai_1 _0919_ (.B1(_0200_),
    .Y(_0201_),
    .A1(_0184_),
    .A2(_0195_));
 sg13g2_o21ai_1 _0920_ (.B1(_0192_),
    .Y(_0202_),
    .A1(_0198_),
    .A2(_0201_));
 sg13g2_or3_1 _0921_ (.A(_0192_),
    .B(_0198_),
    .C(_0201_),
    .X(_0203_));
 sg13g2_and2_1 _0922_ (.A(_0202_),
    .B(_0203_),
    .X(_0204_));
 sg13g2_and2_1 _0923_ (.A(_0191_),
    .B(_0202_),
    .X(_0205_));
 sg13g2_nand2_1 _0924_ (.Y(_0206_),
    .A(_0191_),
    .B(_0202_));
 sg13g2_nand2_1 _0925_ (.Y(_0207_),
    .A(\counter[9] ),
    .B(\hvsync_gen.hpos[9] ));
 sg13g2_nor3_2 _0926_ (.A(_0204_),
    .B(_0205_),
    .C(_0207_),
    .Y(_0208_));
 sg13g2_xnor2_1 _0927_ (.Y(_0209_),
    .A(\counter[9] ),
    .B(\hvsync_gen.hpos[9] ));
 sg13g2_a21o_1 _0928_ (.A2(_0202_),
    .A1(_0191_),
    .B1(_0209_),
    .X(_0210_));
 sg13g2_nand3_1 _0929_ (.B(_0207_),
    .C(_0210_),
    .A(_0204_),
    .Y(_0211_));
 sg13g2_nor2b_1 _0930_ (.A(_0208_),
    .B_N(_0211_),
    .Y(_0212_));
 sg13g2_o21ai_1 _0931_ (.B1(_0176_),
    .Y(_0213_),
    .A1(_0178_),
    .A2(_0185_));
 sg13g2_xnor2_1 _0932_ (.Y(_0214_),
    .A(_0194_),
    .B(_0213_));
 sg13g2_or2_1 _0933_ (.X(_0215_),
    .B(_0209_),
    .A(_0206_));
 sg13g2_nand2_1 _0934_ (.Y(_0216_),
    .A(_0206_),
    .B(_0209_));
 sg13g2_xnor2_1 _0935_ (.Y(_0217_),
    .A(_0206_),
    .B(_0209_));
 sg13g2_a221oi_1 _0936_ (.B2(_0210_),
    .C1(_0217_),
    .B1(_0207_),
    .A1(_0202_),
    .Y(_0218_),
    .A2(_0203_));
 sg13g2_nor2b_1 _0937_ (.A(_0208_),
    .B_N(_0217_),
    .Y(_0219_));
 sg13g2_nand3b_1 _0938_ (.B(_0211_),
    .C(_0214_),
    .Y(_0220_),
    .A_N(_0208_));
 sg13g2_a221oi_1 _0939_ (.B2(_0216_),
    .C1(_0208_),
    .B1(_0215_),
    .A1(_0211_),
    .Y(_0221_),
    .A2(_0214_));
 sg13g2_o21ai_1 _0940_ (.B1(_0214_),
    .Y(_0222_),
    .A1(_0218_),
    .A2(_0221_));
 sg13g2_xnor2_1 _0941_ (.Y(_0223_),
    .A(_0212_),
    .B(_0222_));
 sg13g2_a21oi_1 _0942_ (.A1(net185),
    .A2(_0223_),
    .Y(_0224_),
    .B1(_0190_));
 sg13g2_or3_1 _0943_ (.A(_0214_),
    .B(_0218_),
    .C(_0221_),
    .X(_0225_));
 sg13g2_a21oi_1 _0944_ (.A1(_0222_),
    .A2(_0225_),
    .Y(_0226_),
    .B1(_0060_));
 sg13g2_nor2_1 _0945_ (.A(net185),
    .B(_0007_),
    .Y(_0227_));
 sg13g2_nand2_1 _0946_ (.Y(_0228_),
    .A(_0060_),
    .B(_0007_));
 sg13g2_nand3_1 _0947_ (.B(_0222_),
    .C(_0225_),
    .A(net185),
    .Y(_0229_));
 sg13g2_a21o_1 _0948_ (.A2(_0220_),
    .A1(_0218_),
    .B1(_0219_),
    .X(_0230_));
 sg13g2_nor2_1 _0949_ (.A(_0060_),
    .B(_0221_),
    .Y(_0231_));
 sg13g2_a22oi_1 _0950_ (.Y(_0232_),
    .B1(_0230_),
    .B2(_0231_),
    .A2(_0068_),
    .A1(_0060_));
 sg13g2_nor3_1 _0951_ (.A(_0226_),
    .B(_0227_),
    .C(_0232_),
    .Y(_0233_));
 sg13g2_or3_1 _0952_ (.A(_0226_),
    .B(_0227_),
    .C(_0232_),
    .X(_0234_));
 sg13g2_nor2_1 _0953_ (.A(_0224_),
    .B(_0234_),
    .Y(_0235_));
 sg13g2_and3_1 _0954_ (.X(_0236_),
    .A(_0228_),
    .B(_0229_),
    .C(_0232_));
 sg13g2_a21oi_1 _0955_ (.A1(_0224_),
    .A2(_0233_),
    .Y(_0237_),
    .B1(_0236_));
 sg13g2_nand2_1 _0956_ (.Y(_0238_),
    .A(_0189_),
    .B(_0237_));
 sg13g2_nand2_1 _0957_ (.Y(_0239_),
    .A(_0224_),
    .B(_0234_));
 sg13g2_inv_1 _0958_ (.Y(_0240_),
    .A(_0239_));
 sg13g2_a21oi_1 _0959_ (.A1(_0238_),
    .A2(_0240_),
    .Y(_0241_),
    .B1(_0235_));
 sg13g2_inv_4 _0960_ (.A(net155),
    .Y(uio_out[3]));
 sg13g2_nand2_1 _0961_ (.Y(_0242_),
    .A(_0189_),
    .B(_0235_));
 sg13g2_a21o_1 _0962_ (.A2(uio_out[3]),
    .A1(_0189_),
    .B1(_0237_),
    .X(_0243_));
 sg13g2_nand2_1 _0963_ (.Y(_0244_),
    .A(_0242_),
    .B(_0243_));
 sg13g2_xnor2_1 _0964_ (.Y(_0245_),
    .A(_0188_),
    .B(uio_out[3]));
 sg13g2_xnor2_1 _0965_ (.Y(_0246_),
    .A(_0183_),
    .B(_0196_));
 sg13g2_nor2_1 _0966_ (.A(net185),
    .B(_0008_),
    .Y(_0247_));
 sg13g2_a21oi_2 _0967_ (.B1(_0247_),
    .Y(_0248_),
    .A2(_0246_),
    .A1(net186));
 sg13g2_nand2_1 _0968_ (.Y(_0249_),
    .A(_0245_),
    .B(_0248_));
 sg13g2_a22oi_1 _0969_ (.Y(_0250_),
    .B1(_0245_),
    .B2(_0248_),
    .A2(_0243_),
    .A1(_0242_));
 sg13g2_nand2_1 _0970_ (.Y(_0251_),
    .A(_0188_),
    .B(_0235_));
 sg13g2_o21ai_1 _0971_ (.B1(_0251_),
    .Y(_0252_),
    .A1(_0238_),
    .A2(_0239_));
 sg13g2_nor2_2 _0972_ (.A(_0250_),
    .B(_0252_),
    .Y(_0253_));
 sg13g2_inv_1 _0973_ (.Y(net154),
    .A(_0253_));
 sg13g2_a21oi_1 _0974_ (.A1(_0249_),
    .A2(_0252_),
    .Y(_0254_),
    .B1(_0244_));
 sg13g2_nor2_1 _0975_ (.A(_0250_),
    .B(_0254_),
    .Y(_0255_));
 sg13g2_o21ai_1 _0976_ (.B1(_0248_),
    .Y(_0256_),
    .A1(_0250_),
    .A2(_0252_));
 sg13g2_or3_1 _0977_ (.A(_0244_),
    .B(_0248_),
    .C(_0252_),
    .X(_0257_));
 sg13g2_and2_1 _0978_ (.A(_0256_),
    .B(_0257_),
    .X(_0258_));
 sg13g2_nand3_1 _0979_ (.B(_0256_),
    .C(_0257_),
    .A(_0174_),
    .Y(_0259_));
 sg13g2_xor2_1 _0980_ (.B(_0256_),
    .A(_0245_),
    .X(_0260_));
 sg13g2_a21oi_2 _0981_ (.B1(_0255_),
    .Y(_0261_),
    .A2(_0260_),
    .A1(_0259_));
 sg13g2_inv_2 _0982_ (.Y(uio_out[1]),
    .A(_0261_));
 sg13g2_xnor2_1 _0983_ (.Y(_0262_),
    .A(_0174_),
    .B(_0261_));
 sg13g2_nor2_1 _0984_ (.A(net186),
    .B(_0010_),
    .Y(_0263_));
 sg13g2_xor2_1 _0985_ (.B(net178),
    .A(\counter[3] ),
    .X(_0264_));
 sg13g2_xnor2_1 _0986_ (.Y(_0265_),
    .A(_0167_),
    .B(_0264_));
 sg13g2_a21oi_2 _0987_ (.B1(_0263_),
    .Y(_0266_),
    .A2(_0265_),
    .A1(net186));
 sg13g2_nand2_1 _0988_ (.Y(_0267_),
    .A(_0262_),
    .B(_0266_));
 sg13g2_a21o_1 _0989_ (.A2(uio_out[1]),
    .A1(_0174_),
    .B1(_0258_),
    .X(_0268_));
 sg13g2_nand3_1 _0990_ (.B(_0255_),
    .C(_0258_),
    .A(_0174_),
    .Y(_0269_));
 sg13g2_nand2_1 _0991_ (.Y(_0270_),
    .A(_0268_),
    .B(_0269_));
 sg13g2_a22oi_1 _0992_ (.Y(_0271_),
    .B1(_0268_),
    .B2(_0269_),
    .A2(_0266_),
    .A1(_0262_));
 sg13g2_and3_1 _0993_ (.X(_0272_),
    .A(_0174_),
    .B(_0245_),
    .C(_0258_));
 sg13g2_nor2b_1 _0994_ (.A(_0272_),
    .B_N(_0255_),
    .Y(_0273_));
 sg13g2_a21o_2 _0995_ (.A2(_0261_),
    .A1(_0260_),
    .B1(_0273_),
    .X(_0274_));
 sg13g2_nor2_2 _0996_ (.A(net148),
    .B(_0274_),
    .Y(_0275_));
 sg13g2_inv_1 _0997_ (.Y(uio_out[0]),
    .A(_0275_));
 sg13g2_nand2b_1 _0998_ (.Y(_0276_),
    .B(net59),
    .A_N(net162));
 sg13g2_nor2_1 _0999_ (.A(_0079_),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_nor2b_1 _1000_ (.A(\hvsync_gen.vpos[2] ),
    .B_N(net167),
    .Y(_0278_));
 sg13g2_nand4_1 _1001_ (.B(_0057_),
    .C(net55),
    .A(net165),
    .Y(_0279_),
    .D(_0278_));
 sg13g2_nor3_1 _1002_ (.A(_0079_),
    .B(_0276_),
    .C(_0279_),
    .Y(_0001_));
 sg13g2_nor2_1 _1003_ (.A(\hvsync_gen.hpos[8] ),
    .B(net169),
    .Y(_0280_));
 sg13g2_nor2_2 _1004_ (.A(net71),
    .B(_0280_),
    .Y(_0281_));
 sg13g2_nand2_1 _1005_ (.Y(_0282_),
    .A(net171),
    .B(net175));
 sg13g2_nand3_1 _1006_ (.B(net174),
    .C(net175),
    .A(net171),
    .Y(_0283_));
 sg13g2_nand2_1 _1007_ (.Y(_0284_),
    .A(_0062_),
    .B(_0283_));
 sg13g2_nand2_1 _1008_ (.Y(_0285_),
    .A(net169),
    .B(net171));
 sg13g2_nand3_1 _1009_ (.B(net171),
    .C(net173),
    .A(net170),
    .Y(_0286_));
 sg13g2_nor2_1 _1010_ (.A(net173),
    .B(net176),
    .Y(_0287_));
 sg13g2_o21ai_1 _1011_ (.B1(net169),
    .Y(_0288_),
    .A1(net173),
    .A2(net175));
 sg13g2_and2_1 _1012_ (.A(_0285_),
    .B(_0288_),
    .X(_0289_));
 sg13g2_a221oi_1 _1013_ (.B2(_0062_),
    .C1(_0061_),
    .B1(_0289_),
    .A1(_0281_),
    .Y(_0000_),
    .A2(_0284_));
 sg13g2_nand2_1 _1014_ (.Y(_0290_),
    .A(_0054_),
    .B(net164));
 sg13g2_nor3_1 _1015_ (.A(_0056_),
    .B(net166),
    .C(_0290_),
    .Y(_0291_));
 sg13g2_nor2_1 _1016_ (.A(\hvsync_gen.vpos[0] ),
    .B(\hvsync_gen.vpos[1] ),
    .Y(_0292_));
 sg13g2_and2_1 _1017_ (.A(_0278_),
    .B(_0292_),
    .X(_0293_));
 sg13g2_nand2_1 _1018_ (.Y(_0294_),
    .A(_0278_),
    .B(_0292_));
 sg13g2_o21ai_1 _1019_ (.B1(_0291_),
    .Y(_0295_),
    .A1(_0004_),
    .A2(_0293_));
 sg13g2_o21ai_1 _1020_ (.B1(\hvsync_gen.vpos[8] ),
    .Y(_0296_),
    .A1(\hvsync_gen.vpos[7] ),
    .A2(\hvsync_gen.vpos[6] ));
 sg13g2_a21oi_1 _1021_ (.A1(_0054_),
    .A2(_0003_),
    .Y(_0297_),
    .B1(_0296_));
 sg13g2_nor2_1 _1022_ (.A(_0276_),
    .B(_0294_),
    .Y(_0298_));
 sg13g2_a221oi_1 _1023_ (.B2(_0291_),
    .C1(net162),
    .B1(_0298_),
    .A1(_0295_),
    .Y(_0299_),
    .A2(_0297_));
 sg13g2_nor2_1 _1024_ (.A(net179),
    .B(net180),
    .Y(_0300_));
 sg13g2_a21oi_1 _1025_ (.A1(net181),
    .A2(_0061_),
    .Y(_0301_),
    .B1(\hvsync_gen.hpos[3] ));
 sg13g2_a21oi_1 _1026_ (.A1(_0300_),
    .A2(_0301_),
    .Y(_0302_),
    .B1(_0283_));
 sg13g2_nor4_1 _1027_ (.A(\hvsync_gen.hpos[8] ),
    .B(net169),
    .C(_0068_),
    .D(_0302_),
    .Y(_0303_));
 sg13g2_nor2_2 _1028_ (.A(_0299_),
    .B(_0303_),
    .Y(_0304_));
 sg13g2_nor3_1 _1029_ (.A(net176),
    .B(net178),
    .C(net179),
    .Y(_0305_));
 sg13g2_o21ai_1 _1030_ (.B1(_0061_),
    .Y(_0306_),
    .A1(_0286_),
    .A2(_0305_));
 sg13g2_nor2_2 _1031_ (.A(\hvsync_gen.hpos[8] ),
    .B(_0306_),
    .Y(_0307_));
 sg13g2_nand2_1 _1032_ (.Y(_0308_),
    .A(_0304_),
    .B(_0307_));
 sg13g2_nor3_2 _1033_ (.A(_0055_),
    .B(_0056_),
    .C(_0079_),
    .Y(_0309_));
 sg13g2_nor3_2 _1034_ (.A(net163),
    .B(_0281_),
    .C(_0309_),
    .Y(_0310_));
 sg13g2_nand3_1 _1035_ (.B(_0307_),
    .C(_0310_),
    .A(_0304_),
    .Y(_0311_));
 sg13g2_inv_1 _1036_ (.Y(uo_out[5]),
    .A(_0311_));
 sg13g2_nand2_1 _1037_ (.Y(_0312_),
    .A(net153),
    .B(uio_out[1]));
 sg13g2_o21ai_1 _1038_ (.B1(net153),
    .Y(_0313_),
    .A1(net148),
    .A2(_0274_));
 sg13g2_nand2b_1 _1039_ (.Y(_0314_),
    .B(uio_out[1]),
    .A_N(_0313_));
 sg13g2_o21ai_1 _1040_ (.B1(uio_out[1]),
    .Y(_0315_),
    .A1(net148),
    .A2(_0273_));
 sg13g2_inv_1 _1041_ (.Y(_0316_),
    .A(_0315_));
 sg13g2_or3_1 _1042_ (.A(uio_out[1]),
    .B(net148),
    .C(_0274_),
    .X(_0317_));
 sg13g2_and2_1 _1043_ (.A(_0253_),
    .B(_0317_),
    .X(_0318_));
 sg13g2_o21ai_1 _1044_ (.B1(_0261_),
    .Y(_0319_),
    .A1(net148),
    .A2(_0274_));
 sg13g2_or3_1 _1045_ (.A(_0261_),
    .B(net148),
    .C(_0273_),
    .X(_0320_));
 sg13g2_a21oi_1 _1046_ (.A1(_0319_),
    .A2(net145),
    .Y(_0321_),
    .B1(net153));
 sg13g2_inv_1 _1047_ (.Y(_0322_),
    .A(_0321_));
 sg13g2_nor3_1 _1048_ (.A(net149),
    .B(net156),
    .C(_0321_),
    .Y(_0323_));
 sg13g2_nand2_2 _1049_ (.Y(_0324_),
    .A(net155),
    .B(_0253_));
 sg13g2_nand2_1 _1050_ (.Y(_0325_),
    .A(_0253_),
    .B(_0261_));
 sg13g2_nor2_1 _1051_ (.A(uio_out[3]),
    .B(_0275_),
    .Y(_0326_));
 sg13g2_nor2_2 _1052_ (.A(_0319_),
    .B(_0324_),
    .Y(_0327_));
 sg13g2_or2_1 _1053_ (.X(_0328_),
    .B(_0324_),
    .A(_0319_));
 sg13g2_nor2_1 _1054_ (.A(_0253_),
    .B(uio_out[1]),
    .Y(_0329_));
 sg13g2_nand2_1 _1055_ (.Y(_0330_),
    .A(net153),
    .B(_0261_));
 sg13g2_nand2_1 _1056_ (.Y(_0331_),
    .A(net153),
    .B(net145));
 sg13g2_a21oi_1 _1057_ (.A1(_0253_),
    .A2(_0317_),
    .Y(_0332_),
    .B1(net155));
 sg13g2_a21o_1 _1058_ (.A2(_0332_),
    .A1(_0331_),
    .B1(_0327_),
    .X(_0333_));
 sg13g2_nor2_1 _1059_ (.A(_0148_),
    .B(net149),
    .Y(_0334_));
 sg13g2_a221oi_1 _1060_ (.B2(net149),
    .C1(_0148_),
    .B1(_0333_),
    .A1(_0314_),
    .Y(_0335_),
    .A2(_0323_));
 sg13g2_nor2_1 _1061_ (.A(net146),
    .B(_0329_),
    .Y(_0336_));
 sg13g2_a21oi_1 _1062_ (.A1(net156),
    .A2(_0275_),
    .Y(_0337_),
    .B1(_0316_));
 sg13g2_nor2_2 _1063_ (.A(uio_out[5]),
    .B(net146),
    .Y(_0338_));
 sg13g2_a221oi_1 _1064_ (.B2(_0337_),
    .C1(uio_out[5]),
    .B1(_0336_),
    .A1(net146),
    .Y(_0339_),
    .A2(_0333_));
 sg13g2_nor3_1 _1065_ (.A(uio_out[6]),
    .B(_0335_),
    .C(_0339_),
    .Y(_0340_));
 sg13g2_nand4_1 _1066_ (.B(net152),
    .C(net150),
    .A(uio_out[6]),
    .Y(_0341_),
    .D(_0327_));
 sg13g2_nand2_2 _1067_ (.Y(_0342_),
    .A(uio_out[6]),
    .B(_0148_));
 sg13g2_nor2_1 _1068_ (.A(uio_out[2]),
    .B(net145),
    .Y(_0343_));
 sg13g2_or2_1 _1069_ (.X(_0344_),
    .B(_0320_),
    .A(net153));
 sg13g2_nor2_1 _1070_ (.A(net145),
    .B(_0324_),
    .Y(_0345_));
 sg13g2_inv_1 _1071_ (.Y(_0346_),
    .A(_0345_));
 sg13g2_o21ai_1 _1072_ (.B1(_0341_),
    .Y(_0347_),
    .A1(_0342_),
    .A2(_0346_));
 sg13g2_o21ai_1 _1073_ (.B1(uio_out[7]),
    .Y(_0348_),
    .A1(_0340_),
    .A2(_0347_));
 sg13g2_o21ai_1 _1074_ (.B1(_0266_),
    .Y(_0349_),
    .A1(_0271_),
    .A2(_0274_));
 sg13g2_or3_1 _1075_ (.A(_0266_),
    .B(net148),
    .C(_0274_),
    .X(_0350_));
 sg13g2_nand2_1 _1076_ (.Y(_0351_),
    .A(_0159_),
    .B(_0164_));
 sg13g2_nor2_1 _1077_ (.A(_0060_),
    .B(_0165_),
    .Y(_0352_));
 sg13g2_a22oi_1 _1078_ (.Y(_0353_),
    .B1(_0351_),
    .B2(_0352_),
    .A2(_0065_),
    .A1(_0060_));
 sg13g2_and3_1 _1079_ (.X(_0354_),
    .A(_0349_),
    .B(_0350_),
    .C(_0353_));
 sg13g2_xnor2_1 _1080_ (.Y(_0355_),
    .A(_0262_),
    .B(_0349_));
 sg13g2_a21oi_1 _1081_ (.A1(_0267_),
    .A2(_0274_),
    .Y(_0356_),
    .B1(_0270_));
 sg13g2_or2_1 _1082_ (.X(_0357_),
    .B(_0356_),
    .A(net148));
 sg13g2_o21ai_1 _1083_ (.B1(_0357_),
    .Y(_0358_),
    .A1(_0354_),
    .A2(_0355_));
 sg13g2_inv_1 _1084_ (.Y(_0359_),
    .A(_0358_));
 sg13g2_xnor2_1 _1085_ (.Y(_0360_),
    .A(_0161_),
    .B(_0163_));
 sg13g2_nor2_1 _1086_ (.A(net186),
    .B(_0012_),
    .Y(_0361_));
 sg13g2_a21oi_2 _1087_ (.B1(_0361_),
    .Y(_0362_),
    .A2(_0360_),
    .A1(net186));
 sg13g2_o21ai_1 _1088_ (.B1(_0362_),
    .Y(_0363_),
    .A1(_0353_),
    .A2(_0358_));
 sg13g2_a22oi_1 _1089_ (.Y(_0364_),
    .B1(_0353_),
    .B2(_0358_),
    .A2(_0350_),
    .A1(_0349_));
 sg13g2_o21ai_1 _1090_ (.B1(_0357_),
    .Y(_0365_),
    .A1(_0355_),
    .A2(_0358_));
 sg13g2_a21oi_2 _1091_ (.B1(_0365_),
    .Y(_0366_),
    .A2(_0364_),
    .A1(_0363_));
 sg13g2_nor2_2 _1092_ (.A(net152),
    .B(net150),
    .Y(_0367_));
 sg13g2_a21oi_1 _1093_ (.A1(_0327_),
    .A2(_0367_),
    .Y(_0368_),
    .B1(uio_out[6]));
 sg13g2_nand2b_1 _1094_ (.Y(_0369_),
    .B(_0128_),
    .A_N(_0368_));
 sg13g2_nand2_1 _1095_ (.Y(_0370_),
    .A(net152),
    .B(_0345_));
 sg13g2_a21oi_1 _1096_ (.A1(_0368_),
    .A2(_0370_),
    .Y(_0371_),
    .B1(uio_out[7]));
 sg13g2_a221oi_1 _1097_ (.B2(net149),
    .C1(_0148_),
    .B1(_0333_),
    .A1(_0323_),
    .Y(_0372_),
    .A2(_0331_));
 sg13g2_nor2_1 _1098_ (.A(net146),
    .B(net156),
    .Y(_0373_));
 sg13g2_a221oi_1 _1099_ (.B2(_0313_),
    .C1(uio_out[5]),
    .B1(_0373_),
    .A1(uio_out[4]),
    .Y(_0374_),
    .A2(_0333_));
 sg13g2_nor2_1 _1100_ (.A(_0148_),
    .B(_0328_),
    .Y(_0375_));
 sg13g2_a21oi_1 _1101_ (.A1(net146),
    .A2(_0375_),
    .Y(_0376_),
    .B1(_0138_));
 sg13g2_o21ai_1 _1102_ (.B1(_0376_),
    .Y(_0377_),
    .A1(_0372_),
    .A2(_0374_));
 sg13g2_nand2_1 _1103_ (.Y(_0378_),
    .A(_0371_),
    .B(_0377_));
 sg13g2_nand3_1 _1104_ (.B(_0366_),
    .C(_0378_),
    .A(_0348_),
    .Y(_0379_));
 sg13g2_a21oi_2 _1105_ (.B1(uio_out[3]),
    .Y(_0380_),
    .A2(net145),
    .A1(_0319_));
 sg13g2_nand3_1 _1106_ (.B(_0325_),
    .C(_0380_),
    .A(net150),
    .Y(_0381_));
 sg13g2_and2_1 _1107_ (.A(_0319_),
    .B(_0330_),
    .X(_0382_));
 sg13g2_a21o_1 _1108_ (.A2(_0330_),
    .A1(_0319_),
    .B1(net155),
    .X(_0383_));
 sg13g2_o21ai_1 _1109_ (.B1(_0383_),
    .Y(_0384_),
    .A1(net155),
    .A2(_0344_));
 sg13g2_nand2_1 _1110_ (.Y(_0385_),
    .A(net155),
    .B(_0325_));
 sg13g2_nor2b_1 _1111_ (.A(_0385_),
    .B_N(_0312_),
    .Y(_0386_));
 sg13g2_nand2_1 _1112_ (.Y(_0387_),
    .A(_0315_),
    .B(_0386_));
 sg13g2_nand3_1 _1113_ (.B(_0317_),
    .C(_0386_),
    .A(_0315_),
    .Y(_0388_));
 sg13g2_nand2b_1 _1114_ (.Y(_0389_),
    .B(uio_out[4]),
    .A_N(_0388_));
 sg13g2_nor2b_1 _1115_ (.A(_0385_),
    .B_N(_0314_),
    .Y(_0390_));
 sg13g2_a21oi_1 _1116_ (.A1(_0315_),
    .A2(_0317_),
    .Y(_0391_),
    .B1(_0253_));
 sg13g2_nor3_1 _1117_ (.A(net155),
    .B(_0321_),
    .C(_0391_),
    .Y(_0392_));
 sg13g2_o21ai_1 _1118_ (.B1(_0338_),
    .Y(_0393_),
    .A1(_0390_),
    .A2(_0392_));
 sg13g2_o21ai_1 _1119_ (.B1(_0367_),
    .Y(_0394_),
    .A1(_0380_),
    .A2(_0384_));
 sg13g2_and2_1 _1120_ (.A(_0393_),
    .B(_0394_),
    .X(_0395_));
 sg13g2_nand3_1 _1121_ (.B(_0381_),
    .C(_0389_),
    .A(uio_out[6]),
    .Y(_0396_));
 sg13g2_o21ai_1 _1122_ (.B1(_0342_),
    .Y(_0397_),
    .A1(_0384_),
    .A2(_0396_));
 sg13g2_a21o_1 _1123_ (.A2(_0397_),
    .A1(_0395_),
    .B1(_0369_),
    .X(_0398_));
 sg13g2_nand3_1 _1124_ (.B(_0312_),
    .C(_0380_),
    .A(net150),
    .Y(_0399_));
 sg13g2_and4_1 _1125_ (.A(_0148_),
    .B(_0383_),
    .C(_0389_),
    .D(_0399_),
    .X(_0400_));
 sg13g2_nand4_1 _1126_ (.B(net149),
    .C(_0383_),
    .A(net152),
    .Y(_0401_),
    .D(_0388_));
 sg13g2_or3_1 _1127_ (.A(net155),
    .B(net153),
    .C(_0275_),
    .X(_0402_));
 sg13g2_nand4_1 _1128_ (.B(net146),
    .C(_0387_),
    .A(uio_out[5]),
    .Y(_0403_),
    .D(_0402_));
 sg13g2_nand3_1 _1129_ (.B(_0401_),
    .C(_0403_),
    .A(_0138_),
    .Y(_0404_));
 sg13g2_o21ai_1 _1130_ (.B1(_0341_),
    .Y(_0405_),
    .A1(_0400_),
    .A2(_0404_));
 sg13g2_a21oi_1 _1131_ (.A1(uio_out[7]),
    .A2(_0405_),
    .Y(_0406_),
    .B1(_0366_));
 sg13g2_a21oi_1 _1132_ (.A1(_0398_),
    .A2(_0406_),
    .Y(_0407_),
    .B1(_0359_));
 sg13g2_o21ai_1 _1133_ (.B1(uio_out[3]),
    .Y(_0408_),
    .A1(_0318_),
    .A2(_0329_));
 sg13g2_nand3_1 _1134_ (.B(net153),
    .C(uio_out[1]),
    .A(net156),
    .Y(_0409_));
 sg13g2_a21o_1 _1135_ (.A2(_0409_),
    .A1(_0408_),
    .B1(_0338_),
    .X(_0410_));
 sg13g2_a22oi_1 _1136_ (.Y(_0411_),
    .B1(net145),
    .B2(uio_out[2]),
    .A2(_0319_),
    .A1(uio_out[3]));
 sg13g2_nand4_1 _1137_ (.B(uio_out[2]),
    .C(_0319_),
    .A(uio_out[3]),
    .Y(_0412_),
    .D(net145));
 sg13g2_nor3_1 _1138_ (.A(uio_out[5]),
    .B(net146),
    .C(_0411_),
    .Y(_0413_));
 sg13g2_a22oi_1 _1139_ (.Y(_0414_),
    .B1(_0412_),
    .B2(_0413_),
    .A2(_0367_),
    .A1(_0327_));
 sg13g2_a22oi_1 _1140_ (.Y(_0415_),
    .B1(_0410_),
    .B2(_0414_),
    .A2(_0334_),
    .A1(_0326_));
 sg13g2_a21oi_1 _1141_ (.A1(_0345_),
    .A2(_0367_),
    .Y(_0416_),
    .B1(_0375_));
 sg13g2_a21oi_1 _1142_ (.A1(_0138_),
    .A2(_0416_),
    .Y(_0417_),
    .B1(uio_out[7]));
 sg13g2_o21ai_1 _1143_ (.B1(_0417_),
    .Y(_0418_),
    .A1(_0138_),
    .A2(_0415_));
 sg13g2_nor2_1 _1144_ (.A(_0328_),
    .B(_0342_),
    .Y(_0419_));
 sg13g2_a21o_1 _1145_ (.A2(_0409_),
    .A1(_0408_),
    .B1(_0326_),
    .X(_0420_));
 sg13g2_nor2_1 _1146_ (.A(_0334_),
    .B(_0338_),
    .Y(_0421_));
 sg13g2_o21ai_1 _1147_ (.B1(_0324_),
    .Y(_0422_),
    .A1(_0318_),
    .A2(_0380_));
 sg13g2_nor2_1 _1148_ (.A(uio_out[3]),
    .B(net145),
    .Y(_0423_));
 sg13g2_nor3_1 _1149_ (.A(net152),
    .B(uio_out[4]),
    .C(_0423_),
    .Y(_0424_));
 sg13g2_a21o_1 _1150_ (.A2(_0424_),
    .A1(_0408_),
    .B1(uio_out[6]),
    .X(_0425_));
 sg13g2_a221oi_1 _1151_ (.B2(_0334_),
    .C1(_0425_),
    .B1(_0422_),
    .A1(_0420_),
    .Y(_0426_),
    .A2(_0421_));
 sg13g2_o21ai_1 _1152_ (.B1(uio_out[7]),
    .Y(_0427_),
    .A1(_0419_),
    .A2(_0426_));
 sg13g2_nand3b_1 _1153_ (.B(_0418_),
    .C(_0427_),
    .Y(_0428_),
    .A_N(_0366_));
 sg13g2_and3_1 _1154_ (.X(_0429_),
    .A(uio_out[5]),
    .B(net146),
    .C(_0313_));
 sg13g2_nor2_1 _1155_ (.A(net149),
    .B(_0342_),
    .Y(_0430_));
 sg13g2_o21ai_1 _1156_ (.B1(_0382_),
    .Y(_0431_),
    .A1(_0429_),
    .A2(_0430_));
 sg13g2_a21o_1 _1157_ (.A2(_0367_),
    .A1(_0343_),
    .B1(uio_out[6]),
    .X(_0432_));
 sg13g2_o21ai_1 _1158_ (.B1(_0315_),
    .Y(_0433_),
    .A1(uio_out[2]),
    .A2(uio_out[0]));
 sg13g2_a22oi_1 _1159_ (.Y(_0434_),
    .B1(_0338_),
    .B2(_0433_),
    .A2(_0336_),
    .A1(uio_out[5]));
 sg13g2_nand3_1 _1160_ (.B(_0432_),
    .C(_0434_),
    .A(_0431_),
    .Y(_0435_));
 sg13g2_o21ai_1 _1161_ (.B1(_0343_),
    .Y(_0436_),
    .A1(_0148_),
    .A2(net149));
 sg13g2_a22oi_1 _1162_ (.Y(_0437_),
    .B1(_0436_),
    .B2(uio_out[6]),
    .A2(_0331_),
    .A1(_0322_));
 sg13g2_o21ai_1 _1163_ (.B1(net156),
    .Y(_0438_),
    .A1(_0128_),
    .A2(_0437_));
 sg13g2_a21o_1 _1164_ (.A2(_0435_),
    .A1(_0128_),
    .B1(_0438_),
    .X(_0439_));
 sg13g2_a21oi_1 _1165_ (.A1(_0366_),
    .A2(_0439_),
    .Y(_0440_),
    .B1(_0358_));
 sg13g2_a221oi_1 _1166_ (.B2(_0440_),
    .C1(net2),
    .B1(_0428_),
    .A1(_0379_),
    .Y(_0441_),
    .A2(_0407_));
 sg13g2_nor4_2 _1167_ (.A(\hvsync_gen.vpos[7] ),
    .B(net164),
    .C(net165),
    .Y(_0442_),
    .D(_0057_));
 sg13g2_o21ai_1 _1168_ (.B1(_0442_),
    .Y(_0443_),
    .A1(_0004_),
    .A2(_0293_));
 sg13g2_nor4_2 _1169_ (.A(\hvsync_gen.vpos[7] ),
    .B(\hvsync_gen.vpos[6] ),
    .C(net165),
    .Y(_0444_),
    .D(net166));
 sg13g2_nand2_1 _1170_ (.Y(_0445_),
    .A(\hvsync_gen.vpos[8] ),
    .B(_0443_));
 sg13g2_nand2b_1 _1171_ (.Y(_0446_),
    .B(net1),
    .A_N(net163));
 sg13g2_a21oi_1 _1172_ (.A1(_0298_),
    .A2(_0442_),
    .Y(_0447_),
    .B1(_0446_));
 sg13g2_o21ai_1 _1173_ (.B1(_0447_),
    .Y(_0448_),
    .A1(_0444_),
    .A2(_0445_));
 sg13g2_mux4_1 _1174_ (.S0(_0366_),
    .A0(net4),
    .A1(net3),
    .A2(net6),
    .A3(net5),
    .S1(_0358_),
    .X(_0449_));
 sg13g2_nand2b_1 _1175_ (.Y(_0450_),
    .B(net2),
    .A_N(_0449_));
 sg13g2_nand2b_1 _1176_ (.Y(_0451_),
    .B(_0450_),
    .A_N(_0448_));
 sg13g2_and3_1 _1177_ (.X(_0452_),
    .A(_0056_),
    .B(_0057_),
    .C(_0004_));
 sg13g2_a21oi_1 _1178_ (.A1(_0294_),
    .A2(_0452_),
    .Y(_0453_),
    .B1(_0079_));
 sg13g2_nor3_2 _1179_ (.A(net163),
    .B(\hvsync_gen.vpos[8] ),
    .C(_0453_),
    .Y(_0454_));
 sg13g2_or3_1 _1180_ (.A(net163),
    .B(\hvsync_gen.vpos[8] ),
    .C(_0453_),
    .X(_0455_));
 sg13g2_nand2b_1 _1181_ (.Y(_0456_),
    .B(_0013_),
    .A_N(net182));
 sg13g2_nor2_1 _1182_ (.A(net159),
    .B(net160),
    .Y(_0457_));
 sg13g2_or3_2 _1183_ (.A(net159),
    .B(net160),
    .C(\counter[2] ),
    .X(_0458_));
 sg13g2_nor2_1 _1184_ (.A(\counter[3] ),
    .B(_0458_),
    .Y(_0459_));
 sg13g2_nor3_2 _1185_ (.A(\counter[3] ),
    .B(\counter[4] ),
    .C(_0458_),
    .Y(_0460_));
 sg13g2_nor2b_1 _1186_ (.A(\counter[5] ),
    .B_N(_0460_),
    .Y(_0461_));
 sg13g2_nor2b_1 _1187_ (.A(\counter[6] ),
    .B_N(_0461_),
    .Y(_0462_));
 sg13g2_xnor2_1 _1188_ (.Y(_0463_),
    .A(_0016_),
    .B(_0462_));
 sg13g2_nand2_1 _1189_ (.Y(_0464_),
    .A(net170),
    .B(_0463_));
 sg13g2_xnor2_1 _1190_ (.Y(_0465_),
    .A(net170),
    .B(_0463_));
 sg13g2_xnor2_1 _1191_ (.Y(_0466_),
    .A(\counter[5] ),
    .B(_0460_));
 sg13g2_nand2b_1 _1192_ (.Y(_0467_),
    .B(_0466_),
    .A_N(_0008_));
 sg13g2_xor2_1 _1193_ (.B(net160),
    .A(net159),
    .X(_0468_));
 sg13g2_a22oi_1 _1194_ (.Y(_0469_),
    .B1(_0468_),
    .B2(_0066_),
    .A2(_0163_),
    .A1(_0161_));
 sg13g2_xnor2_1 _1195_ (.Y(_0470_),
    .A(_0159_),
    .B(_0457_));
 sg13g2_o21ai_1 _1196_ (.B1(\counter[2] ),
    .Y(_0471_),
    .A1(net159),
    .A2(net160));
 sg13g2_nand3_1 _1197_ (.B(_0458_),
    .C(_0471_),
    .A(_0065_),
    .Y(_0472_));
 sg13g2_o21ai_1 _1198_ (.B1(_0472_),
    .Y(_0473_),
    .A1(_0469_),
    .A2(_0470_));
 sg13g2_xnor2_1 _1199_ (.Y(_0474_),
    .A(_0264_),
    .B(_0458_));
 sg13g2_inv_1 _1200_ (.Y(_0475_),
    .A(_0474_));
 sg13g2_or2_1 _1201_ (.X(_0476_),
    .B(_0459_),
    .A(_0010_));
 sg13g2_a21oi_1 _1202_ (.A1(\counter[3] ),
    .A2(_0458_),
    .Y(_0477_),
    .B1(_0476_));
 sg13g2_a21o_1 _1203_ (.A2(_0475_),
    .A1(_0473_),
    .B1(_0477_),
    .X(_0478_));
 sg13g2_xnor2_1 _1204_ (.Y(_0479_),
    .A(_0157_),
    .B(_0459_));
 sg13g2_xnor2_1 _1205_ (.Y(_0480_),
    .A(\counter[4] ),
    .B(_0459_));
 sg13g2_a22oi_1 _1206_ (.Y(_0481_),
    .B1(_0480_),
    .B2(_0064_),
    .A2(_0479_),
    .A1(_0478_));
 sg13g2_nor2b_1 _1207_ (.A(_0466_),
    .B_N(_0008_),
    .Y(_0482_));
 sg13g2_xnor2_1 _1208_ (.Y(_0483_),
    .A(_0008_),
    .B(_0466_));
 sg13g2_o21ai_1 _1209_ (.B1(_0467_),
    .Y(_0484_),
    .A1(_0481_),
    .A2(_0482_));
 sg13g2_xnor2_1 _1210_ (.Y(_0485_),
    .A(_0178_),
    .B(_0461_));
 sg13g2_inv_1 _1211_ (.Y(_0486_),
    .A(_0485_));
 sg13g2_nand2b_1 _1212_ (.Y(_0487_),
    .B(\counter[6] ),
    .A_N(_0461_));
 sg13g2_nor2_1 _1213_ (.A(_0002_),
    .B(_0462_),
    .Y(_0488_));
 sg13g2_a22oi_1 _1214_ (.Y(_0489_),
    .B1(_0487_),
    .B2(_0488_),
    .A2(_0486_),
    .A1(_0484_));
 sg13g2_o21ai_1 _1215_ (.B1(_0464_),
    .Y(_0490_),
    .A1(_0465_),
    .A2(_0489_));
 sg13g2_nand2b_1 _1216_ (.Y(_0491_),
    .B(\counter[7] ),
    .A_N(_0462_));
 sg13g2_nand2_1 _1217_ (.Y(_0492_),
    .A(_0018_),
    .B(_0491_));
 sg13g2_xor2_1 _1218_ (.B(_0491_),
    .A(_0018_),
    .X(_0493_));
 sg13g2_xnor2_1 _1219_ (.Y(_0494_),
    .A(_0062_),
    .B(_0493_));
 sg13g2_a22oi_1 _1220_ (.Y(_0495_),
    .B1(_0494_),
    .B2(_0490_),
    .A2(_0493_),
    .A1(_0069_));
 sg13g2_xor2_1 _1221_ (.B(_0492_),
    .A(_0015_),
    .X(_0496_));
 sg13g2_xnor2_1 _1222_ (.Y(_0497_),
    .A(\hvsync_gen.hpos[9] ),
    .B(_0496_));
 sg13g2_nand2_1 _1223_ (.Y(_0498_),
    .A(_0495_),
    .B(_0497_));
 sg13g2_nor2b_1 _1224_ (.A(\counter[8] ),
    .B_N(\counter[9] ),
    .Y(_0499_));
 sg13g2_a21oi_1 _1225_ (.A1(_0491_),
    .A2(_0499_),
    .Y(_0500_),
    .B1(_0015_));
 sg13g2_nor2_1 _1226_ (.A(_0495_),
    .B(_0497_),
    .Y(_0501_));
 sg13g2_a21oi_1 _1227_ (.A1(_0068_),
    .A2(_0496_),
    .Y(_0502_),
    .B1(_0501_));
 sg13g2_a21oi_1 _1228_ (.A1(_0500_),
    .A2(_0502_),
    .Y(_0503_),
    .B1(_0498_));
 sg13g2_nand3_1 _1229_ (.B(_0500_),
    .C(_0502_),
    .A(_0498_),
    .Y(_0504_));
 sg13g2_nor2_1 _1230_ (.A(_0501_),
    .B(_0503_),
    .Y(_0505_));
 sg13g2_and2_1 _1231_ (.A(_0504_),
    .B(_0505_),
    .X(_0506_));
 sg13g2_xnor2_1 _1232_ (.Y(_0507_),
    .A(_0490_),
    .B(_0494_));
 sg13g2_o21ai_1 _1233_ (.B1(_0504_),
    .Y(_0508_),
    .A1(_0500_),
    .A2(_0502_));
 sg13g2_and2_1 _1234_ (.A(_0507_),
    .B(_0508_),
    .X(_0509_));
 sg13g2_nand2b_1 _1235_ (.Y(_0510_),
    .B(_0506_),
    .A_N(_0509_));
 sg13g2_xnor2_1 _1236_ (.Y(_0511_),
    .A(_0465_),
    .B(_0489_));
 sg13g2_inv_1 _1237_ (.Y(_0512_),
    .A(_0511_));
 sg13g2_nor2_1 _1238_ (.A(_0507_),
    .B(_0508_),
    .Y(_0513_));
 sg13g2_a21oi_1 _1239_ (.A1(_0506_),
    .A2(_0509_),
    .Y(_0514_),
    .B1(_0513_));
 sg13g2_and2_1 _1240_ (.A(_0511_),
    .B(_0514_),
    .X(_0515_));
 sg13g2_nor2b_1 _1241_ (.A(_0510_),
    .B_N(_0515_),
    .Y(_0516_));
 sg13g2_nand2b_1 _1242_ (.Y(_0517_),
    .B(_0509_),
    .A_N(_0506_));
 sg13g2_o21ai_1 _1243_ (.B1(net182),
    .Y(_0518_),
    .A1(_0511_),
    .A2(_0517_));
 sg13g2_o21ai_1 _1244_ (.B1(_0456_),
    .Y(_0519_),
    .A1(_0516_),
    .A2(_0518_));
 sg13g2_nand2b_1 _1245_ (.Y(_0520_),
    .B(_0019_),
    .A_N(net182));
 sg13g2_o21ai_1 _1246_ (.B1(_0517_),
    .Y(_0521_),
    .A1(_0510_),
    .A2(_0515_));
 sg13g2_a21oi_1 _1247_ (.A1(_0511_),
    .A2(_0521_),
    .Y(_0522_),
    .B1(_0514_));
 sg13g2_o21ai_1 _1248_ (.B1(net182),
    .Y(_0523_),
    .A1(_0512_),
    .A2(_0517_));
 sg13g2_o21ai_1 _1249_ (.B1(_0520_),
    .Y(_0524_),
    .A1(_0522_),
    .A2(_0523_));
 sg13g2_nand2_1 _1250_ (.Y(_0525_),
    .A(_0519_),
    .B(_0524_));
 sg13g2_nor2_1 _1251_ (.A(net169),
    .B(net182),
    .Y(_0526_));
 sg13g2_xnor2_1 _1252_ (.Y(_0527_),
    .A(_0512_),
    .B(_0521_));
 sg13g2_a21oi_2 _1253_ (.B1(_0526_),
    .Y(_0528_),
    .A2(_0527_),
    .A1(net184));
 sg13g2_xnor2_1 _1254_ (.Y(_0529_),
    .A(_0484_),
    .B(_0486_));
 sg13g2_nor2_1 _1255_ (.A(net171),
    .B(net182),
    .Y(_0530_));
 sg13g2_a21oi_2 _1256_ (.B1(_0530_),
    .Y(_0531_),
    .A2(_0529_),
    .A1(net182));
 sg13g2_inv_1 _1257_ (.Y(_0532_),
    .A(_0531_));
 sg13g2_nor2_1 _1258_ (.A(_0528_),
    .B(_0531_),
    .Y(_0533_));
 sg13g2_xnor2_1 _1259_ (.Y(_0534_),
    .A(_0473_),
    .B(_0475_));
 sg13g2_nor2b_1 _1260_ (.A(net183),
    .B_N(_0010_),
    .Y(_0535_));
 sg13g2_a21oi_2 _1261_ (.B1(_0535_),
    .Y(_0536_),
    .A2(_0534_),
    .A1(net183));
 sg13g2_xnor2_1 _1262_ (.Y(_0537_),
    .A(_0469_),
    .B(_0470_));
 sg13g2_nand2_1 _1263_ (.Y(_0538_),
    .A(net184),
    .B(_0537_));
 sg13g2_o21ai_1 _1264_ (.B1(_0538_),
    .Y(_0539_),
    .A1(_0065_),
    .A2(net183));
 sg13g2_nor2_1 _1265_ (.A(_0012_),
    .B(net183),
    .Y(_0540_));
 sg13g2_nor2b_1 _1266_ (.A(net181),
    .B_N(net160),
    .Y(_0541_));
 sg13g2_xnor2_1 _1267_ (.Y(_0542_),
    .A(_0163_),
    .B(_0541_));
 sg13g2_a21oi_1 _1268_ (.A1(net183),
    .A2(_0542_),
    .Y(_0543_),
    .B1(_0540_));
 sg13g2_nand2_1 _1269_ (.Y(_0544_),
    .A(_0539_),
    .B(_0543_));
 sg13g2_nor2_1 _1270_ (.A(_0009_),
    .B(net184),
    .Y(_0545_));
 sg13g2_xor2_1 _1271_ (.B(_0479_),
    .A(_0478_),
    .X(_0546_));
 sg13g2_a21oi_2 _1272_ (.B1(_0545_),
    .Y(_0547_),
    .A2(_0546_),
    .A1(net183));
 sg13g2_inv_1 _1273_ (.Y(_0548_),
    .A(_0547_));
 sg13g2_o21ai_1 _1274_ (.B1(_0548_),
    .Y(_0549_),
    .A1(_0536_),
    .A2(_0544_));
 sg13g2_nor2_1 _1275_ (.A(_0008_),
    .B(net182),
    .Y(_0550_));
 sg13g2_xnor2_1 _1276_ (.Y(_0551_),
    .A(_0481_),
    .B(_0483_));
 sg13g2_a21oi_2 _1277_ (.B1(_0550_),
    .Y(_0552_),
    .A2(_0551_),
    .A1(net184));
 sg13g2_inv_1 _1278_ (.Y(_0553_),
    .A(_0552_));
 sg13g2_nand4_1 _1279_ (.B(_0533_),
    .C(_0549_),
    .A(_0519_),
    .Y(_0554_),
    .D(_0552_));
 sg13g2_and2_1 _1280_ (.A(_0525_),
    .B(_0554_),
    .X(_0555_));
 sg13g2_nand2_1 _1281_ (.Y(_0556_),
    .A(_0525_),
    .B(_0554_));
 sg13g2_nand2_1 _1282_ (.Y(_0557_),
    .A(_0536_),
    .B(_0544_));
 sg13g2_nor2_1 _1283_ (.A(\hvsync_gen.hpos[0] ),
    .B(net160),
    .Y(_0558_));
 sg13g2_o21ai_1 _1284_ (.B1(net183),
    .Y(_0559_),
    .A1(_0161_),
    .A2(_0558_));
 sg13g2_o21ai_1 _1285_ (.B1(_0559_),
    .Y(_0560_),
    .A1(_0067_),
    .A2(net183));
 sg13g2_nand2_1 _1286_ (.Y(_0561_),
    .A(_0539_),
    .B(_0560_));
 sg13g2_inv_1 _1287_ (.Y(_0562_),
    .A(_0561_));
 sg13g2_nor2_1 _1288_ (.A(_0543_),
    .B(_0561_),
    .Y(_0563_));
 sg13g2_nand2_1 _1289_ (.Y(_0564_),
    .A(_0536_),
    .B(_0563_));
 sg13g2_nand3_1 _1290_ (.B(_0552_),
    .C(_0557_),
    .A(_0547_),
    .Y(_0565_));
 sg13g2_nand3_1 _1291_ (.B(_0531_),
    .C(_0565_),
    .A(_0528_),
    .Y(_0566_));
 sg13g2_nor2b_1 _1292_ (.A(_0524_),
    .B_N(_0519_),
    .Y(_0567_));
 sg13g2_o21ai_1 _1293_ (.B1(_0519_),
    .Y(_0568_),
    .A1(_0524_),
    .A2(_0566_));
 sg13g2_nor2_1 _1294_ (.A(_0539_),
    .B(_0543_),
    .Y(_0569_));
 sg13g2_nand2_1 _1295_ (.Y(_0570_),
    .A(_0536_),
    .B(_0569_));
 sg13g2_a21oi_1 _1296_ (.A1(_0547_),
    .A2(_0570_),
    .Y(_0571_),
    .B1(_0552_));
 sg13g2_a21o_1 _1297_ (.A2(_0571_),
    .A1(_0531_),
    .B1(_0528_),
    .X(_0572_));
 sg13g2_nand3_1 _1298_ (.B(_0567_),
    .C(_0572_),
    .A(_0566_),
    .Y(_0573_));
 sg13g2_o21ai_1 _1299_ (.B1(_0553_),
    .Y(_0574_),
    .A1(_0536_),
    .A2(_0569_));
 sg13g2_o21ai_1 _1300_ (.B1(_0574_),
    .Y(_0575_),
    .A1(_0547_),
    .A2(_0552_));
 sg13g2_nor2b_1 _1301_ (.A(_0575_),
    .B_N(_0524_),
    .Y(_0576_));
 sg13g2_a21o_1 _1302_ (.A2(_0576_),
    .A1(_0533_),
    .B1(_0519_),
    .X(_0577_));
 sg13g2_and2_1 _1303_ (.A(_0573_),
    .B(_0577_),
    .X(_0578_));
 sg13g2_o21ai_1 _1304_ (.B1(_0532_),
    .Y(_0579_),
    .A1(_0547_),
    .A2(_0574_));
 sg13g2_a21oi_1 _1305_ (.A1(_0528_),
    .A2(_0579_),
    .Y(_0580_),
    .B1(_0525_));
 sg13g2_or4_1 _1306_ (.A(_0533_),
    .B(_0547_),
    .C(_0557_),
    .D(_0562_),
    .X(_0581_));
 sg13g2_o21ai_1 _1307_ (.B1(_0552_),
    .Y(_0582_),
    .A1(_0547_),
    .A2(_0564_));
 sg13g2_a21oi_1 _1308_ (.A1(_0531_),
    .A2(_0582_),
    .Y(_0583_),
    .B1(_0528_));
 sg13g2_nand4_1 _1309_ (.B(_0524_),
    .C(_0581_),
    .A(_0519_),
    .Y(_0584_),
    .D(_0583_));
 sg13g2_a22oi_1 _1310_ (.Y(_0585_),
    .B1(_0580_),
    .B2(_0584_),
    .A2(_0578_),
    .A1(_0555_));
 sg13g2_nand2_1 _1311_ (.Y(_0586_),
    .A(_0299_),
    .B(_0585_));
 sg13g2_nor2b_2 _1312_ (.A(net163),
    .B_N(_0296_),
    .Y(_0587_));
 sg13g2_nand2b_1 _1313_ (.Y(_0588_),
    .B(_0296_),
    .A_N(net163));
 sg13g2_nand3_1 _1314_ (.B(_0586_),
    .C(_0588_),
    .A(_0308_),
    .Y(_0589_));
 sg13g2_a21oi_1 _1315_ (.A1(_0448_),
    .A2(_0589_),
    .Y(_0590_),
    .B1(_0454_));
 sg13g2_o21ai_1 _1316_ (.B1(_0590_),
    .Y(_0591_),
    .A1(_0441_),
    .A2(_0451_));
 sg13g2_a21oi_1 _1317_ (.A1(net181),
    .A2(net180),
    .Y(_0592_),
    .B1(net179));
 sg13g2_o21ai_1 _1318_ (.B1(_0287_),
    .Y(_0593_),
    .A1(_0063_),
    .A2(_0592_));
 sg13g2_nand2b_1 _1319_ (.Y(_0594_),
    .B(net180),
    .A_N(net181));
 sg13g2_nand2b_1 _1320_ (.Y(_0595_),
    .B(net178),
    .A_N(net179));
 sg13g2_nor2_1 _1321_ (.A(_0594_),
    .B(_0595_),
    .Y(_0596_));
 sg13g2_a22oi_1 _1322_ (.Y(_0597_),
    .B1(_0596_),
    .B2(_0287_),
    .A2(_0593_),
    .A1(net168));
 sg13g2_o21ai_1 _1323_ (.B1(_0061_),
    .Y(_0598_),
    .A1(_0285_),
    .A2(_0597_));
 sg13g2_nand2_1 _1324_ (.Y(_0599_),
    .A(net179),
    .B(net180));
 sg13g2_nand3_1 _1325_ (.B(net179),
    .C(net180),
    .A(net181),
    .Y(_0600_));
 sg13g2_nor2_1 _1326_ (.A(net178),
    .B(_0600_),
    .Y(_0601_));
 sg13g2_nand2_1 _1327_ (.Y(_0602_),
    .A(_0061_),
    .B(net168));
 sg13g2_nor4_1 _1328_ (.A(net169),
    .B(net173),
    .C(_0282_),
    .D(_0602_),
    .Y(_0603_));
 sg13g2_a21oi_1 _1329_ (.A1(_0601_),
    .A2(_0603_),
    .Y(_0604_),
    .B1(_0068_));
 sg13g2_a21o_1 _1330_ (.A2(net178),
    .A1(net176),
    .B1(net173),
    .X(_0605_));
 sg13g2_a21oi_1 _1331_ (.A1(net171),
    .A2(_0605_),
    .Y(_0606_),
    .B1(net169));
 sg13g2_o21ai_1 _1332_ (.B1(_0604_),
    .Y(_0607_),
    .A1(_0062_),
    .A2(_0606_));
 sg13g2_nand2b_1 _1333_ (.Y(_0608_),
    .B(net181),
    .A_N(net180));
 sg13g2_or4_1 _1334_ (.A(net176),
    .B(_0595_),
    .C(_0602_),
    .D(_0608_),
    .X(_0609_));
 sg13g2_nor3_1 _1335_ (.A(net175),
    .B(net179),
    .C(net180),
    .Y(_0610_));
 sg13g2_o21ai_1 _1336_ (.B1(net168),
    .Y(_0611_),
    .A1(net175),
    .A2(net178));
 sg13g2_o21ai_1 _1337_ (.B1(_0609_),
    .Y(_0612_),
    .A1(_0610_),
    .A2(_0611_));
 sg13g2_nand2b_1 _1338_ (.Y(_0613_),
    .B(_0612_),
    .A_N(_0286_));
 sg13g2_and4_1 _1339_ (.A(_0013_),
    .B(_0598_),
    .C(_0607_),
    .D(_0613_),
    .X(_0614_));
 sg13g2_inv_1 _1340_ (.Y(_0615_),
    .A(_0614_));
 sg13g2_and2_1 _1341_ (.A(_0299_),
    .B(_0573_),
    .X(_0616_));
 sg13g2_a22oi_1 _1342_ (.Y(_0617_),
    .B1(_0616_),
    .B2(_0584_),
    .A2(_0615_),
    .A1(_0304_));
 sg13g2_o21ai_1 _1343_ (.B1(_0448_),
    .Y(_0618_),
    .A1(_0587_),
    .A2(_0617_));
 sg13g2_o21ai_1 _1344_ (.B1(_0584_),
    .Y(_0619_),
    .A1(_0556_),
    .A2(_0568_));
 sg13g2_a22oi_1 _1345_ (.Y(_0620_),
    .B1(_0619_),
    .B2(_0587_),
    .A2(_0618_),
    .A1(_0455_));
 sg13g2_nand2_1 _1346_ (.Y(_0621_),
    .A(_0010_),
    .B(_0287_));
 sg13g2_nor4_1 _1347_ (.A(net169),
    .B(net172),
    .C(_0601_),
    .D(_0621_),
    .Y(_0622_));
 sg13g2_nand3b_1 _1348_ (.B(_0063_),
    .C(_0599_),
    .Y(_0623_),
    .A_N(net176));
 sg13g2_nand3b_1 _1349_ (.B(net173),
    .C(_0623_),
    .Y(_0624_),
    .A_N(net171));
 sg13g2_nand4_1 _1350_ (.B(_0002_),
    .C(_0280_),
    .A(\hvsync_gen.hpos[9] ),
    .Y(_0625_),
    .D(_0624_));
 sg13g2_nor3_1 _1351_ (.A(_0604_),
    .B(_0622_),
    .C(_0625_),
    .Y(_0626_));
 sg13g2_or2_1 _1352_ (.X(_0627_),
    .B(_0626_),
    .A(_0307_));
 sg13g2_o21ai_1 _1353_ (.B1(_0304_),
    .Y(_0628_),
    .A1(_0614_),
    .A2(_0627_));
 sg13g2_nand2_1 _1354_ (.Y(_0629_),
    .A(_0588_),
    .B(_0628_));
 sg13g2_a21oi_1 _1355_ (.A1(_0448_),
    .A2(_0629_),
    .Y(_0630_),
    .B1(_0454_));
 sg13g2_or2_1 _1356_ (.X(_0631_),
    .B(_0630_),
    .A(_0585_));
 sg13g2_and2_1 _1357_ (.A(_0628_),
    .B(_0631_),
    .X(_0632_));
 sg13g2_nand2_1 _1358_ (.Y(_0633_),
    .A(_0620_),
    .B(_0632_));
 sg13g2_or2_1 _1359_ (.X(_0634_),
    .B(_0632_),
    .A(_0620_));
 sg13g2_inv_1 _1360_ (.Y(_0635_),
    .A(_0634_));
 sg13g2_nor2_1 _1361_ (.A(_0299_),
    .B(_0307_),
    .Y(_0636_));
 sg13g2_a22oi_1 _1362_ (.Y(_0637_),
    .B1(_0607_),
    .B2(_0636_),
    .A2(_0578_),
    .A1(_0299_));
 sg13g2_or2_1 _1363_ (.X(_0638_),
    .B(_0637_),
    .A(_0587_));
 sg13g2_a21oi_1 _1364_ (.A1(_0555_),
    .A2(_0587_),
    .Y(_0639_),
    .B1(_0454_));
 sg13g2_and3_1 _1365_ (.X(_0640_),
    .A(_0448_),
    .B(_0638_),
    .C(_0639_));
 sg13g2_nand4_1 _1366_ (.B(_0633_),
    .C(_0634_),
    .A(_0310_),
    .Y(_0641_),
    .D(_0640_));
 sg13g2_o21ai_1 _1367_ (.B1(_0311_),
    .Y(uo_out[4]),
    .A1(_0591_),
    .A2(_0641_));
 sg13g2_nor3_1 _1368_ (.A(_0441_),
    .B(_0451_),
    .C(_0454_),
    .Y(_0642_));
 sg13g2_nor2_1 _1369_ (.A(_0455_),
    .B(_0555_),
    .Y(_0643_));
 sg13g2_nor3_2 _1370_ (.A(_0640_),
    .B(_0642_),
    .C(_0643_),
    .Y(_0644_));
 sg13g2_nand2_1 _1371_ (.Y(_0645_),
    .A(_0310_),
    .B(_0591_));
 sg13g2_nand3_1 _1372_ (.B(_0591_),
    .C(_0633_),
    .A(_0310_),
    .Y(_0646_));
 sg13g2_a21oi_2 _1373_ (.B1(_0646_),
    .Y(uo_out[0]),
    .A2(_0644_),
    .A1(_0635_));
 sg13g2_a21oi_2 _1374_ (.B1(_0645_),
    .Y(uo_out[1]),
    .A2(_0644_),
    .A1(_0634_));
 sg13g2_nand3_1 _1375_ (.B(_0620_),
    .C(_0632_),
    .A(_0310_),
    .Y(_0647_));
 sg13g2_o21ai_1 _1376_ (.B1(_0311_),
    .Y(uo_out[6]),
    .A1(_0591_),
    .A2(_0647_));
 sg13g2_nand2b_1 _1377_ (.Y(_0648_),
    .B(_0310_),
    .A_N(_0620_));
 sg13g2_nand3_1 _1378_ (.B(_0591_),
    .C(_0632_),
    .A(_0310_),
    .Y(_0649_));
 sg13g2_o21ai_1 _1379_ (.B1(_0649_),
    .Y(uo_out[2]),
    .A1(_0644_),
    .A2(_0648_));
 sg13g2_and2_1 _1380_ (.A(net187),
    .B(_0022_),
    .X(_0023_));
 sg13g2_and2_1 _1381_ (.A(net187),
    .B(_0468_),
    .X(_0024_));
 sg13g2_a21oi_2 _1382_ (.B1(\counter[2] ),
    .Y(_0650_),
    .A2(net160),
    .A1(net159));
 sg13g2_nand3_1 _1383_ (.B(net160),
    .C(\counter[2] ),
    .A(net159),
    .Y(_0651_));
 sg13g2_nand2b_1 _1384_ (.Y(_0652_),
    .B(_0651_),
    .A_N(_0650_));
 sg13g2_and2_1 _1385_ (.A(net187),
    .B(_0652_),
    .X(_0025_));
 sg13g2_nor2_1 _1386_ (.A(_0053_),
    .B(_0650_),
    .Y(_0653_));
 sg13g2_o21ai_1 _1387_ (.B1(net187),
    .Y(_0654_),
    .A1(_0053_),
    .A2(_0650_));
 sg13g2_a21oi_1 _1388_ (.A1(_0053_),
    .A2(_0650_),
    .Y(_0026_),
    .B1(_0654_));
 sg13g2_xor2_1 _1389_ (.B(_0653_),
    .A(\counter[4] ),
    .X(_0655_));
 sg13g2_and2_1 _1390_ (.A(net189),
    .B(_0655_),
    .X(_0027_));
 sg13g2_a21oi_1 _1391_ (.A1(\counter[4] ),
    .A2(_0653_),
    .Y(_0656_),
    .B1(\counter[5] ));
 sg13g2_nand3_1 _1392_ (.B(\counter[4] ),
    .C(_0653_),
    .A(\counter[5] ),
    .Y(_0657_));
 sg13g2_nand2_1 _1393_ (.Y(_0658_),
    .A(net189),
    .B(_0657_));
 sg13g2_nor2_1 _1394_ (.A(_0656_),
    .B(_0658_),
    .Y(_0028_));
 sg13g2_nor2_1 _1395_ (.A(_0017_),
    .B(_0657_),
    .Y(_0659_));
 sg13g2_o21ai_1 _1396_ (.B1(net189),
    .Y(_0660_),
    .A1(_0017_),
    .A2(_0657_));
 sg13g2_a21oi_1 _1397_ (.A1(_0017_),
    .A2(_0657_),
    .Y(_0029_),
    .B1(_0660_));
 sg13g2_nand2_1 _1398_ (.Y(_0661_),
    .A(\counter[7] ),
    .B(\counter[6] ));
 sg13g2_nor2_1 _1399_ (.A(_0657_),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_nand2_1 _1400_ (.Y(_0663_),
    .A(\counter[8] ),
    .B(_0662_));
 sg13g2_or2_1 _1401_ (.X(_0664_),
    .B(_0663_),
    .A(\counter[9] ));
 sg13g2_o21ai_1 _1402_ (.B1(_0664_),
    .Y(_0665_),
    .A1(\counter[8] ),
    .A2(_0662_));
 sg13g2_xnor2_1 _1403_ (.Y(_0666_),
    .A(_0016_),
    .B(_0659_));
 sg13g2_or3_1 _1404_ (.A(_0015_),
    .B(_0665_),
    .C(_0666_),
    .X(_0667_));
 sg13g2_nor2_1 _1405_ (.A(_0015_),
    .B(_0663_),
    .Y(_0668_));
 sg13g2_a21oi_1 _1406_ (.A1(_0015_),
    .A2(_0664_),
    .Y(_0669_),
    .B1(_0668_));
 sg13g2_nand2_1 _1407_ (.Y(_0670_),
    .A(\counter[9] ),
    .B(_0668_));
 sg13g2_nand2_1 _1408_ (.Y(_0671_),
    .A(_0666_),
    .B(_0670_));
 sg13g2_o21ai_1 _1409_ (.B1(_0667_),
    .Y(_0672_),
    .A1(_0669_),
    .A2(_0671_));
 sg13g2_and2_1 _1410_ (.A(net189),
    .B(_0672_),
    .X(_0030_));
 sg13g2_nor2_1 _1411_ (.A(_0665_),
    .B(_0668_),
    .Y(_0673_));
 sg13g2_nand2_1 _1412_ (.Y(_0674_),
    .A(_0667_),
    .B(_0673_));
 sg13g2_o21ai_1 _1413_ (.B1(_0674_),
    .Y(_0675_),
    .A1(_0666_),
    .A2(_0670_));
 sg13g2_and2_1 _1414_ (.A(net189),
    .B(_0675_),
    .X(_0031_));
 sg13g2_a21o_1 _1415_ (.A2(_0669_),
    .A1(_0665_),
    .B1(_0666_),
    .X(_0676_));
 sg13g2_and3_1 _1416_ (.X(_0032_),
    .A(net189),
    .B(_0671_),
    .C(_0676_));
 sg13g2_nor2_1 _1417_ (.A(_0063_),
    .B(_0600_),
    .Y(_0677_));
 sg13g2_and2_1 _1418_ (.A(net175),
    .B(_0677_),
    .X(_0678_));
 sg13g2_nor3_1 _1419_ (.A(\hvsync_gen.hpos[7] ),
    .B(net171),
    .C(net173),
    .Y(_0679_));
 sg13g2_and4_2 _1420_ (.A(\hvsync_gen.hpos[9] ),
    .B(net168),
    .C(_0678_),
    .D(_0679_),
    .X(_0680_));
 sg13g2_nor2b_2 _1421_ (.A(_0680_),
    .B_N(net188),
    .Y(_0681_));
 sg13g2_nand2b_2 _1422_ (.Y(_0682_),
    .B(net188),
    .A_N(_0680_));
 sg13g2_and2_1 _1423_ (.A(net47),
    .B(_0681_),
    .X(_0033_));
 sg13g2_a21oi_1 _1424_ (.A1(_0594_),
    .A2(_0608_),
    .Y(_0034_),
    .B1(_0682_));
 sg13g2_nand2_1 _1425_ (.Y(_0683_),
    .A(net187),
    .B(_0600_));
 sg13g2_nor2_1 _1426_ (.A(net74),
    .B(_0683_),
    .Y(_0035_));
 sg13g2_nand3_1 _1427_ (.B(net180),
    .C(_0065_),
    .A(net181),
    .Y(_0684_));
 sg13g2_xnor2_1 _1428_ (.Y(_0685_),
    .A(_0063_),
    .B(_0684_));
 sg13g2_nor2_1 _1429_ (.A(_0682_),
    .B(_0685_),
    .Y(_0036_));
 sg13g2_o21ai_1 _1430_ (.B1(net189),
    .Y(_0686_),
    .A1(net175),
    .A2(_0677_));
 sg13g2_nor2_1 _1431_ (.A(_0678_),
    .B(_0686_),
    .Y(_0037_));
 sg13g2_nor3_1 _1432_ (.A(_0063_),
    .B(net63),
    .C(_0600_),
    .Y(_0687_));
 sg13g2_xnor2_1 _1433_ (.Y(_0688_),
    .A(net174),
    .B(_0687_));
 sg13g2_nor2_1 _1434_ (.A(_0682_),
    .B(net64),
    .Y(_0038_));
 sg13g2_nand2_1 _1435_ (.Y(_0689_),
    .A(net173),
    .B(_0678_));
 sg13g2_xor2_1 _1436_ (.B(_0689_),
    .A(net172),
    .X(_0690_));
 sg13g2_nor2_1 _1437_ (.A(_0682_),
    .B(_0690_),
    .Y(_0039_));
 sg13g2_nor2_1 _1438_ (.A(net66),
    .B(_0689_),
    .Y(_0691_));
 sg13g2_o21ai_1 _1439_ (.B1(_0681_),
    .Y(_0692_),
    .A1(net170),
    .A2(_0691_));
 sg13g2_a21oi_1 _1440_ (.A1(net170),
    .A2(_0691_),
    .Y(_0040_),
    .B1(_0692_));
 sg13g2_nand2b_1 _1441_ (.Y(_0693_),
    .B(_0678_),
    .A_N(_0286_));
 sg13g2_xnor2_1 _1442_ (.Y(_0694_),
    .A(_0062_),
    .B(_0693_));
 sg13g2_nor2_1 _1443_ (.A(_0682_),
    .B(_0694_),
    .Y(_0041_));
 sg13g2_nor2_1 _1444_ (.A(net61),
    .B(_0693_),
    .Y(_0695_));
 sg13g2_o21ai_1 _1445_ (.B1(_0681_),
    .Y(_0696_),
    .A1(\hvsync_gen.hpos[9] ),
    .A2(_0695_));
 sg13g2_a21oi_1 _1446_ (.A1(\hvsync_gen.hpos[9] ),
    .A2(_0695_),
    .Y(_0042_),
    .B1(_0696_));
 sg13g2_nand2_1 _1447_ (.Y(_0697_),
    .A(\hvsync_gen.vpos[0] ),
    .B(_0681_));
 sg13g2_nand4_1 _1448_ (.B(_0055_),
    .C(net167),
    .A(net162),
    .Y(_0698_),
    .D(\hvsync_gen.vpos[2] ));
 sg13g2_nand2_1 _1449_ (.Y(_0699_),
    .A(_0292_),
    .B(_0444_));
 sg13g2_o21ai_1 _1450_ (.B1(net188),
    .Y(_0700_),
    .A1(_0698_),
    .A2(_0699_));
 sg13g2_nand2_1 _1451_ (.Y(_0701_),
    .A(net48),
    .B(_0680_));
 sg13g2_o21ai_1 _1452_ (.B1(_0697_),
    .Y(_0043_),
    .A1(_0700_),
    .A2(_0701_));
 sg13g2_nand2_1 _1453_ (.Y(_0702_),
    .A(\hvsync_gen.vpos[0] ),
    .B(net55));
 sg13g2_a21oi_1 _1454_ (.A1(\hvsync_gen.vpos[0] ),
    .A2(_0680_),
    .Y(_0703_),
    .B1(net55));
 sg13g2_nand2_1 _1455_ (.Y(_0704_),
    .A(net188),
    .B(_0702_));
 sg13g2_a21oi_1 _1456_ (.A1(_0682_),
    .A2(_0704_),
    .Y(_0044_),
    .B1(net56));
 sg13g2_nor2_1 _1457_ (.A(_0681_),
    .B(_0702_),
    .Y(_0705_));
 sg13g2_and2_2 _1458_ (.A(_0682_),
    .B(_0700_),
    .X(_0706_));
 sg13g2_xnor2_1 _1459_ (.Y(_0707_),
    .A(net65),
    .B(_0705_));
 sg13g2_nor2_1 _1460_ (.A(_0706_),
    .B(_0707_),
    .Y(_0045_));
 sg13g2_nor3_1 _1461_ (.A(net52),
    .B(_0681_),
    .C(_0702_),
    .Y(_0708_));
 sg13g2_xnor2_1 _1462_ (.Y(_0709_),
    .A(net167),
    .B(net53));
 sg13g2_nor2_1 _1463_ (.A(_0706_),
    .B(net54),
    .Y(_0046_));
 sg13g2_and3_1 _1464_ (.X(_0710_),
    .A(net167),
    .B(net65),
    .C(_0705_));
 sg13g2_and2_1 _1465_ (.A(net166),
    .B(_0710_),
    .X(_0711_));
 sg13g2_nor2_1 _1466_ (.A(net166),
    .B(_0710_),
    .Y(_0712_));
 sg13g2_nor3_1 _1467_ (.A(_0706_),
    .B(net158),
    .C(_0712_),
    .Y(_0047_));
 sg13g2_nor3_1 _1468_ (.A(_0056_),
    .B(_0706_),
    .C(net158),
    .Y(_0713_));
 sg13g2_nand4_1 _1469_ (.B(net166),
    .C(net187),
    .A(_0056_),
    .Y(_0714_),
    .D(_0710_));
 sg13g2_nand2b_1 _1470_ (.Y(_0048_),
    .B(_0714_),
    .A_N(_0713_));
 sg13g2_a21oi_1 _1471_ (.A1(net50),
    .A2(net158),
    .Y(_0715_),
    .B1(net164));
 sg13g2_nand3_1 _1472_ (.B(net50),
    .C(net158),
    .A(net164),
    .Y(_0716_));
 sg13g2_inv_1 _1473_ (.Y(_0717_),
    .A(_0716_));
 sg13g2_nor3_1 _1474_ (.A(_0706_),
    .B(_0715_),
    .C(_0717_),
    .Y(_0049_));
 sg13g2_nand3b_1 _1475_ (.B(_0716_),
    .C(\hvsync_gen.vpos[7] ),
    .Y(_0718_),
    .A_N(_0706_));
 sg13g2_nand3_1 _1476_ (.B(net187),
    .C(net158),
    .A(net50),
    .Y(_0719_));
 sg13g2_o21ai_1 _1477_ (.B1(_0718_),
    .Y(_0050_),
    .A1(_0290_),
    .A2(_0719_));
 sg13g2_a21oi_1 _1478_ (.A1(_0309_),
    .A2(_0711_),
    .Y(_0720_),
    .B1(_0706_));
 sg13g2_nand3_1 _1479_ (.B(_0078_),
    .C(net158),
    .A(net165),
    .Y(_0721_));
 sg13g2_a221oi_1 _1480_ (.B2(_0055_),
    .C1(_0706_),
    .B1(_0721_),
    .A1(_0309_),
    .Y(_0051_),
    .A2(net158));
 sg13g2_nand2_1 _1481_ (.Y(_0722_),
    .A(net163),
    .B(_0720_));
 sg13g2_nand4_1 _1482_ (.B(net187),
    .C(_0277_),
    .A(net165),
    .Y(_0723_),
    .D(net158));
 sg13g2_nand2_1 _1483_ (.Y(_0052_),
    .A(_0722_),
    .B(_0723_));
 sg13g2_dfrbp_1 _1484_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net27),
    .D(_0023_),
    .Q_N(_0022_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _1485_ (.CLK(net161),
    .RESET_B(net12),
    .D(_0024_),
    .Q_N(_0734_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _1486_ (.CLK(net161),
    .RESET_B(net11),
    .D(_0025_),
    .Q_N(_0733_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _1487_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net10),
    .D(_0026_),
    .Q_N(_0732_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _1488_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net9),
    .D(_0027_),
    .Q_N(_0731_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _1489_ (.CLK(net161),
    .RESET_B(net8),
    .D(_0028_),
    .Q_N(_0730_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _1490_ (.CLK(net161),
    .RESET_B(net7),
    .D(_0029_),
    .Q_N(_0017_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _1491_ (.CLK(net161),
    .RESET_B(net37),
    .D(_0030_),
    .Q_N(_0016_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _1492_ (.CLK(net161),
    .RESET_B(net36),
    .D(_0031_),
    .Q_N(_0018_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _1493_ (.CLK(net161),
    .RESET_B(net35),
    .D(_0032_),
    .Q_N(_0015_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 _1494_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net34),
    .D(_0033_),
    .Q_N(_0021_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 _1495_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net33),
    .D(net77),
    .Q_N(_0012_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _1496_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net32),
    .D(_0035_),
    .Q_N(_0011_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _1497_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net31),
    .D(_0036_),
    .Q_N(_0010_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _1498_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net30),
    .D(_0037_),
    .Q_N(_0009_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _1499_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net29),
    .D(_0038_),
    .Q_N(_0008_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _1500_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net28),
    .D(_0039_),
    .Q_N(_0002_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _1501_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net26),
    .D(net67),
    .Q_N(_0007_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _1502_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net25),
    .D(_0041_),
    .Q_N(_0019_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _1503_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net38),
    .D(net62),
    .Q_N(_0013_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _1504_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net24),
    .D(net72),
    .Q_N(_0729_),
    .Q(hsync));
 sg13g2_dfrbp_1 _1505_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net23),
    .D(net49),
    .Q_N(_0020_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _1506_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net21),
    .D(net57),
    .Q_N(_0006_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _1507_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net19),
    .D(_0045_),
    .Q_N(_0005_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _1508_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net17),
    .D(_0046_),
    .Q_N(_0004_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _1509_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net15),
    .D(_0047_),
    .Q_N(_0728_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _1510_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net13),
    .D(_0048_),
    .Q_N(_0003_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _1511_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net20),
    .D(_0049_),
    .Q_N(_0727_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _1512_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net16),
    .D(net51),
    .Q_N(_0726_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _1513_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net22),
    .D(_0051_),
    .Q_N(_0725_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _1514_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net18),
    .D(_0052_),
    .Q_N(_0014_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _1515_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net14),
    .D(net60),
    .Q_N(_0724_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_tiehi _1489__8 (.L_HI(net8));
 sg13g2_tiehi _1488__9 (.L_HI(net9));
 sg13g2_tiehi _1487__10 (.L_HI(net10));
 sg13g2_tiehi _1486__11 (.L_HI(net11));
 sg13g2_tiehi _1485__12 (.L_HI(net12));
 sg13g2_tiehi _1510__13 (.L_HI(net13));
 sg13g2_tiehi _1515__14 (.L_HI(net14));
 sg13g2_tiehi _1509__15 (.L_HI(net15));
 sg13g2_tiehi _1512__16 (.L_HI(net16));
 sg13g2_tiehi _1508__17 (.L_HI(net17));
 sg13g2_tiehi _1514__18 (.L_HI(net18));
 sg13g2_tiehi _1507__19 (.L_HI(net19));
 sg13g2_tiehi _1511__20 (.L_HI(net20));
 sg13g2_tiehi _1506__21 (.L_HI(net21));
 sg13g2_tiehi _1513__22 (.L_HI(net22));
 sg13g2_tiehi _1505__23 (.L_HI(net23));
 sg13g2_tiehi _1504__24 (.L_HI(net24));
 sg13g2_tiehi _1502__25 (.L_HI(net25));
 sg13g2_tiehi _1501__26 (.L_HI(net26));
 sg13g2_tiehi _1484__27 (.L_HI(net27));
 sg13g2_tiehi _1500__28 (.L_HI(net28));
 sg13g2_tiehi _1499__29 (.L_HI(net29));
 sg13g2_tiehi _1498__30 (.L_HI(net30));
 sg13g2_tiehi _1497__31 (.L_HI(net31));
 sg13g2_tiehi _1496__32 (.L_HI(net32));
 sg13g2_tiehi _1495__33 (.L_HI(net33));
 sg13g2_tiehi _1494__34 (.L_HI(net34));
 sg13g2_tiehi _1493__35 (.L_HI(net35));
 sg13g2_tiehi _1492__36 (.L_HI(net36));
 sg13g2_tiehi _1491__37 (.L_HI(net37));
 sg13g2_tiehi _1503__38 (.L_HI(net38));
 sg13g2_tiehi tt_um_rebeccargb_colorbars_39 (.L_HI(net39));
 sg13g2_tiehi tt_um_rebeccargb_colorbars_40 (.L_HI(net40));
 sg13g2_tiehi tt_um_rebeccargb_colorbars_41 (.L_HI(net41));
 sg13g2_tiehi tt_um_rebeccargb_colorbars_42 (.L_HI(net42));
 sg13g2_tiehi tt_um_rebeccargb_colorbars_43 (.L_HI(net43));
 sg13g2_tiehi tt_um_rebeccargb_colorbars_44 (.L_HI(net44));
 sg13g2_tiehi tt_um_rebeccargb_colorbars_45 (.L_HI(net45));
 sg13g2_tiehi tt_um_rebeccargb_colorbars_46 (.L_HI(net46));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 _1556_ (.A(net161),
    .X(uo_out[3]));
 sg13g2_buf_1 _1557_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout145 (.A(_0320_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(uio_out[4]),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(net147),
    .X(uio_out[4]));
 sg13g2_buf_2 fanout148 (.A(_0271_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_0156_),
    .X(net149));
 sg13g2_buf_1 fanout150 (.A(_0156_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(net152),
    .X(uio_out[5]));
 sg13g2_buf_2 fanout152 (.A(net151),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(net154),
    .X(uio_out[2]));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(_0241_));
 sg13g2_buf_2 fanout156 (.A(_0241_),
    .X(net156));
 sg13g2_buf_4 fanout157 (.X(uio_out[7]),
    .A(net157));
 sg13g2_buf_2 fanout158 (.A(_0711_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(\counter[1] ),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(\counter[0] ),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(\hvsync_gen.vsync ),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(net163),
    .X(net162));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(net69));
 sg13g2_buf_2 fanout164 (.A(net58),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(net50),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(net75),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(\hvsync_gen.vpos[3] ),
    .X(net167));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(\hvsync_gen.hpos[8] ));
 sg13g2_buf_2 fanout169 (.A(\hvsync_gen.hpos[7] ),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(\hvsync_gen.hpos[7] ),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(net70));
 sg13g2_buf_2 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(\hvsync_gen.hpos[5] ),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(net177),
    .X(net175));
 sg13g2_buf_1 fanout176 (.A(net177),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(\hvsync_gen.hpos[4] ),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(\hvsync_gen.hpos[3] ),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(net73),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(\hvsync_gen.hpos[1] ),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(net76),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(net184),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(net184),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(ui_in[3]),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(ui_in[2]),
    .X(net186));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(rst_n));
 sg13g2_buf_2 fanout188 (.A(net189),
    .X(net188));
 sg13g2_buf_4 fanout189 (.X(net189),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_tiehi _1490__7 (.L_HI(net7));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0021_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0020_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0043_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold4 (.A(\hvsync_gen.vpos[5] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0050_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0005_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0708_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0709_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold9 (.A(\hvsync_gen.vpos[1] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0703_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0044_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold12 (.A(\hvsync_gen.vpos[6] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold13 (.A(\hvsync_gen.vpos[8] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0001_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0019_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0042_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0009_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0688_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold19 (.A(\hvsync_gen.vpos[2] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0002_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0040_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0011_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold23 (.A(\hvsync_gen.vpos[9] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold24 (.A(\hvsync_gen.hpos[6] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0013_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0000_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold27 (.A(\hvsync_gen.hpos[2] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0592_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold29 (.A(\hvsync_gen.vpos[4] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold30 (.A(\hvsync_gen.hpos[0] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0034_),
    .X(net77));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_fill_2 FILLER_13_105 ();
 sg13g2_fill_1 FILLER_13_107 ();
 sg13g2_decap_8 FILLER_13_113 ();
 sg13g2_decap_8 FILLER_13_120 ();
 sg13g2_decap_8 FILLER_13_127 ();
 sg13g2_decap_8 FILLER_13_138 ();
 sg13g2_decap_8 FILLER_13_145 ();
 sg13g2_decap_8 FILLER_13_152 ();
 sg13g2_decap_8 FILLER_13_159 ();
 sg13g2_decap_8 FILLER_13_166 ();
 sg13g2_decap_8 FILLER_13_173 ();
 sg13g2_decap_8 FILLER_13_180 ();
 sg13g2_decap_8 FILLER_13_187 ();
 sg13g2_decap_8 FILLER_13_194 ();
 sg13g2_decap_8 FILLER_13_201 ();
 sg13g2_decap_8 FILLER_13_208 ();
 sg13g2_decap_8 FILLER_13_215 ();
 sg13g2_decap_8 FILLER_13_222 ();
 sg13g2_decap_8 FILLER_13_229 ();
 sg13g2_decap_8 FILLER_13_236 ();
 sg13g2_decap_8 FILLER_13_243 ();
 sg13g2_decap_8 FILLER_13_250 ();
 sg13g2_decap_8 FILLER_13_257 ();
 sg13g2_decap_8 FILLER_13_264 ();
 sg13g2_decap_8 FILLER_13_271 ();
 sg13g2_decap_8 FILLER_13_278 ();
 sg13g2_decap_8 FILLER_13_285 ();
 sg13g2_decap_8 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_299 ();
 sg13g2_decap_8 FILLER_13_306 ();
 sg13g2_decap_8 FILLER_13_313 ();
 sg13g2_decap_8 FILLER_13_320 ();
 sg13g2_decap_8 FILLER_13_327 ();
 sg13g2_decap_8 FILLER_13_334 ();
 sg13g2_decap_8 FILLER_13_341 ();
 sg13g2_decap_8 FILLER_13_348 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_decap_8 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_fill_1 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_76 ();
 sg13g2_decap_8 FILLER_14_87 ();
 sg13g2_decap_4 FILLER_14_94 ();
 sg13g2_fill_2 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_162 ();
 sg13g2_fill_2 FILLER_14_169 ();
 sg13g2_fill_1 FILLER_14_171 ();
 sg13g2_fill_2 FILLER_14_229 ();
 sg13g2_fill_2 FILLER_14_278 ();
 sg13g2_fill_1 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_286 ();
 sg13g2_decap_8 FILLER_14_293 ();
 sg13g2_decap_8 FILLER_14_300 ();
 sg13g2_decap_8 FILLER_14_307 ();
 sg13g2_decap_8 FILLER_14_314 ();
 sg13g2_decap_8 FILLER_14_321 ();
 sg13g2_decap_8 FILLER_14_328 ();
 sg13g2_decap_8 FILLER_14_335 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_356 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_fill_1 FILLER_15_56 ();
 sg13g2_fill_1 FILLER_15_65 ();
 sg13g2_fill_1 FILLER_15_71 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_fill_2 FILLER_15_113 ();
 sg13g2_fill_1 FILLER_15_115 ();
 sg13g2_decap_8 FILLER_15_120 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_decap_4 FILLER_15_138 ();
 sg13g2_fill_2 FILLER_15_146 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_fill_2 FILLER_15_154 ();
 sg13g2_fill_2 FILLER_15_166 ();
 sg13g2_decap_4 FILLER_15_176 ();
 sg13g2_fill_1 FILLER_15_180 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_187 ();
 sg13g2_decap_8 FILLER_15_192 ();
 sg13g2_fill_1 FILLER_15_199 ();
 sg13g2_decap_8 FILLER_15_218 ();
 sg13g2_decap_4 FILLER_15_225 ();
 sg13g2_fill_1 FILLER_15_229 ();
 sg13g2_decap_8 FILLER_15_237 ();
 sg13g2_fill_1 FILLER_15_262 ();
 sg13g2_decap_8 FILLER_15_267 ();
 sg13g2_decap_8 FILLER_15_274 ();
 sg13g2_decap_4 FILLER_15_291 ();
 sg13g2_decap_8 FILLER_15_299 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_313 ();
 sg13g2_decap_8 FILLER_15_320 ();
 sg13g2_decap_8 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_decap_8 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_decap_8 FILLER_15_369 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_79 ();
 sg13g2_fill_2 FILLER_16_86 ();
 sg13g2_decap_4 FILLER_16_96 ();
 sg13g2_fill_2 FILLER_16_100 ();
 sg13g2_decap_4 FILLER_16_106 ();
 sg13g2_fill_1 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_125 ();
 sg13g2_fill_1 FILLER_16_127 ();
 sg13g2_decap_4 FILLER_16_133 ();
 sg13g2_fill_2 FILLER_16_137 ();
 sg13g2_fill_1 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_167 ();
 sg13g2_decap_4 FILLER_16_174 ();
 sg13g2_fill_1 FILLER_16_178 ();
 sg13g2_decap_8 FILLER_16_187 ();
 sg13g2_fill_2 FILLER_16_207 ();
 sg13g2_fill_1 FILLER_16_225 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_fill_1 FILLER_16_252 ();
 sg13g2_decap_4 FILLER_16_271 ();
 sg13g2_fill_2 FILLER_16_275 ();
 sg13g2_decap_8 FILLER_16_311 ();
 sg13g2_decap_8 FILLER_16_318 ();
 sg13g2_decap_8 FILLER_16_325 ();
 sg13g2_decap_8 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_4 FILLER_17_49 ();
 sg13g2_fill_2 FILLER_17_62 ();
 sg13g2_fill_1 FILLER_17_64 ();
 sg13g2_fill_1 FILLER_17_100 ();
 sg13g2_fill_2 FILLER_17_123 ();
 sg13g2_fill_1 FILLER_17_137 ();
 sg13g2_fill_1 FILLER_17_143 ();
 sg13g2_fill_1 FILLER_17_149 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_fill_1 FILLER_17_172 ();
 sg13g2_decap_4 FILLER_17_214 ();
 sg13g2_fill_2 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_228 ();
 sg13g2_fill_2 FILLER_17_242 ();
 sg13g2_fill_1 FILLER_17_244 ();
 sg13g2_decap_4 FILLER_17_249 ();
 sg13g2_fill_2 FILLER_17_253 ();
 sg13g2_decap_8 FILLER_17_272 ();
 sg13g2_fill_2 FILLER_17_279 ();
 sg13g2_fill_1 FILLER_17_281 ();
 sg13g2_decap_8 FILLER_17_290 ();
 sg13g2_fill_1 FILLER_17_297 ();
 sg13g2_decap_8 FILLER_17_303 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_316 ();
 sg13g2_decap_8 FILLER_17_323 ();
 sg13g2_decap_8 FILLER_17_330 ();
 sg13g2_decap_8 FILLER_17_337 ();
 sg13g2_decap_8 FILLER_17_344 ();
 sg13g2_decap_8 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_358 ();
 sg13g2_decap_8 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_4 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_58 ();
 sg13g2_fill_1 FILLER_18_71 ();
 sg13g2_decap_4 FILLER_18_97 ();
 sg13g2_fill_2 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_107 ();
 sg13g2_fill_2 FILLER_18_112 ();
 sg13g2_fill_1 FILLER_18_114 ();
 sg13g2_fill_2 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_135 ();
 sg13g2_fill_1 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_4 FILLER_18_175 ();
 sg13g2_fill_2 FILLER_18_179 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_4 FILLER_18_196 ();
 sg13g2_fill_2 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_215 ();
 sg13g2_fill_1 FILLER_18_222 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_fill_1 FILLER_18_277 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_decap_8 FILLER_18_332 ();
 sg13g2_decap_8 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_4 FILLER_19_49 ();
 sg13g2_fill_2 FILLER_19_84 ();
 sg13g2_fill_1 FILLER_19_115 ();
 sg13g2_decap_8 FILLER_19_134 ();
 sg13g2_fill_1 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_155 ();
 sg13g2_fill_2 FILLER_19_161 ();
 sg13g2_fill_2 FILLER_19_189 ();
 sg13g2_fill_1 FILLER_19_191 ();
 sg13g2_fill_1 FILLER_19_218 ();
 sg13g2_fill_1 FILLER_19_261 ();
 sg13g2_decap_4 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_fill_2 FILLER_20_70 ();
 sg13g2_fill_1 FILLER_20_72 ();
 sg13g2_fill_1 FILLER_20_78 ();
 sg13g2_decap_8 FILLER_20_87 ();
 sg13g2_decap_4 FILLER_20_94 ();
 sg13g2_fill_2 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_106 ();
 sg13g2_decap_8 FILLER_20_113 ();
 sg13g2_fill_1 FILLER_20_120 ();
 sg13g2_decap_4 FILLER_20_124 ();
 sg13g2_fill_1 FILLER_20_128 ();
 sg13g2_decap_8 FILLER_20_167 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_211 ();
 sg13g2_decap_8 FILLER_20_218 ();
 sg13g2_decap_4 FILLER_20_225 ();
 sg13g2_fill_1 FILLER_20_229 ();
 sg13g2_fill_1 FILLER_20_234 ();
 sg13g2_decap_4 FILLER_20_240 ();
 sg13g2_fill_1 FILLER_20_244 ();
 sg13g2_fill_2 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_279 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_decap_8 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_314 ();
 sg13g2_decap_8 FILLER_20_321 ();
 sg13g2_decap_8 FILLER_20_328 ();
 sg13g2_decap_8 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_342 ();
 sg13g2_decap_8 FILLER_20_349 ();
 sg13g2_decap_8 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_fill_2 FILLER_21_63 ();
 sg13g2_fill_1 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_79 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_111 ();
 sg13g2_decap_8 FILLER_21_146 ();
 sg13g2_fill_2 FILLER_21_153 ();
 sg13g2_fill_2 FILLER_21_159 ();
 sg13g2_fill_2 FILLER_21_166 ();
 sg13g2_fill_1 FILLER_21_172 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_fill_1 FILLER_21_186 ();
 sg13g2_fill_1 FILLER_21_195 ();
 sg13g2_decap_8 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_221 ();
 sg13g2_fill_2 FILLER_21_259 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_278 ();
 sg13g2_fill_1 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_303 ();
 sg13g2_decap_8 FILLER_21_310 ();
 sg13g2_decap_8 FILLER_21_317 ();
 sg13g2_decap_8 FILLER_21_324 ();
 sg13g2_decap_8 FILLER_21_331 ();
 sg13g2_decap_8 FILLER_21_338 ();
 sg13g2_decap_8 FILLER_21_345 ();
 sg13g2_decap_8 FILLER_21_352 ();
 sg13g2_decap_8 FILLER_21_359 ();
 sg13g2_decap_8 FILLER_21_366 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_4 FILLER_22_56 ();
 sg13g2_fill_1 FILLER_22_60 ();
 sg13g2_fill_2 FILLER_22_76 ();
 sg13g2_fill_1 FILLER_22_78 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_decap_4 FILLER_22_109 ();
 sg13g2_fill_1 FILLER_22_125 ();
 sg13g2_fill_1 FILLER_22_144 ();
 sg13g2_fill_2 FILLER_22_158 ();
 sg13g2_fill_1 FILLER_22_160 ();
 sg13g2_decap_4 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_192 ();
 sg13g2_fill_2 FILLER_22_200 ();
 sg13g2_fill_2 FILLER_22_206 ();
 sg13g2_decap_4 FILLER_22_230 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_fill_2 FILLER_22_245 ();
 sg13g2_fill_1 FILLER_22_247 ();
 sg13g2_fill_1 FILLER_22_266 ();
 sg13g2_decap_4 FILLER_22_288 ();
 sg13g2_decap_8 FILLER_22_300 ();
 sg13g2_decap_8 FILLER_22_307 ();
 sg13g2_decap_8 FILLER_22_314 ();
 sg13g2_decap_8 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_4 FILLER_23_56 ();
 sg13g2_fill_2 FILLER_23_60 ();
 sg13g2_fill_2 FILLER_23_78 ();
 sg13g2_fill_1 FILLER_23_80 ();
 sg13g2_decap_8 FILLER_23_86 ();
 sg13g2_fill_2 FILLER_23_93 ();
 sg13g2_fill_2 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_163 ();
 sg13g2_decap_8 FILLER_23_173 ();
 sg13g2_decap_8 FILLER_23_180 ();
 sg13g2_fill_2 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_203 ();
 sg13g2_fill_2 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_230 ();
 sg13g2_fill_1 FILLER_23_232 ();
 sg13g2_decap_8 FILLER_23_253 ();
 sg13g2_fill_1 FILLER_23_260 ();
 sg13g2_decap_4 FILLER_23_280 ();
 sg13g2_fill_1 FILLER_23_284 ();
 sg13g2_fill_1 FILLER_23_289 ();
 sg13g2_decap_8 FILLER_23_316 ();
 sg13g2_decap_8 FILLER_23_323 ();
 sg13g2_decap_8 FILLER_23_330 ();
 sg13g2_decap_8 FILLER_23_337 ();
 sg13g2_decap_8 FILLER_23_344 ();
 sg13g2_decap_8 FILLER_23_351 ();
 sg13g2_decap_8 FILLER_23_358 ();
 sg13g2_decap_8 FILLER_23_365 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_68 ();
 sg13g2_decap_4 FILLER_24_90 ();
 sg13g2_fill_1 FILLER_24_94 ();
 sg13g2_decap_4 FILLER_24_115 ();
 sg13g2_fill_2 FILLER_24_124 ();
 sg13g2_fill_2 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_138 ();
 sg13g2_decap_4 FILLER_24_148 ();
 sg13g2_fill_1 FILLER_24_152 ();
 sg13g2_fill_1 FILLER_24_158 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_fill_1 FILLER_24_175 ();
 sg13g2_fill_2 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_191 ();
 sg13g2_decap_8 FILLER_24_233 ();
 sg13g2_fill_1 FILLER_24_240 ();
 sg13g2_fill_2 FILLER_24_258 ();
 sg13g2_decap_8 FILLER_24_326 ();
 sg13g2_decap_8 FILLER_24_333 ();
 sg13g2_decap_8 FILLER_24_340 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_decap_8 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_361 ();
 sg13g2_decap_8 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_fill_2 FILLER_25_56 ();
 sg13g2_fill_1 FILLER_25_58 ();
 sg13g2_fill_2 FILLER_25_67 ();
 sg13g2_fill_1 FILLER_25_69 ();
 sg13g2_decap_8 FILLER_25_92 ();
 sg13g2_decap_4 FILLER_25_99 ();
 sg13g2_fill_1 FILLER_25_103 ();
 sg13g2_fill_1 FILLER_25_108 ();
 sg13g2_fill_2 FILLER_25_123 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_fill_2 FILLER_25_172 ();
 sg13g2_decap_8 FILLER_25_179 ();
 sg13g2_fill_2 FILLER_25_186 ();
 sg13g2_fill_1 FILLER_25_188 ();
 sg13g2_decap_4 FILLER_25_204 ();
 sg13g2_fill_1 FILLER_25_208 ();
 sg13g2_decap_8 FILLER_25_228 ();
 sg13g2_decap_4 FILLER_25_235 ();
 sg13g2_fill_2 FILLER_25_239 ();
 sg13g2_fill_2 FILLER_25_256 ();
 sg13g2_fill_1 FILLER_25_258 ();
 sg13g2_decap_4 FILLER_25_280 ();
 sg13g2_fill_2 FILLER_25_284 ();
 sg13g2_decap_4 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_8 FILLER_25_338 ();
 sg13g2_decap_8 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_352 ();
 sg13g2_decap_8 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_366 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_380 ();
 sg13g2_decap_8 FILLER_25_387 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_fill_2 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_58 ();
 sg13g2_fill_2 FILLER_26_83 ();
 sg13g2_decap_4 FILLER_26_97 ();
 sg13g2_fill_1 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_110 ();
 sg13g2_decap_8 FILLER_26_121 ();
 sg13g2_fill_2 FILLER_26_128 ();
 sg13g2_fill_1 FILLER_26_130 ();
 sg13g2_fill_2 FILLER_26_153 ();
 sg13g2_fill_1 FILLER_26_155 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_168 ();
 sg13g2_fill_2 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_209 ();
 sg13g2_fill_2 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_228 ();
 sg13g2_fill_1 FILLER_26_230 ();
 sg13g2_decap_8 FILLER_26_248 ();
 sg13g2_fill_2 FILLER_26_260 ();
 sg13g2_fill_1 FILLER_26_262 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_70 ();
 sg13g2_fill_1 FILLER_27_72 ();
 sg13g2_decap_4 FILLER_27_78 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_decap_4 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_95 ();
 sg13g2_fill_1 FILLER_27_120 ();
 sg13g2_fill_2 FILLER_27_133 ();
 sg13g2_fill_1 FILLER_27_135 ();
 sg13g2_decap_4 FILLER_27_140 ();
 sg13g2_decap_4 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_184 ();
 sg13g2_decap_4 FILLER_27_212 ();
 sg13g2_fill_1 FILLER_27_216 ();
 sg13g2_fill_1 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_254 ();
 sg13g2_fill_1 FILLER_27_256 ();
 sg13g2_decap_8 FILLER_27_269 ();
 sg13g2_fill_2 FILLER_27_276 ();
 sg13g2_fill_1 FILLER_27_278 ();
 sg13g2_fill_2 FILLER_27_324 ();
 sg13g2_fill_1 FILLER_27_326 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_fill_1 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_117 ();
 sg13g2_fill_1 FILLER_28_124 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_fill_2 FILLER_28_178 ();
 sg13g2_decap_8 FILLER_28_223 ();
 sg13g2_fill_2 FILLER_28_230 ();
 sg13g2_fill_1 FILLER_28_237 ();
 sg13g2_decap_4 FILLER_28_246 ();
 sg13g2_fill_2 FILLER_28_250 ();
 sg13g2_fill_1 FILLER_28_257 ();
 sg13g2_decap_4 FILLER_28_263 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_fill_2 FILLER_28_294 ();
 sg13g2_decap_4 FILLER_28_302 ();
 sg13g2_fill_2 FILLER_28_306 ();
 sg13g2_fill_2 FILLER_28_313 ();
 sg13g2_fill_2 FILLER_28_352 ();
 sg13g2_decap_4 FILLER_28_374 ();
 sg13g2_fill_1 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_4 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_124 ();
 sg13g2_decap_4 FILLER_29_131 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_192 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_decap_8 FILLER_29_209 ();
 sg13g2_decap_4 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_220 ();
 sg13g2_fill_2 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_229 ();
 sg13g2_fill_1 FILLER_29_254 ();
 sg13g2_fill_2 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_295 ();
 sg13g2_fill_2 FILLER_29_301 ();
 sg13g2_fill_1 FILLER_29_313 ();
 sg13g2_decap_4 FILLER_29_348 ();
 sg13g2_fill_1 FILLER_29_352 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_4 FILLER_30_98 ();
 sg13g2_fill_1 FILLER_30_129 ();
 sg13g2_fill_2 FILLER_30_138 ();
 sg13g2_fill_2 FILLER_30_200 ();
 sg13g2_decap_4 FILLER_30_215 ();
 sg13g2_decap_4 FILLER_30_237 ();
 sg13g2_decap_8 FILLER_30_246 ();
 sg13g2_fill_1 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_fill_1 FILLER_30_261 ();
 sg13g2_fill_2 FILLER_30_282 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_fill_1 FILLER_30_294 ();
 sg13g2_fill_1 FILLER_30_299 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_decap_4 FILLER_30_327 ();
 sg13g2_fill_2 FILLER_30_331 ();
 sg13g2_fill_2 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_1 FILLER_30_377 ();
 sg13g2_fill_1 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_fill_1 FILLER_31_116 ();
 sg13g2_decap_8 FILLER_31_122 ();
 sg13g2_decap_4 FILLER_31_129 ();
 sg13g2_fill_2 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_139 ();
 sg13g2_decap_8 FILLER_31_149 ();
 sg13g2_decap_4 FILLER_31_156 ();
 sg13g2_fill_1 FILLER_31_165 ();
 sg13g2_decap_4 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_183 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_fill_2 FILLER_31_200 ();
 sg13g2_fill_1 FILLER_31_202 ();
 sg13g2_fill_2 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_209 ();
 sg13g2_decap_8 FILLER_31_235 ();
 sg13g2_decap_8 FILLER_31_242 ();
 sg13g2_fill_2 FILLER_31_249 ();
 sg13g2_fill_1 FILLER_31_251 ();
 sg13g2_fill_2 FILLER_31_280 ();
 sg13g2_fill_1 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_fill_1 FILLER_31_312 ();
 sg13g2_fill_1 FILLER_31_319 ();
 sg13g2_fill_2 FILLER_31_334 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_fill_2 FILLER_32_112 ();
 sg13g2_fill_1 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_151 ();
 sg13g2_decap_4 FILLER_32_158 ();
 sg13g2_fill_2 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_182 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_decap_8 FILLER_32_205 ();
 sg13g2_decap_4 FILLER_32_212 ();
 sg13g2_fill_2 FILLER_32_216 ();
 sg13g2_fill_2 FILLER_32_254 ();
 sg13g2_fill_2 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_280 ();
 sg13g2_fill_1 FILLER_32_304 ();
 sg13g2_fill_2 FILLER_32_323 ();
 sg13g2_fill_2 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_346 ();
 sg13g2_decap_8 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_375 ();
 sg13g2_decap_8 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_fill_2 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_114 ();
 sg13g2_fill_2 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_133 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_fill_2 FILLER_33_164 ();
 sg13g2_fill_1 FILLER_33_176 ();
 sg13g2_fill_2 FILLER_33_182 ();
 sg13g2_fill_2 FILLER_33_192 ();
 sg13g2_decap_4 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_225 ();
 sg13g2_decap_4 FILLER_33_232 ();
 sg13g2_fill_1 FILLER_33_236 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_fill_2 FILLER_33_252 ();
 sg13g2_fill_1 FILLER_33_254 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_decap_4 FILLER_33_268 ();
 sg13g2_fill_1 FILLER_33_272 ();
 sg13g2_fill_1 FILLER_33_282 ();
 sg13g2_fill_2 FILLER_33_309 ();
 sg13g2_decap_4 FILLER_33_336 ();
 sg13g2_fill_1 FILLER_33_340 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_decap_8 FILLER_33_356 ();
 sg13g2_fill_1 FILLER_33_363 ();
 sg13g2_fill_2 FILLER_33_376 ();
 sg13g2_fill_1 FILLER_33_378 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_fill_2 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_132 ();
 sg13g2_decap_4 FILLER_34_143 ();
 sg13g2_decap_4 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_157 ();
 sg13g2_fill_1 FILLER_34_171 ();
 sg13g2_fill_1 FILLER_34_182 ();
 sg13g2_fill_2 FILLER_34_193 ();
 sg13g2_fill_2 FILLER_34_230 ();
 sg13g2_fill_2 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_252 ();
 sg13g2_fill_1 FILLER_34_348 ();
 sg13g2_decap_4 FILLER_34_358 ();
 sg13g2_fill_1 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_fill_1 FILLER_35_137 ();
 sg13g2_fill_2 FILLER_35_150 ();
 sg13g2_fill_1 FILLER_35_152 ();
 sg13g2_decap_8 FILLER_35_159 ();
 sg13g2_fill_1 FILLER_35_166 ();
 sg13g2_decap_4 FILLER_35_181 ();
 sg13g2_fill_2 FILLER_35_191 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_fill_1 FILLER_35_206 ();
 sg13g2_fill_1 FILLER_35_215 ();
 sg13g2_fill_2 FILLER_35_226 ();
 sg13g2_fill_1 FILLER_35_228 ();
 sg13g2_decap_4 FILLER_35_234 ();
 sg13g2_decap_4 FILLER_35_255 ();
 sg13g2_fill_2 FILLER_35_259 ();
 sg13g2_fill_2 FILLER_35_275 ();
 sg13g2_fill_2 FILLER_35_280 ();
 sg13g2_fill_2 FILLER_35_290 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_326 ();
 sg13g2_fill_2 FILLER_35_333 ();
 sg13g2_fill_1 FILLER_35_335 ();
 sg13g2_fill_2 FILLER_35_349 ();
 sg13g2_decap_8 FILLER_35_359 ();
 sg13g2_decap_8 FILLER_35_366 ();
 sg13g2_fill_1 FILLER_35_373 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_fill_1 FILLER_35_391 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_4 FILLER_36_112 ();
 sg13g2_fill_2 FILLER_36_116 ();
 sg13g2_fill_2 FILLER_36_129 ();
 sg13g2_decap_4 FILLER_36_140 ();
 sg13g2_fill_1 FILLER_36_144 ();
 sg13g2_decap_8 FILLER_36_159 ();
 sg13g2_decap_8 FILLER_36_176 ();
 sg13g2_fill_2 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_189 ();
 sg13g2_decap_4 FILLER_36_204 ();
 sg13g2_fill_1 FILLER_36_212 ();
 sg13g2_decap_8 FILLER_36_223 ();
 sg13g2_fill_2 FILLER_36_230 ();
 sg13g2_fill_2 FILLER_36_237 ();
 sg13g2_fill_1 FILLER_36_239 ();
 sg13g2_decap_8 FILLER_36_250 ();
 sg13g2_fill_2 FILLER_36_257 ();
 sg13g2_fill_2 FILLER_36_272 ();
 sg13g2_fill_1 FILLER_36_281 ();
 sg13g2_fill_1 FILLER_36_303 ();
 sg13g2_decap_4 FILLER_36_340 ();
 sg13g2_fill_1 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_358 ();
 sg13g2_fill_1 FILLER_36_360 ();
 sg13g2_fill_1 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_377 ();
 sg13g2_decap_4 FILLER_36_384 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_137 ();
 sg13g2_fill_1 FILLER_37_139 ();
 sg13g2_fill_2 FILLER_37_243 ();
 sg13g2_decap_4 FILLER_37_263 ();
 sg13g2_decap_4 FILLER_37_288 ();
 sg13g2_fill_1 FILLER_37_292 ();
 sg13g2_fill_2 FILLER_37_308 ();
 sg13g2_fill_2 FILLER_37_317 ();
 sg13g2_fill_1 FILLER_37_319 ();
 sg13g2_fill_2 FILLER_37_335 ();
 sg13g2_fill_1 FILLER_37_337 ();
 sg13g2_fill_1 FILLER_37_344 ();
 sg13g2_fill_1 FILLER_37_359 ();
 sg13g2_fill_1 FILLER_37_387 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_130 ();
 sg13g2_decap_4 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_153 ();
 sg13g2_decap_4 FILLER_38_160 ();
 sg13g2_fill_1 FILLER_38_164 ();
 sg13g2_decap_8 FILLER_38_176 ();
 sg13g2_decap_8 FILLER_38_183 ();
 sg13g2_fill_2 FILLER_38_190 ();
 sg13g2_decap_8 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_206 ();
 sg13g2_fill_1 FILLER_38_213 ();
 sg13g2_fill_1 FILLER_38_220 ();
 sg13g2_decap_4 FILLER_38_224 ();
 sg13g2_fill_1 FILLER_38_228 ();
 sg13g2_fill_1 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_241 ();
 sg13g2_decap_8 FILLER_38_253 ();
 sg13g2_decap_8 FILLER_38_260 ();
 sg13g2_fill_1 FILLER_38_267 ();
 sg13g2_decap_8 FILLER_38_284 ();
 sg13g2_fill_1 FILLER_38_291 ();
 sg13g2_fill_2 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_305 ();
 sg13g2_fill_1 FILLER_38_345 ();
 sg13g2_fill_2 FILLER_38_365 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_decap_4 FILLER_38_391 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net39;
 assign uio_oe[1] = net40;
 assign uio_oe[2] = net41;
 assign uio_oe[3] = net42;
 assign uio_oe[4] = net43;
 assign uio_oe[5] = net44;
 assign uio_oe[6] = net45;
 assign uio_oe[7] = net46;
endmodule

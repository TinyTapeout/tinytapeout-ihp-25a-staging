module tt_um_mattvenn_spi_test (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire \config_regs[0] ;
 wire \config_regs[10] ;
 wire \config_regs[11] ;
 wire \config_regs[12] ;
 wire \config_regs[13] ;
 wire \config_regs[14] ;
 wire \config_regs[15] ;
 wire \config_regs[1] ;
 wire \config_regs[2] ;
 wire \config_regs[3] ;
 wire \config_regs[4] ;
 wire \config_regs[5] ;
 wire \config_regs[6] ;
 wire \config_regs[7] ;
 wire \config_regs[8] ;
 wire \config_regs[9] ;
 wire cpha_sync;
 wire cpol_sync;
 wire spi_clk_sync;
 wire spi_cs_n_sync;
 wire spi_miso;
 wire spi_mosi_sync;
 wire \spi_wrapper_i.reg_addr[0] ;
 wire \spi_wrapper_i.reg_addr[1] ;
 wire \spi_wrapper_i.reg_data_o[0] ;
 wire \spi_wrapper_i.reg_data_o[1] ;
 wire \spi_wrapper_i.reg_data_o[2] ;
 wire \spi_wrapper_i.reg_data_o[3] ;
 wire \spi_wrapper_i.reg_data_o[4] ;
 wire \spi_wrapper_i.reg_data_o[5] ;
 wire \spi_wrapper_i.reg_data_o[6] ;
 wire \spi_wrapper_i.reg_data_o[7] ;
 wire \spi_wrapper_i.reg_data_o_vld ;
 wire \spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ;
 wire \spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ;
 wire \spi_wrapper_i.spi_reg_inst.reg_rw ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[0] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[1] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[2] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[3] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[4] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[5] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[6] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[7] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ;
 wire \spi_wrapper_i.spi_reg_inst.state[0] ;
 wire \spi_wrapper_i.spi_reg_inst.state[1] ;
 wire \spi_wrapper_i.spi_reg_inst.state[2] ;
 wire \spi_wrapper_i.spi_reg_inst.state[3] ;
 wire \spi_wrapper_i.spi_reg_inst.state[4] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[0] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[1] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[2] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[3] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[4] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[5] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[6] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ;
 wire \synchronizer_spi_clk_inst.data_sync[1] ;
 wire \synchronizer_spi_cs_n_inst.data_sync[1] ;
 wire \synchronizer_spi_mode_cpha.data_sync[1] ;
 wire \synchronizer_spi_mode_cpol.data_sync[1] ;
 wire \synchronizer_spi_mosi_inst.data_sync[1] ;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_0_clk;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;

 sg13g2_inv_2 _237_ (.Y(_070_),
    .A(net1));
 sg13g2_inv_1 _238_ (.Y(_071_),
    .A(spi_cs_n_sync));
 sg13g2_inv_1 _239_ (.Y(_072_),
    .A(\spi_wrapper_i.spi_reg_inst.reg_rw ));
 sg13g2_inv_1 _240_ (.Y(_073_),
    .A(net69));
 sg13g2_inv_1 _241_ (.Y(_074_),
    .A(spi_clk_sync));
 sg13g2_inv_1 _242_ (.Y(_075_),
    .A(net30));
 sg13g2_inv_1 _243_ (.Y(_076_),
    .A(\spi_wrapper_i.reg_data_o_vld ));
 sg13g2_inv_2 _244_ (.Y(_077_),
    .A(\spi_wrapper_i.reg_addr[1] ));
 sg13g2_nor3_2 _245_ (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ),
    .B(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ),
    .C(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .Y(_078_));
 sg13g2_nand2b_1 _246_ (.Y(_079_),
    .B(net162),
    .A_N(_078_));
 sg13g2_nor3_2 _247_ (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ),
    .B(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ),
    .C(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ),
    .Y(_080_));
 sg13g2_nand2_1 _248_ (.Y(_081_),
    .A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ),
    .B(_080_));
 sg13g2_o21ai_1 _249_ (.B1(_081_),
    .Y(_082_),
    .A1(net76),
    .A2(net120));
 sg13g2_nor2_1 _250_ (.A(net79),
    .B(_071_),
    .Y(_083_));
 sg13g2_nand2_1 _251_ (.Y(_084_),
    .A(net107),
    .B(_083_));
 sg13g2_a21oi_1 _252_ (.A1(_079_),
    .A2(_082_),
    .Y(_085_),
    .B1(_084_));
 sg13g2_nand2_1 _253_ (.Y(_086_),
    .A(net159),
    .B(_078_));
 sg13g2_nand3_1 _254_ (.B(net159),
    .C(_078_),
    .A(net105),
    .Y(_087_));
 sg13g2_nand4_1 _255_ (.B(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ),
    .C(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .A(net105),
    .Y(_088_),
    .D(_078_));
 sg13g2_nand3_1 _256_ (.B(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ),
    .C(_080_),
    .A(net105),
    .Y(_089_));
 sg13g2_nand4_1 _257_ (.B(net105),
    .C(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ),
    .A(net76),
    .Y(_090_),
    .D(_080_));
 sg13g2_nor2b_1 _258_ (.A(spi_cs_n_sync),
    .B_N(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .Y(_091_));
 sg13g2_nand2_1 _259_ (.Y(_092_),
    .A(net107),
    .B(_091_));
 sg13g2_nand2_1 _260_ (.Y(_093_),
    .A(net30),
    .B(_092_));
 sg13g2_nand3_1 _261_ (.B(_090_),
    .C(_093_),
    .A(_088_),
    .Y(_094_));
 sg13g2_nor2_1 _262_ (.A(net121),
    .B(_094_),
    .Y(_005_));
 sg13g2_nand3_1 _263_ (.B(_084_),
    .C(_089_),
    .A(net76),
    .Y(_095_));
 sg13g2_nand3_1 _264_ (.B(\spi_wrapper_i.spi_reg_inst.reg_rw ),
    .C(net69),
    .A(net105),
    .Y(_096_));
 sg13g2_nand2_1 _265_ (.Y(_003_),
    .A(_095_),
    .B(_096_));
 sg13g2_nand2_1 _266_ (.Y(_097_),
    .A(_072_),
    .B(net69));
 sg13g2_o21ai_1 _267_ (.B1(_097_),
    .Y(_098_),
    .A1(_079_),
    .A2(_083_));
 sg13g2_nand2_1 _268_ (.Y(_099_),
    .A(net105),
    .B(_098_));
 sg13g2_nand3b_1 _269_ (.B(net162),
    .C(_078_),
    .Y(_100_),
    .A_N(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ));
 sg13g2_nand2_1 _270_ (.Y(_101_),
    .A(_070_),
    .B(net162));
 sg13g2_nand3_1 _271_ (.B(net88),
    .C(_101_),
    .A(_099_),
    .Y(_000_));
 sg13g2_nand4_1 _272_ (.B(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ),
    .C(net120),
    .A(net105),
    .Y(_102_),
    .D(_080_));
 sg13g2_o21ai_1 _273_ (.B1(_102_),
    .Y(_001_),
    .A1(net105),
    .A2(_073_));
 sg13g2_nand3_1 _274_ (.B(_084_),
    .C(_089_),
    .A(\spi_wrapper_i.spi_reg_inst.state[3] ),
    .Y(_103_));
 sg13g2_o21ai_1 _275_ (.B1(_103_),
    .Y(_002_),
    .A1(_075_),
    .A2(_092_));
 sg13g2_xor2_1 _276_ (.B(cpol_sync),
    .A(cpha_sync),
    .X(_104_));
 sg13g2_nand2b_1 _277_ (.Y(_105_),
    .B(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .A_N(spi_clk_sync));
 sg13g2_o21ai_1 _278_ (.B1(_104_),
    .Y(_106_),
    .A1(spi_cs_n_sync),
    .A2(_105_));
 sg13g2_nor2b_1 _279_ (.A(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .B_N(spi_clk_sync),
    .Y(_107_));
 sg13g2_nor3_1 _280_ (.A(spi_cs_n_sync),
    .B(_074_),
    .C(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .Y(_108_));
 sg13g2_a21o_1 _281_ (.A2(_107_),
    .A1(_071_),
    .B1(_104_),
    .X(_109_));
 sg13g2_and3_1 _282_ (.X(_110_),
    .A(net106),
    .B(_106_),
    .C(_109_));
 sg13g2_mux2_1 _283_ (.A0(net67),
    .A1(net63),
    .S(net84),
    .X(_006_));
 sg13g2_mux2_1 _284_ (.A0(net115),
    .A1(net67),
    .S(net84),
    .X(_007_));
 sg13g2_mux2_1 _285_ (.A0(net138),
    .A1(net115),
    .S(net85),
    .X(_008_));
 sg13g2_mux2_1 _286_ (.A0(net118),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .S(net85),
    .X(_009_));
 sg13g2_mux2_1 _287_ (.A0(net123),
    .A1(net118),
    .S(net85),
    .X(_010_));
 sg13g2_mux2_1 _288_ (.A0(net127),
    .A1(net123),
    .S(net85),
    .X(_011_));
 sg13g2_mux2_1 _289_ (.A0(net111),
    .A1(net127),
    .S(net85),
    .X(_012_));
 sg13g2_mux2_1 _290_ (.A0(net50),
    .A1(net111),
    .S(net85),
    .X(_013_));
 sg13g2_nor2_1 _291_ (.A(net107),
    .B(net79),
    .Y(_111_));
 sg13g2_a21oi_1 _292_ (.A1(net107),
    .A2(_071_),
    .Y(_014_),
    .B1(_111_));
 sg13g2_nor3_2 _293_ (.A(_070_),
    .B(_076_),
    .C(net91),
    .Y(_112_));
 sg13g2_mux2_1 _294_ (.A0(net74),
    .A1(\spi_wrapper_i.reg_data_o[0] ),
    .S(_112_),
    .X(_015_));
 sg13g2_mux2_1 _295_ (.A0(net71),
    .A1(\spi_wrapper_i.reg_data_o[1] ),
    .S(_112_),
    .X(_016_));
 sg13g2_mux2_1 _296_ (.A0(net40),
    .A1(\spi_wrapper_i.reg_data_o[2] ),
    .S(_112_),
    .X(_017_));
 sg13g2_mux2_1 _297_ (.A0(net46),
    .A1(\spi_wrapper_i.reg_data_o[3] ),
    .S(_112_),
    .X(_018_));
 sg13g2_mux2_1 _298_ (.A0(net65),
    .A1(\spi_wrapper_i.reg_data_o[4] ),
    .S(_112_),
    .X(_019_));
 sg13g2_mux2_1 _299_ (.A0(net38),
    .A1(\spi_wrapper_i.reg_data_o[5] ),
    .S(_112_),
    .X(_020_));
 sg13g2_mux2_1 _300_ (.A0(net36),
    .A1(\spi_wrapper_i.reg_data_o[6] ),
    .S(_112_),
    .X(_021_));
 sg13g2_mux2_1 _301_ (.A0(net42),
    .A1(\spi_wrapper_i.reg_data_o[7] ),
    .S(_112_),
    .X(_022_));
 sg13g2_mux2_1 _302_ (.A0(net32),
    .A1(net4),
    .S(net106),
    .X(_023_));
 sg13g2_nand2_1 _303_ (.Y(_113_),
    .A(net107),
    .B(net34));
 sg13g2_o21ai_1 _304_ (.B1(_113_),
    .Y(_024_),
    .A1(net106),
    .A2(_074_));
 sg13g2_mux2_1 _305_ (.A0(net34),
    .A1(net5),
    .S(net106),
    .X(_025_));
 sg13g2_nor2_1 _306_ (.A(net108),
    .B(net157),
    .Y(_114_));
 sg13g2_a21oi_1 _307_ (.A1(net108),
    .A2(_074_),
    .Y(_026_),
    .B1(_114_));
 sg13g2_mux2_1 _308_ (.A0(net81),
    .A1(net6),
    .S(net106),
    .X(_027_));
 sg13g2_mux2_1 _309_ (.A0(net112),
    .A1(net62),
    .S(net108),
    .X(_028_));
 sg13g2_mux2_1 _310_ (.A0(net62),
    .A1(net2),
    .S(net108),
    .X(_029_));
 sg13g2_mux2_1 _311_ (.A0(net82),
    .A1(net68),
    .S(net108),
    .X(_030_));
 sg13g2_mux2_1 _312_ (.A0(net68),
    .A1(net3),
    .S(net108),
    .X(_031_));
 sg13g2_nand2_1 _313_ (.Y(_115_),
    .A(net106),
    .B(net32));
 sg13g2_o21ai_1 _314_ (.B1(_115_),
    .Y(_032_),
    .A1(net106),
    .A2(_071_));
 sg13g2_mux2_1 _315_ (.A0(net63),
    .A1(\synchronizer_spi_mosi_inst.data_sync[1] ),
    .S(net106),
    .X(_033_));
 sg13g2_a21oi_1 _316_ (.A1(_081_),
    .A2(net83),
    .Y(_116_),
    .B1(net153));
 sg13g2_a21oi_1 _317_ (.A1(net153),
    .A2(net83),
    .Y(_034_),
    .B1(net154));
 sg13g2_and3_1 _318_ (.X(_117_),
    .A(net143),
    .B(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ),
    .C(net83));
 sg13g2_a21oi_1 _319_ (.A1(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ),
    .A2(net83),
    .Y(_118_),
    .B1(net143));
 sg13g2_nor2_1 _320_ (.A(_117_),
    .B(net144),
    .Y(_035_));
 sg13g2_xor2_1 _321_ (.B(_117_),
    .A(net109),
    .X(_036_));
 sg13g2_nand3b_1 _322_ (.B(net164),
    .C(_089_),
    .Y(_119_),
    .A_N(net84));
 sg13g2_nand3_1 _323_ (.B(net153),
    .C(net109),
    .A(net143),
    .Y(_120_));
 sg13g2_xnor2_1 _324_ (.Y(_121_),
    .A(net164),
    .B(_120_));
 sg13g2_nand3_1 _325_ (.B(net83),
    .C(_121_),
    .A(_081_),
    .Y(_122_));
 sg13g2_nand2_1 _326_ (.Y(_037_),
    .A(net165),
    .B(_122_));
 sg13g2_nor2_1 _327_ (.A(net50),
    .B(_102_),
    .Y(_123_));
 sg13g2_a21oi_1 _328_ (.A1(_072_),
    .A2(_102_),
    .Y(_038_),
    .B1(net51));
 sg13g2_mux2_1 _329_ (.A0(net67),
    .A1(net91),
    .S(_102_),
    .X(_039_));
 sg13g2_nor2_1 _330_ (.A(net115),
    .B(_102_),
    .Y(_124_));
 sg13g2_a21oi_1 _331_ (.A1(_077_),
    .A2(_102_),
    .Y(_040_),
    .B1(net116));
 sg13g2_nand2_1 _332_ (.Y(_125_),
    .A(_070_),
    .B(net59));
 sg13g2_o21ai_1 _333_ (.B1(_125_),
    .Y(_041_),
    .A1(_072_),
    .A2(net89));
 sg13g2_mux2_1 _334_ (.A0(net67),
    .A1(net151),
    .S(_090_),
    .X(_042_));
 sg13g2_mux2_1 _335_ (.A0(net115),
    .A1(net148),
    .S(net89),
    .X(_043_));
 sg13g2_mux2_1 _336_ (.A0(net138),
    .A1(\spi_wrapper_i.reg_data_o[2] ),
    .S(net89),
    .X(_044_));
 sg13g2_mux2_1 _337_ (.A0(net118),
    .A1(net136),
    .S(net89),
    .X(_045_));
 sg13g2_mux2_1 _338_ (.A0(net123),
    .A1(net124),
    .S(net89),
    .X(_046_));
 sg13g2_mux2_1 _339_ (.A0(net127),
    .A1(net137),
    .S(net89),
    .X(_047_));
 sg13g2_mux2_1 _340_ (.A0(net111),
    .A1(net130),
    .S(net89),
    .X(_048_));
 sg13g2_mux2_1 _341_ (.A0(net50),
    .A1(net131),
    .S(net89),
    .X(_049_));
 sg13g2_a21oi_1 _342_ (.A1(_086_),
    .A2(net83),
    .Y(_126_),
    .B1(net149));
 sg13g2_a21oi_1 _343_ (.A1(net149),
    .A2(net83),
    .Y(_050_),
    .B1(net150));
 sg13g2_and3_1 _344_ (.X(_127_),
    .A(net155),
    .B(net149),
    .C(net85));
 sg13g2_a21oi_1 _345_ (.A1(net149),
    .A2(net85),
    .Y(_128_),
    .B1(net155));
 sg13g2_nor2_1 _346_ (.A(_127_),
    .B(_128_),
    .Y(_051_));
 sg13g2_xor2_1 _347_ (.B(_127_),
    .A(net140),
    .X(_052_));
 sg13g2_nand3b_1 _348_ (.B(net159),
    .C(_087_),
    .Y(_129_),
    .A_N(net84));
 sg13g2_nand3_1 _349_ (.B(net149),
    .C(net140),
    .A(net155),
    .Y(_130_));
 sg13g2_xnor2_1 _350_ (.Y(_131_),
    .A(net159),
    .B(_130_));
 sg13g2_nand3_1 _351_ (.B(net83),
    .C(_131_),
    .A(_086_),
    .Y(_132_));
 sg13g2_nand2_1 _352_ (.Y(_053_),
    .A(net160),
    .B(_132_));
 sg13g2_nand3_1 _353_ (.B(\spi_wrapper_i.reg_data_o_vld ),
    .C(net91),
    .A(net108),
    .Y(_133_));
 sg13g2_mux2_1 _354_ (.A0(\spi_wrapper_i.reg_data_o[0] ),
    .A1(net134),
    .S(_133_),
    .X(_054_));
 sg13g2_mux2_1 _355_ (.A0(\spi_wrapper_i.reg_data_o[1] ),
    .A1(net125),
    .S(_133_),
    .X(_055_));
 sg13g2_mux2_1 _356_ (.A0(\spi_wrapper_i.reg_data_o[2] ),
    .A1(net128),
    .S(_133_),
    .X(_056_));
 sg13g2_mux2_1 _357_ (.A0(\spi_wrapper_i.reg_data_o[3] ),
    .A1(net113),
    .S(_133_),
    .X(_057_));
 sg13g2_mux2_1 _358_ (.A0(net124),
    .A1(net142),
    .S(_133_),
    .X(_058_));
 sg13g2_mux2_1 _359_ (.A0(\spi_wrapper_i.reg_data_o[5] ),
    .A1(net132),
    .S(_133_),
    .X(_059_));
 sg13g2_mux2_1 _360_ (.A0(net130),
    .A1(net147),
    .S(_133_),
    .X(_060_));
 sg13g2_mux2_1 _361_ (.A0(net131),
    .A1(net146),
    .S(_133_),
    .X(_061_));
 sg13g2_nor3_1 _362_ (.A(spi_cs_n_sync),
    .B(_104_),
    .C(_105_),
    .Y(_134_));
 sg13g2_a21oi_1 _363_ (.A1(_104_),
    .A2(_108_),
    .Y(_135_),
    .B1(_134_));
 sg13g2_nor2b_1 _364_ (.A(net90),
    .B_N(net88),
    .Y(_136_));
 sg13g2_a21oi_2 _365_ (.B1(_070_),
    .Y(_137_),
    .A2(_136_),
    .A1(_135_));
 sg13g2_nand2b_1 _366_ (.Y(_138_),
    .B(net91),
    .A_N(\config_regs[8] ));
 sg13g2_o21ai_1 _367_ (.B1(_138_),
    .Y(_139_),
    .A1(net91),
    .A2(\config_regs[0] ));
 sg13g2_nor4_1 _368_ (.A(\spi_wrapper_i.reg_addr[1] ),
    .B(net90),
    .C(net87),
    .D(_139_),
    .Y(_140_));
 sg13g2_mux2_1 _369_ (.A0(net53),
    .A1(_140_),
    .S(_137_),
    .X(_062_));
 sg13g2_mux2_1 _370_ (.A0(\config_regs[1] ),
    .A1(\config_regs[9] ),
    .S(net92),
    .X(_141_));
 sg13g2_a21oi_1 _371_ (.A1(_077_),
    .A2(_141_),
    .Y(_142_),
    .B1(net86));
 sg13g2_nor2b_1 _372_ (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[0] ),
    .B_N(net86),
    .Y(_143_));
 sg13g2_nor3_1 _373_ (.A(net90),
    .B(_142_),
    .C(_143_),
    .Y(_144_));
 sg13g2_mux2_1 _374_ (.A0(net48),
    .A1(_144_),
    .S(_137_),
    .X(_063_));
 sg13g2_mux2_1 _375_ (.A0(\config_regs[2] ),
    .A1(\config_regs[10] ),
    .S(net92),
    .X(_145_));
 sg13g2_a21oi_1 _376_ (.A1(_077_),
    .A2(_145_),
    .Y(_146_),
    .B1(net86));
 sg13g2_nor2b_1 _377_ (.A(net48),
    .B_N(net87),
    .Y(_147_));
 sg13g2_nor3_1 _378_ (.A(net90),
    .B(_146_),
    .C(_147_),
    .Y(_148_));
 sg13g2_mux2_1 _379_ (.A0(net73),
    .A1(_148_),
    .S(_137_),
    .X(_064_));
 sg13g2_nor2b_1 _380_ (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[2] ),
    .B_N(net87),
    .Y(_149_));
 sg13g2_mux2_1 _381_ (.A0(\config_regs[3] ),
    .A1(\config_regs[11] ),
    .S(net92),
    .X(_150_));
 sg13g2_a21oi_1 _382_ (.A1(_077_),
    .A2(_150_),
    .Y(_151_),
    .B1(net86));
 sg13g2_nor3_1 _383_ (.A(net90),
    .B(_149_),
    .C(_151_),
    .Y(_152_));
 sg13g2_mux2_1 _384_ (.A0(net44),
    .A1(_152_),
    .S(_137_),
    .X(_065_));
 sg13g2_nor2b_1 _385_ (.A(net44),
    .B_N(net87),
    .Y(_153_));
 sg13g2_mux2_1 _386_ (.A0(\config_regs[4] ),
    .A1(\config_regs[12] ),
    .S(net92),
    .X(_154_));
 sg13g2_a21oi_1 _387_ (.A1(_077_),
    .A2(_154_),
    .Y(_155_),
    .B1(net86));
 sg13g2_nor3_1 _388_ (.A(net90),
    .B(_153_),
    .C(_155_),
    .Y(_156_));
 sg13g2_mux2_1 _389_ (.A0(net78),
    .A1(_156_),
    .S(_137_),
    .X(_066_));
 sg13g2_mux2_1 _390_ (.A0(\config_regs[5] ),
    .A1(\config_regs[13] ),
    .S(net91),
    .X(_157_));
 sg13g2_a21oi_1 _391_ (.A1(_077_),
    .A2(_157_),
    .Y(_158_),
    .B1(net86));
 sg13g2_nor2b_1 _392_ (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[4] ),
    .B_N(net87),
    .Y(_159_));
 sg13g2_nor3_1 _393_ (.A(net90),
    .B(_158_),
    .C(_159_),
    .Y(_160_));
 sg13g2_mux2_1 _394_ (.A0(net57),
    .A1(_160_),
    .S(_137_),
    .X(_067_));
 sg13g2_nor2b_1 _395_ (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[5] ),
    .B_N(net86),
    .Y(_161_));
 sg13g2_mux2_1 _396_ (.A0(\config_regs[6] ),
    .A1(\config_regs[14] ),
    .S(net91),
    .X(_162_));
 sg13g2_a21oi_1 _397_ (.A1(_077_),
    .A2(_162_),
    .Y(_163_),
    .B1(net86));
 sg13g2_nor3_1 _398_ (.A(_091_),
    .B(_161_),
    .C(_163_),
    .Y(_164_));
 sg13g2_mux2_1 _399_ (.A0(net55),
    .A1(_164_),
    .S(_137_),
    .X(_068_));
 sg13g2_mux2_1 _400_ (.A0(\config_regs[7] ),
    .A1(\config_regs[15] ),
    .S(net91),
    .X(_165_));
 sg13g2_a21oi_1 _401_ (.A1(_077_),
    .A2(_165_),
    .Y(_166_),
    .B1(net88));
 sg13g2_nor2b_1 _402_ (.A(net55),
    .B_N(net87),
    .Y(_167_));
 sg13g2_nor3_1 _403_ (.A(net90),
    .B(_166_),
    .C(_167_),
    .Y(_168_));
 sg13g2_mux2_1 _404_ (.A0(net61),
    .A1(_168_),
    .S(_137_),
    .X(_069_));
 sg13g2_dfrbp_1 _405_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net96),
    .D(net122),
    .Q_N(\spi_wrapper_i.spi_reg_inst.state[0] ),
    .Q(_004_));
 sg13g2_dfrbp_1 _406_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net96),
    .D(net163),
    .Q_N(_234_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[1] ));
 sg13g2_dfrbp_1 _407_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net96),
    .D(net70),
    .Q_N(_235_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[2] ));
 sg13g2_dfrbp_1 _408_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net96),
    .D(net31),
    .Q_N(_236_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[3] ));
 sg13g2_dfrbp_1 _409_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net95),
    .D(net77),
    .Q_N(_233_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[4] ));
 sg13g2_dfrbp_1 _410_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net96),
    .D(_006_),
    .Q_N(_232_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ));
 sg13g2_dfrbp_1 _411_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net93),
    .D(_007_),
    .Q_N(_231_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[1] ));
 sg13g2_dfrbp_1 _412_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net94),
    .D(_008_),
    .Q_N(_230_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ));
 sg13g2_dfrbp_1 _413_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net94),
    .D(net119),
    .Q_N(_229_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ));
 sg13g2_dfrbp_1 _414_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net94),
    .D(_010_),
    .Q_N(_228_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[4] ));
 sg13g2_dfrbp_1 _415_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net93),
    .D(_011_),
    .Q_N(_227_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[5] ));
 sg13g2_dfrbp_1 _416_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net93),
    .D(_012_),
    .Q_N(_226_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[6] ));
 sg13g2_dfrbp_1 _417_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net94),
    .D(_013_),
    .Q_N(_225_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[7] ));
 sg13g2_dfrbp_1 _418_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net104),
    .D(net80),
    .Q_N(_224_),
    .Q(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ));
 sg13g2_dfrbp_1 _419_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net100),
    .D(net75),
    .Q_N(_223_),
    .Q(\config_regs[0] ));
 sg13g2_dfrbp_1 _420_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net100),
    .D(net72),
    .Q_N(_222_),
    .Q(\config_regs[1] ));
 sg13g2_dfrbp_1 _421_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net99),
    .D(net41),
    .Q_N(_221_),
    .Q(\config_regs[2] ));
 sg13g2_dfrbp_1 _422_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net99),
    .D(net47),
    .Q_N(_220_),
    .Q(\config_regs[3] ));
 sg13g2_dfrbp_1 _423_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net99),
    .D(net66),
    .Q_N(_219_),
    .Q(\config_regs[4] ));
 sg13g2_dfrbp_1 _424_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net99),
    .D(net39),
    .Q_N(_218_),
    .Q(\config_regs[5] ));
 sg13g2_dfrbp_1 _425_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net99),
    .D(net37),
    .Q_N(_217_),
    .Q(\config_regs[6] ));
 sg13g2_dfrbp_1 _426_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net101),
    .D(net43),
    .Q_N(_216_),
    .Q(\config_regs[7] ));
 sg13g2_dfrbp_1 _427_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net96),
    .D(_023_),
    .Q_N(_215_),
    .Q(\synchronizer_spi_cs_n_inst.data_sync[1] ));
 sg13g2_dfrbp_1 _428_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net104),
    .D(net35),
    .Q_N(_214_),
    .Q(spi_clk_sync));
 sg13g2_dfrbp_1 _429_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net95),
    .D(_025_),
    .Q_N(_213_),
    .Q(\synchronizer_spi_clk_inst.data_sync[1] ));
 sg13g2_dfrbp_1 _430_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net104),
    .D(net158),
    .Q_N(_212_),
    .Q(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ));
 sg13g2_dfrbp_1 _431_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net95),
    .D(_027_),
    .Q_N(_211_),
    .Q(\synchronizer_spi_mosi_inst.data_sync[1] ));
 sg13g2_dfrbp_1 _432_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net103),
    .D(_028_),
    .Q_N(_210_),
    .Q(cpol_sync));
 sg13g2_dfrbp_1 _433_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net102),
    .D(_029_),
    .Q_N(_209_),
    .Q(\synchronizer_spi_mode_cpol.data_sync[1] ));
 sg13g2_dfrbp_1 _434_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net103),
    .D(_030_),
    .Q_N(_208_),
    .Q(cpha_sync));
 sg13g2_dfrbp_1 _435_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net103),
    .D(_031_),
    .Q_N(_207_),
    .Q(\synchronizer_spi_mode_cpha.data_sync[1] ));
 sg13g2_dfrbp_1 _436_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net104),
    .D(net33),
    .Q_N(_206_),
    .Q(spi_cs_n_sync));
 sg13g2_dfrbp_1 _437_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net95),
    .D(net64),
    .Q_N(_205_),
    .Q(spi_mosi_sync));
 sg13g2_dfrbp_1 _438_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net95),
    .D(_034_),
    .Q_N(_204_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ));
 sg13g2_dfrbp_1 _439_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net95),
    .D(net145),
    .Q_N(_203_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ));
 sg13g2_dfrbp_1 _440_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net95),
    .D(net110),
    .Q_N(_202_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ));
 sg13g2_dfrbp_1 _441_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net95),
    .D(net166),
    .Q_N(_201_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ));
 sg13g2_dfrbp_1 _442_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net96),
    .D(net52),
    .Q_N(_200_),
    .Q(\spi_wrapper_i.spi_reg_inst.reg_rw ));
 sg13g2_dfrbp_1 _443_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net98),
    .D(_039_),
    .Q_N(_199_),
    .Q(\spi_wrapper_i.reg_addr[0] ));
 sg13g2_dfrbp_1 _444_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net104),
    .D(net117),
    .Q_N(_198_),
    .Q(\spi_wrapper_i.reg_addr[1] ));
 sg13g2_dfrbp_1 _445_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net104),
    .D(net60),
    .Q_N(_197_),
    .Q(\spi_wrapper_i.reg_data_o_vld ));
 sg13g2_dfrbp_1 _446_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net98),
    .D(net152),
    .Q_N(_196_),
    .Q(\spi_wrapper_i.reg_data_o[0] ));
 sg13g2_dfrbp_1 _447_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net101),
    .D(_043_),
    .Q_N(_195_),
    .Q(\spi_wrapper_i.reg_data_o[1] ));
 sg13g2_dfrbp_1 _448_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net98),
    .D(net139),
    .Q_N(_194_),
    .Q(\spi_wrapper_i.reg_data_o[2] ));
 sg13g2_dfrbp_1 _449_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net98),
    .D(_045_),
    .Q_N(_193_),
    .Q(\spi_wrapper_i.reg_data_o[3] ));
 sg13g2_dfrbp_1 _450_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net98),
    .D(_046_),
    .Q_N(_192_),
    .Q(\spi_wrapper_i.reg_data_o[4] ));
 sg13g2_dfrbp_1 _451_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net94),
    .D(_047_),
    .Q_N(_191_),
    .Q(\spi_wrapper_i.reg_data_o[5] ));
 sg13g2_dfrbp_1 _452_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net98),
    .D(_048_),
    .Q_N(_190_),
    .Q(\spi_wrapper_i.reg_data_o[6] ));
 sg13g2_dfrbp_1 _453_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net93),
    .D(_049_),
    .Q_N(_189_),
    .Q(\spi_wrapper_i.reg_data_o[7] ));
 sg13g2_dfrbp_1 _454_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net93),
    .D(_050_),
    .Q_N(_188_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ));
 sg13g2_dfrbp_1 _455_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net93),
    .D(_051_),
    .Q_N(_187_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ));
 sg13g2_dfrbp_1 _456_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net93),
    .D(net141),
    .Q_N(_186_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ));
 sg13g2_dfrbp_1 _457_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net93),
    .D(net161),
    .Q_N(_185_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ));
 sg13g2_dfrbp_1 _458_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net100),
    .D(net135),
    .Q_N(_184_),
    .Q(\config_regs[8] ));
 sg13g2_dfrbp_1 _459_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net100),
    .D(net126),
    .Q_N(_183_),
    .Q(\config_regs[9] ));
 sg13g2_dfrbp_1 _460_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net100),
    .D(net129),
    .Q_N(_182_),
    .Q(\config_regs[10] ));
 sg13g2_dfrbp_1 _461_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net99),
    .D(net114),
    .Q_N(_181_),
    .Q(\config_regs[11] ));
 sg13g2_dfrbp_1 _462_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net99),
    .D(_058_),
    .Q_N(_180_),
    .Q(\config_regs[12] ));
 sg13g2_dfrbp_1 _463_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net98),
    .D(net133),
    .Q_N(_179_),
    .Q(\config_regs[13] ));
 sg13g2_dfrbp_1 _464_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net99),
    .D(_060_),
    .Q_N(_178_),
    .Q(\config_regs[14] ));
 sg13g2_dfrbp_1 _465_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net98),
    .D(_061_),
    .Q_N(_177_),
    .Q(\config_regs[15] ));
 sg13g2_dfrbp_1 _466_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net102),
    .D(net54),
    .Q_N(_176_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[0] ));
 sg13g2_dfrbp_1 _467_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net102),
    .D(net49),
    .Q_N(_175_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[1] ));
 sg13g2_dfrbp_1 _468_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net102),
    .D(_064_),
    .Q_N(_174_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[2] ));
 sg13g2_dfrbp_1 _469_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net102),
    .D(net45),
    .Q_N(_173_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[3] ));
 sg13g2_dfrbp_1 _470_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net102),
    .D(_066_),
    .Q_N(_172_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[4] ));
 sg13g2_dfrbp_1 _471_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net102),
    .D(net58),
    .Q_N(_171_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[5] ));
 sg13g2_dfrbp_1 _472_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net102),
    .D(net56),
    .Q_N(_170_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[6] ));
 sg13g2_dfrbp_1 _473_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net103),
    .D(_069_),
    .Q_N(_169_),
    .Q(spi_miso));
 sg13g2_tiehi tt_um_mattvenn_spi_test_26 (.L_HI(net26));
 sg13g2_tiehi tt_um_mattvenn_spi_test_27 (.L_HI(net27));
 sg13g2_tiehi tt_um_mattvenn_spi_test_28 (.L_HI(net28));
 sg13g2_tiehi tt_um_mattvenn_spi_test_29 (.L_HI(net29));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_mattvenn_spi_test_8 (.L_LO(net8));
 sg13g2_tielo tt_um_mattvenn_spi_test_9 (.L_LO(net9));
 sg13g2_tielo tt_um_mattvenn_spi_test_10 (.L_LO(net10));
 sg13g2_tielo tt_um_mattvenn_spi_test_11 (.L_LO(net11));
 sg13g2_tielo tt_um_mattvenn_spi_test_12 (.L_LO(net12));
 sg13g2_tielo tt_um_mattvenn_spi_test_13 (.L_LO(net13));
 sg13g2_tielo tt_um_mattvenn_spi_test_14 (.L_LO(net14));
 sg13g2_tielo tt_um_mattvenn_spi_test_15 (.L_LO(net15));
 sg13g2_tielo tt_um_mattvenn_spi_test_16 (.L_LO(net16));
 sg13g2_tielo tt_um_mattvenn_spi_test_17 (.L_LO(net17));
 sg13g2_tielo tt_um_mattvenn_spi_test_18 (.L_LO(net18));
 sg13g2_tielo tt_um_mattvenn_spi_test_19 (.L_LO(net19));
 sg13g2_tielo tt_um_mattvenn_spi_test_20 (.L_LO(net20));
 sg13g2_tielo tt_um_mattvenn_spi_test_21 (.L_LO(net21));
 sg13g2_tielo tt_um_mattvenn_spi_test_22 (.L_LO(net22));
 sg13g2_tielo tt_um_mattvenn_spi_test_23 (.L_LO(net23));
 sg13g2_tielo tt_um_mattvenn_spi_test_24 (.L_LO(net24));
 sg13g2_tiehi tt_um_mattvenn_spi_test_25 (.L_HI(net25));
 sg13g2_buf_1 _497_ (.A(spi_miso),
    .X(uio_out[3]));
 sg13g2_buf_2 fanout83 (.A(_110_),
    .X(net83));
 sg13g2_buf_1 fanout84 (.A(_110_),
    .X(net84));
 sg13g2_buf_4 fanout85 (.X(net85),
    .A(_110_));
 sg13g2_buf_2 fanout86 (.A(net88),
    .X(net86));
 sg13g2_buf_1 fanout87 (.A(net88),
    .X(net87));
 sg13g2_buf_1 fanout88 (.A(_100_),
    .X(net88));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(_090_));
 sg13g2_buf_2 fanout90 (.A(_091_),
    .X(net90));
 sg13g2_buf_4 fanout91 (.X(net91),
    .A(net156));
 sg13g2_buf_2 fanout92 (.A(\spi_wrapper_i.reg_addr[0] ),
    .X(net92));
 sg13g2_buf_4 fanout93 (.X(net93),
    .A(net97));
 sg13g2_buf_2 fanout94 (.A(net97),
    .X(net94));
 sg13g2_buf_4 fanout95 (.X(net95),
    .A(net97));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(net97));
 sg13g2_buf_2 fanout97 (.A(rst_n),
    .X(net97));
 sg13g2_buf_4 fanout98 (.X(net98),
    .A(net101));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(net100));
 sg13g2_buf_2 fanout100 (.A(net101),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(rst_n),
    .X(net101));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(net104));
 sg13g2_buf_2 fanout103 (.A(net104),
    .X(net103));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(rst_n));
 sg13g2_buf_2 fanout105 (.A(net107),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(net107),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(net108),
    .X(net107));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(net1));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[4]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[5]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[6]),
    .X(net6));
 sg13g2_tielo tt_um_mattvenn_spi_test_7 (.L_LO(net7));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\spi_wrapper_i.spi_reg_inst.state[0] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold2 (.A(_002_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold3 (.A(\synchronizer_spi_cs_n_inst.data_sync[1] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold4 (.A(_032_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold5 (.A(\synchronizer_spi_clk_inst.data_sync[1] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold6 (.A(_024_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold7 (.A(\config_regs[6] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold8 (.A(_021_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold9 (.A(\config_regs[5] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold10 (.A(_020_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold11 (.A(\config_regs[2] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold12 (.A(_017_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold13 (.A(\config_regs[7] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold14 (.A(_022_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold15 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[3] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold16 (.A(_065_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold17 (.A(\config_regs[3] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold18 (.A(_018_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold19 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[1] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold20 (.A(_063_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold21 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[7] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold22 (.A(_123_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold23 (.A(_038_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold24 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[0] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold25 (.A(_062_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold26 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[6] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold27 (.A(_068_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold28 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[5] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold29 (.A(_067_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold30 (.A(\spi_wrapper_i.reg_data_o_vld ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold31 (.A(_041_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold32 (.A(spi_miso),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold33 (.A(\synchronizer_spi_mode_cpol.data_sync[1] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold34 (.A(spi_mosi_sync),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold35 (.A(_033_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold36 (.A(\config_regs[4] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold37 (.A(_019_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold38 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold39 (.A(\synchronizer_spi_mode_cpha.data_sync[1] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold40 (.A(\spi_wrapper_i.spi_reg_inst.state[2] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold41 (.A(_001_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold42 (.A(\config_regs[1] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold43 (.A(_016_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold44 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[2] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold45 (.A(\config_regs[0] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold46 (.A(_015_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold47 (.A(\spi_wrapper_i.spi_reg_inst.state[4] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold48 (.A(_003_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold49 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer[4] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold50 (.A(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold51 (.A(_014_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold52 (.A(\synchronizer_spi_mosi_inst.data_sync[1] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold53 (.A(cpha_sync),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold54 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold55 (.A(_036_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold56 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[6] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold57 (.A(cpol_sync),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold58 (.A(\config_regs[11] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold59 (.A(_057_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold60 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold61 (.A(_124_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold62 (.A(_040_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold63 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold64 (.A(_009_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold65 (.A(\spi_wrapper_i.spi_reg_inst.state[3] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold66 (.A(_085_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold67 (.A(_005_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold68 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[4] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold69 (.A(\spi_wrapper_i.reg_data_o[4] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold70 (.A(\config_regs[9] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold71 (.A(_055_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold72 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[5] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold73 (.A(\config_regs[10] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold74 (.A(_056_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold75 (.A(\spi_wrapper_i.reg_data_o[6] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold76 (.A(\spi_wrapper_i.reg_data_o[7] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold77 (.A(\config_regs[13] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold78 (.A(_059_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold79 (.A(\config_regs[8] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold80 (.A(_054_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold81 (.A(\spi_wrapper_i.reg_data_o[3] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold82 (.A(\spi_wrapper_i.reg_data_o[5] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold83 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold84 (.A(_044_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold85 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold86 (.A(_052_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold87 (.A(\config_regs[12] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold88 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold89 (.A(_118_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold90 (.A(_035_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold91 (.A(\config_regs[15] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold92 (.A(\config_regs[14] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold93 (.A(\spi_wrapper_i.reg_data_o[1] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold94 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold95 (.A(_126_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold96 (.A(\spi_wrapper_i.reg_data_o[0] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold97 (.A(_042_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold98 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold99 (.A(_116_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold100 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold101 (.A(\spi_wrapper_i.reg_addr[0] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold102 (.A(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold103 (.A(_026_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold104 (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold105 (.A(_129_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold106 (.A(_053_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold107 (.A(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold108 (.A(_000_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold109 (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold110 (.A(_119_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold111 (.A(_037_),
    .X(net166));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_4 FILLER_19_224 ();
 sg13g2_fill_1 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_325 ();
 sg13g2_decap_8 FILLER_19_332 ();
 sg13g2_decap_8 FILLER_19_339 ();
 sg13g2_decap_8 FILLER_19_346 ();
 sg13g2_decap_8 FILLER_19_353 ();
 sg13g2_decap_8 FILLER_19_360 ();
 sg13g2_decap_8 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_374 ();
 sg13g2_decap_8 FILLER_19_381 ();
 sg13g2_fill_2 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_4 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_4 FILLER_20_273 ();
 sg13g2_fill_1 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_fill_2 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_fill_1 FILLER_20_370 ();
 sg13g2_fill_2 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_4 FILLER_21_262 ();
 sg13g2_fill_2 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_4 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_356 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_fill_1 FILLER_22_196 ();
 sg13g2_fill_2 FILLER_22_223 ();
 sg13g2_fill_1 FILLER_22_225 ();
 sg13g2_decap_4 FILLER_22_252 ();
 sg13g2_fill_2 FILLER_22_256 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_fill_1 FILLER_22_301 ();
 sg13g2_fill_2 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_fill_2 FILLER_23_189 ();
 sg13g2_fill_1 FILLER_23_191 ();
 sg13g2_decap_4 FILLER_23_227 ();
 sg13g2_fill_2 FILLER_23_231 ();
 sg13g2_fill_1 FILLER_23_259 ();
 sg13g2_fill_2 FILLER_23_296 ();
 sg13g2_fill_2 FILLER_23_317 ();
 sg13g2_fill_1 FILLER_23_345 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_4 FILLER_24_196 ();
 sg13g2_fill_2 FILLER_24_200 ();
 sg13g2_fill_2 FILLER_24_222 ();
 sg13g2_fill_1 FILLER_24_224 ();
 sg13g2_fill_1 FILLER_24_251 ();
 sg13g2_fill_2 FILLER_24_272 ();
 sg13g2_fill_1 FILLER_24_274 ();
 sg13g2_fill_2 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_299 ();
 sg13g2_fill_1 FILLER_24_356 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_4 FILLER_25_161 ();
 sg13g2_fill_2 FILLER_25_165 ();
 sg13g2_decap_8 FILLER_25_184 ();
 sg13g2_decap_8 FILLER_25_191 ();
 sg13g2_decap_4 FILLER_25_198 ();
 sg13g2_fill_2 FILLER_25_247 ();
 sg13g2_fill_2 FILLER_25_290 ();
 sg13g2_fill_1 FILLER_25_300 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_4 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_191 ();
 sg13g2_decap_4 FILLER_26_198 ();
 sg13g2_decap_4 FILLER_26_210 ();
 sg13g2_fill_1 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_263 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_fill_2 FILLER_27_210 ();
 sg13g2_fill_1 FILLER_27_227 ();
 sg13g2_decap_4 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_285 ();
 sg13g2_fill_1 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_4 FILLER_28_154 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_decap_4 FILLER_28_211 ();
 sg13g2_fill_2 FILLER_28_241 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_268 ();
 sg13g2_fill_2 FILLER_28_279 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_154 ();
 sg13g2_fill_1 FILLER_29_156 ();
 sg13g2_decap_4 FILLER_29_220 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_229 ();
 sg13g2_fill_2 FILLER_29_243 ();
 sg13g2_fill_1 FILLER_29_245 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_fill_1 FILLER_30_191 ();
 sg13g2_fill_1 FILLER_30_197 ();
 sg13g2_fill_1 FILLER_30_234 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_fill_2 FILLER_30_307 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_fill_2 FILLER_31_154 ();
 sg13g2_fill_1 FILLER_31_156 ();
 sg13g2_fill_1 FILLER_31_227 ();
 sg13g2_fill_2 FILLER_31_249 ();
 sg13g2_fill_1 FILLER_31_251 ();
 sg13g2_fill_1 FILLER_31_296 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_fill_2 FILLER_32_147 ();
 sg13g2_fill_2 FILLER_32_184 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_fill_2 FILLER_32_294 ();
 sg13g2_fill_2 FILLER_32_322 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_4 FILLER_33_140 ();
 sg13g2_fill_2 FILLER_33_144 ();
 sg13g2_fill_1 FILLER_33_210 ();
 sg13g2_fill_2 FILLER_33_262 ();
 sg13g2_fill_2 FILLER_33_287 ();
 sg13g2_fill_1 FILLER_33_319 ();
 sg13g2_fill_2 FILLER_33_362 ();
 sg13g2_fill_1 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_4 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_151 ();
 sg13g2_fill_1 FILLER_34_166 ();
 sg13g2_fill_2 FILLER_34_198 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_fill_2 FILLER_34_218 ();
 sg13g2_fill_2 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_4 FILLER_35_154 ();
 sg13g2_fill_2 FILLER_35_158 ();
 sg13g2_fill_2 FILLER_35_181 ();
 sg13g2_fill_1 FILLER_35_209 ();
 sg13g2_fill_2 FILLER_35_313 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_fill_1 FILLER_36_215 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_351 ();
 sg13g2_fill_1 FILLER_36_353 ();
 sg13g2_fill_2 FILLER_36_369 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_fill_2 FILLER_37_161 ();
 sg13g2_fill_1 FILLER_37_207 ();
 sg13g2_fill_2 FILLER_37_218 ();
 sg13g2_fill_2 FILLER_37_301 ();
 sg13g2_fill_1 FILLER_37_334 ();
 sg13g2_fill_2 FILLER_37_349 ();
 sg13g2_fill_1 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_fill_2 FILLER_38_164 ();
 sg13g2_fill_1 FILLER_38_221 ();
 sg13g2_fill_2 FILLER_38_232 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_fill_1 FILLER_38_259 ();
 sg13g2_fill_1 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_331 ();
 sg13g2_fill_2 FILLER_38_340 ();
 sg13g2_fill_1 FILLER_38_342 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net25;
 assign uio_oe[1] = net26;
 assign uio_oe[2] = net27;
 assign uio_oe[3] = net28;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net29;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
 assign uio_out[7] = net16;
 assign uo_out[0] = net17;
 assign uo_out[1] = net18;
 assign uo_out[2] = net19;
 assign uo_out[3] = net20;
 assign uo_out[4] = net21;
 assign uo_out[5] = net22;
 assign uo_out[6] = net23;
 assign uo_out[7] = net24;
endmodule

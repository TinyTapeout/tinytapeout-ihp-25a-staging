module tt_um_comm_ic_bhavuk (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire \comm_ic0.MOSI ;
 wire \comm_ic0.SCL ;
 wire \comm_ic0.SCLK ;
 wire \comm_ic0.SDA_op ;
 wire \comm_ic0.SDA_op_en ;
 wire \comm_ic0.SEN ;
 wire \comm_ic0.UART_TX ;
 wire \comm_ic0.busy_i2c ;
 wire \comm_ic0.busy_spi ;
 wire \comm_ic0.busy_uart ;
 wire \comm_ic0.comm_sel[0] ;
 wire \comm_ic0.comm_sel[1] ;
 wire \comm_ic0.curr_st[0] ;
 wire \comm_ic0.curr_st[1] ;
 wire \comm_ic0.curr_st[2] ;
 wire \comm_ic0.curr_st[3] ;
 wire \comm_ic0.error_i2c ;
 wire \comm_ic0.i2c0.addr_ind[0] ;
 wire \comm_ic0.i2c0.addr_ind[1] ;
 wire \comm_ic0.i2c0.addr_ind[2] ;
 wire \comm_ic0.i2c0.addr_wr[0] ;
 wire \comm_ic0.i2c0.addr_wr[1] ;
 wire \comm_ic0.i2c0.addr_wr[2] ;
 wire \comm_ic0.i2c0.addr_wr[3] ;
 wire \comm_ic0.i2c0.addr_wr[4] ;
 wire \comm_ic0.i2c0.addr_wr[5] ;
 wire \comm_ic0.i2c0.addr_wr[6] ;
 wire \comm_ic0.i2c0.addr_wr[7] ;
 wire \comm_ic0.i2c0.address[0] ;
 wire \comm_ic0.i2c0.address[1] ;
 wire \comm_ic0.i2c0.address[2] ;
 wire \comm_ic0.i2c0.address[3] ;
 wire \comm_ic0.i2c0.address[4] ;
 wire \comm_ic0.i2c0.address[5] ;
 wire \comm_ic0.i2c0.address[6] ;
 wire \comm_ic0.i2c0.bits16 ;
 wire \comm_ic0.i2c0.clk_cnt[0] ;
 wire \comm_ic0.i2c0.clk_cnt[1] ;
 wire \comm_ic0.i2c0.clk_cnt[2] ;
 wire \comm_ic0.i2c0.clk_cnt[3] ;
 wire \comm_ic0.i2c0.clk_cnt[4] ;
 wire \comm_ic0.i2c0.clk_cnt[5] ;
 wire \comm_ic0.i2c0.clk_cnt[6] ;
 wire \comm_ic0.i2c0.clk_cnt[7] ;
 wire \comm_ic0.i2c0.clk_cnt_reg[0] ;
 wire \comm_ic0.i2c0.clk_cnt_reg[1] ;
 wire \comm_ic0.i2c0.clk_cnt_reg[2] ;
 wire \comm_ic0.i2c0.clk_cnt_reg[3] ;
 wire \comm_ic0.i2c0.clk_cnt_reg[4] ;
 wire \comm_ic0.i2c0.clk_cnt_reg[5] ;
 wire \comm_ic0.i2c0.clk_cnt_reg[6] ;
 wire \comm_ic0.i2c0.clk_cnt_reg[7] ;
 wire \comm_ic0.i2c0.curr_st[0] ;
 wire \comm_ic0.i2c0.curr_st[1] ;
 wire \comm_ic0.i2c0.curr_st[2] ;
 wire \comm_ic0.i2c0.curr_st[3] ;
 wire \comm_ic0.i2c0.curr_st[4] ;
 wire \comm_ic0.i2c0.curr_st[5] ;
 wire \comm_ic0.i2c0.curr_st[6] ;
 wire \comm_ic0.i2c0.curr_st[7] ;
 wire \comm_ic0.i2c0.data_in[0] ;
 wire \comm_ic0.i2c0.data_in[10] ;
 wire \comm_ic0.i2c0.data_in[11] ;
 wire \comm_ic0.i2c0.data_in[12] ;
 wire \comm_ic0.i2c0.data_in[13] ;
 wire \comm_ic0.i2c0.data_in[14] ;
 wire \comm_ic0.i2c0.data_in[15] ;
 wire \comm_ic0.i2c0.data_in[1] ;
 wire \comm_ic0.i2c0.data_in[2] ;
 wire \comm_ic0.i2c0.data_in[3] ;
 wire \comm_ic0.i2c0.data_in[4] ;
 wire \comm_ic0.i2c0.data_in[5] ;
 wire \comm_ic0.i2c0.data_in[6] ;
 wire \comm_ic0.i2c0.data_in[7] ;
 wire \comm_ic0.i2c0.data_in[8] ;
 wire \comm_ic0.i2c0.data_in[9] ;
 wire \comm_ic0.i2c0.data_ind[0] ;
 wire \comm_ic0.i2c0.data_ind[1] ;
 wire \comm_ic0.i2c0.data_ind[2] ;
 wire \comm_ic0.i2c0.data_ind[3] ;
 wire \comm_ic0.i2c0.data_out[0] ;
 wire \comm_ic0.i2c0.data_out[10] ;
 wire \comm_ic0.i2c0.data_out[11] ;
 wire \comm_ic0.i2c0.data_out[12] ;
 wire \comm_ic0.i2c0.data_out[13] ;
 wire \comm_ic0.i2c0.data_out[14] ;
 wire \comm_ic0.i2c0.data_out[15] ;
 wire \comm_ic0.i2c0.data_out[1] ;
 wire \comm_ic0.i2c0.data_out[2] ;
 wire \comm_ic0.i2c0.data_out[3] ;
 wire \comm_ic0.i2c0.data_out[4] ;
 wire \comm_ic0.i2c0.data_out[5] ;
 wire \comm_ic0.i2c0.data_out[6] ;
 wire \comm_ic0.i2c0.data_out[7] ;
 wire \comm_ic0.i2c0.data_out[8] ;
 wire \comm_ic0.i2c0.data_out[9] ;
 wire \comm_ic0.i2c0.data_wr[0] ;
 wire \comm_ic0.i2c0.data_wr[10] ;
 wire \comm_ic0.i2c0.data_wr[11] ;
 wire \comm_ic0.i2c0.data_wr[12] ;
 wire \comm_ic0.i2c0.data_wr[13] ;
 wire \comm_ic0.i2c0.data_wr[14] ;
 wire \comm_ic0.i2c0.data_wr[15] ;
 wire \comm_ic0.i2c0.data_wr[1] ;
 wire \comm_ic0.i2c0.data_wr[2] ;
 wire \comm_ic0.i2c0.data_wr[3] ;
 wire \comm_ic0.i2c0.data_wr[4] ;
 wire \comm_ic0.i2c0.data_wr[5] ;
 wire \comm_ic0.i2c0.data_wr[6] ;
 wire \comm_ic0.i2c0.data_wr[7] ;
 wire \comm_ic0.i2c0.data_wr[8] ;
 wire \comm_ic0.i2c0.data_wr[9] ;
 wire \comm_ic0.i2c0.scl_cnt[0] ;
 wire \comm_ic0.i2c0.scl_cnt[1] ;
 wire \comm_ic0.i2c0.scl_cnt[2] ;
 wire \comm_ic0.i2c0.scl_cnt[3] ;
 wire \comm_ic0.i2c0.scl_cnt[4] ;
 wire \comm_ic0.i2c0.scl_cnt[5] ;
 wire \comm_ic0.i2c0.scl_cnt[6] ;
 wire \comm_ic0.i2c0.scl_cnt[7] ;
 wire \comm_ic0.i2c0.start ;
 wire \comm_ic0.i2c0.write_n ;
 wire \comm_ic0.i2c_addr_en ;
 wire \comm_ic0.new_uart ;
 wire \comm_ic0.parity_en ;
 wire \comm_ic0.parity_odd ;
 wire \comm_ic0.rx_ack ;
 wire \comm_ic0.rx_data[0] ;
 wire \comm_ic0.rx_data[1] ;
 wire \comm_ic0.rx_data[2] ;
 wire \comm_ic0.rx_data[3] ;
 wire \comm_ic0.rx_data[4] ;
 wire \comm_ic0.rx_data[5] ;
 wire \comm_ic0.rx_data[6] ;
 wire \comm_ic0.rx_data[7] ;
 wire \comm_ic0.rx_error ;
 wire \comm_ic0.rx_new ;
 wire \comm_ic0.send_cnt[0] ;
 wire \comm_ic0.send_cnt[1] ;
 wire \comm_ic0.send_cnt[2] ;
 wire \comm_ic0.send_cnt[3] ;
 wire \comm_ic0.spi0.CPHA ;
 wire \comm_ic0.spi0.CPOL ;
 wire \comm_ic0.spi0.bits16 ;
 wire \comm_ic0.spi0.clk_cnt[0] ;
 wire \comm_ic0.spi0.clk_cnt[1] ;
 wire \comm_ic0.spi0.clk_cnt[2] ;
 wire \comm_ic0.spi0.clk_cnt[3] ;
 wire \comm_ic0.spi0.clk_cnt[4] ;
 wire \comm_ic0.spi0.clk_cnt[5] ;
 wire \comm_ic0.spi0.clk_cnt[6] ;
 wire \comm_ic0.spi0.clk_cnt[7] ;
 wire \comm_ic0.spi0.clk_cnt_reg[0] ;
 wire \comm_ic0.spi0.clk_cnt_reg[1] ;
 wire \comm_ic0.spi0.clk_cnt_reg[2] ;
 wire \comm_ic0.spi0.clk_cnt_reg[3] ;
 wire \comm_ic0.spi0.clk_cnt_reg[4] ;
 wire \comm_ic0.spi0.clk_cnt_reg[5] ;
 wire \comm_ic0.spi0.clk_cnt_reg[6] ;
 wire \comm_ic0.spi0.clk_cnt_reg[7] ;
 wire \comm_ic0.spi0.curr_st[0] ;
 wire \comm_ic0.spi0.curr_st[1] ;
 wire \comm_ic0.spi0.curr_st[2] ;
 wire \comm_ic0.spi0.curr_st[3] ;
 wire \comm_ic0.spi0.data_in[0] ;
 wire \comm_ic0.spi0.data_in[10] ;
 wire \comm_ic0.spi0.data_in[11] ;
 wire \comm_ic0.spi0.data_in[12] ;
 wire \comm_ic0.spi0.data_in[13] ;
 wire \comm_ic0.spi0.data_in[14] ;
 wire \comm_ic0.spi0.data_in[15] ;
 wire \comm_ic0.spi0.data_in[1] ;
 wire \comm_ic0.spi0.data_in[2] ;
 wire \comm_ic0.spi0.data_in[3] ;
 wire \comm_ic0.spi0.data_in[4] ;
 wire \comm_ic0.spi0.data_in[5] ;
 wire \comm_ic0.spi0.data_in[6] ;
 wire \comm_ic0.spi0.data_in[7] ;
 wire \comm_ic0.spi0.data_in[8] ;
 wire \comm_ic0.spi0.data_in[9] ;
 wire \comm_ic0.spi0.data_ind[0] ;
 wire \comm_ic0.spi0.data_ind[1] ;
 wire \comm_ic0.spi0.data_ind[2] ;
 wire \comm_ic0.spi0.data_ind[3] ;
 wire \comm_ic0.spi0.data_out[0] ;
 wire \comm_ic0.spi0.data_out[10] ;
 wire \comm_ic0.spi0.data_out[11] ;
 wire \comm_ic0.spi0.data_out[12] ;
 wire \comm_ic0.spi0.data_out[13] ;
 wire \comm_ic0.spi0.data_out[14] ;
 wire \comm_ic0.spi0.data_out[15] ;
 wire \comm_ic0.spi0.data_out[1] ;
 wire \comm_ic0.spi0.data_out[2] ;
 wire \comm_ic0.spi0.data_out[3] ;
 wire \comm_ic0.spi0.data_out[4] ;
 wire \comm_ic0.spi0.data_out[5] ;
 wire \comm_ic0.spi0.data_out[6] ;
 wire \comm_ic0.spi0.data_out[7] ;
 wire \comm_ic0.spi0.data_out[8] ;
 wire \comm_ic0.spi0.data_out[9] ;
 wire \comm_ic0.spi0.data_wr[0] ;
 wire \comm_ic0.spi0.data_wr[10] ;
 wire \comm_ic0.spi0.data_wr[11] ;
 wire \comm_ic0.spi0.data_wr[12] ;
 wire \comm_ic0.spi0.data_wr[13] ;
 wire \comm_ic0.spi0.data_wr[14] ;
 wire \comm_ic0.spi0.data_wr[15] ;
 wire \comm_ic0.spi0.data_wr[1] ;
 wire \comm_ic0.spi0.data_wr[2] ;
 wire \comm_ic0.spi0.data_wr[3] ;
 wire \comm_ic0.spi0.data_wr[4] ;
 wire \comm_ic0.spi0.data_wr[5] ;
 wire \comm_ic0.spi0.data_wr[6] ;
 wire \comm_ic0.spi0.data_wr[7] ;
 wire \comm_ic0.spi0.data_wr[8] ;
 wire \comm_ic0.spi0.data_wr[9] ;
 wire \comm_ic0.spi0.mode[0] ;
 wire \comm_ic0.spi0.mode[1] ;
 wire \comm_ic0.spi0.sclk_cnt[0] ;
 wire \comm_ic0.spi0.sclk_cnt[1] ;
 wire \comm_ic0.spi0.sclk_cnt[2] ;
 wire \comm_ic0.spi0.sclk_cnt[3] ;
 wire \comm_ic0.spi0.sclk_cnt[4] ;
 wire \comm_ic0.spi0.sclk_cnt[5] ;
 wire \comm_ic0.spi0.sclk_cnt[6] ;
 wire \comm_ic0.spi0.sclk_cnt[7] ;
 wire \comm_ic0.spi0.start ;
 wire \comm_ic0.tx_data[0] ;
 wire \comm_ic0.tx_data[1] ;
 wire \comm_ic0.tx_data[2] ;
 wire \comm_ic0.tx_data[3] ;
 wire \comm_ic0.tx_data[4] ;
 wire \comm_ic0.tx_data[5] ;
 wire \comm_ic0.tx_data[6] ;
 wire \comm_ic0.tx_data[7] ;
 wire \comm_ic0.tx_new ;
 wire \comm_ic0.uart0.clk_b ;
 wire \comm_ic0.uart0.clk_cnt[0] ;
 wire \comm_ic0.uart0.clk_cnt[1] ;
 wire \comm_ic0.uart0.clk_cnt[2] ;
 wire \comm_ic0.uart0.clk_cnt[3] ;
 wire \comm_ic0.uart0.clk_cnt[4] ;
 wire \comm_ic0.uart0.clk_cnt[5] ;
 wire \comm_ic0.uart0.clk_cnt[6] ;
 wire \comm_ic0.uart0.clk_cnt[7] ;
 wire \comm_ic0.uart0.clk_cnt_reg[0] ;
 wire \comm_ic0.uart0.clk_cnt_reg[1] ;
 wire \comm_ic0.uart0.clk_cnt_reg[2] ;
 wire \comm_ic0.uart0.clk_cnt_reg[3] ;
 wire \comm_ic0.uart0.clk_cnt_reg[4] ;
 wire \comm_ic0.uart0.clk_cnt_reg[5] ;
 wire \comm_ic0.uart0.clk_cnt_reg[6] ;
 wire \comm_ic0.uart0.clk_cnt_reg[7] ;
 wire \comm_ic0.uart0.curr_st[0] ;
 wire \comm_ic0.uart0.curr_st[1] ;
 wire \comm_ic0.uart0.curr_st[2] ;
 wire \comm_ic0.uart0.enable ;
 wire \comm_ic0.uart0.par_en ;
 wire \comm_ic0.uart0.par_odd ;
 wire \comm_ic0.uart0.rx_data_reg[0] ;
 wire \comm_ic0.uart0.rx_data_reg[10] ;
 wire \comm_ic0.uart0.rx_data_reg[1] ;
 wire \comm_ic0.uart0.rx_data_reg[2] ;
 wire \comm_ic0.uart0.rx_data_reg[3] ;
 wire \comm_ic0.uart0.rx_data_reg[4] ;
 wire \comm_ic0.uart0.rx_data_reg[5] ;
 wire \comm_ic0.uart0.rx_data_reg[6] ;
 wire \comm_ic0.uart0.rx_data_reg[7] ;
 wire \comm_ic0.uart0.rx_data_reg[8] ;
 wire \comm_ic0.uart0.rx_data_reg[9] ;
 wire \comm_ic0.uart0.rx_ind[0] ;
 wire \comm_ic0.uart0.rx_ind[1] ;
 wire \comm_ic0.uart0.rx_ind[2] ;
 wire \comm_ic0.uart0.rx_ind[3] ;
 wire \comm_ic0.uart0.rx_st[0] ;
 wire \comm_ic0.uart0.rx_st[1] ;
 wire \comm_ic0.uart0.rx_st[2] ;
 wire \comm_ic0.uart0.setting ;
 wire \comm_ic0.uart0.tx_data_reg[0] ;
 wire \comm_ic0.uart0.tx_data_reg[1] ;
 wire \comm_ic0.uart0.tx_data_reg[2] ;
 wire \comm_ic0.uart0.tx_data_reg[3] ;
 wire \comm_ic0.uart0.tx_data_reg[4] ;
 wire \comm_ic0.uart0.tx_data_reg[5] ;
 wire \comm_ic0.uart0.tx_data_reg[6] ;
 wire \comm_ic0.uart0.tx_data_reg[7] ;
 wire \comm_ic0.uart0.tx_data_reg[8] ;
 wire \comm_ic0.uart0.tx_data_reg[9] ;
 wire \comm_ic0.uart0.tx_ind[0] ;
 wire \comm_ic0.uart0.tx_ind[1] ;
 wire \comm_ic0.uart0.tx_ind[2] ;
 wire \comm_ic0.uart0.tx_ind[3] ;
 wire \comm_ic0.uart0.tx_st ;
 wire \comm_ic0.uart0.uclk_cnt[0] ;
 wire \comm_ic0.uart0.uclk_cnt[1] ;
 wire \comm_ic0.uart0.uclk_cnt[2] ;
 wire \comm_ic0.uart0.uclk_cnt[3] ;
 wire \comm_ic0.uart0.uclk_cnt[4] ;
 wire \comm_ic0.uart0.uclk_cnt[5] ;
 wire \comm_ic0.uart0.uclk_cnt[6] ;
 wire \comm_ic0.uart0.uclk_cnt[7] ;
 wire net312;
 wire net313;
 wire net314;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;

 sg13g2_inv_1 _2194_ (.Y(_1329_),
    .A(net429));
 sg13g2_inv_4 _2195_ (.A(net661),
    .Y(_1330_));
 sg13g2_inv_1 _2196_ (.Y(_1331_),
    .A(net332));
 sg13g2_inv_4 _2197_ (.A(net664),
    .Y(_1332_));
 sg13g2_inv_1 _2198_ (.Y(_1333_),
    .A(net423));
 sg13g2_inv_1 _2199_ (.Y(_1334_),
    .A(net669));
 sg13g2_inv_4 _2200_ (.A(net672),
    .Y(_1335_));
 sg13g2_inv_2 _2201_ (.Y(_1336_),
    .A(net868));
 sg13g2_inv_1 _2202_ (.Y(_1337_),
    .A(net1068));
 sg13g2_inv_1 _2203_ (.Y(_1338_),
    .A(net917));
 sg13g2_inv_1 _2204_ (.Y(_1339_),
    .A(net850));
 sg13g2_inv_1 _2205_ (.Y(_1340_),
    .A(net821));
 sg13g2_inv_1 _2206_ (.Y(_1341_),
    .A(net395));
 sg13g2_inv_1 _2207_ (.Y(_1342_),
    .A(net711));
 sg13g2_inv_1 _2208_ (.Y(_1343_),
    .A(net780));
 sg13g2_inv_1 _2209_ (.Y(_1344_),
    .A(net398));
 sg13g2_inv_1 _2210_ (.Y(_1345_),
    .A(net767));
 sg13g2_inv_1 _2211_ (.Y(_1346_),
    .A(net353));
 sg13g2_inv_1 _2212_ (.Y(_1347_),
    .A(net438));
 sg13g2_inv_1 _2213_ (.Y(_1348_),
    .A(net350));
 sg13g2_inv_1 _2214_ (.Y(_1349_),
    .A(net380));
 sg13g2_inv_1 _2215_ (.Y(_1350_),
    .A(net441));
 sg13g2_inv_1 _2216_ (.Y(_1351_),
    .A(net432));
 sg13g2_inv_1 _2217_ (.Y(_1352_),
    .A(net356));
 sg13g2_inv_1 _2218_ (.Y(_1353_),
    .A(net404));
 sg13g2_inv_1 _2219_ (.Y(_1354_),
    .A(net347));
 sg13g2_inv_1 _2220_ (.Y(_1355_),
    .A(net469));
 sg13g2_inv_1 _2221_ (.Y(_1356_),
    .A(net478));
 sg13g2_inv_1 _2222_ (.Y(_1357_),
    .A(net401));
 sg13g2_inv_1 _2223_ (.Y(_1358_),
    .A(net865));
 sg13g2_inv_1 _2224_ (.Y(_1359_),
    .A(net792));
 sg13g2_inv_1 _2225_ (.Y(_1360_),
    .A(net750));
 sg13g2_inv_1 _2226_ (.Y(_1361_),
    .A(net523));
 sg13g2_inv_1 _2227_ (.Y(_1362_),
    .A(net383));
 sg13g2_inv_1 _2228_ (.Y(_1363_),
    .A(net726));
 sg13g2_inv_1 _2229_ (.Y(_1364_),
    .A(net486));
 sg13g2_inv_1 _2230_ (.Y(_1365_),
    .A(net326));
 sg13g2_inv_1 _2231_ (.Y(_1366_),
    .A(net374));
 sg13g2_inv_1 _2232_ (.Y(_1367_),
    .A(net368));
 sg13g2_inv_1 _2233_ (.Y(_1368_),
    .A(net481));
 sg13g2_inv_1 _2234_ (.Y(_1369_),
    .A(net806));
 sg13g2_inv_1 _2235_ (.Y(_1370_),
    .A(net702));
 sg13g2_inv_1 _2236_ (.Y(_1371_),
    .A(net752));
 sg13g2_inv_1 _2237_ (.Y(_1372_),
    .A(net1112));
 sg13g2_inv_4 _2238_ (.A(net623),
    .Y(_1373_));
 sg13g2_inv_1 _2239_ (.Y(_1374_),
    .A(net980));
 sg13g2_inv_1 _2240_ (.Y(_1375_),
    .A(net892));
 sg13g2_inv_1 _2241_ (.Y(_1376_),
    .A(net902));
 sg13g2_inv_1 _2242_ (.Y(_1377_),
    .A(net927));
 sg13g2_inv_1 _2243_ (.Y(_1378_),
    .A(net783));
 sg13g2_inv_1 _2244_ (.Y(_1379_),
    .A(net466));
 sg13g2_inv_1 _2245_ (.Y(_1380_),
    .A(net747));
 sg13g2_inv_1 _2246_ (.Y(_1381_),
    .A(net863));
 sg13g2_inv_2 _2247_ (.Y(_1382_),
    .A(net1074));
 sg13g2_inv_1 _2248_ (.Y(_1383_),
    .A(net942));
 sg13g2_inv_1 _2249_ (.Y(_1384_),
    .A(net1304));
 sg13g2_inv_1 _2250_ (.Y(_1385_),
    .A(net983));
 sg13g2_inv_1 _2251_ (.Y(_1386_),
    .A(net844));
 sg13g2_inv_1 _2252_ (.Y(_1387_),
    .A(net930));
 sg13g2_inv_1 _2253_ (.Y(_1388_),
    .A(net962));
 sg13g2_inv_1 _2254_ (.Y(_1389_),
    .A(net738));
 sg13g2_inv_4 _2255_ (.A(net1213),
    .Y(_1390_));
 sg13g2_inv_1 _2256_ (.Y(_1391_),
    .A(net410));
 sg13g2_inv_1 _2257_ (.Y(_1392_),
    .A(net460));
 sg13g2_inv_1 _2258_ (.Y(_1393_),
    .A(net344));
 sg13g2_inv_1 _2259_ (.Y(_1394_),
    .A(net475));
 sg13g2_inv_1 _2260_ (.Y(_1395_),
    .A(net452));
 sg13g2_inv_1 _2261_ (.Y(_1396_),
    .A(net389));
 sg13g2_inv_1 _2262_ (.Y(_1397_),
    .A(net708));
 sg13g2_inv_1 _2263_ (.Y(_1398_),
    .A(net498));
 sg13g2_inv_1 _2264_ (.Y(_1399_),
    .A(net413));
 sg13g2_inv_1 _2265_ (.Y(_1400_),
    .A(\comm_ic0.spi0.CPHA ));
 sg13g2_inv_2 _2266_ (.Y(_1401_),
    .A(net585));
 sg13g2_inv_1 _2267_ (.Y(_1402_),
    .A(net1251));
 sg13g2_inv_1 _2268_ (.Y(_1403_),
    .A(net911));
 sg13g2_inv_1 _2269_ (.Y(_1404_),
    .A(\comm_ic0.spi0.clk_cnt_reg[0] ));
 sg13g2_inv_1 _2270_ (.Y(_1405_),
    .A(net871));
 sg13g2_inv_1 _2271_ (.Y(_1406_),
    .A(net1031));
 sg13g2_inv_1 _2272_ (.Y(_1407_),
    .A(net1303));
 sg13g2_inv_2 _2273_ (.Y(_1408_),
    .A(net1348));
 sg13g2_inv_1 _2274_ (.Y(_1409_),
    .A(net314));
 sg13g2_inv_1 _2275_ (.Y(_1410_),
    .A(net1190));
 sg13g2_inv_2 _2276_ (.Y(_1411_),
    .A(net1038));
 sg13g2_inv_1 _2277_ (.Y(_1412_),
    .A(\comm_ic0.uart0.tx_st ));
 sg13g2_inv_2 _2278_ (.Y(_1413_),
    .A(\comm_ic0.uart0.rx_ind[3] ));
 sg13g2_inv_1 _2279_ (.Y(_1414_),
    .A(\comm_ic0.uart0.rx_data_reg[0] ));
 sg13g2_inv_1 _2280_ (.Y(_1415_),
    .A(\comm_ic0.rx_error ));
 sg13g2_inv_1 _2281_ (.Y(_1416_),
    .A(\comm_ic0.uart0.rx_st[1] ));
 sg13g2_inv_1 _2282_ (.Y(_1417_),
    .A(net611));
 sg13g2_inv_1 _2283_ (.Y(_1418_),
    .A(net838));
 sg13g2_inv_1 _2284_ (.Y(_1419_),
    .A(net1149));
 sg13g2_inv_1 _2285_ (.Y(_1420_),
    .A(net1048));
 sg13g2_inv_2 _2286_ (.Y(_1421_),
    .A(net678));
 sg13g2_inv_1 _2287_ (.Y(_1422_),
    .A(net1234));
 sg13g2_inv_1 _2288_ (.Y(_1423_),
    .A(net1221));
 sg13g2_inv_1 _2289_ (.Y(_1424_),
    .A(\comm_ic0.spi0.sclk_cnt[6] ));
 sg13g2_inv_2 _2290_ (.Y(_1425_),
    .A(net621));
 sg13g2_inv_1 _2291_ (.Y(_1426_),
    .A(net1182));
 sg13g2_inv_1 _2292_ (.Y(_1427_),
    .A(net1071));
 sg13g2_inv_1 _2293_ (.Y(_1428_),
    .A(net595));
 sg13g2_inv_1 _2294_ (.Y(_1429_),
    .A(net589));
 sg13g2_inv_1 _2295_ (.Y(_1430_),
    .A(net591));
 sg13g2_inv_2 _2296_ (.Y(_1431_),
    .A(net4));
 sg13g2_inv_1 _2297_ (.Y(_1432_),
    .A(net599));
 sg13g2_inv_1 _2298_ (.Y(_1433_),
    .A(\comm_ic0.uart0.tx_ind[3] ));
 sg13g2_inv_2 _2299_ (.Y(_1434_),
    .A(net638));
 sg13g2_inv_1 _2300_ (.Y(_1435_),
    .A(_0030_));
 sg13g2_inv_1 _2301_ (.Y(_1436_),
    .A(_0036_));
 sg13g2_inv_1 _2302_ (.Y(_1437_),
    .A(_0043_));
 sg13g2_inv_1 _2303_ (.Y(_1438_),
    .A(_0050_));
 sg13g2_inv_1 _2304_ (.Y(_1439_),
    .A(_0064_));
 sg13g2_inv_1 _2305_ (.Y(_1440_),
    .A(net1196));
 sg13g2_nor2b_1 _2306_ (.A(net1333),
    .B_N(net911),
    .Y(_1441_));
 sg13g2_xnor2_1 _2307_ (.Y(_1442_),
    .A(net828),
    .B(\comm_ic0.spi0.sclk_cnt[3] ));
 sg13g2_nor2b_1 _2308_ (.A(net744),
    .B_N(net1221),
    .Y(_1443_));
 sg13g2_a221oi_1 _2309_ (.B2(_1402_),
    .C1(_1443_),
    .B1(\comm_ic0.spi0.sclk_cnt[6] ),
    .A1(_1403_),
    .Y(_1444_),
    .A2(net1333));
 sg13g2_xor2_1 _2310_ (.B(\comm_ic0.spi0.sclk_cnt[2] ),
    .A(net992),
    .X(_1445_));
 sg13g2_a221oi_1 _2311_ (.B2(net1251),
    .C1(_1445_),
    .B1(_1424_),
    .A1(net744),
    .Y(_1446_),
    .A2(_1423_));
 sg13g2_xor2_1 _2312_ (.B(net1234),
    .A(\comm_ic0.spi0.clk_cnt_reg[1] ),
    .X(_1447_));
 sg13g2_xor2_1 _2313_ (.B(net1265),
    .A(net880),
    .X(_1448_));
 sg13g2_nor4_1 _2314_ (.A(net1328),
    .B(_1441_),
    .C(_1447_),
    .D(_1448_),
    .Y(_1449_));
 sg13g2_and4_2 _2315_ (.A(_1442_),
    .B(net1334),
    .C(_1446_),
    .D(_1449_),
    .X(_1450_));
 sg13g2_nand4_1 _2316_ (.B(_1444_),
    .C(_1446_),
    .A(_1442_),
    .Y(_1451_),
    .D(_1449_));
 sg13g2_nor2_1 _2317_ (.A(net1234),
    .B(\comm_ic0.spi0.sclk_cnt[1] ),
    .Y(_1452_));
 sg13g2_or4_2 _2318_ (.A(net1234),
    .B(net1265),
    .C(\comm_ic0.spi0.sclk_cnt[2] ),
    .D(\comm_ic0.spi0.sclk_cnt[3] ),
    .X(_1453_));
 sg13g2_or2_1 _2319_ (.X(_1454_),
    .B(net1221),
    .A(\comm_ic0.spi0.sclk_cnt[4] ));
 sg13g2_nor3_1 _2320_ (.A(\comm_ic0.spi0.sclk_cnt[6] ),
    .B(_1453_),
    .C(_1454_),
    .Y(_1455_));
 sg13g2_nor4_2 _2321_ (.A(\comm_ic0.spi0.sclk_cnt[6] ),
    .B(net1328),
    .C(_1453_),
    .Y(_1456_),
    .D(_1454_));
 sg13g2_nor2_1 _2322_ (.A(_1450_),
    .B(_1456_),
    .Y(_1457_));
 sg13g2_o21ai_1 _2323_ (.B1(net1106),
    .Y(_1458_),
    .A1(_1450_),
    .A2(net1329));
 sg13g2_nand2_2 _2324_ (.Y(_1459_),
    .A(_1384_),
    .B(net1193));
 sg13g2_nand3_1 _2325_ (.B(_1458_),
    .C(net1194),
    .A(net683),
    .Y(_0018_));
 sg13g2_and3_1 _2326_ (.X(_1460_),
    .A(\comm_ic0.spi0.start ),
    .B(\comm_ic0.spi0.curr_st[0] ),
    .C(net681));
 sg13g2_inv_1 _2327_ (.Y(_1461_),
    .A(net569));
 sg13g2_nand3_1 _2328_ (.B(net1134),
    .C(_1451_),
    .A(net681),
    .Y(_1462_));
 sg13g2_nand2_1 _2329_ (.Y(_0019_),
    .A(_1461_),
    .B(net1135));
 sg13g2_nor2b_2 _2330_ (.A(net580),
    .B_N(net579),
    .Y(_1463_));
 sg13g2_nand2b_1 _2331_ (.Y(_1464_),
    .B(net771),
    .A_N(net581));
 sg13g2_nor2_2 _2332_ (.A(_1425_),
    .B(net566),
    .Y(_1465_));
 sg13g2_nor2_2 _2333_ (.A(net657),
    .B(_1425_),
    .Y(_1466_));
 sg13g2_nor2b_1 _2334_ (.A(net579),
    .B_N(net580),
    .Y(_1467_));
 sg13g2_nand2b_2 _2335_ (.Y(_1468_),
    .B(net1129),
    .A_N(net579));
 sg13g2_nor2_1 _2336_ (.A(net672),
    .B(_1468_),
    .Y(_1469_));
 sg13g2_a22oi_1 _2337_ (.Y(_1470_),
    .B1(_1466_),
    .B2(_1469_),
    .A2(_1465_),
    .A1(net660));
 sg13g2_nor2_1 _2338_ (.A(net658),
    .B(_1470_),
    .Y(_1471_));
 sg13g2_nor2_2 _2339_ (.A(net1034),
    .B(net658),
    .Y(_1472_));
 sg13g2_nor2_2 _2340_ (.A(net623),
    .B(net621),
    .Y(_1473_));
 sg13g2_nand3b_1 _2341_ (.B(_1472_),
    .C(_1473_),
    .Y(_1474_),
    .A_N(net1168));
 sg13g2_nand2_1 _2342_ (.Y(_1475_),
    .A(net579),
    .B(net580));
 sg13g2_nand3_1 _2343_ (.B(net580),
    .C(_1466_),
    .A(net579),
    .Y(_1476_));
 sg13g2_inv_1 _2344_ (.Y(_1477_),
    .A(_1476_));
 sg13g2_and2_1 _2345_ (.A(net690),
    .B(net1168),
    .X(_1478_));
 sg13g2_nand2_1 _2346_ (.Y(_1479_),
    .A(net694),
    .B(net1168));
 sg13g2_nand2_1 _2347_ (.Y(_1480_),
    .A(net623),
    .B(net690));
 sg13g2_o21ai_1 _2348_ (.B1(net694),
    .Y(_1481_),
    .A1(net623),
    .A2(net1168));
 sg13g2_nand3_1 _2349_ (.B(_1476_),
    .C(_1481_),
    .A(_1474_),
    .Y(_1482_));
 sg13g2_o21ai_1 _2350_ (.B1(net636),
    .Y(_1483_),
    .A1(_1471_),
    .A2(_1482_));
 sg13g2_nand2_1 _2351_ (.Y(_1484_),
    .A(net662),
    .B(net666));
 sg13g2_nor2_2 _2352_ (.A(net579),
    .B(net580),
    .Y(_1485_));
 sg13g2_and3_2 _2353_ (.X(_1486_),
    .A(net636),
    .B(net825),
    .C(_1485_));
 sg13g2_o21ai_1 _2354_ (.B1(net3),
    .Y(_1487_),
    .A1(net662),
    .A2(_1332_));
 sg13g2_a221oi_1 _2355_ (.B2(net625),
    .C1(net657),
    .B1(_1487_),
    .A1(_1484_),
    .Y(_1488_),
    .A2(_1486_));
 sg13g2_nand2_1 _2356_ (.Y(_1489_),
    .A(_1473_),
    .B(_1479_));
 sg13g2_and2_2 _2357_ (.A(net626),
    .B(_1485_),
    .X(_1490_));
 sg13g2_nand2_2 _2358_ (.Y(_1491_),
    .A(net565),
    .B(net563));
 sg13g2_a22oi_1 _2359_ (.Y(_1492_),
    .B1(_1481_),
    .B2(_1425_),
    .A2(net563),
    .A1(net566));
 sg13g2_a22oi_1 _2360_ (.Y(_1493_),
    .B1(_1492_),
    .B2(net626),
    .A2(_1490_),
    .A1(_1489_));
 sg13g2_nand3_1 _2361_ (.B(_1488_),
    .C(_1493_),
    .A(_1483_),
    .Y(_0014_));
 sg13g2_and2_2 _2362_ (.A(net633),
    .B(_1467_),
    .X(_1494_));
 sg13g2_o21ai_1 _2363_ (.B1(_1494_),
    .Y(_1495_),
    .A1(net623),
    .A2(net1168));
 sg13g2_and2_1 _2364_ (.A(net635),
    .B(net1168),
    .X(_1496_));
 sg13g2_nand2b_1 _2365_ (.Y(_1497_),
    .B(net338),
    .A_N(net634));
 sg13g2_nand2_1 _2366_ (.Y(_1498_),
    .A(net634),
    .B(net1116));
 sg13g2_o21ai_1 _2367_ (.B1(_1498_),
    .Y(_1499_),
    .A1(net627),
    .A2(_1497_));
 sg13g2_a21oi_1 _2368_ (.A1(net623),
    .A2(_1499_),
    .Y(_1500_),
    .B1(_1496_));
 sg13g2_o21ai_1 _2369_ (.B1(_1495_),
    .Y(_1501_),
    .A1(net565),
    .A2(_1500_));
 sg13g2_nand2_1 _2370_ (.Y(_1502_),
    .A(net694),
    .B(_1501_));
 sg13g2_or2_1 _2371_ (.X(_1503_),
    .B(_1470_),
    .A(net1182));
 sg13g2_or3_2 _2372_ (.A(net626),
    .B(net634),
    .C(net631),
    .X(_1504_));
 sg13g2_nor3_1 _2373_ (.A(net657),
    .B(_1425_),
    .C(_1504_),
    .Y(_1505_));
 sg13g2_nor3_2 _2374_ (.A(net579),
    .B(net1129),
    .C(net626),
    .Y(_1506_));
 sg13g2_nor2b_1 _2375_ (.A(_1481_),
    .B_N(_1506_),
    .Y(_1507_));
 sg13g2_a21oi_1 _2376_ (.A1(_1475_),
    .A2(_1505_),
    .Y(_1508_),
    .B1(_1507_));
 sg13g2_nand4_1 _2377_ (.B(_1502_),
    .C(_1503_),
    .A(_1488_),
    .Y(_0002_),
    .D(_1508_));
 sg13g2_nand2_1 _2378_ (.Y(_1509_),
    .A(net1116),
    .B(_1463_));
 sg13g2_nand4_1 _2379_ (.B(net694),
    .C(net563),
    .A(net623),
    .Y(_1510_),
    .D(net1117));
 sg13g2_nand3_1 _2380_ (.B(net563),
    .C(_1478_),
    .A(net565),
    .Y(_1511_));
 sg13g2_nand3_1 _2381_ (.B(net1118),
    .C(_1511_),
    .A(_1474_),
    .Y(_1512_));
 sg13g2_o21ai_1 _2382_ (.B1(net631),
    .Y(_1513_),
    .A1(_1477_),
    .A2(net1119));
 sg13g2_nand2_1 _2383_ (.Y(_1514_),
    .A(_1478_),
    .B(_1491_));
 sg13g2_o21ai_1 _2384_ (.B1(_1514_),
    .Y(_1515_),
    .A1(_1480_),
    .A2(net1117));
 sg13g2_nand2_1 _2385_ (.Y(_1516_),
    .A(net444),
    .B(_1515_));
 sg13g2_nor2_2 _2386_ (.A(_1373_),
    .B(_1468_),
    .Y(_1517_));
 sg13g2_and2_1 _2387_ (.A(net444),
    .B(_1517_),
    .X(_1518_));
 sg13g2_nand2_1 _2388_ (.Y(_1519_),
    .A(net687),
    .B(net548));
 sg13g2_and3_2 _2389_ (.X(_1520_),
    .A(net1034),
    .B(net694),
    .C(net3));
 sg13g2_nand2b_1 _2390_ (.Y(_1521_),
    .B(_1520_),
    .A_N(_1484_));
 sg13g2_nand4_1 _2391_ (.B(net1170),
    .C(_1519_),
    .A(_1513_),
    .Y(_0015_),
    .D(_1521_));
 sg13g2_o21ai_1 _2392_ (.B1(net444),
    .Y(_1522_),
    .A1(_1466_),
    .A2(net1119));
 sg13g2_and2_2 _2393_ (.A(net825),
    .B(_1494_),
    .X(_1523_));
 sg13g2_nand4_1 _2394_ (.B(net672),
    .C(net687),
    .A(net670),
    .Y(_1524_),
    .D(_1523_));
 sg13g2_and2_1 _2395_ (.A(_1332_),
    .B(_1520_),
    .X(_1525_));
 sg13g2_nor2_1 _2396_ (.A(net670),
    .B(_1335_),
    .Y(_1526_));
 sg13g2_nor2_1 _2397_ (.A(net660),
    .B(net672),
    .Y(_1527_));
 sg13g2_nor2_1 _2398_ (.A(net662),
    .B(net739),
    .Y(_1528_));
 sg13g2_a22oi_1 _2399_ (.Y(_1529_),
    .B1(_1527_),
    .B2(_1528_),
    .A2(_1526_),
    .A1(net1109));
 sg13g2_nand2b_1 _2400_ (.Y(_1530_),
    .B(_1525_),
    .A_N(_1529_));
 sg13g2_nand3_1 _2401_ (.B(_1524_),
    .C(_1530_),
    .A(net1120),
    .Y(_0017_));
 sg13g2_nand4_1 _2402_ (.B(net666),
    .C(net694),
    .A(net662),
    .Y(_1531_),
    .D(_1486_));
 sg13g2_nand2_2 _2403_ (.Y(_1532_),
    .A(net633),
    .B(_1465_));
 sg13g2_nand4_1 _2404_ (.B(net694),
    .C(net636),
    .A(net670),
    .Y(_1533_),
    .D(_1465_));
 sg13g2_and2_1 _2405_ (.A(_1466_),
    .B(_1526_),
    .X(_1534_));
 sg13g2_a22oi_1 _2406_ (.Y(_1535_),
    .B1(_1534_),
    .B2(_1494_),
    .A2(_1529_),
    .A1(_1525_));
 sg13g2_a21o_1 _2407_ (.A2(net623),
    .A1(net580),
    .B1(net621),
    .X(_1536_));
 sg13g2_nand3_1 _2408_ (.B(_1475_),
    .C(_1536_),
    .A(net694),
    .Y(_1537_));
 sg13g2_nand2b_1 _2409_ (.Y(_1538_),
    .B(_1537_),
    .A_N(_1515_));
 sg13g2_or2_1 _2410_ (.X(_1539_),
    .B(_1481_),
    .A(_1475_));
 sg13g2_nand3_1 _2411_ (.B(_1476_),
    .C(_1539_),
    .A(_1474_),
    .Y(_1540_));
 sg13g2_a22oi_1 _2412_ (.Y(_1541_),
    .B1(_1540_),
    .B2(net626),
    .A2(_1538_),
    .A1(net631));
 sg13g2_nand4_1 _2413_ (.B(_1533_),
    .C(_1535_),
    .A(_1531_),
    .Y(_0016_),
    .D(_1541_));
 sg13g2_nor2_1 _2414_ (.A(\comm_ic0.i2c0.scl_cnt[0] ),
    .B(\comm_ic0.i2c0.scl_cnt[1] ),
    .Y(_1542_));
 sg13g2_or4_2 _2415_ (.A(\comm_ic0.i2c0.scl_cnt[0] ),
    .B(\comm_ic0.i2c0.scl_cnt[1] ),
    .C(\comm_ic0.i2c0.scl_cnt[3] ),
    .D(\comm_ic0.i2c0.scl_cnt[2] ),
    .X(_1543_));
 sg13g2_nor3_2 _2416_ (.A(\comm_ic0.i2c0.scl_cnt[5] ),
    .B(net1313),
    .C(_1543_),
    .Y(_1544_));
 sg13g2_nor2b_1 _2417_ (.A(net1156),
    .B_N(_1544_),
    .Y(_1545_));
 sg13g2_nor2b_2 _2418_ (.A(net1079),
    .B_N(_1545_),
    .Y(_1546_));
 sg13g2_nand2b_1 _2419_ (.Y(_1547_),
    .B(_1545_),
    .A_N(net1079));
 sg13g2_nand3_1 _2420_ (.B(net831),
    .C(net539),
    .A(net690),
    .Y(_1548_));
 sg13g2_nor2b_1 _2421_ (.A(net1270),
    .B_N(\comm_ic0.i2c0.clk_cnt_reg[2] ),
    .Y(_1549_));
 sg13g2_nor2b_1 _2422_ (.A(\comm_ic0.i2c0.clk_cnt_reg[2] ),
    .B_N(net1270),
    .Y(_1550_));
 sg13g2_nor2b_1 _2423_ (.A(\comm_ic0.i2c0.clk_cnt_reg[6] ),
    .B_N(\comm_ic0.i2c0.scl_cnt[5] ),
    .Y(_1551_));
 sg13g2_nor4_2 _2424_ (.A(net1079),
    .B(_1549_),
    .C(_1550_),
    .Y(_1552_),
    .D(_1551_));
 sg13g2_xnor2_1 _2425_ (.Y(_1553_),
    .A(\comm_ic0.i2c0.clk_cnt_reg[5] ),
    .B(net1313));
 sg13g2_xnor2_1 _2426_ (.Y(_1554_),
    .A(net1331),
    .B(net1156));
 sg13g2_nor2b_1 _2427_ (.A(\comm_ic0.i2c0.scl_cnt[5] ),
    .B_N(\comm_ic0.i2c0.clk_cnt_reg[6] ),
    .Y(_1555_));
 sg13g2_nor2b_1 _2428_ (.A(\comm_ic0.i2c0.scl_cnt[2] ),
    .B_N(\comm_ic0.i2c0.clk_cnt_reg[3] ),
    .Y(_1556_));
 sg13g2_nor2b_1 _2429_ (.A(net1246),
    .B_N(\comm_ic0.i2c0.scl_cnt[2] ),
    .Y(_1557_));
 sg13g2_nand2b_1 _2430_ (.Y(_1558_),
    .B(\comm_ic0.i2c0.clk_cnt_reg[4] ),
    .A_N(\comm_ic0.i2c0.scl_cnt[3] ));
 sg13g2_nand2b_1 _2431_ (.Y(_1559_),
    .B(\comm_ic0.i2c0.clk_cnt_reg[1] ),
    .A_N(\comm_ic0.i2c0.scl_cnt[0] ));
 sg13g2_nand2b_1 _2432_ (.Y(_1560_),
    .B(\comm_ic0.i2c0.scl_cnt[3] ),
    .A_N(\comm_ic0.i2c0.clk_cnt_reg[4] ));
 sg13g2_nand2b_1 _2433_ (.Y(_1561_),
    .B(\comm_ic0.i2c0.scl_cnt[0] ),
    .A_N(\comm_ic0.i2c0.clk_cnt_reg[1] ));
 sg13g2_nand4_1 _2434_ (.B(_1559_),
    .C(_1560_),
    .A(_1558_),
    .Y(_1562_),
    .D(_1561_));
 sg13g2_nor4_2 _2435_ (.A(_1555_),
    .B(_1556_),
    .C(_1557_),
    .Y(_1563_),
    .D(_1562_));
 sg13g2_and4_2 _2436_ (.A(_1552_),
    .B(_1553_),
    .C(_1554_),
    .D(_1563_),
    .X(_1564_));
 sg13g2_nand4_1 _2437_ (.B(_1553_),
    .C(_1554_),
    .A(_1552_),
    .Y(_1565_),
    .D(_1563_));
 sg13g2_nand2_2 _2438_ (.Y(_1566_),
    .A(net689),
    .B(net1332));
 sg13g2_o21ai_1 _2439_ (.B1(net832),
    .Y(_0013_),
    .A1(_1427_),
    .A2(_1566_));
 sg13g2_nor2_2 _2440_ (.A(net655),
    .B(_1564_),
    .Y(_1567_));
 sg13g2_nand2_1 _2441_ (.Y(_1568_),
    .A(net590),
    .B(_1567_));
 sg13g2_nor2_1 _2442_ (.A(net1153),
    .B(\comm_ic0.i2c0.addr_ind[0] ),
    .Y(_1569_));
 sg13g2_nand2_1 _2443_ (.Y(_1570_),
    .A(net386),
    .B(_1569_));
 sg13g2_nand2_1 _2444_ (.Y(_1571_),
    .A(net589),
    .B(_1570_));
 sg13g2_a21oi_1 _2445_ (.A1(net589),
    .A2(_1570_),
    .Y(_1572_),
    .B1(net914));
 sg13g2_o21ai_1 _2446_ (.B1(_1568_),
    .Y(_0012_),
    .A1(_1566_),
    .A2(net915));
 sg13g2_nor2_1 _2447_ (.A(net1122),
    .B(net1290),
    .Y(_1573_));
 sg13g2_nor3_2 _2448_ (.A(net604),
    .B(net1122),
    .C(net1290),
    .Y(_1574_));
 sg13g2_and2_2 _2449_ (.A(_1411_),
    .B(_1574_),
    .X(_1575_));
 sg13g2_nand2_2 _2450_ (.Y(_1576_),
    .A(_1411_),
    .B(_1574_));
 sg13g2_nand2_2 _2451_ (.Y(_1577_),
    .A(net592),
    .B(_1576_));
 sg13g2_nand2_1 _2452_ (.Y(_1578_),
    .A(net1190),
    .B(_1431_));
 sg13g2_a21oi_1 _2453_ (.A1(_1577_),
    .A2(_1578_),
    .Y(_1579_),
    .B1(_1566_));
 sg13g2_a21o_1 _2454_ (.A2(_1567_),
    .A1(net1132),
    .B1(_1579_),
    .X(_0011_));
 sg13g2_nor2_1 _2455_ (.A(_1390_),
    .B(net578),
    .Y(_1580_));
 sg13g2_a21oi_1 _2456_ (.A1(net1045),
    .A2(net1081),
    .Y(_1581_),
    .B1(net554));
 sg13g2_nor2_1 _2457_ (.A(net656),
    .B(net1082),
    .Y(_0010_));
 sg13g2_nor2_1 _2458_ (.A(_1382_),
    .B(net1),
    .Y(_1582_));
 sg13g2_o21ai_1 _2459_ (.B1(\comm_ic0.uart0.rx_st[0] ),
    .Y(_1583_),
    .A1(_1382_),
    .A2(net1));
 sg13g2_nand3_1 _2460_ (.B(net693),
    .C(_1583_),
    .A(_1416_),
    .Y(_0024_));
 sg13g2_nand2_1 _2461_ (.Y(_1584_),
    .A(net1071),
    .B(net538));
 sg13g2_nand3_1 _2462_ (.B(net1332),
    .C(_1575_),
    .A(net593),
    .Y(_1585_));
 sg13g2_a21oi_1 _2463_ (.A1(net1072),
    .A2(_1585_),
    .Y(_0009_),
    .B1(net656));
 sg13g2_a22oi_1 _2464_ (.Y(_1586_),
    .B1(net597),
    .B2(_1382_),
    .A2(\comm_ic0.uart0.curr_st[0] ),
    .A1(net942));
 sg13g2_nor2_1 _2465_ (.A(net648),
    .B(net943),
    .Y(_0023_));
 sg13g2_nand3_1 _2466_ (.B(net1045),
    .C(_1546_),
    .A(net689),
    .Y(_1587_));
 sg13g2_nand2_1 _2467_ (.Y(_1588_),
    .A(net595),
    .B(_1567_));
 sg13g2_nand2_1 _2468_ (.Y(_0008_),
    .A(net1046),
    .B(_1588_));
 sg13g2_nand2_1 _2469_ (.Y(_1589_),
    .A(net1190),
    .B(_1567_));
 sg13g2_nand3_1 _2470_ (.B(net589),
    .C(_1569_),
    .A(net386),
    .Y(_1590_));
 sg13g2_o21ai_1 _2471_ (.B1(_1589_),
    .Y(_0007_),
    .A1(_1566_),
    .A2(net387));
 sg13g2_nand3_1 _2472_ (.B(net588),
    .C(_1546_),
    .A(net689),
    .Y(_1591_));
 sg13g2_nand3_1 _2473_ (.B(net4),
    .C(_1564_),
    .A(net1190),
    .Y(_1592_));
 sg13g2_nand2_2 _2474_ (.Y(_1593_),
    .A(_1390_),
    .B(net1312));
 sg13g2_nand4_1 _2475_ (.B(_1591_),
    .C(net1191),
    .A(net689),
    .Y(_0006_),
    .D(_1593_));
 sg13g2_nand2_1 _2476_ (.Y(_1594_),
    .A(net1106),
    .B(_1457_));
 sg13g2_and2_2 _2477_ (.A(\comm_ic0.spi0.CPHA ),
    .B(_1456_),
    .X(_1595_));
 sg13g2_nand2_2 _2478_ (.Y(_1596_),
    .A(_1400_),
    .B(_1450_));
 sg13g2_a21oi_1 _2479_ (.A1(_1400_),
    .A2(_1450_),
    .Y(_1597_),
    .B1(_1595_));
 sg13g2_a21o_2 _2480_ (.A2(_1450_),
    .A1(_1400_),
    .B1(_1595_),
    .X(_1598_));
 sg13g2_nor2_2 _2481_ (.A(net586),
    .B(net587),
    .Y(_1599_));
 sg13g2_nand2_1 _2482_ (.Y(_1600_),
    .A(net532),
    .B(_1599_));
 sg13g2_nor3_2 _2483_ (.A(net583),
    .B(net586),
    .C(net587),
    .Y(_1601_));
 sg13g2_nand2_1 _2484_ (.Y(_1602_),
    .A(net532),
    .B(_1601_));
 sg13g2_nor2b_2 _2485_ (.A(net1146),
    .B_N(_1601_),
    .Y(_1603_));
 sg13g2_or4_2 _2486_ (.A(net1146),
    .B(net583),
    .C(net586),
    .D(net1209),
    .X(_1604_));
 sg13g2_nand3_1 _2487_ (.B(net532),
    .C(_1603_),
    .A(net639),
    .Y(_1605_));
 sg13g2_a21oi_1 _2488_ (.A1(net1107),
    .A2(_1605_),
    .Y(_0021_),
    .B1(net645));
 sg13g2_nor2_1 _2489_ (.A(\comm_ic0.uart0.rx_ind[1] ),
    .B(\comm_ic0.uart0.rx_ind[0] ),
    .Y(_1606_));
 sg13g2_nor3_2 _2490_ (.A(net555),
    .B(\comm_ic0.uart0.rx_ind[1] ),
    .C(\comm_ic0.uart0.rx_ind[0] ),
    .Y(_1607_));
 sg13g2_nand2_2 _2491_ (.Y(_1608_),
    .A(_1413_),
    .B(_1607_));
 sg13g2_nand2_1 _2492_ (.Y(_1609_),
    .A(\comm_ic0.uart0.rx_st[2] ),
    .B(_1608_));
 sg13g2_nand2_1 _2493_ (.Y(_1610_),
    .A(\comm_ic0.uart0.rx_st[0] ),
    .B(_1582_));
 sg13g2_a21oi_1 _2494_ (.A1(_1609_),
    .A2(_1610_),
    .Y(_0025_),
    .B1(net658));
 sg13g2_a21oi_1 _2495_ (.A1(_1383_),
    .A2(net1296),
    .Y(_1611_),
    .B1(net648));
 sg13g2_o21ai_1 _2496_ (.B1(_1611_),
    .Y(_0022_),
    .A1(net1074),
    .A2(_1432_));
 sg13g2_o21ai_1 _2497_ (.B1(_1466_),
    .Y(_1612_),
    .A1(net626),
    .A2(net631));
 sg13g2_nand3_1 _2498_ (.B(_1521_),
    .C(_1612_),
    .A(_1476_),
    .Y(_0005_));
 sg13g2_nand2_1 _2499_ (.Y(_1613_),
    .A(net1134),
    .B(net1335));
 sg13g2_o21ai_1 _2500_ (.B1(net1143),
    .Y(_1614_),
    .A1(net534),
    .A2(_1604_));
 sg13g2_a21oi_1 _2501_ (.A1(_1613_),
    .A2(net1144),
    .Y(_0020_),
    .B1(net645));
 sg13g2_and2_2 _2502_ (.A(_1330_),
    .B(_1525_),
    .X(_1615_));
 sg13g2_nand2b_1 _2503_ (.Y(_1616_),
    .B(net1169),
    .A_N(_1506_));
 sg13g2_a21oi_1 _2504_ (.A1(net520),
    .A2(_1491_),
    .Y(_1617_),
    .B1(_1616_));
 sg13g2_or2_1 _2505_ (.X(_0004_),
    .B(_1617_),
    .A(_1615_));
 sg13g2_o21ai_1 _2506_ (.B1(net1116),
    .Y(_1618_),
    .A1(net338),
    .A2(net634));
 sg13g2_o21ai_1 _2507_ (.B1(_1618_),
    .Y(_1619_),
    .A1(net626),
    .A2(_1497_));
 sg13g2_nor2_1 _2508_ (.A(_1463_),
    .B(_1494_),
    .Y(_1620_));
 sg13g2_o21ai_1 _2509_ (.B1(_1620_),
    .Y(_1621_),
    .A1(net580),
    .A2(net626));
 sg13g2_o21ai_1 _2510_ (.B1(_1621_),
    .Y(_1622_),
    .A1(net565),
    .A2(net1219));
 sg13g2_nand2b_1 _2511_ (.Y(_1623_),
    .B(_1622_),
    .A_N(_1480_));
 sg13g2_nor2_1 _2512_ (.A(_1330_),
    .B(net666),
    .Y(_1624_));
 sg13g2_nand4_1 _2513_ (.B(_1426_),
    .C(_1466_),
    .A(net672),
    .Y(_1625_),
    .D(net564));
 sg13g2_nor3_1 _2514_ (.A(net660),
    .B(net657),
    .C(net1182),
    .Y(_1626_));
 sg13g2_a22oi_1 _2515_ (.Y(_1627_),
    .B1(_1626_),
    .B2(_1465_),
    .A2(_1525_),
    .A1(net663));
 sg13g2_nand4_1 _2516_ (.B(_1623_),
    .C(_1625_),
    .A(_1531_),
    .Y(_0003_),
    .D(_1627_));
 sg13g2_and2_2 _2517_ (.A(net693),
    .B(\comm_ic0.uart0.rx_st[2] ),
    .X(_1628_));
 sg13g2_nand2_2 _2518_ (.Y(_1629_),
    .A(net695),
    .B(\comm_ic0.uart0.rx_st[2] ));
 sg13g2_nor2_1 _2519_ (.A(_1608_),
    .B(_1629_),
    .Y(_0001_));
 sg13g2_nor2_2 _2520_ (.A(net1139),
    .B(net1161),
    .Y(_1630_));
 sg13g2_or2_2 _2521_ (.X(_1631_),
    .B(net596),
    .A(net598));
 sg13g2_nor3_1 _2522_ (.A(_1382_),
    .B(net649),
    .C(_1630_),
    .Y(_0000_));
 sg13g2_nor2b_1 _2523_ (.A(\comm_ic0.rx_error ),
    .B_N(\comm_ic0.rx_new ),
    .Y(\comm_ic0.new_uart ));
 sg13g2_nor4_2 _2524_ (.A(_1372_),
    .B(_1382_),
    .C(\comm_ic0.uart0.tx_st ),
    .Y(_1632_),
    .D(net657));
 sg13g2_nand4_1 _2525_ (.B(\comm_ic0.uart0.enable ),
    .C(_1412_),
    .A(\comm_ic0.tx_new ),
    .Y(_0354_),
    .D(net692));
 sg13g2_nor3_2 _2526_ (.A(\comm_ic0.uart0.tx_ind[0] ),
    .B(\comm_ic0.uart0.tx_ind[1] ),
    .C(\comm_ic0.uart0.tx_ind[2] ),
    .Y(_0355_));
 sg13g2_a21oi_1 _2527_ (.A1(_1433_),
    .A2(_0355_),
    .Y(_0356_),
    .B1(_0028_));
 sg13g2_a21o_1 _2528_ (.A2(_0356_),
    .A1(net693),
    .B1(_1632_),
    .X(_0075_));
 sg13g2_nor2_2 _2529_ (.A(\comm_ic0.uart0.curr_st[0] ),
    .B(net597),
    .Y(_0357_));
 sg13g2_nor2_2 _2530_ (.A(\comm_ic0.uart0.curr_st[0] ),
    .B(_1631_),
    .Y(_0358_));
 sg13g2_nor4_2 _2531_ (.A(net1051),
    .B(net1016),
    .C(net1013),
    .Y(_0359_),
    .D(net1048));
 sg13g2_nor4_2 _2532_ (.A(net965),
    .B(net1149),
    .C(net1084),
    .Y(_0360_),
    .D(net1010));
 sg13g2_nand2_1 _2533_ (.Y(_0361_),
    .A(_0359_),
    .B(_0360_));
 sg13g2_nand3_1 _2534_ (.B(_0359_),
    .C(_0360_),
    .A(net320),
    .Y(_0362_));
 sg13g2_nor2_1 _2535_ (.A(net1048),
    .B(net572),
    .Y(_0363_));
 sg13g2_a22oi_1 _2536_ (.Y(_0364_),
    .B1(_0362_),
    .B2(_0363_),
    .A2(net572),
    .A1(net864));
 sg13g2_nor2_1 _2537_ (.A(_1630_),
    .B(_0364_),
    .Y(_0365_));
 sg13g2_a21oi_1 _2538_ (.A1(net1048),
    .A2(_0358_),
    .Y(_0366_),
    .B1(_0365_));
 sg13g2_nor2_1 _2539_ (.A(net648),
    .B(net1049),
    .Y(_0076_));
 sg13g2_nand3_1 _2540_ (.B(_0359_),
    .C(_0360_),
    .A(\comm_ic0.uart0.clk_cnt_reg[1] ),
    .Y(_0367_));
 sg13g2_nor2_1 _2541_ (.A(net1013),
    .B(net572),
    .Y(_0368_));
 sg13g2_a22oi_1 _2542_ (.Y(_0369_),
    .B1(_0367_),
    .B2(_0368_),
    .A2(net572),
    .A1(_1380_));
 sg13g2_nor2_1 _2543_ (.A(_0364_),
    .B(_0369_),
    .Y(_0370_));
 sg13g2_xnor2_1 _2544_ (.Y(_0371_),
    .A(_0364_),
    .B(_0369_));
 sg13g2_a22oi_1 _2545_ (.Y(_0372_),
    .B1(_0371_),
    .B2(_1631_),
    .A2(_0358_),
    .A1(net1013));
 sg13g2_nor2_1 _2546_ (.A(net648),
    .B(net1014),
    .Y(_0077_));
 sg13g2_and3_2 _2547_ (.X(_0373_),
    .A(net598),
    .B(_0359_),
    .C(_0360_));
 sg13g2_nand2_1 _2548_ (.Y(_0374_),
    .A(net1016),
    .B(net599));
 sg13g2_o21ai_1 _2549_ (.B1(_0374_),
    .Y(_0375_),
    .A1(_1379_),
    .A2(net599));
 sg13g2_a21oi_1 _2550_ (.A1(\comm_ic0.uart0.clk_cnt_reg[2] ),
    .A2(_0373_),
    .Y(_0376_),
    .B1(_0375_));
 sg13g2_a21o_1 _2551_ (.A2(_0373_),
    .A1(\comm_ic0.uart0.clk_cnt_reg[2] ),
    .B1(_0375_),
    .X(_0377_));
 sg13g2_nand2_1 _2552_ (.Y(_0378_),
    .A(_0370_),
    .B(_0376_));
 sg13g2_xnor2_1 _2553_ (.Y(_0379_),
    .A(_0370_),
    .B(_0376_));
 sg13g2_a22oi_1 _2554_ (.Y(_0380_),
    .B1(_0379_),
    .B2(_1631_),
    .A2(_0358_),
    .A1(net1016));
 sg13g2_nor2_1 _2555_ (.A(net648),
    .B(net1017),
    .Y(_0078_));
 sg13g2_nand2_1 _2556_ (.Y(_0381_),
    .A(net1051),
    .B(net598));
 sg13g2_o21ai_1 _2557_ (.B1(_0381_),
    .Y(_0382_),
    .A1(_1378_),
    .A2(net599));
 sg13g2_a21o_1 _2558_ (.A2(_0373_),
    .A1(\comm_ic0.uart0.clk_cnt_reg[3] ),
    .B1(_0382_),
    .X(_0383_));
 sg13g2_nor4_2 _2559_ (.A(_0364_),
    .B(_0369_),
    .C(_0377_),
    .Y(_0384_),
    .D(_0383_));
 sg13g2_xnor2_1 _2560_ (.Y(_0385_),
    .A(_0378_),
    .B(_0383_));
 sg13g2_a22oi_1 _2561_ (.Y(_0386_),
    .B1(_0385_),
    .B2(_1631_),
    .A2(_0358_),
    .A1(net1051));
 sg13g2_nor2_1 _2562_ (.A(net648),
    .B(net1052),
    .Y(_0079_));
 sg13g2_nor2_1 _2563_ (.A(_1343_),
    .B(net598),
    .Y(_0387_));
 sg13g2_a221oi_1 _2564_ (.B2(\comm_ic0.uart0.clk_cnt_reg[4] ),
    .C1(_0387_),
    .B1(_0373_),
    .A1(net1010),
    .Y(_0388_),
    .A2(net598));
 sg13g2_nand2_1 _2565_ (.Y(_0389_),
    .A(_0384_),
    .B(_0388_));
 sg13g2_xnor2_1 _2566_ (.Y(_0390_),
    .A(_0384_),
    .B(_0388_));
 sg13g2_a22oi_1 _2567_ (.Y(_0391_),
    .B1(_0390_),
    .B2(_1631_),
    .A2(_0358_),
    .A1(net1010));
 sg13g2_nor2_1 _2568_ (.A(net646),
    .B(net1011),
    .Y(_0080_));
 sg13g2_nand2_1 _2569_ (.Y(_0392_),
    .A(net1084),
    .B(net598));
 sg13g2_o21ai_1 _2570_ (.B1(_0392_),
    .Y(_0393_),
    .A1(_1342_),
    .A2(net598));
 sg13g2_a21o_1 _2571_ (.A2(_0373_),
    .A1(\comm_ic0.uart0.clk_cnt_reg[5] ),
    .B1(_0393_),
    .X(_0394_));
 sg13g2_inv_1 _2572_ (.Y(_0395_),
    .A(_0394_));
 sg13g2_nand3_1 _2573_ (.B(_0388_),
    .C(_0395_),
    .A(_0384_),
    .Y(_0396_));
 sg13g2_xnor2_1 _2574_ (.Y(_0397_),
    .A(_0389_),
    .B(_0394_));
 sg13g2_a22oi_1 _2575_ (.Y(_0398_),
    .B1(_0397_),
    .B2(_1631_),
    .A2(_0358_),
    .A1(net1084));
 sg13g2_nor2_1 _2576_ (.A(net646),
    .B(net1085),
    .Y(_0081_));
 sg13g2_nand2_1 _2577_ (.Y(_0399_),
    .A(net1149),
    .B(_0358_));
 sg13g2_nand3_1 _2578_ (.B(_0359_),
    .C(_0360_),
    .A(net1324),
    .Y(_0400_));
 sg13g2_a21oi_1 _2579_ (.A1(_0037_),
    .A2(_0361_),
    .Y(_0401_),
    .B1(net572));
 sg13g2_a22oi_1 _2580_ (.Y(_0402_),
    .B1(_0400_),
    .B2(_0401_),
    .A2(_1436_),
    .A1(net572));
 sg13g2_nand4_1 _2581_ (.B(_0388_),
    .C(_0395_),
    .A(_0384_),
    .Y(_0403_),
    .D(net1325));
 sg13g2_xnor2_1 _2582_ (.Y(_0404_),
    .A(_0396_),
    .B(_0402_));
 sg13g2_o21ai_1 _2583_ (.B1(net1150),
    .Y(_0405_),
    .A1(_1630_),
    .A2(_0404_));
 sg13g2_and2_1 _2584_ (.A(net684),
    .B(net1151),
    .X(_0082_));
 sg13g2_nand2_1 _2585_ (.Y(_0406_),
    .A(net965),
    .B(_0358_));
 sg13g2_nor2_1 _2586_ (.A(net965),
    .B(net572),
    .Y(_0407_));
 sg13g2_o21ai_1 _2587_ (.B1(_0407_),
    .Y(_0408_),
    .A1(_1418_),
    .A2(_0361_));
 sg13g2_o21ai_1 _2588_ (.B1(_0408_),
    .Y(_0409_),
    .A1(net821),
    .A2(net598));
 sg13g2_a21oi_1 _2589_ (.A1(net1326),
    .A2(_0409_),
    .Y(_0410_),
    .B1(_1630_));
 sg13g2_o21ai_1 _2590_ (.B1(_0410_),
    .Y(_0411_),
    .A1(_0403_),
    .A2(_0409_));
 sg13g2_a21oi_1 _2591_ (.A1(net966),
    .A2(_0411_),
    .Y(_0083_),
    .B1(net646));
 sg13g2_a22oi_1 _2592_ (.Y(_0412_),
    .B1(net560),
    .B2(net320),
    .A2(net596),
    .A1(net863));
 sg13g2_nor2_1 _2593_ (.A(net648),
    .B(net321),
    .Y(_0084_));
 sg13g2_a22oi_1 _2594_ (.Y(_0413_),
    .B1(net560),
    .B2(net1321),
    .A2(net596),
    .A1(net747));
 sg13g2_nor2_1 _2595_ (.A(net646),
    .B(net748),
    .Y(_0085_));
 sg13g2_a22oi_1 _2596_ (.Y(_0414_),
    .B1(net560),
    .B2(\comm_ic0.uart0.clk_cnt_reg[2] ),
    .A2(net596),
    .A1(net466));
 sg13g2_nor2_1 _2597_ (.A(net648),
    .B(net467),
    .Y(_0086_));
 sg13g2_a22oi_1 _2598_ (.Y(_0415_),
    .B1(_0357_),
    .B2(\comm_ic0.uart0.clk_cnt_reg[3] ),
    .A2(net597),
    .A1(net783));
 sg13g2_nor2_1 _2599_ (.A(net649),
    .B(net784),
    .Y(_0087_));
 sg13g2_a22oi_1 _2600_ (.Y(_0416_),
    .B1(net560),
    .B2(\comm_ic0.uart0.clk_cnt_reg[4] ),
    .A2(net596),
    .A1(net780));
 sg13g2_nor2_1 _2601_ (.A(net646),
    .B(net781),
    .Y(_0088_));
 sg13g2_a22oi_1 _2602_ (.Y(_0417_),
    .B1(net560),
    .B2(\comm_ic0.uart0.clk_cnt_reg[5] ),
    .A2(net596),
    .A1(net711));
 sg13g2_nor2_1 _2603_ (.A(net646),
    .B(net712),
    .Y(_0089_));
 sg13g2_a22oi_1 _2604_ (.Y(_0418_),
    .B1(net560),
    .B2(net456),
    .A2(net596),
    .A1(net395));
 sg13g2_nor2_1 _2605_ (.A(net646),
    .B(net457),
    .Y(_0090_));
 sg13g2_a22oi_1 _2606_ (.Y(_0419_),
    .B1(net560),
    .B2(net838),
    .A2(net596),
    .A1(net821));
 sg13g2_nor2_1 _2607_ (.A(net645),
    .B(net839),
    .Y(_0091_));
 sg13g2_nor2b_1 _2608_ (.A(net1139),
    .B_N(\comm_ic0.uart0.curr_st[0] ),
    .Y(_0420_));
 sg13g2_nor2b_1 _2609_ (.A(net1016),
    .B_N(\comm_ic0.uart0.clk_cnt_reg[3] ),
    .Y(_0421_));
 sg13g2_nor2b_1 _2610_ (.A(\comm_ic0.uart0.clk_cnt_reg[3] ),
    .B_N(net1016),
    .Y(_0422_));
 sg13g2_xor2_1 _2611_ (.B(net1084),
    .A(net456),
    .X(_0423_));
 sg13g2_nand2b_1 _2612_ (.Y(_0424_),
    .B(\comm_ic0.uart0.uclk_cnt[6] ),
    .A_N(net838));
 sg13g2_xor2_1 _2613_ (.B(net1013),
    .A(\comm_ic0.uart0.clk_cnt_reg[2] ),
    .X(_0425_));
 sg13g2_o21ai_1 _2614_ (.B1(_0424_),
    .Y(_0426_),
    .A1(net1321),
    .A2(_1420_));
 sg13g2_nor4_1 _2615_ (.A(_0421_),
    .B(_0423_),
    .C(_0425_),
    .D(_0426_),
    .Y(_0427_));
 sg13g2_a22oi_1 _2616_ (.Y(_0428_),
    .B1(_1420_),
    .B2(net1321),
    .A2(_1419_),
    .A1(net838));
 sg13g2_xnor2_1 _2617_ (.Y(_0429_),
    .A(\comm_ic0.uart0.clk_cnt_reg[4] ),
    .B(net1051));
 sg13g2_xor2_1 _2618_ (.B(net1010),
    .A(\comm_ic0.uart0.clk_cnt_reg[5] ),
    .X(_0430_));
 sg13g2_nor4_1 _2619_ (.A(net965),
    .B(net572),
    .C(_0422_),
    .D(_0430_),
    .Y(_0431_));
 sg13g2_nand4_1 _2620_ (.B(_0428_),
    .C(_0429_),
    .A(_0427_),
    .Y(_0432_),
    .D(_0431_));
 sg13g2_o21ai_1 _2621_ (.B1(net1322),
    .Y(_0433_),
    .A1(net613),
    .A2(_0373_));
 sg13g2_nor3_1 _2622_ (.A(net649),
    .B(net1140),
    .C(net1323),
    .Y(_0092_));
 sg13g2_a22oi_1 _2623_ (.Y(_0434_),
    .B1(net560),
    .B2(\comm_ic0.uart0.par_odd ),
    .A2(net597),
    .A1(net801));
 sg13g2_nor2_1 _2624_ (.A(net658),
    .B(net802),
    .Y(_0093_));
 sg13g2_a22oi_1 _2625_ (.Y(_0435_),
    .B1(_0357_),
    .B2(net612),
    .A2(net597),
    .A1(net760));
 sg13g2_nor2_1 _2626_ (.A(net657),
    .B(net761),
    .Y(_0094_));
 sg13g2_nand2b_1 _2627_ (.Y(_0436_),
    .B(\comm_ic0.uart0.tx_ind[1] ),
    .A_N(\comm_ic0.uart0.tx_ind[0] ));
 sg13g2_nor2_1 _2628_ (.A(\comm_ic0.uart0.tx_data_reg[2] ),
    .B(_0436_),
    .Y(_0437_));
 sg13g2_nand2_1 _2629_ (.Y(_0438_),
    .A(\comm_ic0.uart0.tx_ind[0] ),
    .B(\comm_ic0.uart0.tx_ind[1] ));
 sg13g2_or2_1 _2630_ (.X(_0439_),
    .B(_0438_),
    .A(\comm_ic0.uart0.tx_data_reg[3] ));
 sg13g2_nand2b_1 _2631_ (.Y(_0440_),
    .B(\comm_ic0.uart0.tx_ind[0] ),
    .A_N(\comm_ic0.uart0.tx_ind[1] ));
 sg13g2_nor3_1 _2632_ (.A(\comm_ic0.uart0.tx_data_reg[0] ),
    .B(\comm_ic0.uart0.tx_ind[0] ),
    .C(\comm_ic0.uart0.tx_ind[1] ),
    .Y(_0441_));
 sg13g2_o21ai_1 _2633_ (.B1(_0439_),
    .Y(_0442_),
    .A1(\comm_ic0.uart0.tx_data_reg[1] ),
    .A2(_0440_));
 sg13g2_nor4_1 _2634_ (.A(\comm_ic0.uart0.tx_ind[2] ),
    .B(_0437_),
    .C(_0441_),
    .D(_0442_),
    .Y(_0443_));
 sg13g2_nor3_1 _2635_ (.A(\comm_ic0.uart0.tx_data_reg[4] ),
    .B(\comm_ic0.uart0.tx_ind[0] ),
    .C(\comm_ic0.uart0.tx_ind[1] ),
    .Y(_0444_));
 sg13g2_nor2_1 _2636_ (.A(\comm_ic0.uart0.tx_data_reg[5] ),
    .B(_0440_),
    .Y(_0445_));
 sg13g2_nor2_1 _2637_ (.A(\comm_ic0.uart0.tx_data_reg[6] ),
    .B(_0436_),
    .Y(_0446_));
 sg13g2_o21ai_1 _2638_ (.B1(\comm_ic0.uart0.tx_ind[2] ),
    .Y(_0447_),
    .A1(\comm_ic0.uart0.tx_data_reg[7] ),
    .A2(_0438_));
 sg13g2_nor4_1 _2639_ (.A(_0444_),
    .B(_0445_),
    .C(_0446_),
    .D(_0447_),
    .Y(_0448_));
 sg13g2_o21ai_1 _2640_ (.B1(_1433_),
    .Y(_0449_),
    .A1(_0443_),
    .A2(_0448_));
 sg13g2_mux2_1 _2641_ (.A0(\comm_ic0.uart0.tx_data_reg[8] ),
    .A1(\comm_ic0.uart0.tx_data_reg[9] ),
    .S(\comm_ic0.uart0.tx_ind[0] ),
    .X(_0450_));
 sg13g2_nand4_1 _2642_ (.B(_0060_),
    .C(_0059_),
    .A(\comm_ic0.uart0.tx_ind[3] ),
    .Y(_0451_),
    .D(_0450_));
 sg13g2_nor2_1 _2643_ (.A(_1412_),
    .B(net657),
    .Y(_0452_));
 sg13g2_nand3_1 _2644_ (.B(_0451_),
    .C(net546),
    .A(_0449_),
    .Y(_0095_));
 sg13g2_o21ai_1 _2645_ (.B1(\comm_ic0.uart0.tx_ind[2] ),
    .Y(_0453_),
    .A1(\comm_ic0.uart0.tx_ind[0] ),
    .A2(\comm_ic0.uart0.tx_ind[1] ));
 sg13g2_nand2b_1 _2646_ (.Y(_0454_),
    .B(_0453_),
    .A_N(_0355_));
 sg13g2_and2_1 _2647_ (.A(net546),
    .B(_0454_),
    .X(_0096_));
 sg13g2_nor3_1 _2648_ (.A(_1407_),
    .B(net1106),
    .C(net638),
    .Y(_0455_));
 sg13g2_and2_2 _2649_ (.A(\comm_ic0.spi0.start ),
    .B(net549),
    .X(_0456_));
 sg13g2_nand2_1 _2650_ (.Y(_0457_),
    .A(_1388_),
    .B(_0456_));
 sg13g2_a21oi_1 _2651_ (.A1(net1134),
    .A2(_1451_),
    .Y(_0458_),
    .B1(net1106));
 sg13g2_o21ai_1 _2652_ (.B1(_0458_),
    .Y(_0459_),
    .A1(_1434_),
    .A2(_1456_));
 sg13g2_nand2_1 _2653_ (.Y(_0460_),
    .A(net638),
    .B(_1456_));
 sg13g2_nand2_2 _2654_ (.Y(_0461_),
    .A(_1613_),
    .B(_0460_));
 sg13g2_a22oi_1 _2655_ (.Y(_0462_),
    .B1(_0461_),
    .B2(_1404_),
    .A2(_0459_),
    .A1(net1235));
 sg13g2_o21ai_1 _2656_ (.B1(_0457_),
    .Y(_0463_),
    .A1(net549),
    .A2(net1236));
 sg13g2_and2_1 _2657_ (.A(net685),
    .B(net1237),
    .X(_0097_));
 sg13g2_nor2_1 _2658_ (.A(net930),
    .B(net962),
    .Y(_0464_));
 sg13g2_nor2_1 _2659_ (.A(_1387_),
    .B(_1388_),
    .Y(_0465_));
 sg13g2_o21ai_1 _2660_ (.B1(_0456_),
    .Y(_0466_),
    .A1(_0464_),
    .A2(_0465_));
 sg13g2_xnor2_1 _2661_ (.Y(_0467_),
    .A(net1234),
    .B(net1265));
 sg13g2_xnor2_1 _2662_ (.Y(_0468_),
    .A(\comm_ic0.spi0.clk_cnt_reg[1] ),
    .B(\comm_ic0.spi0.clk_cnt_reg[0] ));
 sg13g2_a22oi_1 _2663_ (.Y(_0469_),
    .B1(_0468_),
    .B2(_0461_),
    .A2(net1266),
    .A1(_0459_));
 sg13g2_o21ai_1 _2664_ (.B1(_0466_),
    .Y(_0470_),
    .A1(net549),
    .A2(net1267));
 sg13g2_and2_1 _2665_ (.A(net685),
    .B(net1268),
    .X(_0098_));
 sg13g2_nand2_1 _2666_ (.Y(_0471_),
    .A(net1172),
    .B(_0464_));
 sg13g2_xnor2_1 _2667_ (.Y(_0472_),
    .A(net1172),
    .B(_0464_));
 sg13g2_nand2_1 _2668_ (.Y(_0473_),
    .A(_0456_),
    .B(net1173));
 sg13g2_nand2_1 _2669_ (.Y(_0474_),
    .A(net1239),
    .B(_1452_));
 sg13g2_xnor2_1 _2670_ (.Y(_0475_),
    .A(_0062_),
    .B(_1452_));
 sg13g2_nor3_1 _2671_ (.A(net880),
    .B(\comm_ic0.spi0.clk_cnt_reg[1] ),
    .C(\comm_ic0.spi0.clk_cnt_reg[0] ),
    .Y(_0476_));
 sg13g2_o21ai_1 _2672_ (.B1(net880),
    .Y(_0477_),
    .A1(\comm_ic0.spi0.clk_cnt_reg[1] ),
    .A2(\comm_ic0.spi0.clk_cnt_reg[0] ));
 sg13g2_nand2b_1 _2673_ (.Y(_0478_),
    .B(_0477_),
    .A_N(_0476_));
 sg13g2_a22oi_1 _2674_ (.Y(_0479_),
    .B1(_0478_),
    .B2(_0461_),
    .A2(_0475_),
    .A1(_0459_));
 sg13g2_o21ai_1 _2675_ (.B1(net1174),
    .Y(_0480_),
    .A1(net549),
    .A2(_0479_));
 sg13g2_and2_1 _2676_ (.A(net682),
    .B(net1175),
    .X(_0099_));
 sg13g2_nor4_2 _2677_ (.A(net992),
    .B(net880),
    .C(\comm_ic0.spi0.clk_cnt_reg[1] ),
    .Y(_0481_),
    .D(\comm_ic0.spi0.clk_cnt_reg[0] ));
 sg13g2_inv_1 _2678_ (.Y(_0482_),
    .A(_0481_));
 sg13g2_xor2_1 _2679_ (.B(_0476_),
    .A(net992),
    .X(_0483_));
 sg13g2_xnor2_1 _2680_ (.Y(_0484_),
    .A(\comm_ic0.spi0.sclk_cnt[3] ),
    .B(net1240));
 sg13g2_a22oi_1 _2681_ (.Y(_0485_),
    .B1(net1241),
    .B2(_0459_),
    .A2(_0483_),
    .A1(_0461_));
 sg13g2_xnor2_1 _2682_ (.Y(_0486_),
    .A(net983),
    .B(_0471_));
 sg13g2_nand2_1 _2683_ (.Y(_0487_),
    .A(_0456_),
    .B(_0486_));
 sg13g2_o21ai_1 _2684_ (.B1(_0487_),
    .Y(_0488_),
    .A1(net549),
    .A2(net1242));
 sg13g2_and2_1 _2685_ (.A(net682),
    .B(net1243),
    .X(_0100_));
 sg13g2_nor4_2 _2686_ (.A(net983),
    .B(net844),
    .C(net930),
    .Y(_0489_),
    .D(net962));
 sg13g2_nand2_1 _2687_ (.Y(_0490_),
    .A(net1163),
    .B(_0489_));
 sg13g2_xnor2_1 _2688_ (.Y(_0491_),
    .A(net1163),
    .B(_0489_));
 sg13g2_nand2_1 _2689_ (.Y(_0492_),
    .A(_0456_),
    .B(net1164));
 sg13g2_nor2_1 _2690_ (.A(_1439_),
    .B(_1453_),
    .Y(_0493_));
 sg13g2_xnor2_1 _2691_ (.Y(_0494_),
    .A(_1439_),
    .B(_1453_));
 sg13g2_xor2_1 _2692_ (.B(_0481_),
    .A(net828),
    .X(_0495_));
 sg13g2_a22oi_1 _2693_ (.Y(_0496_),
    .B1(_0495_),
    .B2(_0461_),
    .A2(_0494_),
    .A1(_0459_));
 sg13g2_o21ai_1 _2694_ (.B1(net1165),
    .Y(_0497_),
    .A1(net549),
    .A2(_0496_));
 sg13g2_and2_1 _2695_ (.A(net682),
    .B(net1166),
    .X(_0101_));
 sg13g2_nor3_2 _2696_ (.A(net911),
    .B(net828),
    .C(_0482_),
    .Y(_0498_));
 sg13g2_o21ai_1 _2697_ (.B1(net911),
    .Y(_0499_),
    .A1(net828),
    .A2(_0482_));
 sg13g2_nand2b_1 _2698_ (.Y(_0500_),
    .B(_0499_),
    .A_N(_0498_));
 sg13g2_xnor2_1 _2699_ (.Y(_0501_),
    .A(net1222),
    .B(_0493_));
 sg13g2_a22oi_1 _2700_ (.Y(_0502_),
    .B1(net1223),
    .B2(_0459_),
    .A2(_0500_),
    .A1(_0461_));
 sg13g2_xnor2_1 _2701_ (.Y(_0503_),
    .A(net865),
    .B(_0490_));
 sg13g2_nand2_1 _2702_ (.Y(_0504_),
    .A(_0456_),
    .B(_0503_));
 sg13g2_o21ai_1 _2703_ (.B1(_0504_),
    .Y(_0505_),
    .A1(_0455_),
    .A2(net1224));
 sg13g2_and2_1 _2704_ (.A(net682),
    .B(net1225),
    .X(_0102_));
 sg13g2_nor2_1 _2705_ (.A(net865),
    .B(net792),
    .Y(_0506_));
 sg13g2_and3_1 _2706_ (.X(_0507_),
    .A(net1177),
    .B(_0489_),
    .C(_0506_));
 sg13g2_a21oi_1 _2707_ (.A1(_0489_),
    .A2(_0506_),
    .Y(_0508_),
    .B1(net1177));
 sg13g2_o21ai_1 _2708_ (.B1(_0456_),
    .Y(_0509_),
    .A1(_0507_),
    .A2(net1178));
 sg13g2_o21ai_1 _2709_ (.B1(\comm_ic0.spi0.sclk_cnt[6] ),
    .Y(_0510_),
    .A1(_1453_),
    .A2(_1454_));
 sg13g2_nand2b_1 _2710_ (.Y(_0511_),
    .B(_0510_),
    .A_N(_1455_));
 sg13g2_nand2b_1 _2711_ (.Y(_0512_),
    .B(_0498_),
    .A_N(net744));
 sg13g2_xor2_1 _2712_ (.B(_0498_),
    .A(net744),
    .X(_0513_));
 sg13g2_a22oi_1 _2713_ (.Y(_0514_),
    .B1(_0513_),
    .B2(_0461_),
    .A2(_0511_),
    .A1(_0459_));
 sg13g2_o21ai_1 _2714_ (.B1(net1179),
    .Y(_0515_),
    .A1(net549),
    .A2(_0514_));
 sg13g2_and2_1 _2715_ (.A(net682),
    .B(net1180),
    .X(_0103_));
 sg13g2_xor2_1 _2716_ (.B(_1455_),
    .A(\comm_ic0.spi0.sclk_cnt[7] ),
    .X(_0516_));
 sg13g2_xnor2_1 _2717_ (.Y(_0517_),
    .A(net1251),
    .B(_0512_));
 sg13g2_a22oi_1 _2718_ (.Y(_0518_),
    .B1(net1252),
    .B2(_0461_),
    .A2(_0516_),
    .A1(_0459_));
 sg13g2_xnor2_1 _2719_ (.Y(_0519_),
    .A(_1356_),
    .B(_0507_));
 sg13g2_nand2_1 _2720_ (.Y(_0520_),
    .A(_0456_),
    .B(_0519_));
 sg13g2_o21ai_1 _2721_ (.B1(_0520_),
    .Y(_0521_),
    .A1(net549),
    .A2(net1253));
 sg13g2_and2_1 _2722_ (.A(net682),
    .B(net1254),
    .X(_0104_));
 sg13g2_nand2b_1 _2723_ (.Y(_0522_),
    .B(\comm_ic0.uart0.rx_data_reg[0] ),
    .A_N(\comm_ic0.uart0.rx_data_reg[9] ));
 sg13g2_nand2_1 _2724_ (.Y(_0523_),
    .A(_0030_),
    .B(_0522_));
 sg13g2_nand3_1 _2725_ (.B(net693),
    .C(_0523_),
    .A(\comm_ic0.uart0.rx_st[1] ),
    .Y(_0524_));
 sg13g2_and2_1 _2726_ (.A(net611),
    .B(\comm_ic0.uart0.par_odd ),
    .X(_0525_));
 sg13g2_nor2_1 _2727_ (.A(\comm_ic0.uart0.rx_data_reg[10] ),
    .B(_1414_),
    .Y(_0526_));
 sg13g2_nand2b_1 _2728_ (.Y(_0527_),
    .B(\comm_ic0.uart0.rx_data_reg[0] ),
    .A_N(\comm_ic0.uart0.rx_data_reg[10] ));
 sg13g2_xnor2_1 _2729_ (.Y(_0528_),
    .A(\comm_ic0.uart0.rx_data_reg[3] ),
    .B(\comm_ic0.uart0.rx_data_reg[2] ));
 sg13g2_xor2_1 _2730_ (.B(\comm_ic0.uart0.rx_data_reg[8] ),
    .A(\comm_ic0.uart0.rx_data_reg[9] ),
    .X(_0529_));
 sg13g2_xnor2_1 _2731_ (.Y(_0530_),
    .A(_0528_),
    .B(_0529_));
 sg13g2_xnor2_1 _2732_ (.Y(_0531_),
    .A(\comm_ic0.uart0.rx_data_reg[7] ),
    .B(\comm_ic0.uart0.rx_data_reg[6] ));
 sg13g2_xnor2_1 _2733_ (.Y(_0532_),
    .A(\comm_ic0.uart0.rx_data_reg[5] ),
    .B(_0531_));
 sg13g2_xnor2_1 _2734_ (.Y(_0533_),
    .A(\comm_ic0.uart0.rx_data_reg[4] ),
    .B(\comm_ic0.uart0.rx_data_reg[1] ));
 sg13g2_xnor2_1 _2735_ (.Y(_0534_),
    .A(_0532_),
    .B(_0533_));
 sg13g2_xor2_1 _2736_ (.B(_0534_),
    .A(_0530_),
    .X(_0535_));
 sg13g2_xnor2_1 _2737_ (.Y(_0536_),
    .A(_0530_),
    .B(_0534_));
 sg13g2_o21ai_1 _2738_ (.B1(_0525_),
    .Y(_0537_),
    .A1(_0527_),
    .A2(_0536_));
 sg13g2_nor2_1 _2739_ (.A(_1417_),
    .B(\comm_ic0.uart0.par_odd ),
    .Y(_0538_));
 sg13g2_o21ai_1 _2740_ (.B1(_0538_),
    .Y(_0539_),
    .A1(_0527_),
    .A2(_0535_));
 sg13g2_a21oi_1 _2741_ (.A1(_0537_),
    .A2(_0539_),
    .Y(_0540_),
    .B1(_0029_));
 sg13g2_nor2_1 _2742_ (.A(\comm_ic0.rx_ack ),
    .B(_1583_),
    .Y(_0541_));
 sg13g2_or3_1 _2743_ (.A(_0524_),
    .B(_0540_),
    .C(_0541_),
    .X(_0542_));
 sg13g2_o21ai_1 _2744_ (.B1(\comm_ic0.uart0.rx_st[0] ),
    .Y(_0543_),
    .A1(_1416_),
    .A2(_0523_));
 sg13g2_nor3_1 _2745_ (.A(_0540_),
    .B(_0541_),
    .C(_0543_),
    .Y(_0544_));
 sg13g2_nand2_1 _2746_ (.Y(_0545_),
    .A(\comm_ic0.rx_new ),
    .B(net693));
 sg13g2_o21ai_1 _2747_ (.B1(_0542_),
    .Y(_0105_),
    .A1(_0544_),
    .A2(_0545_));
 sg13g2_nand3_1 _2748_ (.B(_0536_),
    .C(_0538_),
    .A(_0526_),
    .Y(_0546_));
 sg13g2_nor3_1 _2749_ (.A(_1435_),
    .B(_0029_),
    .C(_0522_),
    .Y(_0547_));
 sg13g2_nand2b_1 _2750_ (.Y(_0548_),
    .B(\comm_ic0.uart0.rx_st[1] ),
    .A_N(\comm_ic0.uart0.rx_st[0] ));
 sg13g2_a21oi_1 _2751_ (.A1(_1610_),
    .A2(_0548_),
    .Y(_0549_),
    .B1(_0547_));
 sg13g2_nand3_1 _2752_ (.B(_0526_),
    .C(_0535_),
    .A(_0525_),
    .Y(_0550_));
 sg13g2_nand3_1 _2753_ (.B(_0549_),
    .C(_0550_),
    .A(_0546_),
    .Y(_0551_));
 sg13g2_a221oi_1 _2754_ (.B2(_1415_),
    .C1(net658),
    .B1(_0551_),
    .A1(_1416_),
    .Y(_0106_),
    .A2(_0549_));
 sg13g2_nor2_1 _2755_ (.A(\comm_ic0.uart0.rx_st[2] ),
    .B(\comm_ic0.uart0.rx_st[0] ),
    .Y(_0552_));
 sg13g2_o21ai_1 _2756_ (.B1(_0033_),
    .Y(_0553_),
    .A1(\comm_ic0.uart0.rx_st[2] ),
    .A2(\comm_ic0.uart0.rx_st[0] ));
 sg13g2_o21ai_1 _2757_ (.B1(_1414_),
    .Y(_0554_),
    .A1(_1608_),
    .A2(_0553_));
 sg13g2_nor2_1 _2758_ (.A(net1),
    .B(_0553_),
    .Y(_0555_));
 sg13g2_and2_1 _2759_ (.A(net693),
    .B(_0552_),
    .X(_0556_));
 sg13g2_o21ai_1 _2760_ (.B1(_0554_),
    .Y(_0557_),
    .A1(_1628_),
    .A2(net544));
 sg13g2_a21oi_1 _2761_ (.A1(_1609_),
    .A2(_0555_),
    .Y(_0107_),
    .B1(_0557_));
 sg13g2_xnor2_1 _2762_ (.Y(_0558_),
    .A(\comm_ic0.uart0.rx_ind[3] ),
    .B(_1607_));
 sg13g2_inv_1 _2763_ (.Y(_0559_),
    .A(_0558_));
 sg13g2_nand2_1 _2764_ (.Y(_0560_),
    .A(\comm_ic0.uart0.rx_ind[1] ),
    .B(\comm_ic0.uart0.rx_ind[0] ));
 sg13g2_nand2b_1 _2765_ (.Y(_0561_),
    .B(_0560_),
    .A_N(_1606_));
 sg13g2_nand2_2 _2766_ (.Y(_0562_),
    .A(net1),
    .B(_1608_));
 sg13g2_nor3_1 _2767_ (.A(_0033_),
    .B(_1629_),
    .C(_0562_),
    .Y(_0563_));
 sg13g2_nand2b_1 _2768_ (.Y(_0564_),
    .B(_0563_),
    .A_N(_0561_));
 sg13g2_or2_1 _2769_ (.X(_0565_),
    .B(_0564_),
    .A(net555));
 sg13g2_nand2b_1 _2770_ (.Y(_0566_),
    .B(\comm_ic0.uart0.rx_ind[0] ),
    .A_N(\comm_ic0.uart0.rx_ind[1] ));
 sg13g2_nor3_1 _2771_ (.A(\comm_ic0.uart0.rx_ind[3] ),
    .B(net555),
    .C(_0566_),
    .Y(_0567_));
 sg13g2_nor2_1 _2772_ (.A(_1629_),
    .B(_0567_),
    .Y(_0568_));
 sg13g2_o21ai_1 _2773_ (.B1(\comm_ic0.uart0.rx_data_reg[1] ),
    .Y(_0569_),
    .A1(net543),
    .A2(_0568_));
 sg13g2_o21ai_1 _2774_ (.B1(_0569_),
    .Y(_0108_),
    .A1(_0559_),
    .A2(_0565_));
 sg13g2_nand2b_2 _2775_ (.Y(_0570_),
    .B(\comm_ic0.uart0.rx_ind[1] ),
    .A_N(\comm_ic0.uart0.rx_ind[0] ));
 sg13g2_nor2_1 _2776_ (.A(net555),
    .B(_0570_),
    .Y(_0571_));
 sg13g2_nor3_1 _2777_ (.A(\comm_ic0.uart0.rx_ind[3] ),
    .B(net555),
    .C(_0570_),
    .Y(_0572_));
 sg13g2_o21ai_1 _2778_ (.B1(_1628_),
    .Y(_0573_),
    .A1(\comm_ic0.uart0.rx_data_reg[2] ),
    .A2(_0572_));
 sg13g2_a21oi_1 _2779_ (.A1(_0562_),
    .A2(_0572_),
    .Y(_0574_),
    .B1(_0573_));
 sg13g2_a21o_1 _2780_ (.A2(net543),
    .A1(\comm_ic0.uart0.rx_data_reg[2] ),
    .B1(_0574_),
    .X(_0109_));
 sg13g2_xnor2_1 _2781_ (.Y(_0575_),
    .A(net555),
    .B(_1606_));
 sg13g2_nand2_1 _2782_ (.Y(_0576_),
    .A(_1413_),
    .B(_0575_));
 sg13g2_nand2_1 _2783_ (.Y(_0577_),
    .A(_0561_),
    .B(_0563_));
 sg13g2_nor2_1 _2784_ (.A(_0560_),
    .B(_0576_),
    .Y(_0578_));
 sg13g2_nor2_1 _2785_ (.A(_1629_),
    .B(_0578_),
    .Y(_0579_));
 sg13g2_o21ai_1 _2786_ (.B1(\comm_ic0.uart0.rx_data_reg[3] ),
    .Y(_0580_),
    .A1(net543),
    .A2(_0579_));
 sg13g2_o21ai_1 _2787_ (.B1(_0580_),
    .Y(_0110_),
    .A1(_0576_),
    .A2(_0577_));
 sg13g2_nor3_1 _2788_ (.A(\comm_ic0.uart0.rx_ind[1] ),
    .B(\comm_ic0.uart0.rx_ind[0] ),
    .C(_0576_),
    .Y(_0581_));
 sg13g2_o21ai_1 _2789_ (.B1(_1628_),
    .Y(_0582_),
    .A1(\comm_ic0.uart0.rx_data_reg[4] ),
    .A2(_0581_));
 sg13g2_a21oi_1 _2790_ (.A1(_0562_),
    .A2(_0581_),
    .Y(_0583_),
    .B1(_0582_));
 sg13g2_a21o_1 _2791_ (.A2(net543),
    .A1(\comm_ic0.uart0.rx_data_reg[4] ),
    .B1(_0583_),
    .X(_0111_));
 sg13g2_nand2b_2 _2792_ (.Y(_0584_),
    .B(_0558_),
    .A_N(_0575_));
 sg13g2_nor2_1 _2793_ (.A(_0566_),
    .B(_0584_),
    .Y(_0585_));
 sg13g2_nor2_1 _2794_ (.A(_1629_),
    .B(_0585_),
    .Y(_0586_));
 sg13g2_o21ai_1 _2795_ (.B1(\comm_ic0.uart0.rx_data_reg[5] ),
    .Y(_0587_),
    .A1(net543),
    .A2(_0586_));
 sg13g2_o21ai_1 _2796_ (.B1(_0587_),
    .Y(_0112_),
    .A1(_0564_),
    .A2(_0584_));
 sg13g2_nor2_1 _2797_ (.A(_0570_),
    .B(_0584_),
    .Y(_0588_));
 sg13g2_o21ai_1 _2798_ (.B1(_1628_),
    .Y(_0589_),
    .A1(\comm_ic0.uart0.rx_data_reg[6] ),
    .A2(_0588_));
 sg13g2_a21oi_1 _2799_ (.A1(_0562_),
    .A2(_0588_),
    .Y(_0590_),
    .B1(_0589_));
 sg13g2_a21o_1 _2800_ (.A2(net543),
    .A1(\comm_ic0.uart0.rx_data_reg[6] ),
    .B1(_0590_),
    .X(_0113_));
 sg13g2_nor2_1 _2801_ (.A(_0560_),
    .B(_0584_),
    .Y(_0591_));
 sg13g2_nor2_1 _2802_ (.A(_1629_),
    .B(_0591_),
    .Y(_0592_));
 sg13g2_o21ai_1 _2803_ (.B1(\comm_ic0.uart0.rx_data_reg[7] ),
    .Y(_0593_),
    .A1(net543),
    .A2(_0592_));
 sg13g2_o21ai_1 _2804_ (.B1(_0593_),
    .Y(_0114_),
    .A1(_0577_),
    .A2(_0584_));
 sg13g2_nand2_1 _2805_ (.Y(_0594_),
    .A(\comm_ic0.uart0.rx_data_reg[8] ),
    .B(net544));
 sg13g2_nand2_1 _2806_ (.Y(_0595_),
    .A(\comm_ic0.uart0.rx_ind[3] ),
    .B(_1607_));
 sg13g2_a21oi_1 _2807_ (.A1(\comm_ic0.uart0.rx_ind[3] ),
    .A2(_1607_),
    .Y(_0596_),
    .B1(\comm_ic0.uart0.rx_data_reg[8] ));
 sg13g2_o21ai_1 _2808_ (.B1(_1628_),
    .Y(_0597_),
    .A1(net1),
    .A2(_0595_));
 sg13g2_o21ai_1 _2809_ (.B1(_0594_),
    .Y(_0115_),
    .A1(_0596_),
    .A2(_0597_));
 sg13g2_nor3_1 _2810_ (.A(_1413_),
    .B(net555),
    .C(_0566_),
    .Y(_0598_));
 sg13g2_nor2_1 _2811_ (.A(_1629_),
    .B(_0598_),
    .Y(_0599_));
 sg13g2_o21ai_1 _2812_ (.B1(\comm_ic0.uart0.rx_data_reg[9] ),
    .Y(_0600_),
    .A1(net543),
    .A2(_0599_));
 sg13g2_o21ai_1 _2813_ (.B1(_0600_),
    .Y(_0116_),
    .A1(_0558_),
    .A2(_0565_));
 sg13g2_nor4_1 _2814_ (.A(_1413_),
    .B(\comm_ic0.uart0.rx_ind[2] ),
    .C(net1),
    .D(_0570_),
    .Y(_0601_));
 sg13g2_a21oi_1 _2815_ (.A1(\comm_ic0.uart0.rx_ind[3] ),
    .A2(_0571_),
    .Y(_0602_),
    .B1(\comm_ic0.uart0.rx_data_reg[10] ));
 sg13g2_nor3_1 _2816_ (.A(_1629_),
    .B(_0601_),
    .C(_0602_),
    .Y(_0603_));
 sg13g2_a21o_1 _2817_ (.A2(net544),
    .A1(\comm_ic0.uart0.rx_data_reg[10] ),
    .B1(_0603_),
    .X(_0117_));
 sg13g2_nand2_1 _2818_ (.Y(_0604_),
    .A(\comm_ic0.uart0.rx_ind[0] ),
    .B(net544));
 sg13g2_nor2_2 _2819_ (.A(\comm_ic0.uart0.rx_st[2] ),
    .B(_1582_),
    .Y(_0605_));
 sg13g2_o21ai_1 _2820_ (.B1(net693),
    .Y(_0606_),
    .A1(\comm_ic0.uart0.rx_st[2] ),
    .A2(\comm_ic0.uart0.rx_st[0] ));
 sg13g2_a21oi_1 _2821_ (.A1(_1435_),
    .A2(_0605_),
    .Y(_0607_),
    .B1(_0606_));
 sg13g2_o21ai_1 _2822_ (.B1(_0607_),
    .Y(_0608_),
    .A1(_0033_),
    .A2(_0605_));
 sg13g2_nand2_1 _2823_ (.Y(_0118_),
    .A(_0604_),
    .B(_0608_));
 sg13g2_nand2_1 _2824_ (.Y(_0609_),
    .A(\comm_ic0.uart0.rx_ind[1] ),
    .B(net544));
 sg13g2_a21oi_1 _2825_ (.A1(_1417_),
    .A2(_0605_),
    .Y(_0610_),
    .B1(_0606_));
 sg13g2_o21ai_1 _2826_ (.B1(_0610_),
    .Y(_0611_),
    .A1(_0561_),
    .A2(_0605_));
 sg13g2_nand2_1 _2827_ (.Y(_0119_),
    .A(_0609_),
    .B(_0611_));
 sg13g2_nand2_1 _2828_ (.Y(_0612_),
    .A(net555),
    .B(net544));
 sg13g2_nor2_1 _2829_ (.A(_0552_),
    .B(_0605_),
    .Y(_0613_));
 sg13g2_xnor2_1 _2830_ (.Y(_0614_),
    .A(_0034_),
    .B(_1606_));
 sg13g2_nand3_1 _2831_ (.B(_0613_),
    .C(_0614_),
    .A(net693),
    .Y(_0615_));
 sg13g2_nand2_1 _2832_ (.Y(_0120_),
    .A(_0612_),
    .B(_0615_));
 sg13g2_a221oi_1 _2833_ (.B2(_0613_),
    .C1(net658),
    .B1(_0558_),
    .A1(_1413_),
    .Y(_0121_),
    .A2(_0552_));
 sg13g2_nand3b_1 _2834_ (.B(_0537_),
    .C(_0539_),
    .Y(_0616_),
    .A_N(_0524_));
 sg13g2_nand2b_1 _2835_ (.Y(_0617_),
    .B(net609),
    .A_N(\comm_ic0.uart0.rx_data_reg[2] ));
 sg13g2_o21ai_1 _2836_ (.B1(_0617_),
    .Y(_0618_),
    .A1(\comm_ic0.uart0.rx_data_reg[1] ),
    .A2(net610));
 sg13g2_nand2_1 _2837_ (.Y(_0619_),
    .A(\comm_ic0.rx_data[0] ),
    .B(net528));
 sg13g2_o21ai_1 _2838_ (.B1(_0619_),
    .Y(_0122_),
    .A1(net528),
    .A2(_0618_));
 sg13g2_nand2b_1 _2839_ (.Y(_0620_),
    .B(net608),
    .A_N(\comm_ic0.uart0.rx_data_reg[3] ));
 sg13g2_o21ai_1 _2840_ (.B1(_0620_),
    .Y(_0621_),
    .A1(\comm_ic0.uart0.rx_data_reg[2] ),
    .A2(net608));
 sg13g2_nand2_1 _2841_ (.Y(_0622_),
    .A(\comm_ic0.rx_data[1] ),
    .B(net527));
 sg13g2_o21ai_1 _2842_ (.B1(_0622_),
    .Y(_0123_),
    .A1(net528),
    .A2(_0621_));
 sg13g2_nand2b_1 _2843_ (.Y(_0623_),
    .B(net608),
    .A_N(\comm_ic0.uart0.rx_data_reg[4] ));
 sg13g2_o21ai_1 _2844_ (.B1(_0623_),
    .Y(_0624_),
    .A1(\comm_ic0.uart0.rx_data_reg[3] ),
    .A2(net608));
 sg13g2_nand2_1 _2845_ (.Y(_0625_),
    .A(\comm_ic0.rx_data[2] ),
    .B(net527));
 sg13g2_o21ai_1 _2846_ (.B1(_0625_),
    .Y(_0124_),
    .A1(net527),
    .A2(_0624_));
 sg13g2_nand2b_1 _2847_ (.Y(_0626_),
    .B(net608),
    .A_N(\comm_ic0.uart0.rx_data_reg[5] ));
 sg13g2_o21ai_1 _2848_ (.B1(_0626_),
    .Y(_0627_),
    .A1(\comm_ic0.uart0.rx_data_reg[4] ),
    .A2(net610));
 sg13g2_nand2_1 _2849_ (.Y(_0628_),
    .A(\comm_ic0.rx_data[3] ),
    .B(net528));
 sg13g2_o21ai_1 _2850_ (.B1(_0628_),
    .Y(_0125_),
    .A1(net528),
    .A2(_0627_));
 sg13g2_nand2b_1 _2851_ (.Y(_0629_),
    .B(net608),
    .A_N(\comm_ic0.uart0.rx_data_reg[6] ));
 sg13g2_o21ai_1 _2852_ (.B1(_0629_),
    .Y(_0630_),
    .A1(\comm_ic0.uart0.rx_data_reg[5] ),
    .A2(net609));
 sg13g2_nand2_1 _2853_ (.Y(_0631_),
    .A(\comm_ic0.rx_data[4] ),
    .B(net527));
 sg13g2_o21ai_1 _2854_ (.B1(_0631_),
    .Y(_0126_),
    .A1(net527),
    .A2(_0630_));
 sg13g2_nand2b_1 _2855_ (.Y(_0632_),
    .B(net608),
    .A_N(\comm_ic0.uart0.rx_data_reg[7] ));
 sg13g2_o21ai_1 _2856_ (.B1(_0632_),
    .Y(_0633_),
    .A1(\comm_ic0.uart0.rx_data_reg[6] ),
    .A2(net609));
 sg13g2_nand2_1 _2857_ (.Y(_0634_),
    .A(\comm_ic0.rx_data[5] ),
    .B(net527));
 sg13g2_o21ai_1 _2858_ (.B1(_0634_),
    .Y(_0127_),
    .A1(net528),
    .A2(_0633_));
 sg13g2_nand2b_1 _2859_ (.Y(_0635_),
    .B(net609),
    .A_N(\comm_ic0.uart0.rx_data_reg[8] ));
 sg13g2_o21ai_1 _2860_ (.B1(_0635_),
    .Y(_0636_),
    .A1(\comm_ic0.uart0.rx_data_reg[7] ),
    .A2(net608));
 sg13g2_nand2_1 _2861_ (.Y(_0637_),
    .A(\comm_ic0.rx_data[6] ),
    .B(net527));
 sg13g2_o21ai_1 _2862_ (.B1(_0637_),
    .Y(_0128_),
    .A1(net527),
    .A2(_0636_));
 sg13g2_nand2b_1 _2863_ (.Y(_0638_),
    .B(net611),
    .A_N(\comm_ic0.uart0.rx_data_reg[9] ));
 sg13g2_o21ai_1 _2864_ (.B1(_0638_),
    .Y(_0639_),
    .A1(\comm_ic0.uart0.rx_data_reg[8] ),
    .A2(net610));
 sg13g2_nand2_1 _2865_ (.Y(_0640_),
    .A(\comm_ic0.rx_data[7] ),
    .B(net528));
 sg13g2_o21ai_1 _2866_ (.B1(_0640_),
    .Y(_0129_),
    .A1(net528),
    .A2(_0639_));
 sg13g2_nand2b_1 _2867_ (.Y(_0641_),
    .B(_0356_),
    .A_N(\comm_ic0.busy_uart ));
 sg13g2_and2_1 _2868_ (.A(_0075_),
    .B(_0641_),
    .X(_0130_));
 sg13g2_a21o_1 _2869_ (.A2(net546),
    .A1(\comm_ic0.uart0.tx_data_reg[0] ),
    .B1(_1632_),
    .X(_0131_));
 sg13g2_xnor2_1 _2870_ (.Y(_0642_),
    .A(\comm_ic0.tx_data[5] ),
    .B(\comm_ic0.tx_data[4] ));
 sg13g2_xnor2_1 _2871_ (.Y(_0643_),
    .A(_1336_),
    .B(_0642_));
 sg13g2_xor2_1 _2872_ (.B(\comm_ic0.uart0.par_odd ),
    .A(\comm_ic0.tx_data[2] ),
    .X(_0644_));
 sg13g2_xnor2_1 _2873_ (.Y(_0645_),
    .A(\comm_ic0.tx_data[7] ),
    .B(\comm_ic0.tx_data[6] ));
 sg13g2_xor2_1 _2874_ (.B(\comm_ic0.tx_data[0] ),
    .A(\comm_ic0.tx_data[1] ),
    .X(_0646_));
 sg13g2_xnor2_1 _2875_ (.Y(_0647_),
    .A(_0645_),
    .B(_0646_));
 sg13g2_xnor2_1 _2876_ (.Y(_0648_),
    .A(_0644_),
    .B(_0647_));
 sg13g2_xnor2_1 _2877_ (.Y(_0649_),
    .A(_0643_),
    .B(_0648_));
 sg13g2_o21ai_1 _2878_ (.B1(_1632_),
    .Y(_0650_),
    .A1(\comm_ic0.tx_data[0] ),
    .A2(net607));
 sg13g2_a21oi_1 _2879_ (.A1(net606),
    .A2(_0649_),
    .Y(_0651_),
    .B1(_0650_));
 sg13g2_a21o_1 _2880_ (.A2(net545),
    .A1(\comm_ic0.uart0.tx_data_reg[1] ),
    .B1(_0651_),
    .X(_0132_));
 sg13g2_nand2_1 _2881_ (.Y(_0652_),
    .A(\comm_ic0.uart0.tx_data_reg[2] ),
    .B(net546));
 sg13g2_mux2_1 _2882_ (.A0(_1338_),
    .A1(_1339_),
    .S(net606),
    .X(_0653_));
 sg13g2_o21ai_1 _2883_ (.B1(_0652_),
    .Y(_0133_),
    .A1(net547),
    .A2(_0653_));
 sg13g2_nand2_1 _2884_ (.Y(_0654_),
    .A(\comm_ic0.uart0.tx_data_reg[3] ),
    .B(net545));
 sg13g2_mux2_1 _2885_ (.A0(_1337_),
    .A1(_1338_),
    .S(net606),
    .X(_0655_));
 sg13g2_o21ai_1 _2886_ (.B1(_0654_),
    .Y(_0134_),
    .A1(net547),
    .A2(_0655_));
 sg13g2_nand2_1 _2887_ (.Y(_0656_),
    .A(\comm_ic0.uart0.tx_data_reg[4] ),
    .B(net545));
 sg13g2_mux2_1 _2888_ (.A0(_1336_),
    .A1(_1337_),
    .S(net606),
    .X(_0657_));
 sg13g2_o21ai_1 _2889_ (.B1(_0656_),
    .Y(_0135_),
    .A1(_0354_),
    .A2(_0657_));
 sg13g2_o21ai_1 _2890_ (.B1(_1632_),
    .Y(_0658_),
    .A1(\comm_ic0.tx_data[4] ),
    .A2(net606));
 sg13g2_a21oi_1 _2891_ (.A1(_1336_),
    .A2(net606),
    .Y(_0659_),
    .B1(_0658_));
 sg13g2_a21o_1 _2892_ (.A2(net546),
    .A1(\comm_ic0.uart0.tx_data_reg[5] ),
    .B1(_0659_),
    .X(_0136_));
 sg13g2_nand2_1 _2893_ (.Y(_0660_),
    .A(\comm_ic0.uart0.tx_data_reg[6] ),
    .B(net545));
 sg13g2_mux2_1 _2894_ (.A0(_1376_),
    .A1(_1377_),
    .S(net606),
    .X(_0661_));
 sg13g2_o21ai_1 _2895_ (.B1(_0660_),
    .Y(_0137_),
    .A1(net547),
    .A2(_0661_));
 sg13g2_nand2_1 _2896_ (.Y(_0662_),
    .A(\comm_ic0.uart0.tx_data_reg[7] ),
    .B(net545));
 sg13g2_mux2_1 _2897_ (.A0(_1375_),
    .A1(_1376_),
    .S(net607),
    .X(_0663_));
 sg13g2_o21ai_1 _2898_ (.B1(_0662_),
    .Y(_0138_),
    .A1(net547),
    .A2(_0663_));
 sg13g2_nand2_1 _2899_ (.Y(_0664_),
    .A(\comm_ic0.uart0.tx_data_reg[8] ),
    .B(net545));
 sg13g2_mux2_1 _2900_ (.A0(_1374_),
    .A1(_1375_),
    .S(net607),
    .X(_0665_));
 sg13g2_o21ai_1 _2901_ (.B1(_0664_),
    .Y(_0139_),
    .A1(net547),
    .A2(_0665_));
 sg13g2_nand2_1 _2902_ (.Y(_0666_),
    .A(\comm_ic0.uart0.tx_data_reg[9] ),
    .B(net545));
 sg13g2_nand2_1 _2903_ (.Y(_0667_),
    .A(\comm_ic0.tx_data[7] ),
    .B(net607));
 sg13g2_o21ai_1 _2904_ (.B1(_0666_),
    .Y(_0140_),
    .A1(net547),
    .A2(_0667_));
 sg13g2_nand2_1 _2905_ (.Y(_0668_),
    .A(net1312),
    .B(net573));
 sg13g2_o21ai_1 _2906_ (.B1(_0668_),
    .Y(_0669_),
    .A1(net538),
    .A2(_1577_));
 sg13g2_nor2_2 _2907_ (.A(_1390_),
    .B(net591),
    .Y(_0670_));
 sg13g2_a21oi_1 _2908_ (.A1(net591),
    .A2(net899),
    .Y(_0671_),
    .B1(_0670_));
 sg13g2_o21ai_1 _2909_ (.B1(net686),
    .Y(_0672_),
    .A1(net1290),
    .A2(_0669_));
 sg13g2_a21oi_1 _2910_ (.A1(_0669_),
    .A2(net900),
    .Y(_0141_),
    .B1(_0672_));
 sg13g2_and2_2 _2911_ (.A(net1122),
    .B(net1290),
    .X(_0673_));
 sg13g2_o21ai_1 _2912_ (.B1(net591),
    .Y(_0674_),
    .A1(_1573_),
    .A2(_0673_));
 sg13g2_nor2b_1 _2913_ (.A(_0670_),
    .B_N(_0674_),
    .Y(_0675_));
 sg13g2_o21ai_1 _2914_ (.B1(net686),
    .Y(_0676_),
    .A1(net1122),
    .A2(_0669_));
 sg13g2_a21oi_1 _2915_ (.A1(_0669_),
    .A2(_0675_),
    .Y(_0142_),
    .B1(net1123));
 sg13g2_o21ai_1 _2916_ (.B1(_0669_),
    .Y(_0677_),
    .A1(net573),
    .A2(net562));
 sg13g2_a21o_1 _2917_ (.A2(_1574_),
    .A1(net591),
    .B1(_0670_),
    .X(_0678_));
 sg13g2_a22oi_1 _2918_ (.Y(_0679_),
    .B1(_0678_),
    .B2(_0669_),
    .A2(_0677_),
    .A1(net604));
 sg13g2_nor2_1 _2919_ (.A(net644),
    .B(net1263),
    .Y(_0143_));
 sg13g2_nand2b_1 _2920_ (.Y(_0680_),
    .B(net600),
    .A_N(_1574_));
 sg13g2_and2_1 _2921_ (.A(net602),
    .B(_1574_),
    .X(_0681_));
 sg13g2_a21oi_2 _2922_ (.B1(net573),
    .Y(_0682_),
    .A2(_0680_),
    .A1(_1576_));
 sg13g2_a21oi_1 _2923_ (.A1(net738),
    .A2(_0670_),
    .Y(_0683_),
    .B1(_0682_));
 sg13g2_o21ai_1 _2924_ (.B1(net686),
    .Y(_0684_),
    .A1(net1039),
    .A2(_0669_));
 sg13g2_a21oi_1 _2925_ (.A1(_0669_),
    .A2(_0683_),
    .Y(_0144_),
    .B1(net1040));
 sg13g2_nand2_1 _2926_ (.Y(_0685_),
    .A(net1312),
    .B(_1429_));
 sg13g2_o21ai_1 _2927_ (.B1(_0685_),
    .Y(_0686_),
    .A1(net538),
    .A2(_1571_));
 sg13g2_nor2_1 _2928_ (.A(_1390_),
    .B(net590),
    .Y(_0687_));
 sg13g2_a21oi_1 _2929_ (.A1(net589),
    .A2(net720),
    .Y(_0688_),
    .B1(_0687_));
 sg13g2_o21ai_1 _2930_ (.B1(net688),
    .Y(_0689_),
    .A1(net1299),
    .A2(_0686_));
 sg13g2_a21oi_1 _2931_ (.A1(_0686_),
    .A2(net721),
    .Y(_0145_),
    .B1(net1300));
 sg13g2_nand2_1 _2932_ (.Y(_0690_),
    .A(net1153),
    .B(net1299));
 sg13g2_o21ai_1 _2933_ (.B1(net589),
    .Y(_0691_),
    .A1(net1153),
    .A2(net1299));
 sg13g2_nand2b_1 _2934_ (.Y(_0692_),
    .B(_0690_),
    .A_N(_0691_));
 sg13g2_o21ai_1 _2935_ (.B1(_0692_),
    .Y(_0693_),
    .A1(net1213),
    .A2(net589));
 sg13g2_o21ai_1 _2936_ (.B1(net689),
    .Y(_0694_),
    .A1(net1153),
    .A2(_0686_));
 sg13g2_a21oi_1 _2937_ (.A1(_0686_),
    .A2(_0693_),
    .Y(_0146_),
    .B1(net1154));
 sg13g2_nand2_1 _2938_ (.Y(_0695_),
    .A(_0686_),
    .B(_0691_));
 sg13g2_a21oi_1 _2939_ (.A1(_0686_),
    .A2(_0691_),
    .Y(_0696_),
    .B1(net971));
 sg13g2_nor2_1 _2940_ (.A(net971),
    .B(_1429_),
    .Y(_0697_));
 sg13g2_nor3_1 _2941_ (.A(_0687_),
    .B(_0695_),
    .C(_0697_),
    .Y(_0698_));
 sg13g2_nor3_1 _2942_ (.A(net655),
    .B(net972),
    .C(_0698_),
    .Y(_0147_));
 sg13g2_a221oi_1 _2943_ (.B2(_1506_),
    .C1(_1479_),
    .B1(net1202),
    .A1(net579),
    .Y(_0699_),
    .A2(net580));
 sg13g2_nor2_1 _2944_ (.A(net986),
    .B(_0699_),
    .Y(_0700_));
 sg13g2_nor2b_1 _2945_ (.A(net636),
    .B_N(\comm_ic0.rx_data[4] ),
    .Y(_0701_));
 sg13g2_a21oi_1 _2946_ (.A1(net635),
    .A2(\comm_ic0.rx_data[0] ),
    .Y(_0702_),
    .B1(_0701_));
 sg13g2_o21ai_1 _2947_ (.B1(_0699_),
    .Y(_0703_),
    .A1(_1491_),
    .A2(_0702_));
 sg13g2_nand2_1 _2948_ (.Y(_0704_),
    .A(net789),
    .B(net633));
 sg13g2_a22oi_1 _2949_ (.Y(_0705_),
    .B1(net630),
    .B2(net516),
    .A2(net628),
    .A1(net495));
 sg13g2_a21oi_2 _2950_ (.B1(net563),
    .Y(_0706_),
    .A2(_0705_),
    .A1(_0704_));
 sg13g2_nand2_1 _2951_ (.Y(_0707_),
    .A(net1057),
    .B(net633));
 sg13g2_a22oi_1 _2952_ (.Y(_0708_),
    .B1(net630),
    .B2(net365),
    .A2(net628),
    .A1(net377));
 sg13g2_a21oi_1 _2953_ (.A1(_0707_),
    .A2(_0708_),
    .Y(_0709_),
    .B1(net566));
 sg13g2_a22oi_1 _2954_ (.Y(_0710_),
    .B1(net564),
    .B2(net795),
    .A2(_1463_),
    .A1(net714));
 sg13g2_nor2_1 _2955_ (.A(_1504_),
    .B(_0710_),
    .Y(_0711_));
 sg13g2_nor4_2 _2956_ (.A(_0703_),
    .B(_0706_),
    .C(_0709_),
    .Y(_0712_),
    .D(_0711_));
 sg13g2_nor2_1 _2957_ (.A(net987),
    .B(_0712_),
    .Y(_0148_));
 sg13g2_nor2_1 _2958_ (.A(net998),
    .B(_0699_),
    .Y(_0713_));
 sg13g2_nor2b_1 _2959_ (.A(net635),
    .B_N(\comm_ic0.rx_data[5] ),
    .Y(_0714_));
 sg13g2_a21oi_1 _2960_ (.A1(net635),
    .A2(\comm_ic0.rx_data[1] ),
    .Y(_0715_),
    .B1(_0714_));
 sg13g2_o21ai_1 _2961_ (.B1(_0699_),
    .Y(_0716_),
    .A1(_1491_),
    .A2(_0715_));
 sg13g2_nand2_1 _2962_ (.Y(_0717_),
    .A(net841),
    .B(net634));
 sg13g2_a22oi_1 _2963_ (.Y(_0718_),
    .B1(net630),
    .B2(net764),
    .A2(net627),
    .A1(net526));
 sg13g2_a21oi_1 _2964_ (.A1(_0717_),
    .A2(_0718_),
    .Y(_0719_),
    .B1(net565));
 sg13g2_nand2_1 _2965_ (.Y(_0720_),
    .A(net1022),
    .B(net637));
 sg13g2_a22oi_1 _2966_ (.Y(_0721_),
    .B1(net632),
    .B2(net860),
    .A2(net629),
    .A1(net874));
 sg13g2_a21oi_2 _2967_ (.B1(net563),
    .Y(_0722_),
    .A2(_0721_),
    .A1(_0720_));
 sg13g2_a22oi_1 _2968_ (.Y(_0723_),
    .B1(net564),
    .B2(net1330),
    .A2(_1463_),
    .A1(net735));
 sg13g2_nor2_1 _2969_ (.A(_1504_),
    .B(_0723_),
    .Y(_0724_));
 sg13g2_nor4_1 _2970_ (.A(_0716_),
    .B(_0719_),
    .C(_0722_),
    .D(_0724_),
    .Y(_0725_));
 sg13g2_nor2_1 _2971_ (.A(net999),
    .B(_0725_),
    .Y(_0149_));
 sg13g2_nor2_1 _2972_ (.A(net1001),
    .B(_0699_),
    .Y(_0726_));
 sg13g2_nor2b_1 _2973_ (.A(net635),
    .B_N(\comm_ic0.rx_data[6] ),
    .Y(_0727_));
 sg13g2_a21oi_1 _2974_ (.A1(net635),
    .A2(\comm_ic0.rx_data[2] ),
    .Y(_0728_),
    .B1(_0727_));
 sg13g2_o21ai_1 _2975_ (.B1(_0699_),
    .Y(_0729_),
    .A1(_1491_),
    .A2(_0728_));
 sg13g2_nand2_1 _2976_ (.Y(_0730_),
    .A(net786),
    .B(net630));
 sg13g2_a22oi_1 _2977_ (.Y(_0731_),
    .B1(net633),
    .B2(net798),
    .A2(net628),
    .A1(net741));
 sg13g2_a21oi_1 _2978_ (.A1(_0730_),
    .A2(_0731_),
    .Y(_0732_),
    .B1(net566));
 sg13g2_nand2_1 _2979_ (.Y(_0733_),
    .A(net895),
    .B(net633));
 sg13g2_a22oi_1 _2980_ (.Y(_0734_),
    .B1(net630),
    .B2(net889),
    .A2(net629),
    .A1(net717));
 sg13g2_a21oi_2 _2981_ (.B1(net563),
    .Y(_0735_),
    .A2(_0734_),
    .A1(_0733_));
 sg13g2_a22oi_1 _2982_ (.Y(_0736_),
    .B1(net564),
    .B2(net871),
    .A2(_1463_),
    .A1(net723));
 sg13g2_nor2_1 _2983_ (.A(_1504_),
    .B(_0736_),
    .Y(_0737_));
 sg13g2_nor4_2 _2984_ (.A(_0729_),
    .B(_0732_),
    .C(_0735_),
    .Y(_0738_),
    .D(_0737_));
 sg13g2_nor2_1 _2985_ (.A(net1002),
    .B(_0738_),
    .Y(_0150_));
 sg13g2_nor2_1 _2986_ (.A(net933),
    .B(_0699_),
    .Y(_0739_));
 sg13g2_nor2b_1 _2987_ (.A(net635),
    .B_N(\comm_ic0.rx_data[7] ),
    .Y(_0740_));
 sg13g2_a21oi_1 _2988_ (.A1(net635),
    .A2(\comm_ic0.rx_data[3] ),
    .Y(_0741_),
    .B1(_0740_));
 sg13g2_o21ai_1 _2989_ (.B1(_0699_),
    .Y(_0742_),
    .A1(_1491_),
    .A2(_0741_));
 sg13g2_nand2_1 _2990_ (.Y(_0743_),
    .A(net886),
    .B(net520));
 sg13g2_a22oi_1 _2991_ (.Y(_0744_),
    .B1(net630),
    .B2(net877),
    .A2(net629),
    .A1(net1087));
 sg13g2_a21oi_2 _2992_ (.B1(net563),
    .Y(_0745_),
    .A2(_0744_),
    .A1(_0743_));
 sg13g2_nand2_1 _2993_ (.Y(_0746_),
    .A(net953),
    .B(net634));
 sg13g2_a22oi_1 _2994_ (.Y(_0747_),
    .B1(net630),
    .B2(net811),
    .A2(net627),
    .A1(net814));
 sg13g2_a21oi_1 _2995_ (.A1(_0746_),
    .A2(_0747_),
    .Y(_0748_),
    .B1(net565));
 sg13g2_a22oi_1 _2996_ (.Y(_0749_),
    .B1(net564),
    .B2(net1285),
    .A2(_1463_),
    .A1(net732));
 sg13g2_nor2_1 _2997_ (.A(_1504_),
    .B(_0749_),
    .Y(_0750_));
 sg13g2_nor4_2 _2998_ (.A(_0742_),
    .B(_0745_),
    .C(_0748_),
    .Y(_0751_),
    .D(_0750_));
 sg13g2_nor2_1 _2999_ (.A(net934),
    .B(_0751_),
    .Y(_0151_));
 sg13g2_a22oi_1 _3000_ (.Y(_0752_),
    .B1(net550),
    .B2(net726),
    .A2(\comm_ic0.i2c0.data_wr[0] ),
    .A1(net574));
 sg13g2_nor2_1 _3001_ (.A(net641),
    .B(net727),
    .Y(_0152_));
 sg13g2_a22oi_1 _3002_ (.Y(_0753_),
    .B1(net550),
    .B2(net383),
    .A2(\comm_ic0.i2c0.data_wr[1] ),
    .A1(net574));
 sg13g2_nor2_1 _3003_ (.A(net641),
    .B(net384),
    .Y(_0153_));
 sg13g2_a22oi_1 _3004_ (.Y(_0754_),
    .B1(net551),
    .B2(net523),
    .A2(\comm_ic0.i2c0.data_wr[2] ),
    .A1(net575));
 sg13g2_nor2_1 _3005_ (.A(net640),
    .B(net524),
    .Y(_0154_));
 sg13g2_a22oi_1 _3006_ (.Y(_0755_),
    .B1(net551),
    .B2(net750),
    .A2(net817),
    .A1(net575));
 sg13g2_nor2_1 _3007_ (.A(net640),
    .B(net818),
    .Y(_0155_));
 sg13g2_a22oi_1 _3008_ (.Y(_0756_),
    .B1(net550),
    .B2(net752),
    .A2(net804),
    .A1(net574));
 sg13g2_nor2_1 _3009_ (.A(net640),
    .B(net805),
    .Y(_0156_));
 sg13g2_a22oi_1 _3010_ (.Y(_0757_),
    .B1(net550),
    .B2(net702),
    .A2(\comm_ic0.i2c0.data_wr[5] ),
    .A1(net574));
 sg13g2_nor2_1 _3011_ (.A(net640),
    .B(net703),
    .Y(_0157_));
 sg13g2_a22oi_1 _3012_ (.Y(_0758_),
    .B1(net550),
    .B2(net806),
    .A2(net855),
    .A1(net574));
 sg13g2_nor2_1 _3013_ (.A(net640),
    .B(net856),
    .Y(_0158_));
 sg13g2_a22oi_1 _3014_ (.Y(_0759_),
    .B1(net550),
    .B2(net481),
    .A2(net819),
    .A1(net574));
 sg13g2_nor2_1 _3015_ (.A(net640),
    .B(net820),
    .Y(_0159_));
 sg13g2_a22oi_1 _3016_ (.Y(_0760_),
    .B1(net550),
    .B2(net368),
    .A2(net1342),
    .A1(net574));
 sg13g2_nor2_1 _3017_ (.A(net640),
    .B(net369),
    .Y(_0160_));
 sg13g2_a22oi_1 _3018_ (.Y(_0761_),
    .B1(net551),
    .B2(net374),
    .A2(\comm_ic0.i2c0.data_wr[9] ),
    .A1(net575));
 sg13g2_nor2_1 _3019_ (.A(net641),
    .B(net375),
    .Y(_0161_));
 sg13g2_a22oi_1 _3020_ (.Y(_0762_),
    .B1(net551),
    .B2(net326),
    .A2(net1344),
    .A1(net575));
 sg13g2_nor2_1 _3021_ (.A(net641),
    .B(net327),
    .Y(_0162_));
 sg13g2_a22oi_1 _3022_ (.Y(_0763_),
    .B1(net550),
    .B2(net486),
    .A2(\comm_ic0.i2c0.data_wr[11] ),
    .A1(net574));
 sg13g2_nor2_1 _3023_ (.A(net640),
    .B(net487),
    .Y(_0163_));
 sg13g2_a22oi_1 _3024_ (.Y(_0764_),
    .B1(net551),
    .B2(net475),
    .A2(net512),
    .A1(net576));
 sg13g2_nor2_1 _3025_ (.A(net644),
    .B(net513),
    .Y(_0164_));
 sg13g2_a22oi_1 _3026_ (.Y(_0765_),
    .B1(net551),
    .B2(net344),
    .A2(net1347),
    .A1(net575));
 sg13g2_nor2_1 _3027_ (.A(net641),
    .B(net345),
    .Y(_0165_));
 sg13g2_a22oi_1 _3028_ (.Y(_0766_),
    .B1(net551),
    .B2(net460),
    .A2(net463),
    .A1(net575));
 sg13g2_nor2_1 _3029_ (.A(net641),
    .B(net464),
    .Y(_0166_));
 sg13g2_a22oi_1 _3030_ (.Y(_0767_),
    .B1(net552),
    .B2(net410),
    .A2(\comm_ic0.i2c0.data_wr[15] ),
    .A1(net576));
 sg13g2_nor2_1 _3031_ (.A(net642),
    .B(net411),
    .Y(_0167_));
 sg13g2_nand2_1 _3032_ (.Y(_0768_),
    .A(net590),
    .B(net539));
 sg13g2_nor2_1 _3033_ (.A(net1327),
    .B(net1071),
    .Y(_0769_));
 sg13g2_or2_2 _3034_ (.X(_0770_),
    .B(net594),
    .A(net1190));
 sg13g2_nor2_1 _3035_ (.A(net1071),
    .B(_0770_),
    .Y(_0771_));
 sg13g2_nor4_2 _3036_ (.A(net1071),
    .B(net590),
    .C(net1045),
    .Y(_0772_),
    .D(_0770_));
 sg13g2_inv_1 _3037_ (.Y(_0773_),
    .A(_0772_));
 sg13g2_a21o_1 _3038_ (.A2(_0771_),
    .A1(_0768_),
    .B1(net538),
    .X(_0774_));
 sg13g2_o21ai_1 _3039_ (.B1(net905),
    .Y(_0775_),
    .A1(net539),
    .A2(_0772_));
 sg13g2_a21oi_1 _3040_ (.A1(net1312),
    .A2(_0772_),
    .Y(_0776_),
    .B1(net656));
 sg13g2_nand3_1 _3041_ (.B(net906),
    .C(_0776_),
    .A(_0774_),
    .Y(_0168_));
 sg13g2_nor4_1 _3042_ (.A(net588),
    .B(net914),
    .C(net590),
    .D(net1045),
    .Y(_0777_));
 sg13g2_inv_1 _3043_ (.Y(_0778_),
    .A(_0777_));
 sg13g2_nor3_1 _3044_ (.A(net1312),
    .B(_0770_),
    .C(_0778_),
    .Y(_0779_));
 sg13g2_a221oi_1 _3045_ (.B2(net588),
    .C1(_0779_),
    .B1(net1080),
    .A1(\comm_ic0.i2c0.addr_wr[0] ),
    .Y(_0780_),
    .A2(net593));
 sg13g2_nand2_1 _3046_ (.Y(_0781_),
    .A(net539),
    .B(_0770_));
 sg13g2_o21ai_1 _3047_ (.B1(_1565_),
    .Y(_0782_),
    .A1(net595),
    .A2(net1045));
 sg13g2_nand4_1 _3048_ (.B(_0780_),
    .C(_0781_),
    .A(_0768_),
    .Y(_0783_),
    .D(_0782_));
 sg13g2_nor2b_2 _3049_ (.A(net1122),
    .B_N(net1290),
    .Y(_0784_));
 sg13g2_nand2_1 _3050_ (.Y(_0785_),
    .A(net804),
    .B(net562));
 sg13g2_nor2b_2 _3051_ (.A(net1290),
    .B_N(net1122),
    .Y(_0786_));
 sg13g2_nand2_1 _3052_ (.Y(_0787_),
    .A(net819),
    .B(_0673_));
 sg13g2_nand2_1 _3053_ (.Y(_0788_),
    .A(net512),
    .B(net562));
 sg13g2_nand2_1 _3054_ (.Y(_0789_),
    .A(\comm_ic0.i2c0.data_wr[15] ),
    .B(_0673_));
 sg13g2_nand2_1 _3055_ (.Y(_0790_),
    .A(\comm_ic0.i2c0.data_wr[0] ),
    .B(net562));
 sg13g2_a22oi_1 _3056_ (.Y(_0791_),
    .B1(_0673_),
    .B2(\comm_ic0.i2c0.data_wr[11] ),
    .A2(net562),
    .A1(\comm_ic0.i2c0.data_wr[8] ));
 sg13g2_a221oi_1 _3057_ (.B2(\comm_ic0.i2c0.data_wr[10] ),
    .C1(net605),
    .B1(_0786_),
    .A1(\comm_ic0.i2c0.data_wr[9] ),
    .Y(_0792_),
    .A2(_0784_));
 sg13g2_nand2_1 _3058_ (.Y(_0793_),
    .A(_0791_),
    .B(_0792_));
 sg13g2_a22oi_1 _3059_ (.Y(_0794_),
    .B1(_0786_),
    .B2(net463),
    .A2(_0784_),
    .A1(\comm_ic0.i2c0.data_wr[13] ));
 sg13g2_nand4_1 _3060_ (.B(_0788_),
    .C(_0789_),
    .A(net605),
    .Y(_0795_),
    .D(_0794_));
 sg13g2_a21oi_1 _3061_ (.A1(_0793_),
    .A2(_0795_),
    .Y(_0796_),
    .B1(_1411_));
 sg13g2_a22oi_1 _3062_ (.Y(_0797_),
    .B1(_0786_),
    .B2(net855),
    .A2(_0784_),
    .A1(\comm_ic0.i2c0.data_wr[5] ));
 sg13g2_nand4_1 _3063_ (.B(_0785_),
    .C(_0787_),
    .A(net605),
    .Y(_0798_),
    .D(_0797_));
 sg13g2_a21oi_1 _3064_ (.A1(\comm_ic0.i2c0.data_wr[1] ),
    .A2(_0784_),
    .Y(_0799_),
    .B1(net605));
 sg13g2_a22oi_1 _3065_ (.Y(_0800_),
    .B1(_0786_),
    .B2(\comm_ic0.i2c0.data_wr[2] ),
    .A2(_0673_),
    .A1(net817));
 sg13g2_nand3_1 _3066_ (.B(_0799_),
    .C(_0800_),
    .A(_0790_),
    .Y(_0801_));
 sg13g2_a21oi_2 _3067_ (.B1(net1038),
    .Y(_0802_),
    .A2(_0801_),
    .A1(_0798_));
 sg13g2_nor3_2 _3068_ (.A(net1318),
    .B(_0796_),
    .C(_0802_),
    .Y(_0803_));
 sg13g2_nand2b_1 _3069_ (.Y(_0804_),
    .B(\comm_ic0.i2c0.addr_ind[0] ),
    .A_N(\comm_ic0.i2c0.addr_ind[1] ));
 sg13g2_nor2_1 _3070_ (.A(\comm_ic0.i2c0.addr_wr[1] ),
    .B(_0804_),
    .Y(_0805_));
 sg13g2_nor3_1 _3071_ (.A(\comm_ic0.i2c0.addr_wr[0] ),
    .B(\comm_ic0.i2c0.addr_ind[1] ),
    .C(\comm_ic0.i2c0.addr_ind[0] ),
    .Y(_0806_));
 sg13g2_nor2b_1 _3072_ (.A(\comm_ic0.i2c0.addr_ind[0] ),
    .B_N(\comm_ic0.i2c0.addr_ind[1] ),
    .Y(_0807_));
 sg13g2_nor2b_1 _3073_ (.A(\comm_ic0.i2c0.addr_wr[2] ),
    .B_N(_0807_),
    .Y(_0808_));
 sg13g2_nor4_1 _3074_ (.A(net971),
    .B(_0805_),
    .C(_0806_),
    .D(_0808_),
    .Y(_0809_));
 sg13g2_o21ai_1 _3075_ (.B1(_0809_),
    .Y(_0810_),
    .A1(net705),
    .A2(_0690_));
 sg13g2_o21ai_1 _3076_ (.B1(net971),
    .Y(_0811_),
    .A1(net504),
    .A2(_0804_));
 sg13g2_nor2_1 _3077_ (.A(net426),
    .B(_0690_),
    .Y(_0812_));
 sg13g2_nor3_1 _3078_ (.A(\comm_ic0.i2c0.addr_wr[4] ),
    .B(\comm_ic0.i2c0.addr_ind[1] ),
    .C(net1314),
    .Y(_0813_));
 sg13g2_nor2b_1 _3079_ (.A(\comm_ic0.i2c0.addr_wr[6] ),
    .B_N(_0807_),
    .Y(_0814_));
 sg13g2_or4_1 _3080_ (.A(_0811_),
    .B(_0812_),
    .C(_0813_),
    .D(_0814_),
    .X(_0815_));
 sg13g2_a22oi_1 _3081_ (.Y(_0816_),
    .B1(_0810_),
    .B2(_0815_),
    .A2(_1429_),
    .A1(_1428_));
 sg13g2_nor4_1 _3082_ (.A(net595),
    .B(net589),
    .C(net1045),
    .D(_0770_),
    .Y(_0817_));
 sg13g2_nor3_1 _3083_ (.A(_0803_),
    .B(_0816_),
    .C(_0817_),
    .Y(_0818_));
 sg13g2_a21oi_1 _3084_ (.A1(net883),
    .A2(_0783_),
    .Y(_0819_),
    .B1(net656));
 sg13g2_o21ai_1 _3085_ (.B1(net884),
    .Y(_0169_),
    .A1(_0783_),
    .A2(net1319));
 sg13g2_nand2b_1 _3086_ (.Y(_0820_),
    .B(net593),
    .A_N(\comm_ic0.i2c0.addr_wr[0] ));
 sg13g2_nand4_1 _3087_ (.B(_0769_),
    .C(_0777_),
    .A(_1593_),
    .Y(_0821_),
    .D(_0820_));
 sg13g2_a21oi_1 _3088_ (.A1(net593),
    .A2(net538),
    .Y(_0822_),
    .B1(_0821_));
 sg13g2_a21o_2 _3089_ (.A2(net538),
    .A1(net593),
    .B1(_0821_),
    .X(_0823_));
 sg13g2_nand2_1 _3090_ (.Y(_0824_),
    .A(_1577_),
    .B(net529));
 sg13g2_nor3_2 _3091_ (.A(net573),
    .B(_1431_),
    .C(_0823_),
    .Y(_0825_));
 sg13g2_a22oi_1 _3092_ (.Y(_0826_),
    .B1(_0825_),
    .B2(_1575_),
    .A2(_0824_),
    .A1(net1057));
 sg13g2_nor2_1 _3093_ (.A(net653),
    .B(net1058),
    .Y(_0170_));
 sg13g2_nor2b_1 _3094_ (.A(net603),
    .B_N(_0784_),
    .Y(_0827_));
 sg13g2_inv_1 _3095_ (.Y(_0828_),
    .A(_0827_));
 sg13g2_o21ai_1 _3096_ (.B1(net593),
    .Y(_0829_),
    .A1(net600),
    .A2(_0828_));
 sg13g2_nand2_1 _3097_ (.Y(_0830_),
    .A(_0822_),
    .B(_0829_));
 sg13g2_and3_1 _3098_ (.X(_0831_),
    .A(net592),
    .B(_0680_),
    .C(net530));
 sg13g2_and4_2 _3099_ (.A(net592),
    .B(_1576_),
    .C(_0680_),
    .D(net529),
    .X(_0832_));
 sg13g2_nor2_1 _3100_ (.A(_1431_),
    .B(_0828_),
    .Y(_0833_));
 sg13g2_a22oi_1 _3101_ (.Y(_0834_),
    .B1(_0832_),
    .B2(_0833_),
    .A2(_0830_),
    .A1(net841));
 sg13g2_nor2_1 _3102_ (.A(net653),
    .B(net842),
    .Y(_0171_));
 sg13g2_nor2b_1 _3103_ (.A(net603),
    .B_N(_0786_),
    .Y(_0835_));
 sg13g2_nand2b_1 _3104_ (.Y(_0836_),
    .B(_0786_),
    .A_N(net604));
 sg13g2_o21ai_1 _3105_ (.B1(net592),
    .Y(_0837_),
    .A1(net600),
    .A2(_0836_));
 sg13g2_nand2_1 _3106_ (.Y(_0838_),
    .A(net530),
    .B(_0837_));
 sg13g2_nor3_1 _3107_ (.A(_1431_),
    .B(_1575_),
    .C(_0836_),
    .Y(_0839_));
 sg13g2_a22oi_1 _3108_ (.Y(_0840_),
    .B1(_0839_),
    .B2(_0831_),
    .A2(_0838_),
    .A1(net798));
 sg13g2_nor2_1 _3109_ (.A(net652),
    .B(net799),
    .Y(_0172_));
 sg13g2_nor2b_1 _3110_ (.A(net604),
    .B_N(_0673_),
    .Y(_0841_));
 sg13g2_inv_1 _3111_ (.Y(_0842_),
    .A(_0841_));
 sg13g2_o21ai_1 _3112_ (.B1(net593),
    .Y(_0843_),
    .A1(net600),
    .A2(_0842_));
 sg13g2_nand2_1 _3113_ (.Y(_0844_),
    .A(_0822_),
    .B(_0843_));
 sg13g2_nor2_1 _3114_ (.A(_1431_),
    .B(_0842_),
    .Y(_0845_));
 sg13g2_a22oi_1 _3115_ (.Y(_0846_),
    .B1(_0845_),
    .B2(_0832_),
    .A2(_0844_),
    .A1(net953));
 sg13g2_nor2_1 _3116_ (.A(net653),
    .B(net954),
    .Y(_0173_));
 sg13g2_and3_1 _3117_ (.X(_0847_),
    .A(_1411_),
    .B(net604),
    .C(net562));
 sg13g2_o21ai_1 _3118_ (.B1(net530),
    .Y(_0848_),
    .A1(net573),
    .A2(_0847_));
 sg13g2_a22oi_1 _3119_ (.Y(_0849_),
    .B1(_0848_),
    .B2(net377),
    .A2(_0847_),
    .A1(_0825_));
 sg13g2_nor2_1 _3120_ (.A(net643),
    .B(net378),
    .Y(_0174_));
 sg13g2_nand2_1 _3121_ (.Y(_0850_),
    .A(net603),
    .B(_0784_));
 sg13g2_o21ai_1 _3122_ (.B1(net594),
    .Y(_0851_),
    .A1(net601),
    .A2(_0850_));
 sg13g2_nand2_1 _3123_ (.Y(_0852_),
    .A(net529),
    .B(_0851_));
 sg13g2_nor2_1 _3124_ (.A(_1431_),
    .B(_0850_),
    .Y(_0853_));
 sg13g2_a22oi_1 _3125_ (.Y(_0854_),
    .B1(_0853_),
    .B2(_0832_),
    .A2(_0852_),
    .A1(net526));
 sg13g2_nor2_1 _3126_ (.A(net654),
    .B(net697),
    .Y(_0175_));
 sg13g2_nand2_1 _3127_ (.Y(_0855_),
    .A(net603),
    .B(_0786_));
 sg13g2_o21ai_1 _3128_ (.B1(net592),
    .Y(_0856_),
    .A1(net600),
    .A2(_0855_));
 sg13g2_nand2_1 _3129_ (.Y(_0857_),
    .A(net530),
    .B(_0856_));
 sg13g2_nor3_1 _3130_ (.A(_1431_),
    .B(_1575_),
    .C(_0855_),
    .Y(_0858_));
 sg13g2_a22oi_1 _3131_ (.Y(_0859_),
    .B1(_0858_),
    .B2(_0831_),
    .A2(_0857_),
    .A1(net741));
 sg13g2_nor2_1 _3132_ (.A(net652),
    .B(net742),
    .Y(_0176_));
 sg13g2_nand2_1 _3133_ (.Y(_0860_),
    .A(net604),
    .B(_0673_));
 sg13g2_o21ai_1 _3134_ (.B1(net592),
    .Y(_0861_),
    .A1(net601),
    .A2(_0860_));
 sg13g2_nand2_1 _3135_ (.Y(_0862_),
    .A(net529),
    .B(_0861_));
 sg13g2_nor2_1 _3136_ (.A(_1431_),
    .B(_0860_),
    .Y(_0863_));
 sg13g2_a22oi_1 _3137_ (.Y(_0864_),
    .B1(_0863_),
    .B2(_0832_),
    .A2(_0862_),
    .A1(net814));
 sg13g2_nor2_1 _3138_ (.A(net653),
    .B(net815),
    .Y(_0177_));
 sg13g2_o21ai_1 _3139_ (.B1(net530),
    .Y(_0865_),
    .A1(net573),
    .A2(_0681_));
 sg13g2_a22oi_1 _3140_ (.Y(_0866_),
    .B1(_0865_),
    .B2(net365),
    .A2(_0825_),
    .A1(_0681_));
 sg13g2_nor2_1 _3141_ (.A(net643),
    .B(net366),
    .Y(_0178_));
 sg13g2_a21oi_1 _3142_ (.A1(net601),
    .A2(_0827_),
    .Y(_0867_),
    .B1(_1430_));
 sg13g2_o21ai_1 _3143_ (.B1(net764),
    .Y(_0868_),
    .A1(_0823_),
    .A2(_0867_));
 sg13g2_nand3_1 _3144_ (.B(net529),
    .C(_0833_),
    .A(_0682_),
    .Y(_0869_));
 sg13g2_a21oi_1 _3145_ (.A1(net765),
    .A2(_0869_),
    .Y(_0179_),
    .B1(net654));
 sg13g2_a21oi_1 _3146_ (.A1(net600),
    .A2(_0835_),
    .Y(_0870_),
    .B1(net573));
 sg13g2_o21ai_1 _3147_ (.B1(net786),
    .Y(_0871_),
    .A1(_0823_),
    .A2(_0870_));
 sg13g2_nand3_1 _3148_ (.B(net530),
    .C(_0839_),
    .A(_0682_),
    .Y(_0872_));
 sg13g2_a21oi_1 _3149_ (.A1(net787),
    .A2(_0872_),
    .Y(_0180_),
    .B1(net653));
 sg13g2_a21oi_1 _3150_ (.A1(net601),
    .A2(_0841_),
    .Y(_0873_),
    .B1(net573));
 sg13g2_o21ai_1 _3151_ (.B1(net811),
    .Y(_0874_),
    .A1(_0823_),
    .A2(_0873_));
 sg13g2_nand3_1 _3152_ (.B(net529),
    .C(_0845_),
    .A(_0682_),
    .Y(_0875_));
 sg13g2_a21oi_1 _3153_ (.A1(net812),
    .A2(_0875_),
    .Y(_0181_),
    .B1(net654));
 sg13g2_nand3_1 _3154_ (.B(net604),
    .C(net562),
    .A(net602),
    .Y(_0876_));
 sg13g2_and2_1 _3155_ (.A(net591),
    .B(_0876_),
    .X(_0877_));
 sg13g2_o21ai_1 _3156_ (.B1(net714),
    .Y(_0878_),
    .A1(_0823_),
    .A2(_0877_));
 sg13g2_nand4_1 _3157_ (.B(net603),
    .C(net562),
    .A(net602),
    .Y(_0879_),
    .D(_0825_));
 sg13g2_a21oi_1 _3158_ (.A1(net715),
    .A2(_0879_),
    .Y(_0182_),
    .B1(net643));
 sg13g2_nand3_1 _3159_ (.B(net603),
    .C(_0784_),
    .A(net600),
    .Y(_0880_));
 sg13g2_and2_1 _3160_ (.A(net592),
    .B(_0880_),
    .X(_0881_));
 sg13g2_o21ai_1 _3161_ (.B1(net735),
    .Y(_0882_),
    .A1(_0823_),
    .A2(_0881_));
 sg13g2_nand3_1 _3162_ (.B(net529),
    .C(_0853_),
    .A(_0682_),
    .Y(_0883_));
 sg13g2_a21oi_1 _3163_ (.A1(net736),
    .A2(_0883_),
    .Y(_0183_),
    .B1(net653));
 sg13g2_nand3_1 _3164_ (.B(net603),
    .C(_0786_),
    .A(net602),
    .Y(_0884_));
 sg13g2_and2_1 _3165_ (.A(net591),
    .B(_0884_),
    .X(_0885_));
 sg13g2_o21ai_1 _3166_ (.B1(net723),
    .Y(_0886_),
    .A1(_0823_),
    .A2(_0885_));
 sg13g2_nand3_1 _3167_ (.B(net530),
    .C(_0858_),
    .A(_0682_),
    .Y(_0887_));
 sg13g2_a21oi_1 _3168_ (.A1(net724),
    .A2(_0887_),
    .Y(_0184_),
    .B1(net653));
 sg13g2_nand3_1 _3169_ (.B(net603),
    .C(_0673_),
    .A(net600),
    .Y(_0888_));
 sg13g2_and2_1 _3170_ (.A(net591),
    .B(_0888_),
    .X(_0889_));
 sg13g2_o21ai_1 _3171_ (.B1(net732),
    .Y(_0890_),
    .A1(_0823_),
    .A2(_0889_));
 sg13g2_nand3_1 _3172_ (.B(net529),
    .C(_0863_),
    .A(_0682_),
    .Y(_0891_));
 sg13g2_a21oi_1 _3173_ (.A1(net733),
    .A2(_0891_),
    .Y(_0185_),
    .B1(net653));
 sg13g2_a21oi_1 _3174_ (.A1(net588),
    .A2(net539),
    .Y(_0892_),
    .B1(net578));
 sg13g2_nor2_1 _3175_ (.A(net1004),
    .B(_0892_),
    .Y(_0893_));
 sg13g2_nand3b_1 _3176_ (.B(_1593_),
    .C(net690),
    .Y(_0894_),
    .A_N(net588));
 sg13g2_a21oi_1 _3177_ (.A1(net832),
    .A2(_0894_),
    .Y(_0186_),
    .B1(net1005));
 sg13g2_nand2_1 _3178_ (.Y(_0895_),
    .A(net577),
    .B(_1410_));
 sg13g2_and4_1 _3179_ (.A(_1564_),
    .B(_1578_),
    .C(_1593_),
    .D(_0895_),
    .X(_0896_));
 sg13g2_o21ai_1 _3180_ (.B1(net689),
    .Y(_0897_),
    .A1(net920),
    .A2(_0896_));
 sg13g2_a21oi_1 _3181_ (.A1(_1410_),
    .A2(net553),
    .Y(_0187_),
    .B1(net921));
 sg13g2_a22oi_1 _3182_ (.Y(_0898_),
    .B1(_0771_),
    .B2(_1408_),
    .A2(net593),
    .A1(\comm_ic0.i2c0.addr_wr[0] ));
 sg13g2_nand3_1 _3183_ (.B(_0781_),
    .C(_0898_),
    .A(_1584_),
    .Y(_0899_));
 sg13g2_a21oi_1 _3184_ (.A1(net1278),
    .A2(_0899_),
    .Y(_0900_),
    .B1(net655));
 sg13g2_o21ai_1 _3185_ (.B1(net1279),
    .Y(_0188_),
    .A1(net315),
    .A2(_0899_));
 sg13g2_a22oi_1 _3186_ (.Y(_0901_),
    .B1(net552),
    .B2(net1054),
    .A2(\comm_ic0.i2c0.clk_cnt_reg[0] ),
    .A1(net576));
 sg13g2_nor2_1 _3187_ (.A(net642),
    .B(net1055),
    .Y(_0189_));
 sg13g2_a22oi_1 _3188_ (.Y(_0902_),
    .B1(net552),
    .B2(net1062),
    .A2(\comm_ic0.i2c0.clk_cnt_reg[1] ),
    .A1(net576));
 sg13g2_nor2_1 _3189_ (.A(net642),
    .B(net1063),
    .Y(_0190_));
 sg13g2_a22oi_1 _3190_ (.Y(_0903_),
    .B1(net552),
    .B2(net857),
    .A2(\comm_ic0.i2c0.clk_cnt_reg[2] ),
    .A1(net576));
 sg13g2_nor2_1 _3191_ (.A(net642),
    .B(net858),
    .Y(_0191_));
 sg13g2_a22oi_1 _3192_ (.Y(_0904_),
    .B1(net552),
    .B2(net1025),
    .A2(\comm_ic0.i2c0.clk_cnt_reg[3] ),
    .A1(net576));
 sg13g2_nor2_1 _3193_ (.A(net642),
    .B(net1026),
    .Y(_0192_));
 sg13g2_a22oi_1 _3194_ (.Y(_0905_),
    .B1(net554),
    .B2(net847),
    .A2(\comm_ic0.i2c0.clk_cnt_reg[4] ),
    .A1(net578));
 sg13g2_nor2_1 _3195_ (.A(net652),
    .B(net848),
    .Y(_0193_));
 sg13g2_a22oi_1 _3196_ (.Y(_0906_),
    .B1(net554),
    .B2(net1028),
    .A2(\comm_ic0.i2c0.clk_cnt_reg[5] ),
    .A1(net578));
 sg13g2_nor2_1 _3197_ (.A(net654),
    .B(net1029),
    .Y(_0194_));
 sg13g2_a22oi_1 _3198_ (.Y(_0907_),
    .B1(net554),
    .B2(net392),
    .A2(\comm_ic0.i2c0.clk_cnt_reg[6] ),
    .A1(net578));
 sg13g2_nor2_1 _3199_ (.A(net654),
    .B(net393),
    .Y(_0195_));
 sg13g2_a22oi_1 _3200_ (.Y(_0908_),
    .B1(net554),
    .B2(net1019),
    .A2(\comm_ic0.i2c0.clk_cnt_reg[7] ),
    .A1(net578));
 sg13g2_nor2_1 _3201_ (.A(net652),
    .B(net1020),
    .Y(_0196_));
 sg13g2_a22oi_1 _3202_ (.Y(_0909_),
    .B1(net554),
    .B2(net452),
    .A2(\comm_ic0.i2c0.addr_wr[0] ),
    .A1(net578));
 sg13g2_nor2_1 _3203_ (.A(net652),
    .B(net453),
    .Y(_0197_));
 sg13g2_a22oi_1 _3204_ (.Y(_0910_),
    .B1(net553),
    .B2(net423),
    .A2(\comm_ic0.i2c0.addr_wr[1] ),
    .A1(net577));
 sg13g2_nor2_1 _3205_ (.A(net655),
    .B(net424),
    .Y(_0198_));
 sg13g2_a22oi_1 _3206_ (.Y(_0911_),
    .B1(net553),
    .B2(net332),
    .A2(net1345),
    .A1(net577));
 sg13g2_nor2_1 _3207_ (.A(net655),
    .B(net333),
    .Y(_0199_));
 sg13g2_a22oi_1 _3208_ (.Y(_0912_),
    .B1(net553),
    .B2(net429),
    .A2(net705),
    .A1(net577));
 sg13g2_nor2_1 _3209_ (.A(net655),
    .B(net706),
    .Y(_0200_));
 sg13g2_a22oi_1 _3210_ (.Y(_0913_),
    .B1(net553),
    .B2(net413),
    .A2(\comm_ic0.i2c0.addr_wr[4] ),
    .A1(net577));
 sg13g2_nor2_1 _3211_ (.A(net655),
    .B(net414),
    .Y(_0201_));
 sg13g2_a22oi_1 _3212_ (.Y(_0914_),
    .B1(net553),
    .B2(net498),
    .A2(net504),
    .A1(net577));
 sg13g2_nor2_1 _3213_ (.A(net656),
    .B(net505),
    .Y(_0202_));
 sg13g2_a22oi_1 _3214_ (.Y(_0915_),
    .B1(net553),
    .B2(net708),
    .A2(\comm_ic0.i2c0.addr_wr[6] ),
    .A1(net577));
 sg13g2_nor2_1 _3215_ (.A(net655),
    .B(net709),
    .Y(_0203_));
 sg13g2_a22oi_1 _3216_ (.Y(_0916_),
    .B1(net553),
    .B2(net389),
    .A2(net577),
    .A1(net426));
 sg13g2_nor2_1 _3217_ (.A(net656),
    .B(net427),
    .Y(_0204_));
 sg13g2_nor2_1 _3218_ (.A(net1106),
    .B(net1134),
    .Y(_0917_));
 sg13g2_or2_1 _3219_ (.X(_0918_),
    .B(net1134),
    .A(net1193));
 sg13g2_o21ai_1 _3220_ (.B1(_1594_),
    .Y(_0919_),
    .A1(net1106),
    .A2(_0918_));
 sg13g2_nor2_1 _3221_ (.A(_0026_),
    .B(_1450_),
    .Y(_0920_));
 sg13g2_o21ai_1 _3222_ (.B1(net757),
    .Y(_0921_),
    .A1(_0919_),
    .A2(_0920_));
 sg13g2_o21ai_1 _3223_ (.B1(net681),
    .Y(_0922_),
    .A1(_1407_),
    .A2(_0919_));
 sg13g2_nand2b_1 _3224_ (.Y(_0205_),
    .B(net758),
    .A_N(_0922_));
 sg13g2_or2_2 _3225_ (.X(_0923_),
    .B(net638),
    .A(net1193));
 sg13g2_nor2_1 _3226_ (.A(net1134),
    .B(_0923_),
    .Y(_0924_));
 sg13g2_a21oi_1 _3227_ (.A1(net638),
    .A2(_1457_),
    .Y(_0925_),
    .B1(_0924_));
 sg13g2_a22oi_1 _3228_ (.Y(_0926_),
    .B1(net638),
    .B2(_1406_),
    .A2(net1134),
    .A1(net699));
 sg13g2_o21ai_1 _3229_ (.B1(net680),
    .Y(_0927_),
    .A1(net1031),
    .A2(_0925_));
 sg13g2_a21oi_1 _3230_ (.A1(_0925_),
    .A2(_0926_),
    .Y(_0206_),
    .B1(net1032));
 sg13g2_nor2_1 _3231_ (.A(_1400_),
    .B(_1450_),
    .Y(_0928_));
 sg13g2_nor2_1 _3232_ (.A(\comm_ic0.spi0.CPHA ),
    .B(_1456_),
    .Y(_0929_));
 sg13g2_o21ai_1 _3233_ (.B1(net638),
    .Y(_0930_),
    .A1(_0928_),
    .A2(_0929_));
 sg13g2_nor2_1 _3234_ (.A(_0920_),
    .B(_0924_),
    .Y(_0931_));
 sg13g2_nand2_1 _3235_ (.Y(_0932_),
    .A(_0930_),
    .B(_0931_));
 sg13g2_and2_2 _3236_ (.A(net586),
    .B(net587),
    .X(_0933_));
 sg13g2_nand2_1 _3237_ (.Y(_0934_),
    .A(net586),
    .B(net1209));
 sg13g2_nor2b_2 _3238_ (.A(net586),
    .B_N(net587),
    .Y(_0935_));
 sg13g2_nor2b_2 _3239_ (.A(net587),
    .B_N(net586),
    .Y(_0936_));
 sg13g2_a22oi_1 _3240_ (.Y(_0937_),
    .B1(_0936_),
    .B2(net329),
    .A2(_0933_),
    .A1(net492));
 sg13g2_a221oi_1 _3241_ (.B2(net317),
    .C1(net585),
    .B1(_0935_),
    .A1(net435),
    .Y(_0938_),
    .A2(net561));
 sg13g2_nand2_1 _3242_ (.Y(_0939_),
    .A(_0937_),
    .B(_0938_));
 sg13g2_a21oi_1 _3243_ (.A1(net362),
    .A2(_0933_),
    .Y(_0940_),
    .B1(_1401_));
 sg13g2_nand2_1 _3244_ (.Y(_0941_),
    .A(net323),
    .B(net561));
 sg13g2_a22oi_1 _3245_ (.Y(_0942_),
    .B1(_0936_),
    .B2(net371),
    .A2(_0935_),
    .A1(net359));
 sg13g2_nand3_1 _3246_ (.B(_0941_),
    .C(_0942_),
    .A(_0940_),
    .Y(_0943_));
 sg13g2_nand3_1 _3247_ (.B(_0939_),
    .C(_0943_),
    .A(\comm_ic0.spi0.data_ind[3] ),
    .Y(_0944_));
 sg13g2_a21oi_1 _3248_ (.A1(net407),
    .A2(_0933_),
    .Y(_0945_),
    .B1(net585));
 sg13g2_nand2_1 _3249_ (.Y(_0946_),
    .A(net416),
    .B(_0935_));
 sg13g2_a22oi_1 _3250_ (.Y(_0947_),
    .B1(_0936_),
    .B2(net335),
    .A2(net561),
    .A1(net341));
 sg13g2_nand3_1 _3251_ (.B(_0946_),
    .C(_0947_),
    .A(_0945_),
    .Y(_0948_));
 sg13g2_a22oi_1 _3252_ (.Y(_0949_),
    .B1(_0935_),
    .B2(net472),
    .A2(net561),
    .A1(net489));
 sg13g2_a221oi_1 _3253_ (.B2(\comm_ic0.spi0.data_wr[6] ),
    .C1(_1401_),
    .B1(_0936_),
    .A1(net501),
    .Y(_0950_),
    .A2(_0933_));
 sg13g2_a21oi_1 _3254_ (.A1(_0949_),
    .A2(_0950_),
    .Y(_0951_),
    .B1(\comm_ic0.spi0.data_ind[3] ));
 sg13g2_nand2_1 _3255_ (.Y(_0952_),
    .A(_0948_),
    .B(_0951_));
 sg13g2_a21oi_1 _3256_ (.A1(_1407_),
    .A2(\comm_ic0.spi0.curr_st[1] ),
    .Y(_0953_),
    .B1(net638));
 sg13g2_nor3_1 _3257_ (.A(_0920_),
    .B(_0928_),
    .C(_0953_),
    .Y(_0954_));
 sg13g2_a22oi_1 _3258_ (.Y(_0955_),
    .B1(_0944_),
    .B2(_0952_),
    .A2(_0929_),
    .A1(_0026_));
 sg13g2_a22oi_1 _3259_ (.Y(_0956_),
    .B1(_0954_),
    .B2(_0955_),
    .A2(_0932_),
    .A1(net777));
 sg13g2_nor2_1 _3260_ (.A(net645),
    .B(net778),
    .Y(_0207_));
 sg13g2_nand2_2 _3261_ (.Y(_0957_),
    .A(_1459_),
    .B(_0917_));
 sg13g2_nor2_2 _3262_ (.A(_1434_),
    .B(net542),
    .Y(_0958_));
 sg13g2_nand3_1 _3263_ (.B(net1194),
    .C(_0917_),
    .A(net639),
    .Y(_0959_));
 sg13g2_xnor2_1 _3264_ (.Y(_0960_),
    .A(net582),
    .B(_1601_));
 sg13g2_xnor2_1 _3265_ (.Y(_0961_),
    .A(_1437_),
    .B(_1601_));
 sg13g2_nor2_1 _3266_ (.A(net533),
    .B(_0961_),
    .Y(_0962_));
 sg13g2_and4_1 _3267_ (.A(_0042_),
    .B(net531),
    .C(_1603_),
    .D(_0960_),
    .X(_0963_));
 sg13g2_nand4_1 _3268_ (.B(_1598_),
    .C(_1603_),
    .A(net2),
    .Y(_0964_),
    .D(_0960_));
 sg13g2_o21ai_1 _3269_ (.B1(_0964_),
    .Y(_0965_),
    .A1(net1346),
    .A2(_0963_));
 sg13g2_a22oi_1 _3270_ (.Y(_0966_),
    .B1(_0958_),
    .B2(_0965_),
    .A2(net542),
    .A1(net789));
 sg13g2_nor2_1 _3271_ (.A(net647),
    .B(net790),
    .Y(_0208_));
 sg13g2_nand2_1 _3272_ (.Y(_0967_),
    .A(net1022),
    .B(net541));
 sg13g2_and2_1 _3273_ (.A(_1401_),
    .B(_0935_),
    .X(_0968_));
 sg13g2_nand2_1 _3274_ (.Y(_0969_),
    .A(net582),
    .B(_0968_));
 sg13g2_o21ai_1 _3275_ (.B1(_0969_),
    .Y(_0970_),
    .A1(net1022),
    .A2(net535));
 sg13g2_nor2_2 _3276_ (.A(_1599_),
    .B(_0933_),
    .Y(_0971_));
 sg13g2_nand2_2 _3277_ (.Y(_0972_),
    .A(net2),
    .B(_1604_));
 sg13g2_nor4_2 _3278_ (.A(_0042_),
    .B(net561),
    .C(_0933_),
    .Y(_0973_),
    .D(_0972_));
 sg13g2_and2_1 _3279_ (.A(_1401_),
    .B(_0973_),
    .X(_0974_));
 sg13g2_a21oi_1 _3280_ (.A1(_0961_),
    .A2(_0974_),
    .Y(_0975_),
    .B1(net534));
 sg13g2_a22oi_1 _3281_ (.Y(_0976_),
    .B1(_0970_),
    .B2(_0975_),
    .A2(net536),
    .A1(net1297));
 sg13g2_nand2_1 _3282_ (.Y(_0977_),
    .A(_1595_),
    .B(_0974_));
 sg13g2_nor2_1 _3283_ (.A(_0960_),
    .B(_0977_),
    .Y(_0978_));
 sg13g2_o21ai_1 _3284_ (.B1(_0958_),
    .Y(_0979_),
    .A1(_0976_),
    .A2(_0978_));
 sg13g2_a21oi_1 _3285_ (.A1(net1023),
    .A2(net1298),
    .Y(_0209_),
    .B1(net647));
 sg13g2_nand2_1 _3286_ (.Y(_0980_),
    .A(net895),
    .B(net542));
 sg13g2_nand2_2 _3287_ (.Y(_0981_),
    .A(net531),
    .B(_0972_));
 sg13g2_and2_1 _3288_ (.A(_1401_),
    .B(_0936_),
    .X(_0982_));
 sg13g2_nand2_1 _3289_ (.Y(_0983_),
    .A(net1309),
    .B(net533));
 sg13g2_nand4_1 _3290_ (.B(_0981_),
    .C(_0982_),
    .A(net582),
    .Y(_0984_),
    .D(_0983_));
 sg13g2_a22oi_1 _3291_ (.Y(_0985_),
    .B1(_0982_),
    .B2(net582),
    .A2(net537),
    .A1(net1309));
 sg13g2_o21ai_1 _3292_ (.B1(_0985_),
    .Y(_0986_),
    .A1(net895),
    .A2(net535));
 sg13g2_a21o_1 _3293_ (.A2(_0986_),
    .A1(net1310),
    .B1(net540),
    .X(_0987_));
 sg13g2_a21oi_1 _3294_ (.A1(net896),
    .A2(net1311),
    .Y(_0210_),
    .B1(net643));
 sg13g2_nand2_1 _3295_ (.Y(_0988_),
    .A(net886),
    .B(_0957_));
 sg13g2_xnor2_1 _3296_ (.Y(_0989_),
    .A(net583),
    .B(net561));
 sg13g2_xnor2_1 _3297_ (.Y(_0990_),
    .A(_1401_),
    .B(net561));
 sg13g2_nor4_1 _3298_ (.A(_0042_),
    .B(_0971_),
    .C(_0972_),
    .D(_0990_),
    .Y(_0991_));
 sg13g2_and2_1 _3299_ (.A(_0961_),
    .B(_0991_),
    .X(_0992_));
 sg13g2_nor2_1 _3300_ (.A(net886),
    .B(net536),
    .Y(_0993_));
 sg13g2_nor3_1 _3301_ (.A(net583),
    .B(net571),
    .C(_0934_),
    .Y(_0994_));
 sg13g2_a221oi_1 _3302_ (.B2(_0994_),
    .C1(_0993_),
    .B1(_1598_),
    .A1(net1283),
    .Y(_0995_),
    .A2(_1596_));
 sg13g2_a21oi_1 _3303_ (.A1(net1283),
    .A2(net533),
    .Y(_0996_),
    .B1(net540));
 sg13g2_o21ai_1 _3304_ (.B1(_0996_),
    .Y(_0997_),
    .A1(_0992_),
    .A2(_0995_));
 sg13g2_a21oi_1 _3305_ (.A1(net887),
    .A2(net1284),
    .Y(_0211_),
    .B1(net647));
 sg13g2_nand2_1 _3306_ (.Y(_0998_),
    .A(net495),
    .B(_0957_));
 sg13g2_nand2_1 _3307_ (.Y(_0999_),
    .A(net1315),
    .B(_1604_));
 sg13g2_nor2_1 _3308_ (.A(_1603_),
    .B(_0971_),
    .Y(_1000_));
 sg13g2_nand2_1 _3309_ (.Y(_1001_),
    .A(_0042_),
    .B(_1000_));
 sg13g2_nor2_1 _3310_ (.A(_0990_),
    .B(_1001_),
    .Y(_1002_));
 sg13g2_nor2_1 _3311_ (.A(net533),
    .B(_0960_),
    .Y(_1003_));
 sg13g2_a21oi_1 _3312_ (.A1(_1002_),
    .A2(_1003_),
    .Y(_1004_),
    .B1(net1288));
 sg13g2_nand4_1 _3313_ (.B(net2),
    .C(net531),
    .A(net583),
    .Y(_1005_),
    .D(net561));
 sg13g2_nor2_1 _3314_ (.A(_0960_),
    .B(_1005_),
    .Y(_1006_));
 sg13g2_o21ai_1 _3315_ (.B1(_0958_),
    .Y(_1007_),
    .A1(_1004_),
    .A2(_1006_));
 sg13g2_a21oi_1 _3316_ (.A1(net496),
    .A2(_1007_),
    .Y(_0212_),
    .B1(net647));
 sg13g2_nand2_1 _3317_ (.Y(_1008_),
    .A(net874),
    .B(net542));
 sg13g2_and3_1 _3318_ (.X(_1009_),
    .A(net584),
    .B(net582),
    .C(_0973_));
 sg13g2_nor2_1 _3319_ (.A(net874),
    .B(net537),
    .Y(_1010_));
 sg13g2_and3_1 _3320_ (.X(_1011_),
    .A(net584),
    .B(net582),
    .C(_0935_));
 sg13g2_a221oi_1 _3321_ (.B2(_1011_),
    .C1(_1010_),
    .B1(net532),
    .A1(net1286),
    .Y(_1012_),
    .A2(net537));
 sg13g2_a21oi_1 _3322_ (.A1(net1286),
    .A2(net534),
    .Y(_1013_),
    .B1(net540));
 sg13g2_o21ai_1 _3323_ (.B1(_1013_),
    .Y(_1014_),
    .A1(_1009_),
    .A2(_1012_));
 sg13g2_a21oi_1 _3324_ (.A1(net875),
    .A2(net1287),
    .Y(_0213_),
    .B1(net647));
 sg13g2_nand2_1 _3325_ (.Y(_1015_),
    .A(net717),
    .B(net542));
 sg13g2_nand2_1 _3326_ (.Y(_1016_),
    .A(net1307),
    .B(net533));
 sg13g2_and3_1 _3327_ (.X(_1017_),
    .A(net584),
    .B(net582),
    .C(_0936_));
 sg13g2_nand3_1 _3328_ (.B(_1016_),
    .C(_1017_),
    .A(_0981_),
    .Y(_1018_));
 sg13g2_a21oi_1 _3329_ (.A1(net1307),
    .A2(net535),
    .Y(_1019_),
    .B1(_1017_));
 sg13g2_o21ai_1 _3330_ (.B1(_1019_),
    .Y(_1020_),
    .A1(net717),
    .A2(net535));
 sg13g2_a21o_1 _3331_ (.A2(_1020_),
    .A1(_1018_),
    .B1(net540),
    .X(_1021_));
 sg13g2_a21oi_1 _3332_ (.A1(net718),
    .A2(_1021_),
    .Y(_0214_),
    .B1(net643));
 sg13g2_nand2_1 _3333_ (.Y(_1022_),
    .A(net1087),
    .B(net541));
 sg13g2_nor4_1 _3334_ (.A(_0042_),
    .B(_0971_),
    .C(_0972_),
    .D(_0989_),
    .Y(_1023_));
 sg13g2_mux2_1 _3335_ (.A0(net1087),
    .A1(_1438_),
    .S(net536),
    .X(_1024_));
 sg13g2_nand4_1 _3336_ (.B(_0043_),
    .C(net531),
    .A(net583),
    .Y(_1025_),
    .D(_0933_));
 sg13g2_a22oi_1 _3337_ (.Y(_1026_),
    .B1(_1024_),
    .B2(_1025_),
    .A2(_1023_),
    .A1(_0961_));
 sg13g2_o21ai_1 _3338_ (.B1(_0958_),
    .Y(_1027_),
    .A1(_1438_),
    .A2(net531));
 sg13g2_o21ai_1 _3339_ (.B1(net1088),
    .Y(_1028_),
    .A1(_1026_),
    .A2(_1027_));
 sg13g2_and2_1 _3340_ (.A(net683),
    .B(net1089),
    .X(_0215_));
 sg13g2_nor4_1 _3341_ (.A(net533),
    .B(_0960_),
    .C(_0989_),
    .D(_1001_),
    .Y(_1029_));
 sg13g2_nand4_1 _3342_ (.B(net571),
    .C(net2),
    .A(\comm_ic0.spi0.data_ind[3] ),
    .Y(_1030_),
    .D(_1601_));
 sg13g2_nand2b_1 _3343_ (.Y(_1031_),
    .B(net531),
    .A_N(_1030_));
 sg13g2_o21ai_1 _3344_ (.B1(_1031_),
    .Y(_1032_),
    .A1(net1340),
    .A2(_1029_));
 sg13g2_a22oi_1 _3345_ (.Y(_1033_),
    .B1(_0958_),
    .B2(_1032_),
    .A2(net541),
    .A1(net516));
 sg13g2_nor2_1 _3346_ (.A(net647),
    .B(net517),
    .Y(_0216_));
 sg13g2_nand2_1 _3347_ (.Y(_1034_),
    .A(net860),
    .B(net541));
 sg13g2_nand2_1 _3348_ (.Y(_1035_),
    .A(net571),
    .B(_0968_));
 sg13g2_o21ai_1 _3349_ (.B1(_1035_),
    .Y(_1036_),
    .A1(net860),
    .A2(net535));
 sg13g2_a21oi_1 _3350_ (.A1(_0960_),
    .A2(_0974_),
    .Y(_1037_),
    .B1(net533));
 sg13g2_a22oi_1 _3351_ (.Y(_1038_),
    .B1(_1036_),
    .B2(_1037_),
    .A2(net536),
    .A1(net1294));
 sg13g2_nor2_1 _3352_ (.A(_0961_),
    .B(_0977_),
    .Y(_1039_));
 sg13g2_o21ai_1 _3353_ (.B1(_0958_),
    .Y(_1040_),
    .A1(_1038_),
    .A2(_1039_));
 sg13g2_a21oi_1 _3354_ (.A1(net861),
    .A2(net1295),
    .Y(_0217_),
    .B1(net647));
 sg13g2_nand2_1 _3355_ (.Y(_1041_),
    .A(net889),
    .B(net541));
 sg13g2_and2_1 _3356_ (.A(net571),
    .B(_0982_),
    .X(_1042_));
 sg13g2_nand2_1 _3357_ (.Y(_1043_),
    .A(net1308),
    .B(net533));
 sg13g2_a21oi_1 _3358_ (.A1(net1308),
    .A2(net535),
    .Y(_1044_),
    .B1(_1042_));
 sg13g2_o21ai_1 _3359_ (.B1(_1044_),
    .Y(_1045_),
    .A1(net889),
    .A2(net535));
 sg13g2_nand3_1 _3360_ (.B(_1042_),
    .C(_1043_),
    .A(_0981_),
    .Y(_1046_));
 sg13g2_a21o_1 _3361_ (.A2(_1046_),
    .A1(_1045_),
    .B1(net540),
    .X(_1047_));
 sg13g2_a21oi_1 _3362_ (.A1(net890),
    .A2(_1047_),
    .Y(_0218_),
    .B1(net643));
 sg13g2_nand2_1 _3363_ (.Y(_1048_),
    .A(net877),
    .B(net542));
 sg13g2_and2_1 _3364_ (.A(net571),
    .B(_0991_),
    .X(_1049_));
 sg13g2_nor2_1 _3365_ (.A(net877),
    .B(net536),
    .Y(_1050_));
 sg13g2_nor3_1 _3366_ (.A(net583),
    .B(net582),
    .C(_0934_),
    .Y(_1051_));
 sg13g2_a221oi_1 _3367_ (.B2(_1051_),
    .C1(_1050_),
    .B1(net531),
    .A1(net1281),
    .Y(_1052_),
    .A2(net537));
 sg13g2_a21oi_1 _3368_ (.A1(net1281),
    .A2(net534),
    .Y(_1053_),
    .B1(_0959_));
 sg13g2_o21ai_1 _3369_ (.B1(_1053_),
    .Y(_1054_),
    .A1(_1049_),
    .A2(_1052_));
 sg13g2_a21oi_1 _3370_ (.A1(net878),
    .A2(net1282),
    .Y(_0219_),
    .B1(net647));
 sg13g2_nand2_1 _3371_ (.Y(_1055_),
    .A(net795),
    .B(net541));
 sg13g2_a21oi_1 _3372_ (.A1(_0962_),
    .A2(_1002_),
    .Y(_1056_),
    .B1(net1289));
 sg13g2_nor2_1 _3373_ (.A(_0961_),
    .B(_1005_),
    .Y(_1057_));
 sg13g2_o21ai_1 _3374_ (.B1(_0958_),
    .Y(_1058_),
    .A1(_1056_),
    .A2(_1057_));
 sg13g2_a21oi_1 _3375_ (.A1(net796),
    .A2(_1058_),
    .Y(_0220_),
    .B1(net650));
 sg13g2_nand3_1 _3376_ (.B(net571),
    .C(_0973_),
    .A(net584),
    .Y(_1059_));
 sg13g2_o21ai_1 _3377_ (.B1(net923),
    .Y(_1060_),
    .A1(\comm_ic0.spi0.CPHA ),
    .A2(_1451_));
 sg13g2_o21ai_1 _3378_ (.B1(_1060_),
    .Y(_1061_),
    .A1(\comm_ic0.spi0.data_out[13] ),
    .A2(net537));
 sg13g2_and4_1 _3379_ (.A(net584),
    .B(net571),
    .C(net532),
    .D(_0935_),
    .X(_1062_));
 sg13g2_o21ai_1 _3380_ (.B1(_1059_),
    .Y(_1063_),
    .A1(_1061_),
    .A2(_1062_));
 sg13g2_a21oi_1 _3381_ (.A1(net923),
    .A2(net534),
    .Y(_1064_),
    .B1(net540));
 sg13g2_a22oi_1 _3382_ (.Y(_1065_),
    .B1(_1063_),
    .B2(net924),
    .A2(net542),
    .A1(\comm_ic0.spi0.data_out[13] ));
 sg13g2_nor2_1 _3383_ (.A(net645),
    .B(net925),
    .Y(_0221_));
 sg13g2_nand2_1 _3384_ (.Y(_1066_),
    .A(net871),
    .B(net541));
 sg13g2_nand3_1 _3385_ (.B(net571),
    .C(_0936_),
    .A(net584),
    .Y(_1067_));
 sg13g2_nand2b_1 _3386_ (.Y(_1068_),
    .B(net531),
    .A_N(_1067_));
 sg13g2_mux2_1 _3387_ (.A0(_1405_),
    .A1(net1302),
    .S(net536),
    .X(_1069_));
 sg13g2_a21oi_1 _3388_ (.A1(_1068_),
    .A2(_1069_),
    .Y(_1070_),
    .B1(net540));
 sg13g2_o21ai_1 _3389_ (.B1(_1070_),
    .Y(_1071_),
    .A1(_0981_),
    .A2(_1067_));
 sg13g2_a21oi_1 _3390_ (.A1(net872),
    .A2(_1071_),
    .Y(_0222_),
    .B1(net650));
 sg13g2_nand2_1 _3391_ (.Y(_1072_),
    .A(net1285),
    .B(net541));
 sg13g2_and2_1 _3392_ (.A(_0960_),
    .B(_1023_),
    .X(_1073_));
 sg13g2_nor2_1 _3393_ (.A(\comm_ic0.spi0.data_out[15] ),
    .B(net535),
    .Y(_1074_));
 sg13g2_nor3_1 _3394_ (.A(_1401_),
    .B(_0043_),
    .C(_0934_),
    .Y(_1075_));
 sg13g2_a221oi_1 _3395_ (.B2(_1075_),
    .C1(_1074_),
    .B1(_1598_),
    .A1(net956),
    .Y(_1076_),
    .A2(net536));
 sg13g2_a21oi_1 _3396_ (.A1(net956),
    .A2(net534),
    .Y(_1077_),
    .B1(net540));
 sg13g2_o21ai_1 _3397_ (.B1(net957),
    .Y(_1078_),
    .A1(_1073_),
    .A2(_1076_));
 sg13g2_a21oi_1 _3398_ (.A1(_1072_),
    .A2(net958),
    .Y(_0223_),
    .B1(net650));
 sg13g2_nand2b_1 _3399_ (.Y(_1079_),
    .B(\comm_ic0.spi0.curr_st[0] ),
    .A_N(\comm_ic0.spi0.curr_st[3] ));
 sg13g2_nand4_1 _3400_ (.B(net683),
    .C(_1458_),
    .A(net974),
    .Y(_1080_),
    .D(_1079_));
 sg13g2_o21ai_1 _3401_ (.B1(net975),
    .Y(_0224_),
    .A1(net1106),
    .A2(_1461_));
 sg13g2_nor2_1 _3402_ (.A(\comm_ic0.spi0.curr_st[0] ),
    .B(net645),
    .Y(_1081_));
 sg13g2_a22oi_1 _3403_ (.Y(_1082_),
    .B1(net558),
    .B2(\comm_ic0.spi0.clk_cnt_reg[0] ),
    .A2(net570),
    .A1(net962));
 sg13g2_inv_1 _3404_ (.Y(_0225_),
    .A(net963));
 sg13g2_a22oi_1 _3405_ (.Y(_1083_),
    .B1(net558),
    .B2(\comm_ic0.spi0.clk_cnt_reg[1] ),
    .A2(net570),
    .A1(net930));
 sg13g2_inv_1 _3406_ (.Y(_0226_),
    .A(net931));
 sg13g2_a22oi_1 _3407_ (.Y(_1084_),
    .B1(net558),
    .B2(net880),
    .A2(net570),
    .A1(net844));
 sg13g2_inv_1 _3408_ (.Y(_0227_),
    .A(net881));
 sg13g2_a22oi_1 _3409_ (.Y(_1085_),
    .B1(net557),
    .B2(net992),
    .A2(net568),
    .A1(net983));
 sg13g2_inv_1 _3410_ (.Y(_0228_),
    .A(net993));
 sg13g2_a22oi_1 _3411_ (.Y(_1086_),
    .B1(net557),
    .B2(net828),
    .A2(net568),
    .A1(net792));
 sg13g2_inv_1 _3412_ (.Y(_0229_),
    .A(net829));
 sg13g2_a22oi_1 _3413_ (.Y(_1087_),
    .B1(net557),
    .B2(net911),
    .A2(net568),
    .A1(net865));
 sg13g2_inv_1 _3414_ (.Y(_0230_),
    .A(net912));
 sg13g2_a22oi_1 _3415_ (.Y(_1088_),
    .B1(net557),
    .B2(net744),
    .A2(net568),
    .A1(net401));
 sg13g2_inv_1 _3416_ (.Y(_0231_),
    .A(net745));
 sg13g2_a22oi_1 _3417_ (.Y(_1089_),
    .B1(net559),
    .B2(net1336),
    .A2(net570),
    .A1(net478));
 sg13g2_inv_1 _3418_ (.Y(_0232_),
    .A(net479));
 sg13g2_a22oi_1 _3419_ (.Y(_1090_),
    .B1(net557),
    .B2(net341),
    .A2(net568),
    .A1(net438));
 sg13g2_inv_1 _3420_ (.Y(_0233_),
    .A(net342));
 sg13g2_a22oi_1 _3421_ (.Y(_1091_),
    .B1(net557),
    .B2(net416),
    .A2(net568),
    .A1(net353));
 sg13g2_inv_1 _3422_ (.Y(_0234_),
    .A(net417));
 sg13g2_a22oi_1 _3423_ (.Y(_1092_),
    .B1(net556),
    .B2(net335),
    .A2(net567),
    .A1(net767));
 sg13g2_inv_1 _3424_ (.Y(_0235_),
    .A(net336));
 sg13g2_a22oi_1 _3425_ (.Y(_1093_),
    .B1(net559),
    .B2(net407),
    .A2(net569),
    .A1(net398));
 sg13g2_inv_1 _3426_ (.Y(_0236_),
    .A(net408));
 sg13g2_a22oi_1 _3427_ (.Y(_1094_),
    .B1(net556),
    .B2(net489),
    .A2(net567),
    .A1(net469));
 sg13g2_inv_1 _3428_ (.Y(_0237_),
    .A(net490));
 sg13g2_a22oi_1 _3429_ (.Y(_1095_),
    .B1(net556),
    .B2(net472),
    .A2(net567),
    .A1(net347));
 sg13g2_inv_1 _3430_ (.Y(_0238_),
    .A(net473));
 sg13g2_a22oi_1 _3431_ (.Y(_1096_),
    .B1(net556),
    .B2(net808),
    .A2(net567),
    .A1(net404));
 sg13g2_inv_1 _3432_ (.Y(_0239_),
    .A(net809));
 sg13g2_a22oi_1 _3433_ (.Y(_1097_),
    .B1(net556),
    .B2(net501),
    .A2(net567),
    .A1(net356));
 sg13g2_inv_1 _3434_ (.Y(_0240_),
    .A(net502));
 sg13g2_a22oi_1 _3435_ (.Y(_1098_),
    .B1(net556),
    .B2(net435),
    .A2(net567),
    .A1(net432));
 sg13g2_inv_1 _3436_ (.Y(_0241_),
    .A(net436));
 sg13g2_a22oi_1 _3437_ (.Y(_1099_),
    .B1(net557),
    .B2(net317),
    .A2(net568),
    .A1(net441));
 sg13g2_inv_1 _3438_ (.Y(_0242_),
    .A(net318));
 sg13g2_a22oi_1 _3439_ (.Y(_1100_),
    .B1(net556),
    .B2(net329),
    .A2(net567),
    .A1(net380));
 sg13g2_inv_1 _3440_ (.Y(_0243_),
    .A(net330));
 sg13g2_a22oi_1 _3441_ (.Y(_1101_),
    .B1(net556),
    .B2(net492),
    .A2(net567),
    .A1(net350));
 sg13g2_inv_1 _3442_ (.Y(_0244_),
    .A(net493));
 sg13g2_a22oi_1 _3443_ (.Y(_1102_),
    .B1(net558),
    .B2(net323),
    .A2(net569),
    .A1(\comm_ic0.spi0.data_in[12] ));
 sg13g2_inv_1 _3444_ (.Y(_0245_),
    .A(net324));
 sg13g2_a22oi_1 _3445_ (.Y(_1103_),
    .B1(net558),
    .B2(net359),
    .A2(net569),
    .A1(net1343));
 sg13g2_inv_1 _3446_ (.Y(_0246_),
    .A(net360));
 sg13g2_a22oi_1 _3447_ (.Y(_1104_),
    .B1(net558),
    .B2(net371),
    .A2(net569),
    .A1(net968));
 sg13g2_inv_1 _3448_ (.Y(_0247_),
    .A(net372));
 sg13g2_a22oi_1 _3449_ (.Y(_1105_),
    .B1(net558),
    .B2(net362),
    .A2(net569),
    .A1(net995));
 sg13g2_inv_1 _3450_ (.Y(_0248_),
    .A(net363));
 sg13g2_nand2_1 _3451_ (.Y(_1106_),
    .A(_1434_),
    .B(net1194));
 sg13g2_nor3_1 _3452_ (.A(net1210),
    .B(net537),
    .C(_1603_),
    .Y(_1107_));
 sg13g2_a21o_1 _3453_ (.A2(net537),
    .A1(net1210),
    .B1(_1107_),
    .X(_1108_));
 sg13g2_a21oi_1 _3454_ (.A1(_1595_),
    .A2(_0999_),
    .Y(_1109_),
    .B1(_1434_));
 sg13g2_o21ai_1 _3455_ (.B1(net1316),
    .Y(_1110_),
    .A1(_1595_),
    .A2(_1108_));
 sg13g2_o21ai_1 _3456_ (.B1(net683),
    .Y(_1111_),
    .A1(net1210),
    .A2(_0923_));
 sg13g2_a21oi_1 _3457_ (.A1(_1106_),
    .A2(net1317),
    .Y(_0249_),
    .B1(net1211));
 sg13g2_nor2_1 _3458_ (.A(net586),
    .B(net532),
    .Y(_1112_));
 sg13g2_o21ai_1 _3459_ (.B1(net639),
    .Y(_1113_),
    .A1(net534),
    .A2(_1000_));
 sg13g2_o21ai_1 _3460_ (.B1(_1106_),
    .Y(_1114_),
    .A1(_1112_),
    .A2(_1113_));
 sg13g2_o21ai_1 _3461_ (.B1(_1114_),
    .Y(_1115_),
    .A1(net908),
    .A2(_0923_));
 sg13g2_nor2_1 _3462_ (.A(net645),
    .B(net909),
    .Y(_0250_));
 sg13g2_nand4_1 _3463_ (.B(net1143),
    .C(net532),
    .A(net1146),
    .Y(_1116_),
    .D(_1601_));
 sg13g2_nand3_1 _3464_ (.B(net1143),
    .C(_1600_),
    .A(net583),
    .Y(_1117_));
 sg13g2_nand3_1 _3465_ (.B(_1116_),
    .C(_1117_),
    .A(_1106_),
    .Y(_1118_));
 sg13g2_o21ai_1 _3466_ (.B1(net683),
    .Y(_1119_),
    .A1(net1187),
    .A2(_0923_));
 sg13g2_nor2b_1 _3467_ (.A(net1188),
    .B_N(_1118_),
    .Y(_0251_));
 sg13g2_nand3_1 _3468_ (.B(net1143),
    .C(_1602_),
    .A(net1146),
    .Y(_1120_));
 sg13g2_nand2b_1 _3469_ (.Y(_1121_),
    .B(net1193),
    .A_N(net1109));
 sg13g2_nand3_1 _3470_ (.B(net1194),
    .C(_1121_),
    .A(_1434_),
    .Y(_1122_));
 sg13g2_o21ai_1 _3471_ (.B1(net683),
    .Y(_1123_),
    .A1(net1146),
    .A2(_0923_));
 sg13g2_a21oi_1 _3472_ (.A1(net1147),
    .A2(_1122_),
    .Y(_0252_),
    .B1(_1123_));
 sg13g2_a22oi_1 _3473_ (.Y(_1124_),
    .B1(net559),
    .B2(net699),
    .A2(net569),
    .A1(net950));
 sg13g2_inv_1 _3474_ (.Y(_0253_),
    .A(net700));
 sg13g2_a22oi_1 _3475_ (.Y(_1125_),
    .B1(net559),
    .B2(\comm_ic0.spi0.CPHA ),
    .A2(net569),
    .A1(net774));
 sg13g2_inv_1 _3476_ (.Y(_0254_),
    .A(net775));
 sg13g2_a21o_1 _3477_ (.A2(net538),
    .A1(net595),
    .B1(net588),
    .X(_1126_));
 sg13g2_a221oi_1 _3478_ (.B2(net539),
    .C1(net588),
    .B1(_0773_),
    .A1(net595),
    .Y(_1127_),
    .A2(net538));
 sg13g2_nor2_1 _3479_ (.A(\comm_ic0.i2c0.scl_cnt[0] ),
    .B(_1127_),
    .Y(_1128_));
 sg13g2_nor3_2 _3480_ (.A(net588),
    .B(net595),
    .C(_0773_),
    .Y(_1129_));
 sg13g2_nand2_2 _3481_ (.Y(_1130_),
    .A(net1213),
    .B(_1129_));
 sg13g2_nor2_1 _3482_ (.A(net1054),
    .B(_1130_),
    .Y(_1131_));
 sg13g2_a22oi_1 _3483_ (.Y(_1132_),
    .B1(_0773_),
    .B2(_1546_),
    .A2(_1564_),
    .A1(net595));
 sg13g2_nor2_1 _3484_ (.A(net1230),
    .B(_1132_),
    .Y(_1133_));
 sg13g2_nor3_1 _3485_ (.A(_1128_),
    .B(_1131_),
    .C(net1231),
    .Y(_1134_));
 sg13g2_nor2_1 _3486_ (.A(net643),
    .B(net1232),
    .Y(_0255_));
 sg13g2_xor2_1 _3487_ (.B(net1270),
    .A(\comm_ic0.i2c0.scl_cnt[0] ),
    .X(_1135_));
 sg13g2_nor2_1 _3488_ (.A(_1127_),
    .B(net1271),
    .Y(_1136_));
 sg13g2_nor2_1 _3489_ (.A(net1062),
    .B(net1054),
    .Y(_1137_));
 sg13g2_xor2_1 _3490_ (.B(net1054),
    .A(net1062),
    .X(_1138_));
 sg13g2_nor2_1 _3491_ (.A(_1130_),
    .B(_1138_),
    .Y(_1139_));
 sg13g2_xor2_1 _3492_ (.B(net1230),
    .A(\comm_ic0.i2c0.clk_cnt_reg[1] ),
    .X(_1140_));
 sg13g2_nor2_1 _3493_ (.A(_1132_),
    .B(_1140_),
    .Y(_1141_));
 sg13g2_nor3_1 _3494_ (.A(net1272),
    .B(_1139_),
    .C(_1141_),
    .Y(_1142_));
 sg13g2_nor2_1 _3495_ (.A(net642),
    .B(net1273),
    .Y(_0256_));
 sg13g2_nand2_1 _3496_ (.Y(_1143_),
    .A(net1204),
    .B(_1542_));
 sg13g2_or2_1 _3497_ (.X(_1144_),
    .B(_1542_),
    .A(net1204));
 sg13g2_a21oi_1 _3498_ (.A1(net1205),
    .A2(_1144_),
    .Y(_1145_),
    .B1(_1127_));
 sg13g2_nand2_1 _3499_ (.Y(_1146_),
    .A(_0066_),
    .B(_1137_));
 sg13g2_or2_1 _3500_ (.X(_1147_),
    .B(_1137_),
    .A(_0066_));
 sg13g2_a21oi_1 _3501_ (.A1(_1146_),
    .A2(_1147_),
    .Y(_1148_),
    .B1(_1130_));
 sg13g2_nor3_1 _3502_ (.A(\comm_ic0.i2c0.clk_cnt_reg[2] ),
    .B(\comm_ic0.i2c0.clk_cnt_reg[1] ),
    .C(net1230),
    .Y(_1149_));
 sg13g2_o21ai_1 _3503_ (.B1(\comm_ic0.i2c0.clk_cnt_reg[2] ),
    .Y(_1150_),
    .A1(\comm_ic0.i2c0.clk_cnt_reg[1] ),
    .A2(\comm_ic0.i2c0.clk_cnt_reg[0] ));
 sg13g2_nor2b_1 _3504_ (.A(_1149_),
    .B_N(_1150_),
    .Y(_1151_));
 sg13g2_nor2_1 _3505_ (.A(_1132_),
    .B(_1151_),
    .Y(_1152_));
 sg13g2_nor3_1 _3506_ (.A(net1206),
    .B(_1148_),
    .C(_1152_),
    .Y(_1153_));
 sg13g2_nor2_1 _3507_ (.A(net642),
    .B(net1207),
    .Y(_0257_));
 sg13g2_xor2_1 _3508_ (.B(net1205),
    .A(\comm_ic0.i2c0.scl_cnt[3] ),
    .X(_1154_));
 sg13g2_nor2_1 _3509_ (.A(_1127_),
    .B(_1154_),
    .Y(_1155_));
 sg13g2_xor2_1 _3510_ (.B(_1146_),
    .A(net1025),
    .X(_1156_));
 sg13g2_nor2_1 _3511_ (.A(_1130_),
    .B(_1156_),
    .Y(_1157_));
 sg13g2_nor4_2 _3512_ (.A(net1246),
    .B(\comm_ic0.i2c0.clk_cnt_reg[2] ),
    .C(\comm_ic0.i2c0.clk_cnt_reg[1] ),
    .Y(_1158_),
    .D(net1230));
 sg13g2_xnor2_1 _3513_ (.Y(_1159_),
    .A(net1246),
    .B(_1149_));
 sg13g2_nor2_1 _3514_ (.A(_1132_),
    .B(net1247),
    .Y(_1160_));
 sg13g2_nor3_1 _3515_ (.A(_1155_),
    .B(_1157_),
    .C(net1248),
    .Y(_1161_));
 sg13g2_nor2_1 _3516_ (.A(net642),
    .B(net1249),
    .Y(_0258_));
 sg13g2_or2_1 _3517_ (.X(_1162_),
    .B(_1543_),
    .A(net1197));
 sg13g2_nand2_1 _3518_ (.Y(_1163_),
    .A(net1197),
    .B(_1543_));
 sg13g2_a21oi_1 _3519_ (.A1(_1162_),
    .A2(net1198),
    .Y(_1164_),
    .B1(_1127_));
 sg13g2_nor4_2 _3520_ (.A(net1025),
    .B(net857),
    .C(net1062),
    .Y(_1165_),
    .D(net1054));
 sg13g2_nand2_1 _3521_ (.Y(_1166_),
    .A(net1256),
    .B(_1165_));
 sg13g2_or2_1 _3522_ (.X(_1167_),
    .B(_1165_),
    .A(_0068_));
 sg13g2_a21oi_1 _3523_ (.A1(_1166_),
    .A2(_1167_),
    .Y(_1168_),
    .B1(_1130_));
 sg13g2_nor2b_1 _3524_ (.A(\comm_ic0.i2c0.clk_cnt_reg[4] ),
    .B_N(_1158_),
    .Y(_1169_));
 sg13g2_xnor2_1 _3525_ (.Y(_1170_),
    .A(\comm_ic0.i2c0.clk_cnt_reg[4] ),
    .B(_1158_));
 sg13g2_nor2_1 _3526_ (.A(_1132_),
    .B(_1170_),
    .Y(_1171_));
 sg13g2_nor3_1 _3527_ (.A(net1199),
    .B(_1168_),
    .C(_1171_),
    .Y(_1172_));
 sg13g2_nor2_1 _3528_ (.A(net652),
    .B(net1200),
    .Y(_0259_));
 sg13g2_xor2_1 _3529_ (.B(_1162_),
    .A(\comm_ic0.i2c0.scl_cnt[5] ),
    .X(_1173_));
 sg13g2_nor2_1 _3530_ (.A(_1127_),
    .B(_1173_),
    .Y(_1174_));
 sg13g2_nor2b_1 _3531_ (.A(\comm_ic0.i2c0.clk_cnt_reg[5] ),
    .B_N(_1169_),
    .Y(_1175_));
 sg13g2_xnor2_1 _3532_ (.Y(_1176_),
    .A(\comm_ic0.i2c0.clk_cnt_reg[5] ),
    .B(_1169_));
 sg13g2_nor2_1 _3533_ (.A(_1132_),
    .B(_1176_),
    .Y(_1177_));
 sg13g2_xor2_1 _3534_ (.B(net1257),
    .A(net1028),
    .X(_1178_));
 sg13g2_nor2_1 _3535_ (.A(_1130_),
    .B(_1178_),
    .Y(_1179_));
 sg13g2_nor3_1 _3536_ (.A(_1174_),
    .B(_1177_),
    .C(net1258),
    .Y(_1180_));
 sg13g2_nor2_1 _3537_ (.A(net652),
    .B(net1259),
    .Y(_0260_));
 sg13g2_xor2_1 _3538_ (.B(_1544_),
    .A(net1156),
    .X(_1181_));
 sg13g2_nand2b_1 _3539_ (.Y(_1182_),
    .B(net1157),
    .A_N(_1127_));
 sg13g2_nor2_1 _3540_ (.A(net1028),
    .B(net847),
    .Y(_1183_));
 sg13g2_nand3_1 _3541_ (.B(_1165_),
    .C(_1183_),
    .A(net1305),
    .Y(_1184_));
 sg13g2_a21o_1 _3542_ (.A2(_1183_),
    .A1(_1165_),
    .B1(net1305),
    .X(_1185_));
 sg13g2_a21oi_1 _3543_ (.A1(_1184_),
    .A2(_1185_),
    .Y(_1186_),
    .B1(_1130_));
 sg13g2_nor2b_1 _3544_ (.A(\comm_ic0.i2c0.clk_cnt_reg[6] ),
    .B_N(_1175_),
    .Y(_1187_));
 sg13g2_xnor2_1 _3545_ (.Y(_1188_),
    .A(\comm_ic0.i2c0.clk_cnt_reg[6] ),
    .B(_1175_));
 sg13g2_nor2_1 _3546_ (.A(_1132_),
    .B(_1188_),
    .Y(_1189_));
 sg13g2_nor2_1 _3547_ (.A(_1186_),
    .B(_1189_),
    .Y(_1190_));
 sg13g2_a21oi_1 _3548_ (.A1(net1158),
    .A2(net1306),
    .Y(_0261_),
    .B1(net652));
 sg13g2_o21ai_1 _3549_ (.B1(net539),
    .Y(_1191_),
    .A1(_1428_),
    .A2(_1565_));
 sg13g2_xor2_1 _3550_ (.B(_1187_),
    .A(\comm_ic0.i2c0.clk_cnt_reg[7] ),
    .X(_1192_));
 sg13g2_nor2b_1 _3551_ (.A(_1545_),
    .B_N(net1079),
    .Y(_1193_));
 sg13g2_a221oi_1 _3552_ (.B2(_1192_),
    .C1(_1193_),
    .B1(_1191_),
    .A1(_1546_),
    .Y(_1194_),
    .A2(_1126_));
 sg13g2_xnor2_1 _3553_ (.Y(_1195_),
    .A(net1019),
    .B(_1184_));
 sg13g2_nand3_1 _3554_ (.B(_1129_),
    .C(_1195_),
    .A(net1213),
    .Y(_1196_));
 sg13g2_o21ai_1 _3555_ (.B1(net1214),
    .Y(_1197_),
    .A1(_1129_),
    .A2(_1194_));
 sg13g2_and2_1 _3556_ (.A(net689),
    .B(net1215),
    .X(_0262_));
 sg13g2_or2_1 _3557_ (.X(_1198_),
    .B(_1473_),
    .A(_1463_));
 sg13g2_o21ai_1 _3558_ (.B1(net621),
    .Y(_1199_),
    .A1(net660),
    .A2(net1182));
 sg13g2_nand4_1 _3559_ (.B(net3),
    .C(_1527_),
    .A(net625),
    .Y(_1200_),
    .D(_1624_));
 sg13g2_o21ai_1 _3560_ (.B1(_1200_),
    .Y(_1201_),
    .A1(net625),
    .A2(_1473_));
 sg13g2_nand4_1 _3561_ (.B(_1198_),
    .C(net1183),
    .A(net447),
    .Y(_1202_),
    .D(_1201_));
 sg13g2_nand4_1 _3562_ (.B(_1198_),
    .C(net1183),
    .A(net634),
    .Y(_1203_),
    .D(_1201_));
 sg13g2_nand2_1 _3563_ (.Y(_1204_),
    .A(net338),
    .B(_1203_));
 sg13g2_a21o_1 _3564_ (.A2(_1204_),
    .A1(net1184),
    .B1(net656),
    .X(_1205_));
 sg13g2_inv_1 _3565_ (.Y(_0263_),
    .A(net1185));
 sg13g2_and2_2 _3566_ (.A(net628),
    .B(_1465_),
    .X(_1206_));
 sg13g2_o21ai_1 _3567_ (.B1(net686),
    .Y(_1207_),
    .A1(net1054),
    .A2(_1206_));
 sg13g2_a21oi_1 _3568_ (.A1(_1335_),
    .A2(_1206_),
    .Y(_0264_),
    .B1(_1207_));
 sg13g2_o21ai_1 _3569_ (.B1(net677),
    .Y(_1208_),
    .A1(net1062),
    .A2(_1206_));
 sg13g2_a21oi_1 _3570_ (.A1(net660),
    .A2(_1206_),
    .Y(_0265_),
    .B1(net1126));
 sg13g2_o21ai_1 _3571_ (.B1(net677),
    .Y(_1209_),
    .A1(net857),
    .A2(_1206_));
 sg13g2_a21oi_1 _3572_ (.A1(_1332_),
    .A2(_1206_),
    .Y(_0266_),
    .B1(net1043));
 sg13g2_o21ai_1 _3573_ (.B1(net686),
    .Y(_1210_),
    .A1(net1025),
    .A2(_1206_));
 sg13g2_a21oi_1 _3574_ (.A1(_1330_),
    .A2(_1206_),
    .Y(_0267_),
    .B1(net1094));
 sg13g2_nor2_1 _3575_ (.A(net447),
    .B(net565),
    .Y(_1211_));
 sg13g2_nand3_1 _3576_ (.B(net627),
    .C(_1211_),
    .A(net338),
    .Y(_1212_));
 sg13g2_o21ai_1 _3577_ (.B1(net688),
    .Y(_1213_),
    .A1(net672),
    .A2(_1212_));
 sg13g2_a21oi_1 _3578_ (.A1(_1399_),
    .A2(_1212_),
    .Y(_0268_),
    .B1(_1213_));
 sg13g2_o21ai_1 _3579_ (.B1(net688),
    .Y(_1214_),
    .A1(net670),
    .A2(_1212_));
 sg13g2_a21oi_1 _3580_ (.A1(net499),
    .A2(_1212_),
    .Y(_0269_),
    .B1(_1214_));
 sg13g2_o21ai_1 _3581_ (.B1(net688),
    .Y(_1215_),
    .A1(net666),
    .A2(_1212_));
 sg13g2_a21oi_1 _3582_ (.A1(_1397_),
    .A2(_1212_),
    .Y(_0270_),
    .B1(_1215_));
 sg13g2_o21ai_1 _3583_ (.B1(net688),
    .Y(_1216_),
    .A1(net663),
    .A2(_1212_));
 sg13g2_a21oi_1 _3584_ (.A1(net390),
    .A2(_1212_),
    .Y(_0271_),
    .B1(_1216_));
 sg13g2_o21ai_1 _3585_ (.B1(net686),
    .Y(_1217_),
    .A1(net662),
    .A2(net521));
 sg13g2_a21oi_1 _3586_ (.A1(_1395_),
    .A2(net521),
    .Y(_0272_),
    .B1(_1217_));
 sg13g2_nor3_2 _3587_ (.A(net338),
    .B(net447),
    .C(net565),
    .Y(_1218_));
 sg13g2_nand2_2 _3588_ (.Y(_1219_),
    .A(net444),
    .B(_1218_));
 sg13g2_o21ai_1 _3589_ (.B1(net677),
    .Y(_1220_),
    .A1(net671),
    .A2(net445));
 sg13g2_a21oi_1 _3590_ (.A1(net476),
    .A2(net445),
    .Y(_0273_),
    .B1(_1220_));
 sg13g2_o21ai_1 _3591_ (.B1(net678),
    .Y(_1221_),
    .A1(net669),
    .A2(net445));
 sg13g2_a21oi_1 _3592_ (.A1(_1393_),
    .A2(net445),
    .Y(_0274_),
    .B1(_1221_));
 sg13g2_o21ai_1 _3593_ (.B1(net678),
    .Y(_1222_),
    .A1(net664),
    .A2(net445));
 sg13g2_a21oi_1 _3594_ (.A1(net461),
    .A2(net445),
    .Y(_0275_),
    .B1(_1222_));
 sg13g2_o21ai_1 _3595_ (.B1(net677),
    .Y(_1223_),
    .A1(net663),
    .A2(net445));
 sg13g2_a21oi_1 _3596_ (.A1(_1391_),
    .A2(net445),
    .Y(_0276_),
    .B1(_1223_));
 sg13g2_nor2_2 _3597_ (.A(net625),
    .B(_1373_),
    .Y(_1224_));
 sg13g2_a21oi_1 _3598_ (.A1(net1035),
    .A2(net1004),
    .Y(_1225_),
    .B1(_1224_));
 sg13g2_a21oi_1 _3599_ (.A1(net1218),
    .A2(_1211_),
    .Y(_1226_),
    .B1(_1225_));
 sg13g2_o21ai_1 _3600_ (.B1(net1228),
    .Y(_1227_),
    .A1(_1373_),
    .A2(_1463_));
 sg13g2_a221oi_1 _3601_ (.B2(_1390_),
    .C1(net659),
    .B1(_1227_),
    .A1(_1373_),
    .Y(_0277_),
    .A2(net1228));
 sg13g2_o21ai_1 _3602_ (.B1(net686),
    .Y(_1228_),
    .A1(net666),
    .A2(net521));
 sg13g2_a21oi_1 _3603_ (.A1(net739),
    .A2(net521),
    .Y(_0278_),
    .B1(_1228_));
 sg13g2_nand3_1 _3604_ (.B(net825),
    .C(net564),
    .A(net730),
    .Y(_1229_));
 sg13g2_o21ai_1 _3605_ (.B1(net680),
    .Y(_1230_),
    .A1(net673),
    .A2(_1229_));
 sg13g2_a21oi_1 _3606_ (.A1(_1388_),
    .A2(_1229_),
    .Y(_0279_),
    .B1(_1230_));
 sg13g2_o21ai_1 _3607_ (.B1(net680),
    .Y(_1231_),
    .A1(net668),
    .A2(_1229_));
 sg13g2_a21oi_1 _3608_ (.A1(_1387_),
    .A2(_1229_),
    .Y(_0280_),
    .B1(_1231_));
 sg13g2_o21ai_1 _3609_ (.B1(net680),
    .Y(_1232_),
    .A1(net665),
    .A2(_1229_));
 sg13g2_a21oi_1 _3610_ (.A1(net845),
    .A2(_1229_),
    .Y(_0281_),
    .B1(_1232_));
 sg13g2_o21ai_1 _3611_ (.B1(net680),
    .Y(_1233_),
    .A1(net661),
    .A2(_1229_));
 sg13g2_a21oi_1 _3612_ (.A1(net984),
    .A2(_1229_),
    .Y(_0282_),
    .B1(_1233_));
 sg13g2_o21ai_1 _3613_ (.B1(net678),
    .Y(_1234_),
    .A1(net774),
    .A2(_1523_));
 sg13g2_a21oi_1 _3614_ (.A1(_1332_),
    .A2(_1523_),
    .Y(_0283_),
    .B1(net990));
 sg13g2_nor2_2 _3615_ (.A(net662),
    .B(_1425_),
    .Y(_1235_));
 sg13g2_o21ai_1 _3616_ (.B1(net679),
    .Y(_1236_),
    .A1(net950),
    .A2(_1523_));
 sg13g2_a21oi_1 _3617_ (.A1(_1330_),
    .A2(_1523_),
    .Y(_0284_),
    .B1(net951));
 sg13g2_a21oi_1 _3618_ (.A1(net1035),
    .A2(net974),
    .Y(_1237_),
    .B1(_1224_));
 sg13g2_a21oi_2 _3619_ (.B1(_1373_),
    .Y(_1238_),
    .A2(net564),
    .A1(_1426_));
 sg13g2_nor2_1 _3620_ (.A(_1237_),
    .B(_1238_),
    .Y(_1239_));
 sg13g2_a21oi_1 _3621_ (.A1(net1065),
    .A2(_1239_),
    .Y(_1240_),
    .B1(net645));
 sg13g2_o21ai_1 _3622_ (.B1(net1066),
    .Y(_0285_),
    .A1(_1384_),
    .A2(_1239_));
 sg13g2_o21ai_1 _3623_ (.B1(net678),
    .Y(_1241_),
    .A1(net1076),
    .A2(_1518_));
 sg13g2_a21oi_1 _3624_ (.A1(_1335_),
    .A2(net548),
    .Y(_0286_),
    .B1(net1077));
 sg13g2_o21ai_1 _3625_ (.B1(net679),
    .Y(_1242_),
    .A1(net1007),
    .A2(net548));
 sg13g2_a21oi_1 _3626_ (.A1(net660),
    .A2(net548),
    .Y(_0287_),
    .B1(net1008));
 sg13g2_o21ai_1 _3627_ (.B1(net678),
    .Y(_1243_),
    .A1(net968),
    .A2(net548));
 sg13g2_a21oi_1 _3628_ (.A1(_1332_),
    .A2(net548),
    .Y(_0288_),
    .B1(net969));
 sg13g2_o21ai_1 _3629_ (.B1(net678),
    .Y(_1244_),
    .A1(net995),
    .A2(net548));
 sg13g2_a21oi_1 _3630_ (.A1(_1330_),
    .A2(net548),
    .Y(_0289_),
    .B1(net996));
 sg13g2_o21ai_1 _3631_ (.B1(net687),
    .Y(_1245_),
    .A1(net1109),
    .A2(_1523_));
 sg13g2_a21oi_1 _3632_ (.A1(net660),
    .A2(_1523_),
    .Y(_0290_),
    .B1(net1110));
 sg13g2_nand2_1 _3633_ (.Y(_1246_),
    .A(_1426_),
    .B(_1485_));
 sg13g2_nand2_1 _3634_ (.Y(_1247_),
    .A(net1035),
    .B(\comm_ic0.busy_uart ));
 sg13g2_nand2b_1 _3635_ (.Y(_1248_),
    .B(net621),
    .A_N(net1035));
 sg13g2_a22oi_1 _3636_ (.Y(_1249_),
    .B1(_1247_),
    .B2(_1248_),
    .A2(_1246_),
    .A1(net621));
 sg13g2_nand2_1 _3637_ (.Y(_1250_),
    .A(net667),
    .B(net621));
 sg13g2_o21ai_1 _3638_ (.B1(net692),
    .Y(_1251_),
    .A1(net942),
    .A2(net1036));
 sg13g2_a21oi_1 _3639_ (.A1(net1036),
    .A2(_1250_),
    .Y(_0291_),
    .B1(_1251_));
 sg13g2_nor2_1 _3640_ (.A(_1373_),
    .B(_1485_),
    .Y(_1252_));
 sg13g2_a221oi_1 _3641_ (.B2(net621),
    .C1(_1252_),
    .B1(_1246_),
    .A1(_1373_),
    .Y(_1253_),
    .A2(net1099));
 sg13g2_o21ai_1 _3642_ (.B1(net692),
    .Y(_1254_),
    .A1(net1074),
    .A2(net1100));
 sg13g2_a21oi_1 _3643_ (.A1(_1235_),
    .A2(net1100),
    .Y(_0292_),
    .B1(net1101));
 sg13g2_nand2_2 _3644_ (.Y(_1255_),
    .A(net825),
    .B(_1490_));
 sg13g2_o21ai_1 _3645_ (.B1(net683),
    .Y(_1256_),
    .A1(net673),
    .A2(net826));
 sg13g2_a21oi_1 _3646_ (.A1(net864),
    .A2(net826),
    .Y(_0293_),
    .B1(_1256_));
 sg13g2_o21ai_1 _3647_ (.B1(net683),
    .Y(_1257_),
    .A1(net669),
    .A2(net826));
 sg13g2_a21oi_1 _3648_ (.A1(_1380_),
    .A2(net826),
    .Y(_0294_),
    .B1(_1257_));
 sg13g2_o21ai_1 _3649_ (.B1(net684),
    .Y(_1258_),
    .A1(net665),
    .A2(net826));
 sg13g2_a21oi_1 _3650_ (.A1(_1379_),
    .A2(net826),
    .Y(_0295_),
    .B1(_1258_));
 sg13g2_a221oi_1 _3651_ (.B2(_1378_),
    .C1(net649),
    .B1(net826),
    .A1(_1490_),
    .Y(_0296_),
    .A2(_1235_));
 sg13g2_nand2_2 _3652_ (.Y(_1259_),
    .A(net624),
    .B(_1490_));
 sg13g2_o21ai_1 _3653_ (.B1(net691),
    .Y(_1260_),
    .A1(net673),
    .A2(_1259_));
 sg13g2_a21oi_1 _3654_ (.A1(net928),
    .A2(_1259_),
    .Y(_0297_),
    .B1(_1260_));
 sg13g2_o21ai_1 _3655_ (.B1(net691),
    .Y(_1261_),
    .A1(net5),
    .A2(_1259_));
 sg13g2_a21oi_1 _3656_ (.A1(net903),
    .A2(_1259_),
    .Y(_0298_),
    .B1(_1261_));
 sg13g2_o21ai_1 _3657_ (.B1(net691),
    .Y(_1262_),
    .A1(net666),
    .A2(_1259_));
 sg13g2_a21oi_1 _3658_ (.A1(net893),
    .A2(_1259_),
    .Y(_0299_),
    .B1(_1262_));
 sg13g2_o21ai_1 _3659_ (.B1(net691),
    .Y(_1263_),
    .A1(net662),
    .A2(_1259_));
 sg13g2_a21oi_1 _3660_ (.A1(net981),
    .A2(_1259_),
    .Y(_0300_),
    .B1(_1263_));
 sg13g2_nor2b_1 _3661_ (.A(_1224_),
    .B_N(_1247_),
    .Y(_1264_));
 sg13g2_o21ai_1 _3662_ (.B1(net1113),
    .Y(_1265_),
    .A1(_1246_),
    .A2(_1264_));
 sg13g2_o21ai_1 _3663_ (.B1(net1114),
    .Y(_1266_),
    .A1(net624),
    .A2(_1247_));
 sg13g2_nor2_1 _3664_ (.A(net657),
    .B(net1115),
    .Y(_0301_));
 sg13g2_o21ai_1 _3665_ (.B1(net692),
    .Y(_1267_),
    .A1(net801),
    .A2(_1486_));
 sg13g2_a21oi_1 _3666_ (.A1(_1335_),
    .A2(_1486_),
    .Y(_0302_),
    .B1(net937));
 sg13g2_o21ai_1 _3667_ (.B1(net692),
    .Y(_1268_),
    .A1(net760),
    .A2(_1486_));
 sg13g2_a21oi_1 _3668_ (.A1(net660),
    .A2(_1486_),
    .Y(_0303_),
    .B1(net940));
 sg13g2_a21oi_1 _3669_ (.A1(_1485_),
    .A2(_1496_),
    .Y(_1269_),
    .B1(net507));
 sg13g2_nor2_1 _3670_ (.A(net658),
    .B(net508),
    .Y(_0304_));
 sg13g2_a22oi_1 _3671_ (.Y(_1270_),
    .B1(_1520_),
    .B2(net672),
    .A2(_1472_),
    .A1(net1129));
 sg13g2_inv_1 _3672_ (.Y(_0305_),
    .A(net1130));
 sg13g2_a22oi_1 _3673_ (.Y(_1271_),
    .B1(_1520_),
    .B2(net670),
    .A2(_1472_),
    .A1(net771));
 sg13g2_inv_1 _3674_ (.Y(_0306_),
    .A(net772));
 sg13g2_a21o_1 _3675_ (.A2(_1472_),
    .A1(net1091),
    .B1(_1615_),
    .X(_0307_));
 sg13g2_nand2_2 _3676_ (.Y(_1272_),
    .A(net730),
    .B(net448));
 sg13g2_o21ai_1 _3677_ (.B1(net676),
    .Y(_1273_),
    .A1(net671),
    .A2(_1272_));
 sg13g2_a21oi_1 _3678_ (.A1(net753),
    .A2(_1272_),
    .Y(_0308_),
    .B1(_1273_));
 sg13g2_o21ai_1 _3679_ (.B1(net676),
    .Y(_1274_),
    .A1(net668),
    .A2(_1272_));
 sg13g2_a21oi_1 _3680_ (.A1(_1370_),
    .A2(_1272_),
    .Y(_0309_),
    .B1(_1274_));
 sg13g2_o21ai_1 _3681_ (.B1(net676),
    .Y(_1275_),
    .A1(net664),
    .A2(_1272_));
 sg13g2_a21oi_1 _3682_ (.A1(net807),
    .A2(_1272_),
    .Y(_0310_),
    .B1(_1275_));
 sg13g2_o21ai_1 _3683_ (.B1(net676),
    .Y(_1276_),
    .A1(net661),
    .A2(_1272_));
 sg13g2_a21oi_1 _3684_ (.A1(net482),
    .A2(_1272_),
    .Y(_0311_),
    .B1(_1276_));
 sg13g2_nand2_2 _3685_ (.Y(_1277_),
    .A(net420),
    .B(_1218_));
 sg13g2_o21ai_1 _3686_ (.B1(net677),
    .Y(_1278_),
    .A1(net671),
    .A2(net421));
 sg13g2_a21oi_1 _3687_ (.A1(_1367_),
    .A2(net421),
    .Y(_0312_),
    .B1(_1278_));
 sg13g2_o21ai_1 _3688_ (.B1(net677),
    .Y(_1279_),
    .A1(net669),
    .A2(net421));
 sg13g2_a21oi_1 _3689_ (.A1(_1366_),
    .A2(net421),
    .Y(_0313_),
    .B1(_1279_));
 sg13g2_o21ai_1 _3690_ (.B1(net677),
    .Y(_1280_),
    .A1(net664),
    .A2(net421));
 sg13g2_a21oi_1 _3691_ (.A1(_1365_),
    .A2(net421),
    .Y(_0314_),
    .B1(_1280_));
 sg13g2_o21ai_1 _3692_ (.B1(net677),
    .Y(_1281_),
    .A1(net663),
    .A2(net421));
 sg13g2_a21oi_1 _3693_ (.A1(_1364_),
    .A2(net421),
    .Y(_0315_),
    .B1(_1281_));
 sg13g2_nand2_2 _3694_ (.Y(_1282_),
    .A(net633),
    .B(net448));
 sg13g2_o21ai_1 _3695_ (.B1(net676),
    .Y(_1283_),
    .A1(net671),
    .A2(net449));
 sg13g2_a21oi_1 _3696_ (.A1(_1363_),
    .A2(net449),
    .Y(_0316_),
    .B1(_1283_));
 sg13g2_o21ai_1 _3697_ (.B1(net676),
    .Y(_1284_),
    .A1(net668),
    .A2(net449));
 sg13g2_a21oi_1 _3698_ (.A1(_1362_),
    .A2(net449),
    .Y(_0317_),
    .B1(_1284_));
 sg13g2_o21ai_1 _3699_ (.B1(net676),
    .Y(_1285_),
    .A1(net664),
    .A2(net449));
 sg13g2_a21oi_1 _3700_ (.A1(_1361_),
    .A2(net449),
    .Y(_0318_),
    .B1(_1285_));
 sg13g2_o21ai_1 _3701_ (.B1(net676),
    .Y(_1286_),
    .A1(net661),
    .A2(net449));
 sg13g2_a21oi_1 _3702_ (.A1(net751),
    .A2(net449),
    .Y(_0319_),
    .B1(_1286_));
 sg13g2_nand3_1 _3703_ (.B(net420),
    .C(net564),
    .A(net825),
    .Y(_1287_));
 sg13g2_o21ai_1 _3704_ (.B1(net680),
    .Y(_1288_),
    .A1(net673),
    .A2(_1287_));
 sg13g2_a21oi_1 _3705_ (.A1(net793),
    .A2(_1287_),
    .Y(_0320_),
    .B1(_1288_));
 sg13g2_o21ai_1 _3706_ (.B1(net680),
    .Y(_1289_),
    .A1(net668),
    .A2(_1287_));
 sg13g2_a21oi_1 _3707_ (.A1(net866),
    .A2(_1287_),
    .Y(_0321_),
    .B1(_1289_));
 sg13g2_o21ai_1 _3708_ (.B1(net680),
    .Y(_1290_),
    .A1(net665),
    .A2(_1287_));
 sg13g2_a21oi_1 _3709_ (.A1(net402),
    .A2(_1287_),
    .Y(_0322_),
    .B1(_1290_));
 sg13g2_o21ai_1 _3710_ (.B1(net681),
    .Y(_1291_),
    .A1(net661),
    .A2(_1287_));
 sg13g2_a21oi_1 _3711_ (.A1(_1356_),
    .A2(_1287_),
    .Y(_0323_),
    .B1(_1291_));
 sg13g2_nand2_2 _3712_ (.Y(_1292_),
    .A(net629),
    .B(_1517_));
 sg13g2_o21ai_1 _3713_ (.B1(net675),
    .Y(_1293_),
    .A1(net671),
    .A2(_1292_));
 sg13g2_a21oi_1 _3714_ (.A1(net470),
    .A2(_1292_),
    .Y(_0324_),
    .B1(_1293_));
 sg13g2_o21ai_1 _3715_ (.B1(net674),
    .Y(_1294_),
    .A1(net668),
    .A2(_1292_));
 sg13g2_a21oi_1 _3716_ (.A1(net348),
    .A2(_1292_),
    .Y(_0325_),
    .B1(_1294_));
 sg13g2_o21ai_1 _3717_ (.B1(net674),
    .Y(_1295_),
    .A1(net664),
    .A2(_1292_));
 sg13g2_a21oi_1 _3718_ (.A1(net405),
    .A2(_1292_),
    .Y(_0326_),
    .B1(_1295_));
 sg13g2_o21ai_1 _3719_ (.B1(net674),
    .Y(_1296_),
    .A1(net661),
    .A2(_1292_));
 sg13g2_a21oi_1 _3720_ (.A1(net357),
    .A2(_1292_),
    .Y(_0327_),
    .B1(_1296_));
 sg13g2_nand2_2 _3721_ (.Y(_1297_),
    .A(net420),
    .B(_1517_));
 sg13g2_o21ai_1 _3722_ (.B1(net675),
    .Y(_1298_),
    .A1(net671),
    .A2(_1297_));
 sg13g2_a21oi_1 _3723_ (.A1(net433),
    .A2(_1297_),
    .Y(_0328_),
    .B1(_1298_));
 sg13g2_o21ai_1 _3724_ (.B1(net675),
    .Y(_1299_),
    .A1(net668),
    .A2(_1297_));
 sg13g2_a21oi_1 _3725_ (.A1(net442),
    .A2(_1297_),
    .Y(_0329_),
    .B1(_1299_));
 sg13g2_o21ai_1 _3726_ (.B1(net674),
    .Y(_1300_),
    .A1(net664),
    .A2(_1297_));
 sg13g2_a21oi_1 _3727_ (.A1(net381),
    .A2(_1297_),
    .Y(_0330_),
    .B1(_1300_));
 sg13g2_o21ai_1 _3728_ (.B1(net674),
    .Y(_1301_),
    .A1(net661),
    .A2(_1297_));
 sg13g2_a21oi_1 _3729_ (.A1(net351),
    .A2(_1297_),
    .Y(_0331_),
    .B1(_1301_));
 sg13g2_nand2_2 _3730_ (.Y(_1302_),
    .A(net1065),
    .B(_1494_));
 sg13g2_o21ai_1 _3731_ (.B1(net674),
    .Y(_1303_),
    .A1(net671),
    .A2(_1302_));
 sg13g2_a21oi_1 _3732_ (.A1(net439),
    .A2(_1302_),
    .Y(_0332_),
    .B1(_1303_));
 sg13g2_o21ai_1 _3733_ (.B1(net674),
    .Y(_1304_),
    .A1(net668),
    .A2(_1302_));
 sg13g2_a21oi_1 _3734_ (.A1(net354),
    .A2(_1302_),
    .Y(_0333_),
    .B1(_1304_));
 sg13g2_o21ai_1 _3735_ (.B1(net674),
    .Y(_1305_),
    .A1(net664),
    .A2(_1302_));
 sg13g2_a21oi_1 _3736_ (.A1(net768),
    .A2(_1302_),
    .Y(_0334_),
    .B1(_1305_));
 sg13g2_o21ai_1 _3737_ (.B1(net675),
    .Y(_1306_),
    .A1(net661),
    .A2(_1302_));
 sg13g2_a21oi_1 _3738_ (.A1(net399),
    .A2(_1302_),
    .Y(_0335_),
    .B1(_1306_));
 sg13g2_nand3_1 _3739_ (.B(net420),
    .C(_1485_),
    .A(net825),
    .Y(_1307_));
 sg13g2_o21ai_1 _3740_ (.B1(net684),
    .Y(_1308_),
    .A1(net671),
    .A2(_1307_));
 sg13g2_a21oi_1 _3741_ (.A1(_1343_),
    .A2(_1307_),
    .Y(_0336_),
    .B1(_1308_));
 sg13g2_o21ai_1 _3742_ (.B1(net684),
    .Y(_1309_),
    .A1(net668),
    .A2(_1307_));
 sg13g2_a21oi_1 _3743_ (.A1(_1342_),
    .A2(_1307_),
    .Y(_0337_),
    .B1(_1309_));
 sg13g2_o21ai_1 _3744_ (.B1(net684),
    .Y(_1310_),
    .A1(net665),
    .A2(_1307_));
 sg13g2_a21oi_1 _3745_ (.A1(net396),
    .A2(_1307_),
    .Y(_0338_),
    .B1(_1310_));
 sg13g2_o21ai_1 _3746_ (.B1(net684),
    .Y(_1311_),
    .A1(net663),
    .A2(_1307_));
 sg13g2_a21oi_1 _3747_ (.A1(net822),
    .A2(_1307_),
    .Y(_0339_),
    .B1(_1311_));
 sg13g2_nand3_1 _3748_ (.B(net633),
    .C(_1485_),
    .A(net624),
    .Y(_1312_));
 sg13g2_o21ai_1 _3749_ (.B1(net691),
    .Y(_1313_),
    .A1(net672),
    .A2(_1312_));
 sg13g2_a21oi_1 _3750_ (.A1(net851),
    .A2(_1312_),
    .Y(_0340_),
    .B1(_1313_));
 sg13g2_o21ai_1 _3751_ (.B1(net691),
    .Y(_1314_),
    .A1(net5),
    .A2(_1312_));
 sg13g2_a21oi_1 _3752_ (.A1(net918),
    .A2(_1312_),
    .Y(_0341_),
    .B1(_1314_));
 sg13g2_o21ai_1 _3753_ (.B1(net691),
    .Y(_1315_),
    .A1(net666),
    .A2(_1312_));
 sg13g2_a21oi_1 _3754_ (.A1(net1069),
    .A2(_1312_),
    .Y(_0342_),
    .B1(_1315_));
 sg13g2_o21ai_1 _3755_ (.B1(net691),
    .Y(_1316_),
    .A1(net662),
    .A2(_1312_));
 sg13g2_a21oi_1 _3756_ (.A1(net869),
    .A2(_1312_),
    .Y(_0343_),
    .B1(_1316_));
 sg13g2_nand2_1 _3757_ (.Y(_1317_),
    .A(_0035_),
    .B(net545));
 sg13g2_o21ai_1 _3758_ (.B1(_1317_),
    .Y(_0344_),
    .A1(net606),
    .A2(net547));
 sg13g2_nand3_1 _3759_ (.B(_0440_),
    .C(net546),
    .A(_0436_),
    .Y(_1318_));
 sg13g2_o21ai_1 _3760_ (.B1(_1318_),
    .Y(_0345_),
    .A1(_0030_),
    .A2(net547));
 sg13g2_xnor2_1 _3761_ (.Y(_1319_),
    .A(_1433_),
    .B(_0355_));
 sg13g2_a21o_1 _3762_ (.A2(_1319_),
    .A1(net546),
    .B1(_1632_),
    .X(_0346_));
 sg13g2_and2_2 _3763_ (.A(net630),
    .B(_1465_),
    .X(_1320_));
 sg13g2_o21ai_1 _3764_ (.B1(net687),
    .Y(_1321_),
    .A1(net847),
    .A2(_1320_));
 sg13g2_a21oi_1 _3765_ (.A1(_1335_),
    .A2(_1320_),
    .Y(_0347_),
    .B1(net978));
 sg13g2_o21ai_1 _3766_ (.B1(net687),
    .Y(_1322_),
    .A1(net1028),
    .A2(_1320_));
 sg13g2_a21oi_1 _3767_ (.A1(_1334_),
    .A2(_1320_),
    .Y(_0348_),
    .B1(net1097));
 sg13g2_o21ai_1 _3768_ (.B1(net687),
    .Y(_1323_),
    .A1(net392),
    .A2(_1320_));
 sg13g2_a21oi_1 _3769_ (.A1(_1332_),
    .A2(_1320_),
    .Y(_0349_),
    .B1(net948));
 sg13g2_o21ai_1 _3770_ (.B1(net686),
    .Y(_1324_),
    .A1(net1019),
    .A2(_1320_));
 sg13g2_a21oi_1 _3771_ (.A1(_1330_),
    .A2(_1320_),
    .Y(_0350_),
    .B1(net1104));
 sg13g2_nand3_1 _3772_ (.B(net634),
    .C(_1211_),
    .A(net338),
    .Y(_1325_));
 sg13g2_o21ai_1 _3773_ (.B1(net688),
    .Y(_1326_),
    .A1(net670),
    .A2(net339));
 sg13g2_a21oi_1 _3774_ (.A1(_1333_),
    .A2(net339),
    .Y(_0351_),
    .B1(_1326_));
 sg13g2_o21ai_1 _3775_ (.B1(net688),
    .Y(_1327_),
    .A1(net666),
    .A2(net339));
 sg13g2_a21oi_1 _3776_ (.A1(_1331_),
    .A2(net339),
    .Y(_0352_),
    .B1(_1327_));
 sg13g2_o21ai_1 _3777_ (.B1(net688),
    .Y(_1328_),
    .A1(net663),
    .A2(net339));
 sg13g2_a21oi_1 _3778_ (.A1(net430),
    .A2(net339),
    .Y(_0353_),
    .B1(_1328_));
 sg13g2_dfrbp_1 _3779_ (.CLK(clk),
    .RESET_B(net8),
    .D(net1195),
    .Q_N(_1870_),
    .Q(\comm_ic0.spi0.curr_st[0] ));
 sg13g2_dfrbp_1 _3780_ (.CLK(clk),
    .RESET_B(net9),
    .D(net1136),
    .Q_N(_0026_),
    .Q(\comm_ic0.spi0.curr_st[1] ));
 sg13g2_dfrbp_1 _3781_ (.CLK(clk),
    .RESET_B(net10),
    .D(net1145),
    .Q_N(_1871_),
    .Q(\comm_ic0.spi0.curr_st[2] ));
 sg13g2_dfrbp_1 _3782_ (.CLK(clk),
    .RESET_B(net11),
    .D(net1108),
    .Q_N(_1872_),
    .Q(\comm_ic0.spi0.curr_st[3] ));
 sg13g2_dfrbp_1 _3783_ (.CLK(clk),
    .RESET_B(net12),
    .D(_0014_),
    .Q_N(_0073_),
    .Q(\comm_ic0.send_cnt[0] ));
 sg13g2_dfrbp_1 _3784_ (.CLK(clk),
    .RESET_B(net13),
    .D(net1171),
    .Q_N(_1873_),
    .Q(\comm_ic0.send_cnt[1] ));
 sg13g2_dfrbp_1 _3785_ (.CLK(clk),
    .RESET_B(net14),
    .D(_0016_),
    .Q_N(_1874_),
    .Q(\comm_ic0.send_cnt[2] ));
 sg13g2_dfrbp_1 _3786_ (.CLK(clk),
    .RESET_B(net15),
    .D(net1121),
    .Q_N(_1875_),
    .Q(\comm_ic0.send_cnt[3] ));
 sg13g2_dfrbp_1 _3787_ (.CLK(clk),
    .RESET_B(net16),
    .D(net1203),
    .Q_N(_1876_),
    .Q(\comm_ic0.curr_st[0] ));
 sg13g2_dfrbp_1 _3788_ (.CLK(clk),
    .RESET_B(net17),
    .D(net1220),
    .Q_N(_0032_),
    .Q(\comm_ic0.curr_st[1] ));
 sg13g2_dfrbp_1 _3789_ (.CLK(clk),
    .RESET_B(net39),
    .D(_0004_),
    .Q_N(_1877_),
    .Q(\comm_ic0.curr_st[2] ));
 sg13g2_dfrbp_1 _3790_ (.CLK(clk),
    .RESET_B(net7),
    .D(_0005_),
    .Q_N(_0071_),
    .Q(\comm_ic0.curr_st[3] ));
 sg13g2_dfrbp_1 _3791_ (.CLK(net617),
    .RESET_B(net49),
    .D(_0075_),
    .Q_N(_0028_),
    .Q(\comm_ic0.uart0.tx_st ));
 sg13g2_dfrbp_1 _3792_ (.CLK(clk),
    .RESET_B(net48),
    .D(net1050),
    .Q_N(_1869_),
    .Q(\comm_ic0.uart0.uclk_cnt[0] ));
 sg13g2_dfrbp_1 _3793_ (.CLK(clk),
    .RESET_B(net46),
    .D(net1015),
    .Q_N(_1868_),
    .Q(\comm_ic0.uart0.uclk_cnt[1] ));
 sg13g2_dfrbp_1 _3794_ (.CLK(clk),
    .RESET_B(net44),
    .D(net1018),
    .Q_N(_1867_),
    .Q(\comm_ic0.uart0.uclk_cnt[2] ));
 sg13g2_dfrbp_1 _3795_ (.CLK(clk),
    .RESET_B(net42),
    .D(net1053),
    .Q_N(_1866_),
    .Q(\comm_ic0.uart0.uclk_cnt[3] ));
 sg13g2_dfrbp_1 _3796_ (.CLK(clk),
    .RESET_B(net37),
    .D(net1012),
    .Q_N(_1865_),
    .Q(\comm_ic0.uart0.uclk_cnt[4] ));
 sg13g2_dfrbp_1 _3797_ (.CLK(clk),
    .RESET_B(net35),
    .D(net1086),
    .Q_N(_1864_),
    .Q(\comm_ic0.uart0.uclk_cnt[5] ));
 sg13g2_dfrbp_1 _3798_ (.CLK(clk),
    .RESET_B(net33),
    .D(net1152),
    .Q_N(_0037_),
    .Q(\comm_ic0.uart0.uclk_cnt[6] ));
 sg13g2_dfrbp_1 _3799_ (.CLK(clk),
    .RESET_B(net31),
    .D(net967),
    .Q_N(_1863_),
    .Q(\comm_ic0.uart0.uclk_cnt[7] ));
 sg13g2_dfrbp_1 _3800_ (.CLK(clk),
    .RESET_B(net29),
    .D(net322),
    .Q_N(_1862_),
    .Q(\comm_ic0.uart0.clk_cnt_reg[0] ));
 sg13g2_dfrbp_1 _3801_ (.CLK(clk),
    .RESET_B(net27),
    .D(net749),
    .Q_N(_1861_),
    .Q(\comm_ic0.uart0.clk_cnt_reg[1] ));
 sg13g2_dfrbp_1 _3802_ (.CLK(clk),
    .RESET_B(net25),
    .D(net468),
    .Q_N(_1860_),
    .Q(\comm_ic0.uart0.clk_cnt_reg[2] ));
 sg13g2_dfrbp_1 _3803_ (.CLK(clk),
    .RESET_B(net23),
    .D(net785),
    .Q_N(_1859_),
    .Q(\comm_ic0.uart0.clk_cnt_reg[3] ));
 sg13g2_dfrbp_1 _3804_ (.CLK(clk),
    .RESET_B(net21),
    .D(net782),
    .Q_N(_1858_),
    .Q(\comm_ic0.uart0.clk_cnt_reg[4] ));
 sg13g2_dfrbp_1 _3805_ (.CLK(clk),
    .RESET_B(net19),
    .D(net713),
    .Q_N(_1857_),
    .Q(\comm_ic0.uart0.clk_cnt_reg[5] ));
 sg13g2_dfrbp_1 _3806_ (.CLK(clk),
    .RESET_B(net6),
    .D(net458),
    .Q_N(_0038_),
    .Q(\comm_ic0.uart0.clk_cnt_reg[6] ));
 sg13g2_dfrbp_1 _3807_ (.CLK(clk),
    .RESET_B(net309),
    .D(net840),
    .Q_N(_1856_),
    .Q(\comm_ic0.uart0.clk_cnt_reg[7] ));
 sg13g2_dfrbp_1 _3808_ (.CLK(clk),
    .RESET_B(net307),
    .D(net1141),
    .Q_N(_1855_),
    .Q(\comm_ic0.uart0.clk_b ));
 sg13g2_dfrbp_1 _3809_ (.CLK(clk),
    .RESET_B(net305),
    .D(net803),
    .Q_N(_1854_),
    .Q(\comm_ic0.uart0.par_odd ));
 sg13g2_dfrbp_1 _3810_ (.CLK(clk),
    .RESET_B(net303),
    .D(net762),
    .Q_N(_0030_),
    .Q(\comm_ic0.uart0.par_en ));
 sg13g2_dfrbp_1 _3811_ (.CLK(net616),
    .RESET_B(net40),
    .D(_0095_),
    .Q_N(_1878_),
    .Q(\comm_ic0.UART_TX ));
 sg13g2_dfrbp_1 _3812_ (.CLK(net617),
    .RESET_B(net41),
    .D(_0024_),
    .Q_N(_1879_),
    .Q(\comm_ic0.uart0.rx_st[0] ));
 sg13g2_dfrbp_1 _3813_ (.CLK(net617),
    .RESET_B(net114),
    .D(_0001_),
    .Q_N(_0029_),
    .Q(\comm_ic0.uart0.rx_st[1] ));
 sg13g2_dfrbp_1 _3814_ (.CLK(net618),
    .RESET_B(net301),
    .D(_0025_),
    .Q_N(_1853_),
    .Q(\comm_ic0.uart0.rx_st[2] ));
 sg13g2_dfrbp_1 _3815_ (.CLK(net617),
    .RESET_B(net300),
    .D(_0096_),
    .Q_N(_0059_),
    .Q(\comm_ic0.uart0.tx_ind[2] ));
 sg13g2_dfrbp_1 _3816_ (.CLK(clk),
    .RESET_B(net299),
    .D(net1238),
    .Q_N(_1852_),
    .Q(\comm_ic0.spi0.sclk_cnt[0] ));
 sg13g2_dfrbp_1 _3817_ (.CLK(clk),
    .RESET_B(net298),
    .D(net1269),
    .Q_N(_1851_),
    .Q(\comm_ic0.spi0.sclk_cnt[1] ));
 sg13g2_dfrbp_1 _3818_ (.CLK(clk),
    .RESET_B(net297),
    .D(net1176),
    .Q_N(_0062_),
    .Q(\comm_ic0.spi0.sclk_cnt[2] ));
 sg13g2_dfrbp_1 _3819_ (.CLK(clk),
    .RESET_B(net296),
    .D(net1244),
    .Q_N(_1850_),
    .Q(\comm_ic0.spi0.sclk_cnt[3] ));
 sg13g2_dfrbp_1 _3820_ (.CLK(clk),
    .RESET_B(net295),
    .D(net1167),
    .Q_N(_0064_),
    .Q(\comm_ic0.spi0.sclk_cnt[4] ));
 sg13g2_dfrbp_1 _3821_ (.CLK(clk),
    .RESET_B(net294),
    .D(net1226),
    .Q_N(_1849_),
    .Q(\comm_ic0.spi0.sclk_cnt[5] ));
 sg13g2_dfrbp_1 _3822_ (.CLK(clk),
    .RESET_B(net293),
    .D(net1181),
    .Q_N(_1848_),
    .Q(\comm_ic0.spi0.sclk_cnt[6] ));
 sg13g2_dfrbp_1 _3823_ (.CLK(clk),
    .RESET_B(net292),
    .D(net1255),
    .Q_N(_1847_),
    .Q(\comm_ic0.spi0.sclk_cnt[7] ));
 sg13g2_dfrbp_1 _3824_ (.CLK(net616),
    .RESET_B(net291),
    .D(_0105_),
    .Q_N(_1846_),
    .Q(\comm_ic0.rx_new ));
 sg13g2_dfrbp_1 _3825_ (.CLK(net616),
    .RESET_B(net289),
    .D(_0106_),
    .Q_N(_1845_),
    .Q(\comm_ic0.rx_error ));
 sg13g2_dfrbp_1 _3826_ (.CLK(net618),
    .RESET_B(net287),
    .D(_0107_),
    .Q_N(_1844_),
    .Q(\comm_ic0.uart0.rx_data_reg[0] ));
 sg13g2_dfrbp_1 _3827_ (.CLK(net615),
    .RESET_B(net285),
    .D(_0108_),
    .Q_N(_1843_),
    .Q(\comm_ic0.uart0.rx_data_reg[1] ));
 sg13g2_dfrbp_1 _3828_ (.CLK(net615),
    .RESET_B(net283),
    .D(_0109_),
    .Q_N(_1842_),
    .Q(\comm_ic0.uart0.rx_data_reg[2] ));
 sg13g2_dfrbp_1 _3829_ (.CLK(net615),
    .RESET_B(net281),
    .D(_0110_),
    .Q_N(_1841_),
    .Q(\comm_ic0.uart0.rx_data_reg[3] ));
 sg13g2_dfrbp_1 _3830_ (.CLK(net615),
    .RESET_B(net279),
    .D(_0111_),
    .Q_N(_1840_),
    .Q(\comm_ic0.uart0.rx_data_reg[4] ));
 sg13g2_dfrbp_1 _3831_ (.CLK(net615),
    .RESET_B(net277),
    .D(_0112_),
    .Q_N(_1839_),
    .Q(\comm_ic0.uart0.rx_data_reg[5] ));
 sg13g2_dfrbp_1 _3832_ (.CLK(net615),
    .RESET_B(net275),
    .D(_0113_),
    .Q_N(_1838_),
    .Q(\comm_ic0.uart0.rx_data_reg[6] ));
 sg13g2_dfrbp_1 _3833_ (.CLK(net615),
    .RESET_B(net273),
    .D(_0114_),
    .Q_N(_1837_),
    .Q(\comm_ic0.uart0.rx_data_reg[7] ));
 sg13g2_dfrbp_1 _3834_ (.CLK(net618),
    .RESET_B(net271),
    .D(_0115_),
    .Q_N(_1836_),
    .Q(\comm_ic0.uart0.rx_data_reg[8] ));
 sg13g2_dfrbp_1 _3835_ (.CLK(net618),
    .RESET_B(net269),
    .D(_0116_),
    .Q_N(_1835_),
    .Q(\comm_ic0.uart0.rx_data_reg[9] ));
 sg13g2_dfrbp_1 _3836_ (.CLK(net618),
    .RESET_B(net267),
    .D(_0117_),
    .Q_N(_1834_),
    .Q(\comm_ic0.uart0.rx_data_reg[10] ));
 sg13g2_dfrbp_1 _3837_ (.CLK(net619),
    .RESET_B(net265),
    .D(_0118_),
    .Q_N(_0033_),
    .Q(\comm_ic0.uart0.rx_ind[0] ));
 sg13g2_dfrbp_1 _3838_ (.CLK(net618),
    .RESET_B(net263),
    .D(_0119_),
    .Q_N(_1833_),
    .Q(\comm_ic0.uart0.rx_ind[1] ));
 sg13g2_dfrbp_1 _3839_ (.CLK(net618),
    .RESET_B(net261),
    .D(_0120_),
    .Q_N(_0034_),
    .Q(\comm_ic0.uart0.rx_ind[2] ));
 sg13g2_dfrbp_1 _3840_ (.CLK(net618),
    .RESET_B(net259),
    .D(_0121_),
    .Q_N(_1832_),
    .Q(\comm_ic0.uart0.rx_ind[3] ));
 sg13g2_dfrbp_1 _3841_ (.CLK(net614),
    .RESET_B(net257),
    .D(_0122_),
    .Q_N(_1831_),
    .Q(\comm_ic0.rx_data[0] ));
 sg13g2_dfrbp_1 _3842_ (.CLK(net614),
    .RESET_B(net256),
    .D(_0123_),
    .Q_N(_1830_),
    .Q(\comm_ic0.rx_data[1] ));
 sg13g2_dfrbp_1 _3843_ (.CLK(net614),
    .RESET_B(net255),
    .D(_0124_),
    .Q_N(_1829_),
    .Q(\comm_ic0.rx_data[2] ));
 sg13g2_dfrbp_1 _3844_ (.CLK(net614),
    .RESET_B(net254),
    .D(_0125_),
    .Q_N(_1828_),
    .Q(\comm_ic0.rx_data[3] ));
 sg13g2_dfrbp_1 _3845_ (.CLK(net614),
    .RESET_B(net253),
    .D(_0126_),
    .Q_N(_1827_),
    .Q(\comm_ic0.rx_data[4] ));
 sg13g2_dfrbp_1 _3846_ (.CLK(net614),
    .RESET_B(net252),
    .D(_0127_),
    .Q_N(_1826_),
    .Q(\comm_ic0.rx_data[5] ));
 sg13g2_dfrbp_1 _3847_ (.CLK(net614),
    .RESET_B(net251),
    .D(_0128_),
    .Q_N(_1825_),
    .Q(\comm_ic0.rx_data[6] ));
 sg13g2_dfrbp_1 _3848_ (.CLK(net614),
    .RESET_B(net250),
    .D(_0129_),
    .Q_N(_1824_),
    .Q(\comm_ic0.rx_data[7] ));
 sg13g2_dfrbp_1 _3849_ (.CLK(net617),
    .RESET_B(net249),
    .D(_0130_),
    .Q_N(_1823_),
    .Q(\comm_ic0.busy_uart ));
 sg13g2_dfrbp_1 _3850_ (.CLK(net617),
    .RESET_B(net247),
    .D(_0131_),
    .Q_N(_1822_),
    .Q(\comm_ic0.uart0.tx_data_reg[0] ));
 sg13g2_dfrbp_1 _3851_ (.CLK(net613),
    .RESET_B(net245),
    .D(_0132_),
    .Q_N(_1821_),
    .Q(\comm_ic0.uart0.tx_data_reg[1] ));
 sg13g2_dfrbp_1 _3852_ (.CLK(net619),
    .RESET_B(net243),
    .D(_0133_),
    .Q_N(_1820_),
    .Q(\comm_ic0.uart0.tx_data_reg[2] ));
 sg13g2_dfrbp_1 _3853_ (.CLK(net613),
    .RESET_B(net241),
    .D(_0134_),
    .Q_N(_1819_),
    .Q(\comm_ic0.uart0.tx_data_reg[3] ));
 sg13g2_dfrbp_1 _3854_ (.CLK(net613),
    .RESET_B(net239),
    .D(_0135_),
    .Q_N(_1818_),
    .Q(\comm_ic0.uart0.tx_data_reg[4] ));
 sg13g2_dfrbp_1 _3855_ (.CLK(net619),
    .RESET_B(net237),
    .D(_0136_),
    .Q_N(_1817_),
    .Q(\comm_ic0.uart0.tx_data_reg[5] ));
 sg13g2_dfrbp_1 _3856_ (.CLK(net613),
    .RESET_B(net235),
    .D(_0137_),
    .Q_N(_1816_),
    .Q(\comm_ic0.uart0.tx_data_reg[6] ));
 sg13g2_dfrbp_1 _3857_ (.CLK(net613),
    .RESET_B(net233),
    .D(_0138_),
    .Q_N(_1815_),
    .Q(\comm_ic0.uart0.tx_data_reg[7] ));
 sg13g2_dfrbp_1 _3858_ (.CLK(net613),
    .RESET_B(net231),
    .D(_0139_),
    .Q_N(_1814_),
    .Q(\comm_ic0.uart0.tx_data_reg[8] ));
 sg13g2_dfrbp_1 _3859_ (.CLK(net620),
    .RESET_B(net229),
    .D(_0140_),
    .Q_N(_1813_),
    .Q(\comm_ic0.uart0.tx_data_reg[9] ));
 sg13g2_dfrbp_1 _3860_ (.CLK(clk),
    .RESET_B(net227),
    .D(net901),
    .Q_N(_0039_),
    .Q(\comm_ic0.i2c0.data_ind[0] ));
 sg13g2_dfrbp_1 _3861_ (.CLK(clk),
    .RESET_B(net225),
    .D(net1124),
    .Q_N(_1812_),
    .Q(\comm_ic0.i2c0.data_ind[1] ));
 sg13g2_dfrbp_1 _3862_ (.CLK(clk),
    .RESET_B(net223),
    .D(net1264),
    .Q_N(_1811_),
    .Q(\comm_ic0.i2c0.data_ind[2] ));
 sg13g2_dfrbp_1 _3863_ (.CLK(clk),
    .RESET_B(net221),
    .D(net1041),
    .Q_N(_1810_),
    .Q(\comm_ic0.i2c0.data_ind[3] ));
 sg13g2_dfrbp_1 _3864_ (.CLK(clk),
    .RESET_B(net219),
    .D(net722),
    .Q_N(_0040_),
    .Q(\comm_ic0.i2c0.addr_ind[0] ));
 sg13g2_dfrbp_1 _3865_ (.CLK(clk),
    .RESET_B(net217),
    .D(net1155),
    .Q_N(_1809_),
    .Q(\comm_ic0.i2c0.addr_ind[1] ));
 sg13g2_dfrbp_1 _3866_ (.CLK(clk),
    .RESET_B(net215),
    .D(net973),
    .Q_N(_0074_),
    .Q(\comm_ic0.i2c0.addr_ind[2] ));
 sg13g2_dfrbp_1 _3867_ (.CLK(clk),
    .RESET_B(net213),
    .D(net988),
    .Q_N(_1808_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _3868_ (.CLK(clk),
    .RESET_B(net212),
    .D(net1000),
    .Q_N(_1807_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _3869_ (.CLK(clk),
    .RESET_B(net211),
    .D(net1003),
    .Q_N(_1806_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _3870_ (.CLK(clk),
    .RESET_B(net210),
    .D(net935),
    .Q_N(_1805_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _3871_ (.CLK(clk),
    .RESET_B(net209),
    .D(net728),
    .Q_N(_1804_),
    .Q(\comm_ic0.i2c0.data_wr[0] ));
 sg13g2_dfrbp_1 _3872_ (.CLK(clk),
    .RESET_B(net207),
    .D(net385),
    .Q_N(_1803_),
    .Q(\comm_ic0.i2c0.data_wr[1] ));
 sg13g2_dfrbp_1 _3873_ (.CLK(clk),
    .RESET_B(net205),
    .D(net525),
    .Q_N(_1802_),
    .Q(\comm_ic0.i2c0.data_wr[2] ));
 sg13g2_dfrbp_1 _3874_ (.CLK(clk),
    .RESET_B(net203),
    .D(_0155_),
    .Q_N(_1801_),
    .Q(\comm_ic0.i2c0.data_wr[3] ));
 sg13g2_dfrbp_1 _3875_ (.CLK(clk),
    .RESET_B(net201),
    .D(_0156_),
    .Q_N(_1800_),
    .Q(\comm_ic0.i2c0.data_wr[4] ));
 sg13g2_dfrbp_1 _3876_ (.CLK(clk),
    .RESET_B(net199),
    .D(net704),
    .Q_N(_1799_),
    .Q(\comm_ic0.i2c0.data_wr[5] ));
 sg13g2_dfrbp_1 _3877_ (.CLK(clk),
    .RESET_B(net197),
    .D(_0158_),
    .Q_N(_1798_),
    .Q(\comm_ic0.i2c0.data_wr[6] ));
 sg13g2_dfrbp_1 _3878_ (.CLK(clk),
    .RESET_B(net195),
    .D(_0159_),
    .Q_N(_1797_),
    .Q(\comm_ic0.i2c0.data_wr[7] ));
 sg13g2_dfrbp_1 _3879_ (.CLK(clk),
    .RESET_B(net193),
    .D(net370),
    .Q_N(_1796_),
    .Q(\comm_ic0.i2c0.data_wr[8] ));
 sg13g2_dfrbp_1 _3880_ (.CLK(clk),
    .RESET_B(net191),
    .D(net376),
    .Q_N(_1795_),
    .Q(\comm_ic0.i2c0.data_wr[9] ));
 sg13g2_dfrbp_1 _3881_ (.CLK(clk),
    .RESET_B(net189),
    .D(net328),
    .Q_N(_1794_),
    .Q(\comm_ic0.i2c0.data_wr[10] ));
 sg13g2_dfrbp_1 _3882_ (.CLK(clk),
    .RESET_B(net187),
    .D(net488),
    .Q_N(_1793_),
    .Q(\comm_ic0.i2c0.data_wr[11] ));
 sg13g2_dfrbp_1 _3883_ (.CLK(clk),
    .RESET_B(net185),
    .D(net514),
    .Q_N(_1792_),
    .Q(\comm_ic0.i2c0.data_wr[12] ));
 sg13g2_dfrbp_1 _3884_ (.CLK(clk),
    .RESET_B(net183),
    .D(net346),
    .Q_N(_1791_),
    .Q(\comm_ic0.i2c0.data_wr[13] ));
 sg13g2_dfrbp_1 _3885_ (.CLK(clk),
    .RESET_B(net181),
    .D(net465),
    .Q_N(_1790_),
    .Q(\comm_ic0.i2c0.data_wr[14] ));
 sg13g2_dfrbp_1 _3886_ (.CLK(clk),
    .RESET_B(net115),
    .D(net412),
    .Q_N(_1880_),
    .Q(\comm_ic0.i2c0.data_wr[15] ));
 sg13g2_dfrbp_1 _3887_ (.CLK(clk),
    .RESET_B(net116),
    .D(net1075),
    .Q_N(_1881_),
    .Q(\comm_ic0.uart0.curr_st[0] ));
 sg13g2_dfrbp_1 _3888_ (.CLK(clk),
    .RESET_B(net154),
    .D(net1162),
    .Q_N(_1882_),
    .Q(\comm_ic0.uart0.curr_st[1] ));
 sg13g2_dfrbp_1 _3889_ (.CLK(clk),
    .RESET_B(net179),
    .D(net944),
    .Q_N(_1789_),
    .Q(\comm_ic0.uart0.curr_st[2] ));
 sg13g2_dfrbp_1 _3890_ (.CLK(clk),
    .RESET_B(net177),
    .D(net907),
    .Q_N(_1788_),
    .Q(\comm_ic0.SCL ));
 sg13g2_dfrbp_1 _3891_ (.CLK(clk),
    .RESET_B(net175),
    .D(net885),
    .Q_N(_1787_),
    .Q(\comm_ic0.SDA_op ));
 sg13g2_dfrbp_1 _3892_ (.CLK(clk),
    .RESET_B(net173),
    .D(net1059),
    .Q_N(_1786_),
    .Q(\comm_ic0.i2c0.data_out[0] ));
 sg13g2_dfrbp_1 _3893_ (.CLK(clk),
    .RESET_B(net171),
    .D(net843),
    .Q_N(_1785_),
    .Q(\comm_ic0.i2c0.data_out[1] ));
 sg13g2_dfrbp_1 _3894_ (.CLK(clk),
    .RESET_B(net169),
    .D(net800),
    .Q_N(_1784_),
    .Q(\comm_ic0.i2c0.data_out[2] ));
 sg13g2_dfrbp_1 _3895_ (.CLK(clk),
    .RESET_B(net167),
    .D(net955),
    .Q_N(_1783_),
    .Q(\comm_ic0.i2c0.data_out[3] ));
 sg13g2_dfrbp_1 _3896_ (.CLK(clk),
    .RESET_B(net165),
    .D(net379),
    .Q_N(_1782_),
    .Q(\comm_ic0.i2c0.data_out[4] ));
 sg13g2_dfrbp_1 _3897_ (.CLK(clk),
    .RESET_B(net163),
    .D(net698),
    .Q_N(_1781_),
    .Q(\comm_ic0.i2c0.data_out[5] ));
 sg13g2_dfrbp_1 _3898_ (.CLK(clk),
    .RESET_B(net153),
    .D(net743),
    .Q_N(_1780_),
    .Q(\comm_ic0.i2c0.data_out[6] ));
 sg13g2_dfrbp_1 _3899_ (.CLK(clk),
    .RESET_B(net151),
    .D(net816),
    .Q_N(_1779_),
    .Q(\comm_ic0.i2c0.data_out[7] ));
 sg13g2_dfrbp_1 _3900_ (.CLK(clk),
    .RESET_B(net149),
    .D(net367),
    .Q_N(_1778_),
    .Q(\comm_ic0.i2c0.data_out[8] ));
 sg13g2_dfrbp_1 _3901_ (.CLK(clk),
    .RESET_B(net147),
    .D(net766),
    .Q_N(_1777_),
    .Q(\comm_ic0.i2c0.data_out[9] ));
 sg13g2_dfrbp_1 _3902_ (.CLK(clk),
    .RESET_B(net145),
    .D(net788),
    .Q_N(_1776_),
    .Q(\comm_ic0.i2c0.data_out[10] ));
 sg13g2_dfrbp_1 _3903_ (.CLK(clk),
    .RESET_B(net143),
    .D(net813),
    .Q_N(_1775_),
    .Q(\comm_ic0.i2c0.data_out[11] ));
 sg13g2_dfrbp_1 _3904_ (.CLK(clk),
    .RESET_B(net141),
    .D(net716),
    .Q_N(_1774_),
    .Q(\comm_ic0.i2c0.data_out[12] ));
 sg13g2_dfrbp_1 _3905_ (.CLK(clk),
    .RESET_B(net139),
    .D(net737),
    .Q_N(_1773_),
    .Q(\comm_ic0.i2c0.data_out[13] ));
 sg13g2_dfrbp_1 _3906_ (.CLK(clk),
    .RESET_B(net137),
    .D(net725),
    .Q_N(_1772_),
    .Q(\comm_ic0.i2c0.data_out[14] ));
 sg13g2_dfrbp_1 _3907_ (.CLK(clk),
    .RESET_B(net135),
    .D(net734),
    .Q_N(_1771_),
    .Q(\comm_ic0.i2c0.data_out[15] ));
 sg13g2_dfrbp_1 _3908_ (.CLK(clk),
    .RESET_B(net133),
    .D(net1006),
    .Q_N(_1770_),
    .Q(\comm_ic0.busy_i2c ));
 sg13g2_dfrbp_1 _3909_ (.CLK(clk),
    .RESET_B(net131),
    .D(net922),
    .Q_N(_1769_),
    .Q(\comm_ic0.error_i2c ));
 sg13g2_dfrbp_1 _3910_ (.CLK(clk),
    .RESET_B(net129),
    .D(net316),
    .Q_N(_1768_),
    .Q(\comm_ic0.SDA_op_en ));
 sg13g2_dfrbp_1 _3911_ (.CLK(clk),
    .RESET_B(net127),
    .D(net1056),
    .Q_N(_1767_),
    .Q(\comm_ic0.i2c0.clk_cnt_reg[0] ));
 sg13g2_dfrbp_1 _3912_ (.CLK(clk),
    .RESET_B(net125),
    .D(net1064),
    .Q_N(_1766_),
    .Q(\comm_ic0.i2c0.clk_cnt_reg[1] ));
 sg13g2_dfrbp_1 _3913_ (.CLK(clk),
    .RESET_B(net123),
    .D(net859),
    .Q_N(_1765_),
    .Q(\comm_ic0.i2c0.clk_cnt_reg[2] ));
 sg13g2_dfrbp_1 _3914_ (.CLK(clk),
    .RESET_B(net121),
    .D(net1027),
    .Q_N(_1764_),
    .Q(\comm_ic0.i2c0.clk_cnt_reg[3] ));
 sg13g2_dfrbp_1 _3915_ (.CLK(clk),
    .RESET_B(net119),
    .D(net849),
    .Q_N(_1763_),
    .Q(\comm_ic0.i2c0.clk_cnt_reg[4] ));
 sg13g2_dfrbp_1 _3916_ (.CLK(clk),
    .RESET_B(net117),
    .D(net1030),
    .Q_N(_1762_),
    .Q(\comm_ic0.i2c0.clk_cnt_reg[5] ));
 sg13g2_dfrbp_1 _3917_ (.CLK(clk),
    .RESET_B(net112),
    .D(net394),
    .Q_N(_1761_),
    .Q(\comm_ic0.i2c0.clk_cnt_reg[6] ));
 sg13g2_dfrbp_1 _3918_ (.CLK(clk),
    .RESET_B(net110),
    .D(net1021),
    .Q_N(_1760_),
    .Q(\comm_ic0.i2c0.clk_cnt_reg[7] ));
 sg13g2_dfrbp_1 _3919_ (.CLK(clk),
    .RESET_B(net108),
    .D(net454),
    .Q_N(_1759_),
    .Q(\comm_ic0.i2c0.addr_wr[0] ));
 sg13g2_dfrbp_1 _3920_ (.CLK(clk),
    .RESET_B(net106),
    .D(net425),
    .Q_N(_1758_),
    .Q(\comm_ic0.i2c0.addr_wr[1] ));
 sg13g2_dfrbp_1 _3921_ (.CLK(clk),
    .RESET_B(net104),
    .D(net334),
    .Q_N(_1757_),
    .Q(\comm_ic0.i2c0.addr_wr[2] ));
 sg13g2_dfrbp_1 _3922_ (.CLK(clk),
    .RESET_B(net102),
    .D(net707),
    .Q_N(_1756_),
    .Q(\comm_ic0.i2c0.addr_wr[3] ));
 sg13g2_dfrbp_1 _3923_ (.CLK(clk),
    .RESET_B(net100),
    .D(net415),
    .Q_N(_1755_),
    .Q(\comm_ic0.i2c0.addr_wr[4] ));
 sg13g2_dfrbp_1 _3924_ (.CLK(clk),
    .RESET_B(net98),
    .D(net506),
    .Q_N(_1754_),
    .Q(\comm_ic0.i2c0.addr_wr[5] ));
 sg13g2_dfrbp_1 _3925_ (.CLK(clk),
    .RESET_B(net96),
    .D(net710),
    .Q_N(_1753_),
    .Q(\comm_ic0.i2c0.addr_wr[6] ));
 sg13g2_dfrbp_1 _3926_ (.CLK(clk),
    .RESET_B(net155),
    .D(net428),
    .Q_N(_1883_),
    .Q(\comm_ic0.i2c0.addr_wr[7] ));
 sg13g2_dfrbp_1 _3927_ (.CLK(clk),
    .RESET_B(net156),
    .D(net1192),
    .Q_N(_1884_),
    .Q(\comm_ic0.i2c0.curr_st[0] ));
 sg13g2_dfrbp_1 _3928_ (.CLK(clk),
    .RESET_B(net157),
    .D(net388),
    .Q_N(_0027_),
    .Q(\comm_ic0.i2c0.curr_st[1] ));
 sg13g2_dfrbp_1 _3929_ (.CLK(clk),
    .RESET_B(net158),
    .D(net1047),
    .Q_N(_1885_),
    .Q(\comm_ic0.i2c0.curr_st[2] ));
 sg13g2_dfrbp_1 _3930_ (.CLK(clk),
    .RESET_B(net159),
    .D(net1073),
    .Q_N(_1886_),
    .Q(\comm_ic0.i2c0.curr_st[3] ));
 sg13g2_dfrbp_1 _3931_ (.CLK(clk),
    .RESET_B(net160),
    .D(net1083),
    .Q_N(_1887_),
    .Q(\comm_ic0.i2c0.curr_st[4] ));
 sg13g2_dfrbp_1 _3932_ (.CLK(clk),
    .RESET_B(net161),
    .D(net1133),
    .Q_N(_0031_),
    .Q(\comm_ic0.i2c0.curr_st[5] ));
 sg13g2_dfrbp_1 _3933_ (.CLK(clk),
    .RESET_B(net172),
    .D(net916),
    .Q_N(_1888_),
    .Q(\comm_ic0.i2c0.curr_st[6] ));
 sg13g2_dfrbp_1 _3934_ (.CLK(clk),
    .RESET_B(net94),
    .D(net833),
    .Q_N(_1752_),
    .Q(\comm_ic0.i2c0.curr_st[7] ));
 sg13g2_dfrbp_1 _3935_ (.CLK(clk),
    .RESET_B(net92),
    .D(net759),
    .Q_N(_1751_),
    .Q(\comm_ic0.SEN ));
 sg13g2_dfrbp_1 _3936_ (.CLK(clk),
    .RESET_B(net90),
    .D(net1033),
    .Q_N(_1750_),
    .Q(\comm_ic0.SCLK ));
 sg13g2_dfrbp_1 _3937_ (.CLK(clk),
    .RESET_B(net88),
    .D(net779),
    .Q_N(_1749_),
    .Q(\comm_ic0.MOSI ));
 sg13g2_dfrbp_1 _3938_ (.CLK(clk),
    .RESET_B(net86),
    .D(net791),
    .Q_N(_0041_),
    .Q(\comm_ic0.spi0.data_out[0] ));
 sg13g2_dfrbp_1 _3939_ (.CLK(clk),
    .RESET_B(net84),
    .D(net1024),
    .Q_N(_0044_),
    .Q(\comm_ic0.spi0.data_out[1] ));
 sg13g2_dfrbp_1 _3940_ (.CLK(clk),
    .RESET_B(net82),
    .D(net897),
    .Q_N(_0045_),
    .Q(\comm_ic0.spi0.data_out[2] ));
 sg13g2_dfrbp_1 _3941_ (.CLK(clk),
    .RESET_B(net80),
    .D(net888),
    .Q_N(_0046_),
    .Q(\comm_ic0.spi0.data_out[3] ));
 sg13g2_dfrbp_1 _3942_ (.CLK(clk),
    .RESET_B(net78),
    .D(net497),
    .Q_N(_0047_),
    .Q(\comm_ic0.spi0.data_out[4] ));
 sg13g2_dfrbp_1 _3943_ (.CLK(clk),
    .RESET_B(net76),
    .D(net876),
    .Q_N(_0048_),
    .Q(\comm_ic0.spi0.data_out[5] ));
 sg13g2_dfrbp_1 _3944_ (.CLK(clk),
    .RESET_B(net74),
    .D(net719),
    .Q_N(_0049_),
    .Q(\comm_ic0.spi0.data_out[6] ));
 sg13g2_dfrbp_1 _3945_ (.CLK(clk),
    .RESET_B(net72),
    .D(net1090),
    .Q_N(_0050_),
    .Q(\comm_ic0.spi0.data_out[7] ));
 sg13g2_dfrbp_1 _3946_ (.CLK(clk),
    .RESET_B(net70),
    .D(net518),
    .Q_N(_0051_),
    .Q(\comm_ic0.spi0.data_out[8] ));
 sg13g2_dfrbp_1 _3947_ (.CLK(clk),
    .RESET_B(net68),
    .D(net862),
    .Q_N(_0052_),
    .Q(\comm_ic0.spi0.data_out[9] ));
 sg13g2_dfrbp_1 _3948_ (.CLK(clk),
    .RESET_B(net66),
    .D(net891),
    .Q_N(_0053_),
    .Q(\comm_ic0.spi0.data_out[10] ));
 sg13g2_dfrbp_1 _3949_ (.CLK(clk),
    .RESET_B(net64),
    .D(net879),
    .Q_N(_0054_),
    .Q(\comm_ic0.spi0.data_out[11] ));
 sg13g2_dfrbp_1 _3950_ (.CLK(clk),
    .RESET_B(net62),
    .D(net797),
    .Q_N(_0055_),
    .Q(\comm_ic0.spi0.data_out[12] ));
 sg13g2_dfrbp_1 _3951_ (.CLK(clk),
    .RESET_B(net60),
    .D(net926),
    .Q_N(_0056_),
    .Q(\comm_ic0.spi0.data_out[13] ));
 sg13g2_dfrbp_1 _3952_ (.CLK(clk),
    .RESET_B(net58),
    .D(net873),
    .Q_N(_0057_),
    .Q(\comm_ic0.spi0.data_out[14] ));
 sg13g2_dfrbp_1 _3953_ (.CLK(clk),
    .RESET_B(net56),
    .D(net959),
    .Q_N(_0058_),
    .Q(\comm_ic0.spi0.data_out[15] ));
 sg13g2_dfrbp_1 _3954_ (.CLK(clk),
    .RESET_B(net54),
    .D(net976),
    .Q_N(_1748_),
    .Q(\comm_ic0.busy_spi ));
 sg13g2_dfrbp_1 _3955_ (.CLK(clk),
    .RESET_B(net52),
    .D(net964),
    .Q_N(_1747_),
    .Q(\comm_ic0.spi0.clk_cnt_reg[0] ));
 sg13g2_dfrbp_1 _3956_ (.CLK(clk),
    .RESET_B(net50),
    .D(net932),
    .Q_N(_1746_),
    .Q(\comm_ic0.spi0.clk_cnt_reg[1] ));
 sg13g2_dfrbp_1 _3957_ (.CLK(clk),
    .RESET_B(net45),
    .D(net882),
    .Q_N(_1745_),
    .Q(\comm_ic0.spi0.clk_cnt_reg[2] ));
 sg13g2_dfrbp_1 _3958_ (.CLK(clk),
    .RESET_B(net38),
    .D(net994),
    .Q_N(_1744_),
    .Q(\comm_ic0.spi0.clk_cnt_reg[3] ));
 sg13g2_dfrbp_1 _3959_ (.CLK(clk),
    .RESET_B(net34),
    .D(net830),
    .Q_N(_1743_),
    .Q(\comm_ic0.spi0.clk_cnt_reg[4] ));
 sg13g2_dfrbp_1 _3960_ (.CLK(clk),
    .RESET_B(net30),
    .D(net913),
    .Q_N(_1742_),
    .Q(\comm_ic0.spi0.clk_cnt_reg[5] ));
 sg13g2_dfrbp_1 _3961_ (.CLK(clk),
    .RESET_B(net26),
    .D(net746),
    .Q_N(_1741_),
    .Q(\comm_ic0.spi0.clk_cnt_reg[6] ));
 sg13g2_dfrbp_1 _3962_ (.CLK(clk),
    .RESET_B(net22),
    .D(net480),
    .Q_N(_1740_),
    .Q(\comm_ic0.spi0.clk_cnt_reg[7] ));
 sg13g2_dfrbp_1 _3963_ (.CLK(clk),
    .RESET_B(net18),
    .D(net343),
    .Q_N(_1739_),
    .Q(\comm_ic0.spi0.data_wr[0] ));
 sg13g2_dfrbp_1 _3964_ (.CLK(clk),
    .RESET_B(net308),
    .D(net418),
    .Q_N(_1738_),
    .Q(\comm_ic0.spi0.data_wr[1] ));
 sg13g2_dfrbp_1 _3965_ (.CLK(clk),
    .RESET_B(net304),
    .D(net337),
    .Q_N(_1737_),
    .Q(\comm_ic0.spi0.data_wr[2] ));
 sg13g2_dfrbp_1 _3966_ (.CLK(clk),
    .RESET_B(net290),
    .D(net409),
    .Q_N(_1736_),
    .Q(\comm_ic0.spi0.data_wr[3] ));
 sg13g2_dfrbp_1 _3967_ (.CLK(clk),
    .RESET_B(net286),
    .D(net491),
    .Q_N(_1735_),
    .Q(\comm_ic0.spi0.data_wr[4] ));
 sg13g2_dfrbp_1 _3968_ (.CLK(clk),
    .RESET_B(net282),
    .D(net474),
    .Q_N(_1734_),
    .Q(\comm_ic0.spi0.data_wr[5] ));
 sg13g2_dfrbp_1 _3969_ (.CLK(clk),
    .RESET_B(net278),
    .D(net810),
    .Q_N(_1733_),
    .Q(\comm_ic0.spi0.data_wr[6] ));
 sg13g2_dfrbp_1 _3970_ (.CLK(clk),
    .RESET_B(net274),
    .D(net503),
    .Q_N(_1732_),
    .Q(\comm_ic0.spi0.data_wr[7] ));
 sg13g2_dfrbp_1 _3971_ (.CLK(clk),
    .RESET_B(net270),
    .D(net437),
    .Q_N(_1731_),
    .Q(\comm_ic0.spi0.data_wr[8] ));
 sg13g2_dfrbp_1 _3972_ (.CLK(clk),
    .RESET_B(net266),
    .D(net319),
    .Q_N(_1730_),
    .Q(\comm_ic0.spi0.data_wr[9] ));
 sg13g2_dfrbp_1 _3973_ (.CLK(clk),
    .RESET_B(net262),
    .D(net331),
    .Q_N(_1729_),
    .Q(\comm_ic0.spi0.data_wr[10] ));
 sg13g2_dfrbp_1 _3974_ (.CLK(clk),
    .RESET_B(net258),
    .D(net494),
    .Q_N(_1728_),
    .Q(\comm_ic0.spi0.data_wr[11] ));
 sg13g2_dfrbp_1 _3975_ (.CLK(clk),
    .RESET_B(net246),
    .D(net325),
    .Q_N(_1727_),
    .Q(\comm_ic0.spi0.data_wr[12] ));
 sg13g2_dfrbp_1 _3976_ (.CLK(clk),
    .RESET_B(net242),
    .D(net361),
    .Q_N(_1726_),
    .Q(\comm_ic0.spi0.data_wr[13] ));
 sg13g2_dfrbp_1 _3977_ (.CLK(clk),
    .RESET_B(net238),
    .D(net373),
    .Q_N(_1725_),
    .Q(\comm_ic0.spi0.data_wr[14] ));
 sg13g2_dfrbp_1 _3978_ (.CLK(clk),
    .RESET_B(net234),
    .D(net364),
    .Q_N(_1724_),
    .Q(\comm_ic0.spi0.data_wr[15] ));
 sg13g2_dfrbp_1 _3979_ (.CLK(clk),
    .RESET_B(net230),
    .D(net1212),
    .Q_N(_0042_),
    .Q(\comm_ic0.spi0.data_ind[0] ));
 sg13g2_dfrbp_1 _3980_ (.CLK(clk),
    .RESET_B(net226),
    .D(net910),
    .Q_N(_1723_),
    .Q(\comm_ic0.spi0.data_ind[1] ));
 sg13g2_dfrbp_1 _3981_ (.CLK(clk),
    .RESET_B(net222),
    .D(net1189),
    .Q_N(_1722_),
    .Q(\comm_ic0.spi0.data_ind[2] ));
 sg13g2_dfrbp_1 _3982_ (.CLK(clk),
    .RESET_B(net218),
    .D(net1148),
    .Q_N(_0043_),
    .Q(\comm_ic0.spi0.data_ind[3] ));
 sg13g2_dfrbp_1 _3983_ (.CLK(clk),
    .RESET_B(net214),
    .D(net701),
    .Q_N(_1721_),
    .Q(\comm_ic0.spi0.CPOL ));
 sg13g2_dfrbp_1 _3984_ (.CLK(clk),
    .RESET_B(net206),
    .D(net776),
    .Q_N(_1720_),
    .Q(\comm_ic0.spi0.CPHA ));
 sg13g2_dfrbp_1 _3985_ (.CLK(clk),
    .RESET_B(net202),
    .D(net1233),
    .Q_N(_1719_),
    .Q(\comm_ic0.i2c0.scl_cnt[0] ));
 sg13g2_dfrbp_1 _3986_ (.CLK(clk),
    .RESET_B(net200),
    .D(net1274),
    .Q_N(_1718_),
    .Q(\comm_ic0.i2c0.scl_cnt[1] ));
 sg13g2_dfrbp_1 _3987_ (.CLK(clk),
    .RESET_B(net198),
    .D(net1208),
    .Q_N(_0067_),
    .Q(\comm_ic0.i2c0.scl_cnt[2] ));
 sg13g2_dfrbp_1 _3988_ (.CLK(clk),
    .RESET_B(net196),
    .D(net1250),
    .Q_N(_1717_),
    .Q(\comm_ic0.i2c0.scl_cnt[3] ));
 sg13g2_dfrbp_1 _3989_ (.CLK(clk),
    .RESET_B(net194),
    .D(net1201),
    .Q_N(_0069_),
    .Q(\comm_ic0.i2c0.scl_cnt[4] ));
 sg13g2_dfrbp_1 _3990_ (.CLK(clk),
    .RESET_B(net192),
    .D(net1260),
    .Q_N(_1716_),
    .Q(\comm_ic0.i2c0.scl_cnt[5] ));
 sg13g2_dfrbp_1 _3991_ (.CLK(clk),
    .RESET_B(net190),
    .D(net1159),
    .Q_N(_1715_),
    .Q(\comm_ic0.i2c0.scl_cnt[6] ));
 sg13g2_dfrbp_1 _3992_ (.CLK(clk),
    .RESET_B(net188),
    .D(net1216),
    .Q_N(_1714_),
    .Q(\comm_ic0.i2c0.scl_cnt[7] ));
 sg13g2_dfrbp_1 _3993_ (.CLK(clk),
    .RESET_B(net186),
    .D(_0263_),
    .Q_N(_0072_),
    .Q(\comm_ic0.i2c_addr_en ));
 sg13g2_dfrbp_1 _3994_ (.CLK(clk),
    .RESET_B(net182),
    .D(_0264_),
    .Q_N(_1713_),
    .Q(\comm_ic0.i2c0.clk_cnt[0] ));
 sg13g2_dfrbp_1 _3995_ (.CLK(clk),
    .RESET_B(net178),
    .D(net1127),
    .Q_N(_1712_),
    .Q(\comm_ic0.i2c0.clk_cnt[1] ));
 sg13g2_dfrbp_1 _3996_ (.CLK(clk),
    .RESET_B(net174),
    .D(net1044),
    .Q_N(_0066_),
    .Q(\comm_ic0.i2c0.clk_cnt[2] ));
 sg13g2_dfrbp_1 _3997_ (.CLK(clk),
    .RESET_B(net170),
    .D(net1095),
    .Q_N(_1711_),
    .Q(\comm_ic0.i2c0.clk_cnt[3] ));
 sg13g2_dfrbp_1 _3998_ (.CLK(clk),
    .RESET_B(net166),
    .D(net485),
    .Q_N(_1710_),
    .Q(\comm_ic0.i2c0.address[3] ));
 sg13g2_dfrbp_1 _3999_ (.CLK(clk),
    .RESET_B(net162),
    .D(net500),
    .Q_N(_1709_),
    .Q(\comm_ic0.i2c0.address[4] ));
 sg13g2_dfrbp_1 _4000_ (.CLK(clk),
    .RESET_B(net150),
    .D(net756),
    .Q_N(_1708_),
    .Q(\comm_ic0.i2c0.address[5] ));
 sg13g2_dfrbp_1 _4001_ (.CLK(clk),
    .RESET_B(net146),
    .D(net391),
    .Q_N(_1707_),
    .Q(\comm_ic0.i2c0.address[6] ));
 sg13g2_dfrbp_1 _4002_ (.CLK(clk),
    .RESET_B(net142),
    .D(net522),
    .Q_N(_1706_),
    .Q(\comm_ic0.i2c0.write_n ));
 sg13g2_dfrbp_1 _4003_ (.CLK(clk),
    .RESET_B(net138),
    .D(net477),
    .Q_N(_1705_),
    .Q(\comm_ic0.i2c0.data_in[12] ));
 sg13g2_dfrbp_1 _4004_ (.CLK(clk),
    .RESET_B(net134),
    .D(_0274_),
    .Q_N(_1704_),
    .Q(\comm_ic0.i2c0.data_in[13] ));
 sg13g2_dfrbp_1 _4005_ (.CLK(clk),
    .RESET_B(net130),
    .D(net462),
    .Q_N(_1703_),
    .Q(\comm_ic0.i2c0.data_in[14] ));
 sg13g2_dfrbp_1 _4006_ (.CLK(clk),
    .RESET_B(net126),
    .D(net446),
    .Q_N(_1702_),
    .Q(\comm_ic0.i2c0.data_in[15] ));
 sg13g2_dfrbp_1 _4007_ (.CLK(clk),
    .RESET_B(net122),
    .D(net1229),
    .Q_N(_1701_),
    .Q(\comm_ic0.i2c0.start ));
 sg13g2_dfrbp_1 _4008_ (.CLK(clk),
    .RESET_B(net118),
    .D(net740),
    .Q_N(_1700_),
    .Q(\comm_ic0.i2c0.bits16 ));
 sg13g2_dfrbp_1 _4009_ (.CLK(clk),
    .RESET_B(net111),
    .D(net1061),
    .Q_N(_1699_),
    .Q(\comm_ic0.spi0.clk_cnt[0] ));
 sg13g2_dfrbp_1 _4010_ (.CLK(clk),
    .RESET_B(net107),
    .D(net946),
    .Q_N(_1698_),
    .Q(\comm_ic0.spi0.clk_cnt[1] ));
 sg13g2_dfrbp_1 _4011_ (.CLK(clk),
    .RESET_B(net103),
    .D(net846),
    .Q_N(_0061_),
    .Q(\comm_ic0.spi0.clk_cnt[2] ));
 sg13g2_dfrbp_1 _4012_ (.CLK(clk),
    .RESET_B(net99),
    .D(net985),
    .Q_N(_1697_),
    .Q(\comm_ic0.spi0.clk_cnt[3] ));
 sg13g2_dfrbp_1 _4013_ (.CLK(clk),
    .RESET_B(net95),
    .D(net991),
    .Q_N(_1696_),
    .Q(\comm_ic0.spi0.mode[0] ));
 sg13g2_dfrbp_1 _4014_ (.CLK(clk),
    .RESET_B(net91),
    .D(net952),
    .Q_N(_1695_),
    .Q(\comm_ic0.spi0.mode[1] ));
 sg13g2_dfrbp_1 _4015_ (.CLK(clk),
    .RESET_B(net87),
    .D(net1067),
    .Q_N(_1694_),
    .Q(\comm_ic0.spi0.start ));
 sg13g2_dfrbp_1 _4016_ (.CLK(clk),
    .RESET_B(net83),
    .D(net1078),
    .Q_N(_1693_),
    .Q(\comm_ic0.spi0.data_in[12] ));
 sg13g2_dfrbp_1 _4017_ (.CLK(clk),
    .RESET_B(net79),
    .D(net1009),
    .Q_N(_1692_),
    .Q(\comm_ic0.spi0.data_in[13] ));
 sg13g2_dfrbp_1 _4018_ (.CLK(clk),
    .RESET_B(net75),
    .D(net970),
    .Q_N(_1691_),
    .Q(\comm_ic0.spi0.data_in[14] ));
 sg13g2_dfrbp_1 _4019_ (.CLK(clk),
    .RESET_B(net71),
    .D(net997),
    .Q_N(_1690_),
    .Q(\comm_ic0.spi0.data_in[15] ));
 sg13g2_dfrbp_1 _4020_ (.CLK(clk),
    .RESET_B(net67),
    .D(net1111),
    .Q_N(_1689_),
    .Q(\comm_ic0.spi0.bits16 ));
 sg13g2_dfrbp_1 _4021_ (.CLK(clk),
    .RESET_B(net63),
    .D(net1037),
    .Q_N(_1688_),
    .Q(\comm_ic0.uart0.setting ));
 sg13g2_dfrbp_1 _4022_ (.CLK(clk),
    .RESET_B(net59),
    .D(net1102),
    .Q_N(_1687_),
    .Q(\comm_ic0.uart0.enable ));
 sg13g2_dfrbp_1 _4023_ (.CLK(clk),
    .RESET_B(net55),
    .D(_0293_),
    .Q_N(_1686_),
    .Q(\comm_ic0.uart0.clk_cnt[0] ));
 sg13g2_dfrbp_1 _4024_ (.CLK(clk),
    .RESET_B(net51),
    .D(_0294_),
    .Q_N(_1685_),
    .Q(\comm_ic0.uart0.clk_cnt[1] ));
 sg13g2_dfrbp_1 _4025_ (.CLK(clk),
    .RESET_B(net43),
    .D(net827),
    .Q_N(_1684_),
    .Q(\comm_ic0.uart0.clk_cnt[2] ));
 sg13g2_dfrbp_1 _4026_ (.CLK(clk),
    .RESET_B(net32),
    .D(net961),
    .Q_N(_1683_),
    .Q(\comm_ic0.uart0.clk_cnt[3] ));
 sg13g2_dfrbp_1 _4027_ (.CLK(clk),
    .RESET_B(net24),
    .D(net929),
    .Q_N(_1682_),
    .Q(\comm_ic0.tx_data[4] ));
 sg13g2_dfrbp_1 _4028_ (.CLK(clk),
    .RESET_B(net310),
    .D(net904),
    .Q_N(_1681_),
    .Q(\comm_ic0.tx_data[5] ));
 sg13g2_dfrbp_1 _4029_ (.CLK(clk),
    .RESET_B(net302),
    .D(net894),
    .Q_N(_1680_),
    .Q(\comm_ic0.tx_data[6] ));
 sg13g2_dfrbp_1 _4030_ (.CLK(clk),
    .RESET_B(net284),
    .D(net982),
    .Q_N(_1679_),
    .Q(\comm_ic0.tx_data[7] ));
 sg13g2_dfrbp_1 _4031_ (.CLK(clk),
    .RESET_B(net276),
    .D(_0301_),
    .Q_N(_1678_),
    .Q(\comm_ic0.tx_new ));
 sg13g2_dfrbp_1 _4032_ (.CLK(clk),
    .RESET_B(net268),
    .D(net938),
    .Q_N(_1677_),
    .Q(\comm_ic0.parity_odd ));
 sg13g2_dfrbp_1 _4033_ (.CLK(clk),
    .RESET_B(net260),
    .D(net941),
    .Q_N(_1676_),
    .Q(\comm_ic0.parity_en ));
 sg13g2_dfrbp_1 _4034_ (.CLK(clk),
    .RESET_B(net244),
    .D(net509),
    .Q_N(_1675_),
    .Q(\comm_ic0.rx_ack ));
 sg13g2_dfrbp_1 _4035_ (.CLK(clk),
    .RESET_B(net236),
    .D(_0305_),
    .Q_N(_1674_),
    .Q(\comm_ic0.comm_sel[0] ));
 sg13g2_dfrbp_1 _4036_ (.CLK(clk),
    .RESET_B(net228),
    .D(net773),
    .Q_N(_1673_),
    .Q(\comm_ic0.comm_sel[1] ));
 sg13g2_dfrbp_1 _4037_ (.CLK(clk),
    .RESET_B(net220),
    .D(net1092),
    .Q_N(_1672_),
    .Q(uio_oe[5]));
 sg13g2_dfrbp_1 _4038_ (.CLK(clk),
    .RESET_B(net208),
    .D(net754),
    .Q_N(_1671_),
    .Q(\comm_ic0.i2c0.data_in[4] ));
 sg13g2_dfrbp_1 _4039_ (.CLK(clk),
    .RESET_B(net184),
    .D(net731),
    .Q_N(_1670_),
    .Q(\comm_ic0.i2c0.data_in[5] ));
 sg13g2_dfrbp_1 _4040_ (.CLK(clk),
    .RESET_B(net176),
    .D(_0310_),
    .Q_N(_1669_),
    .Q(\comm_ic0.i2c0.data_in[6] ));
 sg13g2_dfrbp_1 _4041_ (.CLK(clk),
    .RESET_B(net168),
    .D(net483),
    .Q_N(_1668_),
    .Q(\comm_ic0.i2c0.data_in[7] ));
 sg13g2_dfrbp_1 _4042_ (.CLK(clk),
    .RESET_B(net152),
    .D(net422),
    .Q_N(_1667_),
    .Q(\comm_ic0.i2c0.data_in[8] ));
 sg13g2_dfrbp_1 _4043_ (.CLK(clk),
    .RESET_B(net144),
    .D(_0313_),
    .Q_N(_1666_),
    .Q(\comm_ic0.i2c0.data_in[9] ));
 sg13g2_dfrbp_1 _4044_ (.CLK(clk),
    .RESET_B(net136),
    .D(_0314_),
    .Q_N(_1665_),
    .Q(\comm_ic0.i2c0.data_in[10] ));
 sg13g2_dfrbp_1 _4045_ (.CLK(clk),
    .RESET_B(net128),
    .D(_0315_),
    .Q_N(_1664_),
    .Q(\comm_ic0.i2c0.data_in[11] ));
 sg13g2_dfrbp_1 _4046_ (.CLK(clk),
    .RESET_B(net120),
    .D(_0316_),
    .Q_N(_1663_),
    .Q(\comm_ic0.i2c0.data_in[0] ));
 sg13g2_dfrbp_1 _4047_ (.CLK(clk),
    .RESET_B(net109),
    .D(net450),
    .Q_N(_1662_),
    .Q(\comm_ic0.i2c0.data_in[1] ));
 sg13g2_dfrbp_1 _4048_ (.CLK(clk),
    .RESET_B(net101),
    .D(_0318_),
    .Q_N(_1661_),
    .Q(\comm_ic0.i2c0.data_in[2] ));
 sg13g2_dfrbp_1 _4049_ (.CLK(clk),
    .RESET_B(net93),
    .D(_0319_),
    .Q_N(_1660_),
    .Q(\comm_ic0.i2c0.data_in[3] ));
 sg13g2_dfrbp_1 _4050_ (.CLK(clk),
    .RESET_B(net85),
    .D(net794),
    .Q_N(_0063_),
    .Q(\comm_ic0.spi0.clk_cnt[4] ));
 sg13g2_dfrbp_1 _4051_ (.CLK(clk),
    .RESET_B(net77),
    .D(net867),
    .Q_N(_1659_),
    .Q(\comm_ic0.spi0.clk_cnt[5] ));
 sg13g2_dfrbp_1 _4052_ (.CLK(clk),
    .RESET_B(net69),
    .D(net403),
    .Q_N(_0065_),
    .Q(\comm_ic0.spi0.clk_cnt[6] ));
 sg13g2_dfrbp_1 _4053_ (.CLK(clk),
    .RESET_B(net61),
    .D(net835),
    .Q_N(_1658_),
    .Q(\comm_ic0.spi0.clk_cnt[7] ));
 sg13g2_dfrbp_1 _4054_ (.CLK(clk),
    .RESET_B(net53),
    .D(net471),
    .Q_N(_1657_),
    .Q(\comm_ic0.spi0.data_in[4] ));
 sg13g2_dfrbp_1 _4055_ (.CLK(clk),
    .RESET_B(net36),
    .D(net349),
    .Q_N(_1656_),
    .Q(\comm_ic0.spi0.data_in[5] ));
 sg13g2_dfrbp_1 _4056_ (.CLK(clk),
    .RESET_B(net20),
    .D(net406),
    .Q_N(_1655_),
    .Q(\comm_ic0.spi0.data_in[6] ));
 sg13g2_dfrbp_1 _4057_ (.CLK(clk),
    .RESET_B(net288),
    .D(net358),
    .Q_N(_1654_),
    .Q(\comm_ic0.spi0.data_in[7] ));
 sg13g2_dfrbp_1 _4058_ (.CLK(clk),
    .RESET_B(net272),
    .D(net434),
    .Q_N(_1653_),
    .Q(\comm_ic0.spi0.data_in[8] ));
 sg13g2_dfrbp_1 _4059_ (.CLK(clk),
    .RESET_B(net248),
    .D(net443),
    .Q_N(_1652_),
    .Q(\comm_ic0.spi0.data_in[9] ));
 sg13g2_dfrbp_1 _4060_ (.CLK(clk),
    .RESET_B(net232),
    .D(net382),
    .Q_N(_1651_),
    .Q(\comm_ic0.spi0.data_in[10] ));
 sg13g2_dfrbp_1 _4061_ (.CLK(clk),
    .RESET_B(net216),
    .D(net352),
    .Q_N(_1650_),
    .Q(\comm_ic0.spi0.data_in[11] ));
 sg13g2_dfrbp_1 _4062_ (.CLK(clk),
    .RESET_B(net180),
    .D(net440),
    .Q_N(_1649_),
    .Q(\comm_ic0.spi0.data_in[0] ));
 sg13g2_dfrbp_1 _4063_ (.CLK(clk),
    .RESET_B(net164),
    .D(net355),
    .Q_N(_1648_),
    .Q(\comm_ic0.spi0.data_in[1] ));
 sg13g2_dfrbp_1 _4064_ (.CLK(clk),
    .RESET_B(net140),
    .D(net769),
    .Q_N(_1647_),
    .Q(\comm_ic0.spi0.data_in[2] ));
 sg13g2_dfrbp_1 _4065_ (.CLK(clk),
    .RESET_B(net124),
    .D(net400),
    .Q_N(_1646_),
    .Q(\comm_ic0.spi0.data_in[3] ));
 sg13g2_dfrbp_1 _4066_ (.CLK(clk),
    .RESET_B(net105),
    .D(net837),
    .Q_N(_1645_),
    .Q(\comm_ic0.uart0.clk_cnt[4] ));
 sg13g2_dfrbp_1 _4067_ (.CLK(clk),
    .RESET_B(net89),
    .D(net854),
    .Q_N(_1644_),
    .Q(\comm_ic0.uart0.clk_cnt[5] ));
 sg13g2_dfrbp_1 _4068_ (.CLK(clk),
    .RESET_B(net73),
    .D(net397),
    .Q_N(_0036_),
    .Q(\comm_ic0.uart0.clk_cnt[6] ));
 sg13g2_dfrbp_1 _4069_ (.CLK(clk),
    .RESET_B(net57),
    .D(net823),
    .Q_N(_1643_),
    .Q(\comm_ic0.uart0.clk_cnt[7] ));
 sg13g2_dfrbp_1 _4070_ (.CLK(clk),
    .RESET_B(net28),
    .D(net852),
    .Q_N(_1642_),
    .Q(\comm_ic0.tx_data[0] ));
 sg13g2_dfrbp_1 _4071_ (.CLK(clk),
    .RESET_B(net280),
    .D(net919),
    .Q_N(_1641_),
    .Q(\comm_ic0.tx_data[1] ));
 sg13g2_dfrbp_1 _4072_ (.CLK(clk),
    .RESET_B(net240),
    .D(net1070),
    .Q_N(_1640_),
    .Q(\comm_ic0.tx_data[2] ));
 sg13g2_dfrbp_1 _4073_ (.CLK(clk),
    .RESET_B(net204),
    .D(net870),
    .Q_N(_1639_),
    .Q(\comm_ic0.tx_data[3] ));
 sg13g2_dfrbp_1 _4074_ (.CLK(net613),
    .RESET_B(net148),
    .D(_0344_),
    .Q_N(_0035_),
    .Q(\comm_ic0.uart0.tx_ind[0] ));
 sg13g2_dfrbp_1 _4075_ (.CLK(net617),
    .RESET_B(net132),
    .D(_0345_),
    .Q_N(_0060_),
    .Q(\comm_ic0.uart0.tx_ind[1] ));
 sg13g2_dfrbp_1 _4076_ (.CLK(net617),
    .RESET_B(net113),
    .D(_0346_),
    .Q_N(_1638_),
    .Q(\comm_ic0.uart0.tx_ind[3] ));
 sg13g2_dfrbp_1 _4077_ (.CLK(clk),
    .RESET_B(net97),
    .D(net979),
    .Q_N(_0068_),
    .Q(\comm_ic0.i2c0.clk_cnt[4] ));
 sg13g2_dfrbp_1 _4078_ (.CLK(clk),
    .RESET_B(net65),
    .D(net1098),
    .Q_N(_1637_),
    .Q(\comm_ic0.i2c0.clk_cnt[5] ));
 sg13g2_dfrbp_1 _4079_ (.CLK(clk),
    .RESET_B(net306),
    .D(net949),
    .Q_N(_0070_),
    .Q(\comm_ic0.i2c0.clk_cnt[6] ));
 sg13g2_dfrbp_1 _4080_ (.CLK(clk),
    .RESET_B(net224),
    .D(net1105),
    .Q_N(_1636_),
    .Q(\comm_ic0.i2c0.clk_cnt[7] ));
 sg13g2_dfrbp_1 _4081_ (.CLK(clk),
    .RESET_B(net81),
    .D(net511),
    .Q_N(_1635_),
    .Q(\comm_ic0.i2c0.address[0] ));
 sg13g2_dfrbp_1 _4082_ (.CLK(clk),
    .RESET_B(net264),
    .D(net340),
    .Q_N(_1634_),
    .Q(\comm_ic0.i2c0.address[1] ));
 sg13g2_dfrbp_1 _4083_ (.CLK(clk),
    .RESET_B(net47),
    .D(net431),
    .Q_N(_1633_),
    .Q(\comm_ic0.i2c0.address[2] ));
 sg13g2_tiehi _3790__7 (.L_HI(net7));
 sg13g2_tiehi _3779__8 (.L_HI(net8));
 sg13g2_tiehi _3780__9 (.L_HI(net9));
 sg13g2_tiehi _3781__10 (.L_HI(net10));
 sg13g2_tiehi _3782__11 (.L_HI(net11));
 sg13g2_tiehi _3783__12 (.L_HI(net12));
 sg13g2_tiehi _3784__13 (.L_HI(net13));
 sg13g2_tiehi _3785__14 (.L_HI(net14));
 sg13g2_tiehi _3786__15 (.L_HI(net15));
 sg13g2_tiehi _3787__16 (.L_HI(net16));
 sg13g2_tiehi _3788__17 (.L_HI(net17));
 sg13g2_tiehi _3963__18 (.L_HI(net18));
 sg13g2_tiehi _3805__19 (.L_HI(net19));
 sg13g2_tiehi _4056__20 (.L_HI(net20));
 sg13g2_tiehi _3804__21 (.L_HI(net21));
 sg13g2_tiehi _3962__22 (.L_HI(net22));
 sg13g2_tiehi _3803__23 (.L_HI(net23));
 sg13g2_tiehi _4027__24 (.L_HI(net24));
 sg13g2_tiehi _3802__25 (.L_HI(net25));
 sg13g2_tiehi _3961__26 (.L_HI(net26));
 sg13g2_tiehi _3801__27 (.L_HI(net27));
 sg13g2_tiehi _4070__28 (.L_HI(net28));
 sg13g2_tiehi _3800__29 (.L_HI(net29));
 sg13g2_tiehi _3960__30 (.L_HI(net30));
 sg13g2_tiehi _3799__31 (.L_HI(net31));
 sg13g2_tiehi _4026__32 (.L_HI(net32));
 sg13g2_tiehi _3798__33 (.L_HI(net33));
 sg13g2_tiehi _3959__34 (.L_HI(net34));
 sg13g2_tiehi _3797__35 (.L_HI(net35));
 sg13g2_tiehi _4055__36 (.L_HI(net36));
 sg13g2_tiehi _3796__37 (.L_HI(net37));
 sg13g2_tiehi _3958__38 (.L_HI(net38));
 sg13g2_tiehi _3789__39 (.L_HI(net39));
 sg13g2_tiehi _3811__40 (.L_HI(net40));
 sg13g2_tiehi _3812__41 (.L_HI(net41));
 sg13g2_tiehi _3795__42 (.L_HI(net42));
 sg13g2_tiehi _4025__43 (.L_HI(net43));
 sg13g2_tiehi _3794__44 (.L_HI(net44));
 sg13g2_tiehi _3957__45 (.L_HI(net45));
 sg13g2_tiehi _3793__46 (.L_HI(net46));
 sg13g2_tiehi _4083__47 (.L_HI(net47));
 sg13g2_tiehi _3792__48 (.L_HI(net48));
 sg13g2_tiehi _3791__49 (.L_HI(net49));
 sg13g2_tiehi _3956__50 (.L_HI(net50));
 sg13g2_tiehi _4024__51 (.L_HI(net51));
 sg13g2_tiehi _3955__52 (.L_HI(net52));
 sg13g2_tiehi _4054__53 (.L_HI(net53));
 sg13g2_tiehi _3954__54 (.L_HI(net54));
 sg13g2_tiehi _4023__55 (.L_HI(net55));
 sg13g2_tiehi _3953__56 (.L_HI(net56));
 sg13g2_tiehi _4069__57 (.L_HI(net57));
 sg13g2_tiehi _3952__58 (.L_HI(net58));
 sg13g2_tiehi _4022__59 (.L_HI(net59));
 sg13g2_tiehi _3951__60 (.L_HI(net60));
 sg13g2_tiehi _4053__61 (.L_HI(net61));
 sg13g2_tiehi _3950__62 (.L_HI(net62));
 sg13g2_tiehi _4021__63 (.L_HI(net63));
 sg13g2_tiehi _3949__64 (.L_HI(net64));
 sg13g2_tiehi _4078__65 (.L_HI(net65));
 sg13g2_tiehi _3948__66 (.L_HI(net66));
 sg13g2_tiehi _4020__67 (.L_HI(net67));
 sg13g2_tiehi _3947__68 (.L_HI(net68));
 sg13g2_tiehi _4052__69 (.L_HI(net69));
 sg13g2_tiehi _3946__70 (.L_HI(net70));
 sg13g2_tiehi _4019__71 (.L_HI(net71));
 sg13g2_tiehi _3945__72 (.L_HI(net72));
 sg13g2_tiehi _4068__73 (.L_HI(net73));
 sg13g2_tiehi _3944__74 (.L_HI(net74));
 sg13g2_tiehi _4018__75 (.L_HI(net75));
 sg13g2_tiehi _3943__76 (.L_HI(net76));
 sg13g2_tiehi _4051__77 (.L_HI(net77));
 sg13g2_tiehi _3942__78 (.L_HI(net78));
 sg13g2_tiehi _4017__79 (.L_HI(net79));
 sg13g2_tiehi _3941__80 (.L_HI(net80));
 sg13g2_tiehi _4081__81 (.L_HI(net81));
 sg13g2_tiehi _3940__82 (.L_HI(net82));
 sg13g2_tiehi _4016__83 (.L_HI(net83));
 sg13g2_tiehi _3939__84 (.L_HI(net84));
 sg13g2_tiehi _4050__85 (.L_HI(net85));
 sg13g2_tiehi _3938__86 (.L_HI(net86));
 sg13g2_tiehi _4015__87 (.L_HI(net87));
 sg13g2_tiehi _3937__88 (.L_HI(net88));
 sg13g2_tiehi _4067__89 (.L_HI(net89));
 sg13g2_tiehi _3936__90 (.L_HI(net90));
 sg13g2_tiehi _4014__91 (.L_HI(net91));
 sg13g2_tiehi _3935__92 (.L_HI(net92));
 sg13g2_tiehi _4049__93 (.L_HI(net93));
 sg13g2_tiehi _3934__94 (.L_HI(net94));
 sg13g2_tiehi _4013__95 (.L_HI(net95));
 sg13g2_tiehi _3925__96 (.L_HI(net96));
 sg13g2_tiehi _4077__97 (.L_HI(net97));
 sg13g2_tiehi _3924__98 (.L_HI(net98));
 sg13g2_tiehi _4012__99 (.L_HI(net99));
 sg13g2_tiehi _3923__100 (.L_HI(net100));
 sg13g2_tiehi _4048__101 (.L_HI(net101));
 sg13g2_tiehi _3922__102 (.L_HI(net102));
 sg13g2_tiehi _4011__103 (.L_HI(net103));
 sg13g2_tiehi _3921__104 (.L_HI(net104));
 sg13g2_tiehi _4066__105 (.L_HI(net105));
 sg13g2_tiehi _3920__106 (.L_HI(net106));
 sg13g2_tiehi _4010__107 (.L_HI(net107));
 sg13g2_tiehi _3919__108 (.L_HI(net108));
 sg13g2_tiehi _4047__109 (.L_HI(net109));
 sg13g2_tiehi _3918__110 (.L_HI(net110));
 sg13g2_tiehi _4009__111 (.L_HI(net111));
 sg13g2_tiehi _3917__112 (.L_HI(net112));
 sg13g2_tiehi _4076__113 (.L_HI(net113));
 sg13g2_tiehi _3813__114 (.L_HI(net114));
 sg13g2_tiehi _3886__115 (.L_HI(net115));
 sg13g2_tiehi _3887__116 (.L_HI(net116));
 sg13g2_tiehi _3916__117 (.L_HI(net117));
 sg13g2_tiehi _4008__118 (.L_HI(net118));
 sg13g2_tiehi _3915__119 (.L_HI(net119));
 sg13g2_tiehi _4046__120 (.L_HI(net120));
 sg13g2_tiehi _3914__121 (.L_HI(net121));
 sg13g2_tiehi _4007__122 (.L_HI(net122));
 sg13g2_tiehi _3913__123 (.L_HI(net123));
 sg13g2_tiehi _4065__124 (.L_HI(net124));
 sg13g2_tiehi _3912__125 (.L_HI(net125));
 sg13g2_tiehi _4006__126 (.L_HI(net126));
 sg13g2_tiehi _3911__127 (.L_HI(net127));
 sg13g2_tiehi _4045__128 (.L_HI(net128));
 sg13g2_tiehi _3910__129 (.L_HI(net129));
 sg13g2_tiehi _4005__130 (.L_HI(net130));
 sg13g2_tiehi _3909__131 (.L_HI(net131));
 sg13g2_tiehi _4075__132 (.L_HI(net132));
 sg13g2_tiehi _3908__133 (.L_HI(net133));
 sg13g2_tiehi _4004__134 (.L_HI(net134));
 sg13g2_tiehi _3907__135 (.L_HI(net135));
 sg13g2_tiehi _4044__136 (.L_HI(net136));
 sg13g2_tiehi _3906__137 (.L_HI(net137));
 sg13g2_tiehi _4003__138 (.L_HI(net138));
 sg13g2_tiehi _3905__139 (.L_HI(net139));
 sg13g2_tiehi _4064__140 (.L_HI(net140));
 sg13g2_tiehi _3904__141 (.L_HI(net141));
 sg13g2_tiehi _4002__142 (.L_HI(net142));
 sg13g2_tiehi _3903__143 (.L_HI(net143));
 sg13g2_tiehi _4043__144 (.L_HI(net144));
 sg13g2_tiehi _3902__145 (.L_HI(net145));
 sg13g2_tiehi _4001__146 (.L_HI(net146));
 sg13g2_tiehi _3901__147 (.L_HI(net147));
 sg13g2_tiehi _4074__148 (.L_HI(net148));
 sg13g2_tiehi _3900__149 (.L_HI(net149));
 sg13g2_tiehi _4000__150 (.L_HI(net150));
 sg13g2_tiehi _3899__151 (.L_HI(net151));
 sg13g2_tiehi _4042__152 (.L_HI(net152));
 sg13g2_tiehi _3898__153 (.L_HI(net153));
 sg13g2_tiehi _3888__154 (.L_HI(net154));
 sg13g2_tiehi _3926__155 (.L_HI(net155));
 sg13g2_tiehi _3927__156 (.L_HI(net156));
 sg13g2_tiehi _3928__157 (.L_HI(net157));
 sg13g2_tiehi _3929__158 (.L_HI(net158));
 sg13g2_tiehi _3930__159 (.L_HI(net159));
 sg13g2_tiehi _3931__160 (.L_HI(net160));
 sg13g2_tiehi _3932__161 (.L_HI(net161));
 sg13g2_tiehi _3999__162 (.L_HI(net162));
 sg13g2_tiehi _3897__163 (.L_HI(net163));
 sg13g2_tiehi _4063__164 (.L_HI(net164));
 sg13g2_tiehi _3896__165 (.L_HI(net165));
 sg13g2_tiehi _3998__166 (.L_HI(net166));
 sg13g2_tiehi _3895__167 (.L_HI(net167));
 sg13g2_tiehi _4041__168 (.L_HI(net168));
 sg13g2_tiehi _3894__169 (.L_HI(net169));
 sg13g2_tiehi _3997__170 (.L_HI(net170));
 sg13g2_tiehi _3893__171 (.L_HI(net171));
 sg13g2_tiehi _3933__172 (.L_HI(net172));
 sg13g2_tiehi _3892__173 (.L_HI(net173));
 sg13g2_tiehi _3996__174 (.L_HI(net174));
 sg13g2_tiehi _3891__175 (.L_HI(net175));
 sg13g2_tiehi _4040__176 (.L_HI(net176));
 sg13g2_tiehi _3890__177 (.L_HI(net177));
 sg13g2_tiehi _3995__178 (.L_HI(net178));
 sg13g2_tiehi _3889__179 (.L_HI(net179));
 sg13g2_tiehi _4062__180 (.L_HI(net180));
 sg13g2_tiehi _3885__181 (.L_HI(net181));
 sg13g2_tiehi _3994__182 (.L_HI(net182));
 sg13g2_tiehi _3884__183 (.L_HI(net183));
 sg13g2_tiehi _4039__184 (.L_HI(net184));
 sg13g2_tiehi _3883__185 (.L_HI(net185));
 sg13g2_tiehi _3993__186 (.L_HI(net186));
 sg13g2_tiehi _3882__187 (.L_HI(net187));
 sg13g2_tiehi _3992__188 (.L_HI(net188));
 sg13g2_tiehi _3881__189 (.L_HI(net189));
 sg13g2_tiehi _3991__190 (.L_HI(net190));
 sg13g2_tiehi _3880__191 (.L_HI(net191));
 sg13g2_tiehi _3990__192 (.L_HI(net192));
 sg13g2_tiehi _3879__193 (.L_HI(net193));
 sg13g2_tiehi _3989__194 (.L_HI(net194));
 sg13g2_tiehi _3878__195 (.L_HI(net195));
 sg13g2_tiehi _3988__196 (.L_HI(net196));
 sg13g2_tiehi _3877__197 (.L_HI(net197));
 sg13g2_tiehi _3987__198 (.L_HI(net198));
 sg13g2_tiehi _3876__199 (.L_HI(net199));
 sg13g2_tiehi _3986__200 (.L_HI(net200));
 sg13g2_tiehi _3875__201 (.L_HI(net201));
 sg13g2_tiehi _3985__202 (.L_HI(net202));
 sg13g2_tiehi _3874__203 (.L_HI(net203));
 sg13g2_tiehi _4073__204 (.L_HI(net204));
 sg13g2_tiehi _3873__205 (.L_HI(net205));
 sg13g2_tiehi _3984__206 (.L_HI(net206));
 sg13g2_tiehi _3872__207 (.L_HI(net207));
 sg13g2_tiehi _4038__208 (.L_HI(net208));
 sg13g2_tiehi _3871__209 (.L_HI(net209));
 sg13g2_tiehi _3870__210 (.L_HI(net210));
 sg13g2_tiehi _3869__211 (.L_HI(net211));
 sg13g2_tiehi _3868__212 (.L_HI(net212));
 sg13g2_tiehi _3867__213 (.L_HI(net213));
 sg13g2_tiehi _3983__214 (.L_HI(net214));
 sg13g2_tiehi _3866__215 (.L_HI(net215));
 sg13g2_tiehi _4061__216 (.L_HI(net216));
 sg13g2_tiehi _3865__217 (.L_HI(net217));
 sg13g2_tiehi _3982__218 (.L_HI(net218));
 sg13g2_tiehi _3864__219 (.L_HI(net219));
 sg13g2_tiehi _4037__220 (.L_HI(net220));
 sg13g2_tiehi _3863__221 (.L_HI(net221));
 sg13g2_tiehi _3981__222 (.L_HI(net222));
 sg13g2_tiehi _3862__223 (.L_HI(net223));
 sg13g2_tiehi _4080__224 (.L_HI(net224));
 sg13g2_tiehi _3861__225 (.L_HI(net225));
 sg13g2_tiehi _3980__226 (.L_HI(net226));
 sg13g2_tiehi _3860__227 (.L_HI(net227));
 sg13g2_tiehi _4036__228 (.L_HI(net228));
 sg13g2_tiehi _3859__229 (.L_HI(net229));
 sg13g2_tiehi _3979__230 (.L_HI(net230));
 sg13g2_tiehi _3858__231 (.L_HI(net231));
 sg13g2_tiehi _4060__232 (.L_HI(net232));
 sg13g2_tiehi _3857__233 (.L_HI(net233));
 sg13g2_tiehi _3978__234 (.L_HI(net234));
 sg13g2_tiehi _3856__235 (.L_HI(net235));
 sg13g2_tiehi _4035__236 (.L_HI(net236));
 sg13g2_tiehi _3855__237 (.L_HI(net237));
 sg13g2_tiehi _3977__238 (.L_HI(net238));
 sg13g2_tiehi _3854__239 (.L_HI(net239));
 sg13g2_tiehi _4072__240 (.L_HI(net240));
 sg13g2_tiehi _3853__241 (.L_HI(net241));
 sg13g2_tiehi _3976__242 (.L_HI(net242));
 sg13g2_tiehi _3852__243 (.L_HI(net243));
 sg13g2_tiehi _4034__244 (.L_HI(net244));
 sg13g2_tiehi _3851__245 (.L_HI(net245));
 sg13g2_tiehi _3975__246 (.L_HI(net246));
 sg13g2_tiehi _3850__247 (.L_HI(net247));
 sg13g2_tiehi _4059__248 (.L_HI(net248));
 sg13g2_tiehi _3849__249 (.L_HI(net249));
 sg13g2_tiehi _3848__250 (.L_HI(net250));
 sg13g2_tiehi _3847__251 (.L_HI(net251));
 sg13g2_tiehi _3846__252 (.L_HI(net252));
 sg13g2_tiehi _3845__253 (.L_HI(net253));
 sg13g2_tiehi _3844__254 (.L_HI(net254));
 sg13g2_tiehi _3843__255 (.L_HI(net255));
 sg13g2_tiehi _3842__256 (.L_HI(net256));
 sg13g2_tiehi _3841__257 (.L_HI(net257));
 sg13g2_tiehi _3974__258 (.L_HI(net258));
 sg13g2_tiehi _3840__259 (.L_HI(net259));
 sg13g2_tiehi _4033__260 (.L_HI(net260));
 sg13g2_tiehi _3839__261 (.L_HI(net261));
 sg13g2_tiehi _3973__262 (.L_HI(net262));
 sg13g2_tiehi _3838__263 (.L_HI(net263));
 sg13g2_tiehi _4082__264 (.L_HI(net264));
 sg13g2_tiehi _3837__265 (.L_HI(net265));
 sg13g2_tiehi _3972__266 (.L_HI(net266));
 sg13g2_tiehi _3836__267 (.L_HI(net267));
 sg13g2_tiehi _4032__268 (.L_HI(net268));
 sg13g2_tiehi _3835__269 (.L_HI(net269));
 sg13g2_tiehi _3971__270 (.L_HI(net270));
 sg13g2_tiehi _3834__271 (.L_HI(net271));
 sg13g2_tiehi _4058__272 (.L_HI(net272));
 sg13g2_tiehi _3833__273 (.L_HI(net273));
 sg13g2_tiehi _3970__274 (.L_HI(net274));
 sg13g2_tiehi _3832__275 (.L_HI(net275));
 sg13g2_tiehi _4031__276 (.L_HI(net276));
 sg13g2_tiehi _3831__277 (.L_HI(net277));
 sg13g2_tiehi _3969__278 (.L_HI(net278));
 sg13g2_tiehi _3830__279 (.L_HI(net279));
 sg13g2_tiehi _4071__280 (.L_HI(net280));
 sg13g2_tiehi _3829__281 (.L_HI(net281));
 sg13g2_tiehi _3968__282 (.L_HI(net282));
 sg13g2_tiehi _3828__283 (.L_HI(net283));
 sg13g2_tiehi _4030__284 (.L_HI(net284));
 sg13g2_tiehi _3827__285 (.L_HI(net285));
 sg13g2_tiehi _3967__286 (.L_HI(net286));
 sg13g2_tiehi _3826__287 (.L_HI(net287));
 sg13g2_tiehi _4057__288 (.L_HI(net288));
 sg13g2_tiehi _3825__289 (.L_HI(net289));
 sg13g2_tiehi _3966__290 (.L_HI(net290));
 sg13g2_tiehi _3824__291 (.L_HI(net291));
 sg13g2_tiehi _3823__292 (.L_HI(net292));
 sg13g2_tiehi _3822__293 (.L_HI(net293));
 sg13g2_tiehi _3821__294 (.L_HI(net294));
 sg13g2_tiehi _3820__295 (.L_HI(net295));
 sg13g2_tiehi _3819__296 (.L_HI(net296));
 sg13g2_tiehi _3818__297 (.L_HI(net297));
 sg13g2_tiehi _3817__298 (.L_HI(net298));
 sg13g2_tiehi _3816__299 (.L_HI(net299));
 sg13g2_tiehi _3815__300 (.L_HI(net300));
 sg13g2_tiehi _3814__301 (.L_HI(net301));
 sg13g2_tiehi _4029__302 (.L_HI(net302));
 sg13g2_tiehi _3810__303 (.L_HI(net303));
 sg13g2_tiehi _3965__304 (.L_HI(net304));
 sg13g2_tiehi _3809__305 (.L_HI(net305));
 sg13g2_tiehi _4079__306 (.L_HI(net306));
 sg13g2_tiehi _3808__307 (.L_HI(net307));
 sg13g2_tiehi _3964__308 (.L_HI(net308));
 sg13g2_tiehi _3807__309 (.L_HI(net309));
 sg13g2_tiehi _4028__310 (.L_HI(net310));
 sg13g2_tiehi tt_um_comm_ic_bhavuk_311 (.L_HI(net311));
 sg13g2_tiehi tt_um_comm_ic_bhavuk_312 (.L_HI(net312));
 sg13g2_tiehi tt_um_comm_ic_bhavuk_313 (.L_HI(net313));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0027_),
    .X(net314));
 sg13g2_buf_1 _4392_ (.A(\comm_ic0.SDA_op_en ),
    .X(uio_oe[0]));
 sg13g2_buf_1 _4393_ (.A(uio_oe[5]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _4394_ (.A(uio_oe[5]),
    .X(uio_oe[3]));
 sg13g2_buf_1 _4395_ (.A(uio_oe[5]),
    .X(uio_oe[4]));
 sg13g2_buf_1 _4396_ (.A(\comm_ic0.SDA_op ),
    .X(uio_out[0]));
 sg13g2_buf_2 _4397_ (.A(\comm_ic0.new_uart ),
    .X(uio_out[1]));
 sg13g2_buf_1 _4398_ (.A(\comm_ic0.error_i2c ),
    .X(uio_out[6]));
 sg13g2_buf_1 _4399_ (.A(clk),
    .X(uio_out[7]));
 sg13g2_buf_2 _4400_ (.A(\comm_ic0.UART_TX ),
    .X(uo_out[0]));
 sg13g2_buf_4 _4401_ (.X(uo_out[1]),
    .A(\comm_ic0.SEN ));
 sg13g2_buf_4 _4402_ (.X(uo_out[2]),
    .A(\comm_ic0.SCLK ));
 sg13g2_buf_4 _4403_ (.X(uo_out[3]),
    .A(\comm_ic0.MOSI ));
 sg13g2_buf_1 _4404_ (.A(\comm_ic0.SCL ),
    .X(uo_out[4]));
 sg13g2_buf_2 _4405_ (.A(\comm_ic0.busy_uart ),
    .X(uo_out[5]));
 sg13g2_buf_2 _4406_ (.A(\comm_ic0.busy_spi ),
    .X(uo_out[6]));
 sg13g2_buf_1 _4407_ (.A(\comm_ic0.busy_i2c ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout527 (.A(_0616_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_0616_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(net530),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_0822_),
    .X(net530));
 sg13g2_buf_4 fanout531 (.X(net531),
    .A(net532));
 sg13g2_buf_2 fanout532 (.A(_1598_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(net534),
    .X(net533));
 sg13g2_buf_4 fanout534 (.X(net534),
    .A(_1597_));
 sg13g2_buf_2 fanout535 (.A(net536),
    .X(net535));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(net537));
 sg13g2_buf_2 fanout537 (.A(_1596_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_1565_),
    .X(net538));
 sg13g2_buf_4 fanout539 (.X(net539),
    .A(net1080));
 sg13g2_buf_2 fanout540 (.A(_0959_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(net542),
    .X(net541));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(_0957_));
 sg13g2_buf_2 fanout543 (.A(_0556_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_0556_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_0452_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_0452_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_0354_),
    .X(net547));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(_1518_));
 sg13g2_buf_2 fanout549 (.A(_0455_),
    .X(net549));
 sg13g2_buf_4 fanout550 (.X(net550),
    .A(net551));
 sg13g2_buf_4 fanout551 (.X(net551),
    .A(net552));
 sg13g2_buf_2 fanout552 (.A(_1580_),
    .X(net552));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(net554));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(_1580_));
 sg13g2_buf_2 fanout555 (.A(\comm_ic0.uart0.rx_ind[2] ),
    .X(net555));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(net557));
 sg13g2_buf_4 fanout557 (.X(net557),
    .A(net558));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(_1081_));
 sg13g2_buf_2 fanout559 (.A(_1081_),
    .X(net559));
 sg13g2_buf_4 fanout560 (.X(net560),
    .A(_0357_));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(_1599_));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(_1573_));
 sg13g2_buf_4 fanout563 (.X(net563),
    .A(_1468_));
 sg13g2_buf_4 fanout564 (.X(net564),
    .A(_1467_));
 sg13g2_buf_2 fanout565 (.A(net566),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_1464_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(net568),
    .X(net567));
 sg13g2_buf_4 fanout568 (.X(net568),
    .A(net570));
 sg13g2_buf_2 fanout569 (.A(net570),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(_1460_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_1437_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_1432_),
    .X(net572));
 sg13g2_buf_4 fanout573 (.X(net573),
    .A(_1430_));
 sg13g2_buf_2 fanout574 (.A(net575),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_1408_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_4 fanout578 (.X(net578),
    .A(_1408_));
 sg13g2_buf_2 fanout579 (.A(net771),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(net1129),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(net1128),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_0043_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(net584),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(net1186),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(net908),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net1209),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(net831),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(net1292),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(net1292),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(net1132),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(net594),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(net1131),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(net914),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(\comm_ic0.uart0.curr_st[2] ),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(net1160),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(net1138),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(net1138),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(net602),
    .X(net600));
 sg13g2_buf_1 fanout601 (.A(net602),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(net1038),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(net604),
    .X(net603));
 sg13g2_buf_4 fanout604 (.X(net604),
    .A(net1262));
 sg13g2_buf_2 fanout605 (.A(net1261),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(net612),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(net612),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(net609),
    .X(net608));
 sg13g2_buf_1 fanout609 (.A(net610),
    .X(net609));
 sg13g2_buf_1 fanout610 (.A(net611),
    .X(net610));
 sg13g2_buf_1 fanout611 (.A(net612),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(\comm_ic0.uart0.par_en ),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net620),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(net616),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(net616),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(net620),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(net619),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(net619),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(\comm_ic0.uart0.clk_b ),
    .X(net620));
 sg13g2_buf_4 fanout621 (.X(net621),
    .A(net825));
 sg13g2_buf_2 fanout622 (.A(net824),
    .X(net622));
 sg13g2_buf_4 fanout623 (.X(net623),
    .A(net624));
 sg13g2_buf_2 fanout624 (.A(net1065),
    .X(net624));
 sg13g2_buf_4 fanout625 (.X(net625),
    .A(net1034));
 sg13g2_buf_4 fanout626 (.X(net626),
    .A(net627));
 sg13g2_buf_2 fanout627 (.A(net628),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(net629),
    .X(net628));
 sg13g2_buf_4 fanout629 (.X(net629),
    .A(net729));
 sg13g2_buf_4 fanout630 (.X(net630),
    .A(net420));
 sg13g2_buf_1 fanout631 (.A(net420),
    .X(net631));
 sg13g2_buf_4 fanout632 (.X(net632),
    .A(net419));
 sg13g2_buf_4 fanout633 (.X(net633),
    .A(net520));
 sg13g2_buf_2 fanout634 (.A(net637),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(net636),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(net520),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(net519),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(net1142),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(net1142),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(net641),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(net644),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(net643),
    .X(net642));
 sg13g2_buf_4 fanout643 (.X(net643),
    .A(net644));
 sg13g2_buf_2 fanout644 (.A(net651),
    .X(net644));
 sg13g2_buf_4 fanout645 (.X(net645),
    .A(net651));
 sg13g2_buf_2 fanout646 (.A(net651),
    .X(net646));
 sg13g2_buf_4 fanout647 (.X(net647),
    .A(net650));
 sg13g2_buf_2 fanout648 (.A(net650),
    .X(net648));
 sg13g2_buf_1 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(net651),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_1421_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(net654),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(net654),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(net659),
    .X(net654));
 sg13g2_buf_4 fanout655 (.X(net655),
    .A(net656));
 sg13g2_buf_4 fanout656 (.X(net656),
    .A(net659));
 sg13g2_buf_4 fanout657 (.X(net657),
    .A(net658));
 sg13g2_buf_4 fanout658 (.X(net658),
    .A(net659));
 sg13g2_buf_2 fanout659 (.A(_1421_),
    .X(net659));
 sg13g2_buf_4 fanout660 (.X(net660),
    .A(_1334_));
 sg13g2_buf_4 fanout661 (.X(net661),
    .A(net663));
 sg13g2_buf_4 fanout662 (.X(net662),
    .A(net663));
 sg13g2_buf_8 fanout663 (.A(uio_in[5]),
    .X(net663));
 sg13g2_buf_4 fanout664 (.X(net664),
    .A(net667));
 sg13g2_buf_2 fanout665 (.A(net667),
    .X(net665));
 sg13g2_buf_4 fanout666 (.X(net666),
    .A(net667));
 sg13g2_buf_2 fanout667 (.A(uio_in[4]),
    .X(net667));
 sg13g2_buf_4 fanout668 (.X(net668),
    .A(net670));
 sg13g2_buf_2 fanout669 (.A(net670),
    .X(net669));
 sg13g2_buf_8 fanout670 (.A(net5),
    .X(net670));
 sg13g2_buf_4 fanout671 (.X(net671),
    .A(net673));
 sg13g2_buf_4 fanout672 (.X(net672),
    .A(net673));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(uio_in[2]));
 sg13g2_buf_2 fanout674 (.A(net675),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(net679),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(net679),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(net679),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(net696),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(net682),
    .X(net680));
 sg13g2_buf_1 fanout681 (.A(net682),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(net685),
    .X(net682));
 sg13g2_buf_4 fanout683 (.X(net683),
    .A(net685));
 sg13g2_buf_2 fanout684 (.A(net685),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(net696),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(net696),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(net689),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(net690),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(net696),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net695),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(net695),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(net695),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_4 fanout696 (.X(net696),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[1]));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(uio_in[0]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(uio_in[3]),
    .X(net5));
 sg13g2_tiehi _3806__6 (.L_HI(net6));
 sg13g2_dlygate4sd3_1 hold2 (.A(_1409_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold3 (.A(net1280),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold4 (.A(\comm_ic0.spi0.data_wr[9] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold5 (.A(_1099_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0242_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold7 (.A(\comm_ic0.uart0.clk_cnt_reg[0] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0412_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0084_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold10 (.A(\comm_ic0.spi0.data_wr[12] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold11 (.A(_1102_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0245_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold13 (.A(net455),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0762_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0162_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold16 (.A(\comm_ic0.spi0.data_wr[10] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold17 (.A(_1100_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0243_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold19 (.A(net1337),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0911_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0199_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold22 (.A(\comm_ic0.spi0.data_wr[2] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold23 (.A(_1092_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0235_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold25 (.A(\comm_ic0.i2c_addr_en ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold26 (.A(_1325_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0352_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold28 (.A(\comm_ic0.spi0.data_wr[0] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold29 (.A(_1090_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0233_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold31 (.A(net459),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0765_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0165_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold34 (.A(\comm_ic0.spi0.data_in[5] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold35 (.A(_1354_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0325_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold37 (.A(\comm_ic0.spi0.data_in[11] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold38 (.A(_1348_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0331_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold40 (.A(\comm_ic0.spi0.data_in[1] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold41 (.A(_1346_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0333_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold43 (.A(\comm_ic0.spi0.data_in[7] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold44 (.A(_1352_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0327_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold46 (.A(\comm_ic0.spi0.data_wr[13] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold47 (.A(_1103_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0246_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold49 (.A(\comm_ic0.spi0.data_wr[15] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold50 (.A(_1105_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0248_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold52 (.A(\comm_ic0.i2c0.data_out[8] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0866_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0178_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold55 (.A(net1339),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0760_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0160_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold58 (.A(\comm_ic0.spi0.data_wr[14] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold59 (.A(_1104_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0247_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold61 (.A(net451),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0761_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0161_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold64 (.A(\comm_ic0.i2c0.data_out[4] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0849_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0174_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold67 (.A(\comm_ic0.spi0.data_in[10] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold68 (.A(_1349_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0330_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold70 (.A(net1338),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0753_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0153_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0074_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold74 (.A(_1590_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0007_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold76 (.A(\comm_ic0.i2c0.address[6] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold77 (.A(_1396_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0271_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold79 (.A(net947),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0907_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0195_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold82 (.A(\comm_ic0.uart0.clk_cnt[6] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold83 (.A(_1341_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0338_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold85 (.A(\comm_ic0.spi0.data_in[3] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold86 (.A(_1344_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0335_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold88 (.A(\comm_ic0.spi0.clk_cnt[6] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold89 (.A(_1357_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0322_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold91 (.A(\comm_ic0.spi0.data_in[6] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold92 (.A(_1353_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0326_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold94 (.A(\comm_ic0.spi0.data_wr[3] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold95 (.A(_1093_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0236_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold97 (.A(net1341),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0767_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0167_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold100 (.A(net484),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0913_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0201_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold103 (.A(\comm_ic0.spi0.data_wr[1] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold104 (.A(_1091_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0234_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold106 (.A(\comm_ic0.send_cnt[1] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold107 (.A(net632),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold108 (.A(_1277_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0312_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold110 (.A(net510),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0910_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0198_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold113 (.A(\comm_ic0.i2c0.addr_wr[7] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0916_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0204_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold116 (.A(\comm_ic0.i2c0.address[2] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold117 (.A(_1329_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0353_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold119 (.A(\comm_ic0.spi0.data_in[8] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold120 (.A(_1351_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0328_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold122 (.A(\comm_ic0.spi0.data_wr[8] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold123 (.A(_1098_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0241_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold125 (.A(\comm_ic0.spi0.data_in[0] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold126 (.A(_1347_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0332_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold128 (.A(\comm_ic0.spi0.data_in[9] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold129 (.A(_1350_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0329_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold131 (.A(\comm_ic0.send_cnt[3] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold132 (.A(_1219_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0276_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0032_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold135 (.A(_1218_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold136 (.A(_1282_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0317_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold138 (.A(\comm_ic0.i2c0.data_in[9] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold139 (.A(\comm_ic0.i2c0.write_n ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0909_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0197_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold142 (.A(\comm_ic0.i2c0.data_in[10] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold143 (.A(\comm_ic0.uart0.clk_cnt_reg[6] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0418_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0090_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold146 (.A(\comm_ic0.i2c0.data_in[13] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold147 (.A(\comm_ic0.i2c0.data_in[14] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold148 (.A(_1392_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0275_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold150 (.A(\comm_ic0.i2c0.data_wr[14] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0766_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0166_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold153 (.A(\comm_ic0.uart0.clk_cnt[2] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0414_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0086_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold156 (.A(\comm_ic0.spi0.data_in[4] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold157 (.A(_1355_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0324_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold159 (.A(\comm_ic0.spi0.data_wr[5] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold160 (.A(_1095_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0238_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold162 (.A(\comm_ic0.i2c0.data_in[12] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold163 (.A(_1394_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0273_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold165 (.A(net834),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold166 (.A(_1089_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0232_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold168 (.A(\comm_ic0.i2c0.data_in[7] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold169 (.A(_1368_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0311_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold171 (.A(\comm_ic0.i2c0.address[3] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0268_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold173 (.A(net515),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0763_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0163_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold176 (.A(\comm_ic0.spi0.data_wr[4] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold177 (.A(_1094_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0237_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold179 (.A(\comm_ic0.spi0.data_wr[11] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold180 (.A(_1101_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0244_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold182 (.A(\comm_ic0.spi0.data_out[4] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0998_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0212_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold185 (.A(\comm_ic0.i2c0.address[4] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold186 (.A(_1398_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0269_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold188 (.A(\comm_ic0.spi0.data_wr[7] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold189 (.A(_1097_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0240_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold191 (.A(\comm_ic0.i2c0.addr_wr[5] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0914_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0202_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold194 (.A(\comm_ic0.rx_ack ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold195 (.A(_1269_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0304_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold197 (.A(\comm_ic0.i2c0.address[0] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0351_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold199 (.A(\comm_ic0.i2c0.data_wr[12] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0764_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0164_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold202 (.A(\comm_ic0.i2c0.data_in[11] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold203 (.A(\comm_ic0.spi0.data_out[8] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold204 (.A(_1033_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0216_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold206 (.A(\comm_ic0.send_cnt[0] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold207 (.A(net637),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold208 (.A(_1532_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0272_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold210 (.A(net763),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0754_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0154_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold213 (.A(\comm_ic0.i2c0.data_out[5] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0854_),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0175_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold216 (.A(\comm_ic0.spi0.CPOL ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold217 (.A(_1124_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0253_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold219 (.A(\comm_ic0.i2c0.data_in[5] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0757_),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0157_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold222 (.A(\comm_ic0.i2c0.addr_wr[3] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0912_),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0200_),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold225 (.A(net755),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0915_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0203_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold228 (.A(net853),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0417_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0089_),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold231 (.A(\comm_ic0.i2c0.data_out[12] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0878_),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0182_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold234 (.A(\comm_ic0.spi0.data_out[6] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold235 (.A(_1015_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0214_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0040_),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0688_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold239 (.A(net1301),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold240 (.A(\comm_ic0.i2c0.data_out[14] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0886_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0184_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold243 (.A(net770),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0752_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0152_),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold246 (.A(\comm_ic0.send_cnt[2] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold247 (.A(net629),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0309_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold249 (.A(\comm_ic0.i2c0.data_out[15] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0890_),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0185_),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold252 (.A(\comm_ic0.i2c0.data_out[13] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0882_),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0183_),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold255 (.A(\comm_ic0.i2c0.bits16 ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold256 (.A(_1389_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0278_),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold258 (.A(\comm_ic0.i2c0.data_out[6] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0859_),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0176_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold261 (.A(\comm_ic0.spi0.clk_cnt_reg[6] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold262 (.A(_1088_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0231_),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold264 (.A(net898),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0413_),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0085_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold267 (.A(\comm_ic0.i2c0.data_in[3] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold268 (.A(_1360_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold269 (.A(\comm_ic0.i2c0.data_in[4] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold270 (.A(_1371_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0308_),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold272 (.A(\comm_ic0.i2c0.address[5] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0270_),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold274 (.A(\comm_ic0.SEN ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0921_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0205_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold277 (.A(net939),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0435_),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0094_),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold280 (.A(\comm_ic0.i2c0.data_in[2] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold281 (.A(\comm_ic0.i2c0.data_out[9] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0868_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0179_),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold284 (.A(\comm_ic0.spi0.data_in[2] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold285 (.A(_1345_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0334_),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold287 (.A(\comm_ic0.i2c0.data_in[0] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold288 (.A(net1245),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold289 (.A(_1271_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0306_),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold291 (.A(net989),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold292 (.A(_1125_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0254_),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold294 (.A(\comm_ic0.MOSI ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0956_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0207_),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold297 (.A(net836),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0416_),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0088_),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold300 (.A(net960),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0415_),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0087_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold303 (.A(\comm_ic0.i2c0.data_out[10] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0871_),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0180_),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold306 (.A(\comm_ic0.spi0.data_out[0] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0966_),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0208_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold309 (.A(\comm_ic0.spi0.clk_cnt[4] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold310 (.A(_1359_),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0320_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold312 (.A(\comm_ic0.spi0.data_out[12] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold313 (.A(_1055_),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0220_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold315 (.A(\comm_ic0.i2c0.data_out[2] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0840_),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0172_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold318 (.A(net936),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0434_),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0093_),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold321 (.A(\comm_ic0.i2c0.data_wr[4] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0756_),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold323 (.A(\comm_ic0.i2c0.data_in[6] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold324 (.A(_1369_),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold325 (.A(\comm_ic0.spi0.data_wr[6] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold326 (.A(_1096_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0239_),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold328 (.A(\comm_ic0.i2c0.data_out[11] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0874_),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0181_),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold331 (.A(\comm_ic0.i2c0.data_out[7] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0864_),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0177_),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold334 (.A(\comm_ic0.i2c0.data_wr[3] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0755_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold336 (.A(\comm_ic0.i2c0.data_wr[7] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0759_),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold338 (.A(\comm_ic0.uart0.clk_cnt[7] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold339 (.A(_1340_),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0339_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold341 (.A(\comm_ic0.curr_st[3] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold342 (.A(net622),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold343 (.A(_1255_),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0295_),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold345 (.A(\comm_ic0.spi0.clk_cnt_reg[4] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold346 (.A(_1086_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0229_),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold348 (.A(\comm_ic0.i2c0.curr_st[7] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold349 (.A(_1548_),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0013_),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold351 (.A(\comm_ic0.spi0.clk_cnt[7] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0323_),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold353 (.A(\comm_ic0.uart0.clk_cnt[4] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0336_),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold355 (.A(\comm_ic0.uart0.clk_cnt_reg[7] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0419_),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0091_),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold358 (.A(\comm_ic0.i2c0.data_out[1] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0834_),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0171_),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold361 (.A(\comm_ic0.spi0.clk_cnt[2] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold362 (.A(_1386_),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0281_),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold364 (.A(net977),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0905_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0193_),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold367 (.A(\comm_ic0.tx_data[0] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold368 (.A(_1339_),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold369 (.A(_0340_),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold370 (.A(\comm_ic0.uart0.clk_cnt[5] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0337_),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold372 (.A(\comm_ic0.i2c0.data_wr[6] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0758_),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold374 (.A(net1042),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0903_),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0191_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold377 (.A(\comm_ic0.spi0.data_out[9] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold378 (.A(_1034_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0217_),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold380 (.A(\comm_ic0.uart0.clk_cnt[0] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold381 (.A(_1381_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold382 (.A(\comm_ic0.spi0.clk_cnt[5] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold383 (.A(_1358_),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0321_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold385 (.A(\comm_ic0.tx_data[3] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold386 (.A(_1336_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold387 (.A(_0343_),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold388 (.A(\comm_ic0.spi0.data_out[14] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold389 (.A(_1066_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0222_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold391 (.A(\comm_ic0.spi0.data_out[5] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold392 (.A(_1008_),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0213_),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold394 (.A(\comm_ic0.spi0.data_out[11] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold395 (.A(_1048_),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0219_),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold397 (.A(\comm_ic0.spi0.clk_cnt_reg[2] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold398 (.A(_1084_),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0227_),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold400 (.A(\comm_ic0.SDA_op ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0819_),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold402 (.A(net1320),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold403 (.A(\comm_ic0.spi0.data_out[3] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0988_),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0211_),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold406 (.A(\comm_ic0.spi0.data_out[10] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold407 (.A(_1041_),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold408 (.A(_0218_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold409 (.A(\comm_ic0.tx_data[6] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold410 (.A(_1375_),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0299_),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold412 (.A(\comm_ic0.spi0.data_out[2] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0980_),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold414 (.A(_0210_),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold415 (.A(\comm_ic0.uart0.clk_cnt[1] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0039_),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0671_),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold418 (.A(net1291),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold419 (.A(\comm_ic0.tx_data[5] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold420 (.A(_1376_),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0298_),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold422 (.A(\comm_ic0.SCL ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0775_),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold424 (.A(_0168_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold425 (.A(\comm_ic0.spi0.data_ind[1] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold426 (.A(_1115_),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0250_),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold428 (.A(\comm_ic0.spi0.clk_cnt_reg[5] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold429 (.A(_1087_),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0230_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold431 (.A(\comm_ic0.i2c0.curr_st[2] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold432 (.A(_1572_),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold433 (.A(net1293),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold434 (.A(\comm_ic0.tx_data[1] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold435 (.A(_1338_),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0341_),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold437 (.A(\comm_ic0.error_i2c ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold438 (.A(_0897_),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold439 (.A(_0187_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold440 (.A(_0056_),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold441 (.A(_1064_),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold442 (.A(_1065_),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold443 (.A(_0221_),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold444 (.A(\comm_ic0.tx_data[4] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold445 (.A(_1377_),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0297_),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold447 (.A(net945),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold448 (.A(_1083_),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold449 (.A(_0226_),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold450 (.A(uio_out[5]),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold451 (.A(_0739_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0151_),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold453 (.A(\comm_ic0.parity_odd ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold454 (.A(_1267_),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold455 (.A(_0302_),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold456 (.A(\comm_ic0.parity_en ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold457 (.A(_1268_),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0303_),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold459 (.A(\comm_ic0.uart0.setting ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold460 (.A(_1586_),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0023_),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold462 (.A(\comm_ic0.spi0.clk_cnt[1] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold463 (.A(_0280_),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold464 (.A(\comm_ic0.i2c0.clk_cnt[6] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold465 (.A(_1323_),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0349_),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold467 (.A(\comm_ic0.spi0.mode[1] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold468 (.A(_1236_),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold469 (.A(_0284_),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold470 (.A(\comm_ic0.i2c0.data_out[3] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold471 (.A(_0846_),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold472 (.A(_0173_),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold473 (.A(_0058_),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold474 (.A(_1077_),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold475 (.A(_1078_),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold476 (.A(_0223_),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold477 (.A(\comm_ic0.uart0.clk_cnt[3] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold478 (.A(_0296_),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold479 (.A(net1060),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold480 (.A(_1082_),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold481 (.A(_0225_),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold482 (.A(\comm_ic0.uart0.uclk_cnt[7] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold483 (.A(_0406_),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0083_),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold485 (.A(\comm_ic0.spi0.data_in[14] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold486 (.A(_1243_),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold487 (.A(_0288_),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold488 (.A(\comm_ic0.i2c0.addr_ind[2] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold489 (.A(_0696_),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold490 (.A(_0147_),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold491 (.A(\comm_ic0.busy_spi ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold492 (.A(_1080_),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0224_),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold494 (.A(\comm_ic0.i2c0.clk_cnt[4] ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold495 (.A(_1321_),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold496 (.A(_0347_),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold497 (.A(\comm_ic0.tx_data[7] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold498 (.A(_1374_),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0300_),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold500 (.A(\comm_ic0.spi0.clk_cnt[3] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold501 (.A(_1385_),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold502 (.A(_0282_),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold503 (.A(uio_out[2]),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold504 (.A(_0700_),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold505 (.A(_0148_),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold506 (.A(\comm_ic0.spi0.mode[0] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold507 (.A(_1234_),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold508 (.A(_0283_),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold509 (.A(\comm_ic0.spi0.clk_cnt_reg[3] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold510 (.A(_1085_),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold511 (.A(_0228_),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold512 (.A(\comm_ic0.spi0.data_in[15] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold513 (.A(_1244_),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold514 (.A(_0289_),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold515 (.A(uio_out[3]),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold516 (.A(_0713_),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold517 (.A(_0149_),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold518 (.A(uio_out[4]),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold519 (.A(_0726_),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold520 (.A(_0150_),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold521 (.A(net1227),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold522 (.A(_0893_),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold523 (.A(_0186_),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold524 (.A(\comm_ic0.spi0.data_in[13] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold525 (.A(_1242_),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold526 (.A(_0287_),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold527 (.A(\comm_ic0.uart0.uclk_cnt[4] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold528 (.A(_0391_),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold529 (.A(_0080_),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold530 (.A(\comm_ic0.uart0.uclk_cnt[1] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold531 (.A(_0372_),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold532 (.A(_0077_),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold533 (.A(\comm_ic0.uart0.uclk_cnt[2] ),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold534 (.A(_0380_),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold535 (.A(_0078_),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold536 (.A(net1103),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0908_),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold538 (.A(_0196_),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold539 (.A(\comm_ic0.spi0.data_out[1] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold540 (.A(_0967_),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold541 (.A(_0209_),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold542 (.A(net1093),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold543 (.A(_0904_),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold544 (.A(_0192_),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold545 (.A(net1096),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold546 (.A(_0906_),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold547 (.A(_0194_),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold548 (.A(\comm_ic0.SCLK ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold549 (.A(_0927_),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold550 (.A(_0206_),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold551 (.A(net1275),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold552 (.A(net625),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold553 (.A(_1249_),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold554 (.A(_0291_),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold555 (.A(\comm_ic0.i2c0.data_ind[3] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold556 (.A(net602),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold557 (.A(_0684_),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold558 (.A(_0144_),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold559 (.A(\comm_ic0.i2c0.clk_cnt[2] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold560 (.A(_1209_),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold561 (.A(_0266_),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold562 (.A(\comm_ic0.i2c0.curr_st[4] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold563 (.A(_1587_),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold564 (.A(_0008_),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold565 (.A(\comm_ic0.uart0.uclk_cnt[0] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold566 (.A(_0366_),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold567 (.A(_0076_),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold568 (.A(\comm_ic0.uart0.uclk_cnt[3] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold569 (.A(_0386_),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold570 (.A(_0079_),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold571 (.A(net1137),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold572 (.A(_0901_),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold573 (.A(_0189_),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold574 (.A(\comm_ic0.i2c0.data_out[0] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold575 (.A(_0826_),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold576 (.A(_0170_),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold577 (.A(\comm_ic0.spi0.clk_cnt[0] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold578 (.A(_0279_),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold579 (.A(net1125),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold580 (.A(_0902_),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold581 (.A(_0190_),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold582 (.A(\comm_ic0.curr_st[1] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold583 (.A(_1240_),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold584 (.A(_0285_),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold585 (.A(\comm_ic0.tx_data[2] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold586 (.A(_1337_),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold587 (.A(_0342_),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold588 (.A(\comm_ic0.i2c0.curr_st[3] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold589 (.A(_1584_),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold590 (.A(_0009_),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold591 (.A(\comm_ic0.uart0.enable ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold592 (.A(_0022_),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold593 (.A(\comm_ic0.spi0.data_in[12] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold594 (.A(_1241_),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold595 (.A(_0286_),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold596 (.A(\comm_ic0.i2c0.scl_cnt[7] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold597 (.A(_1547_),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold598 (.A(net539),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold599 (.A(_1581_),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold600 (.A(_0010_),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold601 (.A(\comm_ic0.uart0.uclk_cnt[5] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold602 (.A(_0398_),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold603 (.A(_0081_),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold604 (.A(\comm_ic0.spi0.data_out[7] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold605 (.A(_1022_),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold606 (.A(_1028_),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold607 (.A(_0215_),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold608 (.A(uio_oe[5]),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold609 (.A(_0307_),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold610 (.A(\comm_ic0.i2c0.clk_cnt[3] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold611 (.A(_1210_),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold612 (.A(_0267_),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold613 (.A(\comm_ic0.i2c0.clk_cnt[5] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold614 (.A(_1322_),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold615 (.A(_0348_),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold616 (.A(_0071_),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold617 (.A(_1253_),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold618 (.A(_1254_),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold619 (.A(_0292_),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold620 (.A(\comm_ic0.i2c0.clk_cnt[7] ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold621 (.A(_1324_),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold622 (.A(_0350_),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold623 (.A(\comm_ic0.spi0.curr_st[3] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold624 (.A(_1594_),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold625 (.A(_0021_),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold626 (.A(net1277),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold627 (.A(_1245_),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold628 (.A(_0290_),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold629 (.A(\comm_ic0.tx_new ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold630 (.A(_1372_),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold631 (.A(_1265_),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold632 (.A(_1266_),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold633 (.A(net1217),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold634 (.A(_1509_),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold635 (.A(_1510_),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold636 (.A(_1512_),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold637 (.A(_1522_),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold638 (.A(_0017_),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold639 (.A(\comm_ic0.i2c0.data_ind[1] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold640 (.A(_0676_),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold641 (.A(_0142_),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold642 (.A(\comm_ic0.i2c0.clk_cnt[1] ),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold643 (.A(_1208_),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold644 (.A(_0265_),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold645 (.A(\comm_ic0.comm_sel[0] ),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold646 (.A(net581),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold647 (.A(_1270_),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold648 (.A(\comm_ic0.i2c0.curr_st[5] ),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold649 (.A(net594),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold650 (.A(_0011_),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold651 (.A(\comm_ic0.spi0.curr_st[1] ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold652 (.A(_1462_),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold653 (.A(_0019_),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold654 (.A(\comm_ic0.i2c0.clk_cnt[0] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold655 (.A(\comm_ic0.uart0.curr_st[1] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold656 (.A(net599),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold657 (.A(_0420_),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold658 (.A(_0092_),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold659 (.A(\comm_ic0.spi0.curr_st[2] ),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold660 (.A(net639),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold661 (.A(_1614_),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold662 (.A(_0020_),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold663 (.A(\comm_ic0.spi0.data_ind[3] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold664 (.A(_1120_),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold665 (.A(_0252_),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold666 (.A(\comm_ic0.uart0.uclk_cnt[6] ),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold667 (.A(_0399_),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold668 (.A(_0405_),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold669 (.A(_0082_),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold670 (.A(\comm_ic0.i2c0.addr_ind[1] ),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold671 (.A(_0694_),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold672 (.A(_0146_),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold673 (.A(\comm_ic0.i2c0.scl_cnt[6] ),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold674 (.A(_1181_),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold675 (.A(_1182_),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold676 (.A(_0261_),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold677 (.A(\comm_ic0.uart0.curr_st[2] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold678 (.A(net597),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold679 (.A(_0000_),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold680 (.A(_0063_),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold681 (.A(_0491_),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold682 (.A(_0492_),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold683 (.A(_0497_),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold684 (.A(_0101_),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold685 (.A(net1276),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold686 (.A(_1478_),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold687 (.A(_1516_),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold688 (.A(_0015_),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold689 (.A(_0061_),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold690 (.A(_0472_),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold691 (.A(_0473_),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold692 (.A(_0480_),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold693 (.A(_0099_),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold694 (.A(_0065_),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold695 (.A(_0508_),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold696 (.A(_0509_),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold697 (.A(_0515_),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold698 (.A(_0103_),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold699 (.A(net1202),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold700 (.A(_1199_),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold701 (.A(_1202_),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold702 (.A(_1205_),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold703 (.A(\comm_ic0.spi0.data_ind[2] ),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold704 (.A(net585),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold705 (.A(_1119_),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold706 (.A(_0251_),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold707 (.A(\comm_ic0.i2c0.curr_st[1] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold708 (.A(_1592_),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold709 (.A(_0006_),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold710 (.A(\comm_ic0.spi0.curr_st[0] ),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold711 (.A(_1459_),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold712 (.A(_0018_),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold713 (.A(_0069_),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold714 (.A(_1440_),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold715 (.A(_1163_),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold716 (.A(_1164_),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold717 (.A(_1172_),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold718 (.A(_0259_),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold719 (.A(_0073_),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold720 (.A(_0002_),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold721 (.A(_0067_),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold722 (.A(_1143_),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold723 (.A(_1145_),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold724 (.A(_1153_),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold725 (.A(_0257_),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold726 (.A(\comm_ic0.spi0.data_ind[0] ),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold727 (.A(net587),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold728 (.A(_1111_),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold729 (.A(_0249_),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold730 (.A(\comm_ic0.i2c0.start ),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold731 (.A(_1196_),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold732 (.A(_1197_),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold733 (.A(_0262_),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold734 (.A(_0072_),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold735 (.A(_1618_),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold736 (.A(_1619_),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold737 (.A(_0003_),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold738 (.A(\comm_ic0.spi0.sclk_cnt[5] ),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold739 (.A(_1423_),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold740 (.A(_0501_),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold741 (.A(_0502_),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold742 (.A(_0505_),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold743 (.A(_0102_),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold744 (.A(\comm_ic0.busy_i2c ),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold745 (.A(_1226_),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold746 (.A(_0277_),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold747 (.A(\comm_ic0.i2c0.clk_cnt_reg[0] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold748 (.A(_1133_),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold749 (.A(_1134_),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold750 (.A(_0255_),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold751 (.A(\comm_ic0.spi0.sclk_cnt[0] ),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold752 (.A(_1422_),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold753 (.A(_0462_),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold754 (.A(_0463_),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold755 (.A(_0097_),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold756 (.A(_0062_),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold757 (.A(_0474_),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold758 (.A(_0484_),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold759 (.A(_0485_),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold760 (.A(_0488_),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold761 (.A(_0100_),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold762 (.A(\comm_ic0.comm_sel[1] ),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold763 (.A(\comm_ic0.i2c0.clk_cnt_reg[3] ),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold764 (.A(_1159_),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold765 (.A(_1160_),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold766 (.A(_1161_),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold767 (.A(_0258_),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold768 (.A(\comm_ic0.spi0.clk_cnt_reg[7] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold769 (.A(_0517_),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold770 (.A(_0518_),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold771 (.A(_0521_),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold772 (.A(_0104_),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold773 (.A(_0068_),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold774 (.A(_1166_),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold775 (.A(_1179_),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold776 (.A(_1180_),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold777 (.A(_0260_),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold778 (.A(\comm_ic0.i2c0.data_ind[2] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold779 (.A(net605),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold780 (.A(_0679_),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold781 (.A(_0143_),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold782 (.A(\comm_ic0.spi0.sclk_cnt[1] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold783 (.A(_0467_),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold784 (.A(_0469_),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold785 (.A(_0470_),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold786 (.A(_0098_),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold787 (.A(\comm_ic0.i2c0.scl_cnt[1] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold788 (.A(_1135_),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold789 (.A(_1136_),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold790 (.A(_1142_),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold791 (.A(_0256_),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold792 (.A(\comm_ic0.curr_st[0] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold793 (.A(\comm_ic0.curr_st[2] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold794 (.A(\comm_ic0.spi0.bits16 ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold795 (.A(\comm_ic0.SDA_op_en ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold796 (.A(_0900_),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold797 (.A(_0188_),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold798 (.A(_0054_),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold799 (.A(_1054_),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold800 (.A(_0046_),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold801 (.A(_0997_),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold802 (.A(\comm_ic0.spi0.data_out[15] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold803 (.A(_0048_),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold804 (.A(_1014_),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold805 (.A(_0047_),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold806 (.A(_0055_),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold807 (.A(\comm_ic0.i2c0.data_ind[0] ),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold808 (.A(_0141_),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold809 (.A(\comm_ic0.i2c0.curr_st[6] ),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold810 (.A(_0012_),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold811 (.A(_0052_),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold812 (.A(_1040_),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold813 (.A(\comm_ic0.uart0.curr_st[0] ),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold814 (.A(_0044_),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold815 (.A(_0979_),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold816 (.A(\comm_ic0.i2c0.addr_ind[0] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold817 (.A(_0689_),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold818 (.A(_0145_),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold819 (.A(_0057_),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold820 (.A(_0026_),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold821 (.A(\comm_ic0.spi0.start ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold822 (.A(_0070_),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold823 (.A(_1190_),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold824 (.A(_0049_),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold825 (.A(_0053_),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold826 (.A(_0045_),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold827 (.A(_0984_),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold828 (.A(_0987_),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold829 (.A(\comm_ic0.i2c0.curr_st[0] ),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold830 (.A(\comm_ic0.i2c0.scl_cnt[4] ),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold831 (.A(\comm_ic0.i2c0.addr_ind[0] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold832 (.A(_0042_),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold833 (.A(_1109_),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold834 (.A(_1110_),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold835 (.A(_0031_),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold836 (.A(_0818_),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold837 (.A(_0169_),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold838 (.A(\comm_ic0.uart0.clk_cnt_reg[1] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold839 (.A(_0432_),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold840 (.A(_0433_),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold841 (.A(_0038_),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold842 (.A(_0402_),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold843 (.A(_0403_),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold844 (.A(\comm_ic0.i2c0.curr_st[1] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold845 (.A(\comm_ic0.spi0.sclk_cnt[7] ),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold846 (.A(_1456_),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold847 (.A(\comm_ic0.spi0.data_out[13] ),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold848 (.A(\comm_ic0.i2c0.clk_cnt_reg[7] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold849 (.A(_1564_),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold850 (.A(\comm_ic0.spi0.sclk_cnt[4] ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold851 (.A(_1444_),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold852 (.A(_1450_),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold853 (.A(\comm_ic0.spi0.clk_cnt_reg[7] ),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold854 (.A(\comm_ic0.i2c0.address[1] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold855 (.A(\comm_ic0.i2c0.data_in[1] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold856 (.A(\comm_ic0.i2c0.data_in[8] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold857 (.A(_0051_),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold858 (.A(\comm_ic0.i2c0.data_in[15] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold859 (.A(\comm_ic0.i2c0.data_wr[8] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold860 (.A(\comm_ic0.spi0.data_in[13] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold861 (.A(\comm_ic0.i2c0.data_wr[10] ),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold862 (.A(\comm_ic0.i2c0.addr_wr[2] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold863 (.A(_0041_),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold864 (.A(\comm_ic0.i2c0.data_wr[13] ),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold865 (.A(\comm_ic0.i2c0.curr_st[0] ),
    .X(net1348));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_fill_2 FILLER_0_140 ();
 sg13g2_fill_2 FILLER_0_157 ();
 sg13g2_fill_2 FILLER_0_165 ();
 sg13g2_fill_1 FILLER_0_206 ();
 sg13g2_fill_2 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_236 ();
 sg13g2_decap_8 FILLER_0_243 ();
 sg13g2_decap_8 FILLER_0_250 ();
 sg13g2_decap_8 FILLER_0_257 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_fill_1 FILLER_0_271 ();
 sg13g2_fill_1 FILLER_0_295 ();
 sg13g2_fill_2 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_4 FILLER_1_126 ();
 sg13g2_fill_2 FILLER_1_130 ();
 sg13g2_decap_8 FILLER_1_244 ();
 sg13g2_decap_8 FILLER_1_251 ();
 sg13g2_decap_8 FILLER_1_258 ();
 sg13g2_fill_1 FILLER_1_298 ();
 sg13g2_fill_2 FILLER_1_334 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_fill_2 FILLER_2_126 ();
 sg13g2_fill_2 FILLER_2_217 ();
 sg13g2_fill_1 FILLER_2_252 ();
 sg13g2_fill_1 FILLER_2_271 ();
 sg13g2_fill_1 FILLER_2_298 ();
 sg13g2_fill_2 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_379 ();
 sg13g2_decap_8 FILLER_2_386 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_fill_2 FILLER_3_105 ();
 sg13g2_fill_1 FILLER_3_111 ();
 sg13g2_fill_2 FILLER_3_117 ();
 sg13g2_fill_1 FILLER_3_119 ();
 sg13g2_fill_1 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_4 FILLER_4_91 ();
 sg13g2_fill_1 FILLER_4_95 ();
 sg13g2_fill_1 FILLER_4_238 ();
 sg13g2_fill_1 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_fill_2 FILLER_5_84 ();
 sg13g2_fill_1 FILLER_5_86 ();
 sg13g2_fill_2 FILLER_5_145 ();
 sg13g2_fill_1 FILLER_5_171 ();
 sg13g2_fill_1 FILLER_5_199 ();
 sg13g2_fill_1 FILLER_5_284 ();
 sg13g2_fill_2 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_4 FILLER_5_403 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_4 FILLER_6_77 ();
 sg13g2_fill_2 FILLER_6_81 ();
 sg13g2_fill_2 FILLER_6_101 ();
 sg13g2_fill_2 FILLER_6_230 ();
 sg13g2_fill_1 FILLER_6_344 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_4 FILLER_7_70 ();
 sg13g2_fill_1 FILLER_7_74 ();
 sg13g2_fill_1 FILLER_7_101 ();
 sg13g2_fill_1 FILLER_7_121 ();
 sg13g2_fill_1 FILLER_7_266 ();
 sg13g2_fill_2 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_387 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_4 FILLER_8_70 ();
 sg13g2_fill_1 FILLER_8_132 ();
 sg13g2_fill_1 FILLER_8_175 ();
 sg13g2_fill_1 FILLER_8_220 ();
 sg13g2_fill_2 FILLER_8_240 ();
 sg13g2_fill_1 FILLER_8_255 ();
 sg13g2_fill_1 FILLER_8_261 ();
 sg13g2_fill_2 FILLER_8_271 ();
 sg13g2_decap_8 FILLER_8_387 ();
 sg13g2_decap_8 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_fill_2 FILLER_9_77 ();
 sg13g2_fill_1 FILLER_9_143 ();
 sg13g2_fill_1 FILLER_9_182 ();
 sg13g2_fill_1 FILLER_9_235 ();
 sg13g2_fill_1 FILLER_9_305 ();
 sg13g2_fill_1 FILLER_9_341 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_fill_1 FILLER_10_160 ();
 sg13g2_fill_1 FILLER_10_204 ();
 sg13g2_fill_2 FILLER_10_226 ();
 sg13g2_fill_2 FILLER_10_236 ();
 sg13g2_fill_1 FILLER_10_238 ();
 sg13g2_fill_1 FILLER_10_324 ();
 sg13g2_fill_2 FILLER_10_334 ();
 sg13g2_fill_2 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_4 FILLER_10_403 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_fill_2 FILLER_11_84 ();
 sg13g2_fill_1 FILLER_11_105 ();
 sg13g2_fill_2 FILLER_11_115 ();
 sg13g2_fill_1 FILLER_11_171 ();
 sg13g2_fill_1 FILLER_11_176 ();
 sg13g2_fill_2 FILLER_11_220 ();
 sg13g2_fill_1 FILLER_11_222 ();
 sg13g2_fill_1 FILLER_11_232 ();
 sg13g2_fill_1 FILLER_11_269 ();
 sg13g2_decap_8 FILLER_11_377 ();
 sg13g2_decap_8 FILLER_11_384 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_fill_2 FILLER_12_77 ();
 sg13g2_fill_1 FILLER_12_79 ();
 sg13g2_fill_2 FILLER_12_139 ();
 sg13g2_fill_1 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_180 ();
 sg13g2_fill_2 FILLER_12_184 ();
 sg13g2_fill_2 FILLER_12_218 ();
 sg13g2_fill_1 FILLER_12_225 ();
 sg13g2_fill_2 FILLER_12_240 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_fill_2 FILLER_13_70 ();
 sg13g2_fill_1 FILLER_13_72 ();
 sg13g2_decap_8 FILLER_13_145 ();
 sg13g2_fill_2 FILLER_13_160 ();
 sg13g2_fill_2 FILLER_13_176 ();
 sg13g2_fill_1 FILLER_13_231 ();
 sg13g2_fill_1 FILLER_13_245 ();
 sg13g2_fill_1 FILLER_13_255 ();
 sg13g2_fill_2 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_fill_1 FILLER_14_70 ();
 sg13g2_fill_2 FILLER_14_153 ();
 sg13g2_fill_2 FILLER_14_278 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_fill_2 FILLER_15_70 ();
 sg13g2_fill_1 FILLER_15_72 ();
 sg13g2_fill_2 FILLER_15_122 ();
 sg13g2_fill_2 FILLER_15_170 ();
 sg13g2_fill_1 FILLER_15_207 ();
 sg13g2_fill_1 FILLER_15_227 ();
 sg13g2_fill_2 FILLER_15_236 ();
 sg13g2_fill_1 FILLER_15_254 ();
 sg13g2_fill_2 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_4 FILLER_16_77 ();
 sg13g2_fill_1 FILLER_16_81 ();
 sg13g2_fill_1 FILLER_16_86 ();
 sg13g2_fill_2 FILLER_16_151 ();
 sg13g2_fill_1 FILLER_16_182 ();
 sg13g2_fill_2 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_325 ();
 sg13g2_fill_2 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_fill_2 FILLER_17_84 ();
 sg13g2_fill_1 FILLER_17_120 ();
 sg13g2_fill_2 FILLER_17_153 ();
 sg13g2_fill_1 FILLER_17_174 ();
 sg13g2_fill_1 FILLER_17_217 ();
 sg13g2_decap_4 FILLER_17_230 ();
 sg13g2_fill_1 FILLER_17_234 ();
 sg13g2_fill_2 FILLER_17_275 ();
 sg13g2_fill_2 FILLER_17_291 ();
 sg13g2_fill_2 FILLER_17_337 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_fill_2 FILLER_18_77 ();
 sg13g2_fill_1 FILLER_18_142 ();
 sg13g2_fill_2 FILLER_18_169 ();
 sg13g2_fill_2 FILLER_18_186 ();
 sg13g2_fill_2 FILLER_18_202 ();
 sg13g2_fill_1 FILLER_18_210 ();
 sg13g2_fill_2 FILLER_18_220 ();
 sg13g2_decap_4 FILLER_18_239 ();
 sg13g2_fill_1 FILLER_18_243 ();
 sg13g2_fill_2 FILLER_18_256 ();
 sg13g2_fill_1 FILLER_18_306 ();
 sg13g2_fill_1 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_383 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_fill_2 FILLER_19_70 ();
 sg13g2_fill_1 FILLER_19_72 ();
 sg13g2_decap_8 FILLER_19_239 ();
 sg13g2_fill_1 FILLER_19_256 ();
 sg13g2_fill_1 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_fill_2 FILLER_20_96 ();
 sg13g2_fill_2 FILLER_20_103 ();
 sg13g2_fill_2 FILLER_20_132 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_fill_2 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_233 ();
 sg13g2_fill_1 FILLER_20_248 ();
 sg13g2_fill_1 FILLER_20_254 ();
 sg13g2_fill_2 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_271 ();
 sg13g2_fill_2 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_fill_2 FILLER_21_56 ();
 sg13g2_fill_2 FILLER_21_97 ();
 sg13g2_decap_4 FILLER_21_225 ();
 sg13g2_decap_8 FILLER_21_275 ();
 sg13g2_decap_8 FILLER_21_282 ();
 sg13g2_decap_8 FILLER_21_289 ();
 sg13g2_fill_2 FILLER_21_320 ();
 sg13g2_fill_2 FILLER_21_338 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_fill_2 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_135 ();
 sg13g2_fill_2 FILLER_22_218 ();
 sg13g2_fill_1 FILLER_22_259 ();
 sg13g2_fill_1 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_290 ();
 sg13g2_decap_4 FILLER_22_297 ();
 sg13g2_fill_1 FILLER_22_353 ();
 sg13g2_decap_8 FILLER_22_360 ();
 sg13g2_decap_8 FILLER_22_367 ();
 sg13g2_decap_8 FILLER_22_374 ();
 sg13g2_decap_8 FILLER_22_381 ();
 sg13g2_decap_8 FILLER_22_388 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_4 FILLER_23_56 ();
 sg13g2_fill_2 FILLER_23_82 ();
 sg13g2_fill_2 FILLER_23_123 ();
 sg13g2_fill_2 FILLER_23_218 ();
 sg13g2_fill_1 FILLER_23_220 ();
 sg13g2_fill_2 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_340 ();
 sg13g2_fill_1 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_91 ();
 sg13g2_fill_2 FILLER_24_201 ();
 sg13g2_fill_1 FILLER_24_252 ();
 sg13g2_fill_1 FILLER_24_288 ();
 sg13g2_fill_1 FILLER_24_315 ();
 sg13g2_fill_1 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_140 ();
 sg13g2_fill_2 FILLER_25_146 ();
 sg13g2_fill_2 FILLER_25_153 ();
 sg13g2_fill_1 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_167 ();
 sg13g2_fill_2 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_265 ();
 sg13g2_fill_1 FILLER_25_275 ();
 sg13g2_fill_2 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_353 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_fill_2 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_155 ();
 sg13g2_fill_1 FILLER_26_177 ();
 sg13g2_decap_4 FILLER_26_222 ();
 sg13g2_fill_1 FILLER_26_226 ();
 sg13g2_fill_2 FILLER_26_255 ();
 sg13g2_fill_2 FILLER_26_283 ();
 sg13g2_fill_1 FILLER_26_308 ();
 sg13g2_fill_1 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_4 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_97 ();
 sg13g2_fill_1 FILLER_27_176 ();
 sg13g2_fill_2 FILLER_27_201 ();
 sg13g2_fill_2 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_228 ();
 sg13g2_fill_1 FILLER_27_313 ();
 sg13g2_fill_1 FILLER_27_332 ();
 sg13g2_fill_1 FILLER_27_344 ();
 sg13g2_fill_2 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_89 ();
 sg13g2_fill_1 FILLER_28_117 ();
 sg13g2_fill_1 FILLER_28_144 ();
 sg13g2_fill_2 FILLER_28_160 ();
 sg13g2_fill_2 FILLER_28_205 ();
 sg13g2_fill_1 FILLER_28_207 ();
 sg13g2_fill_2 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_fill_2 FILLER_28_241 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_278 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_fill_1 FILLER_29_56 ();
 sg13g2_fill_2 FILLER_29_66 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_fill_1 FILLER_29_189 ();
 sg13g2_fill_2 FILLER_29_234 ();
 sg13g2_fill_1 FILLER_29_256 ();
 sg13g2_fill_2 FILLER_29_271 ();
 sg13g2_fill_2 FILLER_29_305 ();
 sg13g2_fill_2 FILLER_29_371 ();
 sg13g2_fill_1 FILLER_29_373 ();
 sg13g2_decap_8 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_4 FILLER_30_42 ();
 sg13g2_fill_1 FILLER_30_46 ();
 sg13g2_fill_2 FILLER_30_73 ();
 sg13g2_fill_2 FILLER_30_84 ();
 sg13g2_fill_1 FILLER_30_122 ();
 sg13g2_fill_2 FILLER_30_157 ();
 sg13g2_fill_2 FILLER_30_214 ();
 sg13g2_fill_1 FILLER_30_216 ();
 sg13g2_fill_1 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_259 ();
 sg13g2_fill_1 FILLER_30_290 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_decap_8 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_35 ();
 sg13g2_fill_2 FILLER_31_41 ();
 sg13g2_fill_1 FILLER_31_43 ();
 sg13g2_fill_2 FILLER_31_166 ();
 sg13g2_fill_2 FILLER_31_196 ();
 sg13g2_decap_4 FILLER_31_222 ();
 sg13g2_fill_1 FILLER_31_255 ();
 sg13g2_fill_1 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_359 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_4 FILLER_32_21 ();
 sg13g2_fill_2 FILLER_32_25 ();
 sg13g2_fill_1 FILLER_32_79 ();
 sg13g2_fill_2 FILLER_32_154 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_fill_2 FILLER_32_196 ();
 sg13g2_fill_1 FILLER_32_218 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_241 ();
 sg13g2_fill_1 FILLER_32_243 ();
 sg13g2_fill_2 FILLER_32_270 ();
 sg13g2_fill_2 FILLER_32_348 ();
 sg13g2_fill_1 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_376 ();
 sg13g2_decap_8 FILLER_32_383 ();
 sg13g2_decap_8 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_397 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_4 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_25 ();
 sg13g2_fill_2 FILLER_33_134 ();
 sg13g2_fill_1 FILLER_33_136 ();
 sg13g2_fill_1 FILLER_33_236 ();
 sg13g2_fill_2 FILLER_33_267 ();
 sg13g2_fill_1 FILLER_33_269 ();
 sg13g2_fill_2 FILLER_33_282 ();
 sg13g2_decap_4 FILLER_33_288 ();
 sg13g2_decap_4 FILLER_33_296 ();
 sg13g2_fill_2 FILLER_33_300 ();
 sg13g2_fill_2 FILLER_33_370 ();
 sg13g2_fill_1 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_25 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_fill_1 FILLER_34_129 ();
 sg13g2_decap_8 FILLER_34_134 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_decap_4 FILLER_34_215 ();
 sg13g2_decap_8 FILLER_34_225 ();
 sg13g2_fill_1 FILLER_34_232 ();
 sg13g2_fill_1 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_252 ();
 sg13g2_fill_1 FILLER_34_254 ();
 sg13g2_decap_4 FILLER_34_263 ();
 sg13g2_fill_1 FILLER_34_276 ();
 sg13g2_decap_4 FILLER_34_282 ();
 sg13g2_fill_1 FILLER_34_286 ();
 sg13g2_fill_2 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_388 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_41 ();
 sg13g2_fill_1 FILLER_35_43 ();
 sg13g2_decap_4 FILLER_35_124 ();
 sg13g2_fill_1 FILLER_35_128 ();
 sg13g2_fill_2 FILLER_35_165 ();
 sg13g2_fill_2 FILLER_35_176 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_decap_8 FILLER_35_214 ();
 sg13g2_fill_2 FILLER_35_221 ();
 sg13g2_fill_2 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_270 ();
 sg13g2_fill_1 FILLER_35_276 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_28 ();
 sg13g2_fill_2 FILLER_36_32 ();
 sg13g2_fill_1 FILLER_36_38 ();
 sg13g2_fill_2 FILLER_36_88 ();
 sg13g2_fill_2 FILLER_36_116 ();
 sg13g2_fill_1 FILLER_36_118 ();
 sg13g2_fill_2 FILLER_36_145 ();
 sg13g2_fill_1 FILLER_36_175 ();
 sg13g2_fill_1 FILLER_36_210 ();
 sg13g2_fill_1 FILLER_36_225 ();
 sg13g2_fill_1 FILLER_36_266 ();
 sg13g2_fill_2 FILLER_36_272 ();
 sg13g2_fill_1 FILLER_36_274 ();
 sg13g2_fill_2 FILLER_36_342 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_44 ();
 sg13g2_fill_2 FILLER_37_68 ();
 sg13g2_fill_1 FILLER_37_96 ();
 sg13g2_fill_2 FILLER_37_140 ();
 sg13g2_fill_1 FILLER_37_142 ();
 sg13g2_fill_1 FILLER_37_176 ();
 sg13g2_fill_2 FILLER_37_192 ();
 sg13g2_fill_1 FILLER_37_194 ();
 sg13g2_fill_1 FILLER_37_274 ();
 sg13g2_fill_1 FILLER_37_285 ();
 sg13g2_decap_4 FILLER_37_294 ();
 sg13g2_fill_2 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_62 ();
 sg13g2_fill_2 FILLER_38_68 ();
 sg13g2_fill_1 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_97 ();
 sg13g2_decap_8 FILLER_38_104 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_fill_2 FILLER_38_225 ();
 sg13g2_fill_1 FILLER_38_227 ();
 sg13g2_fill_1 FILLER_38_274 ();
 sg13g2_decap_4 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_4 FILLER_39_7 ();
 sg13g2_fill_1 FILLER_39_11 ();
 sg13g2_fill_1 FILLER_39_104 ();
 sg13g2_decap_8 FILLER_39_109 ();
 sg13g2_decap_8 FILLER_39_116 ();
 sg13g2_decap_8 FILLER_39_123 ();
 sg13g2_fill_2 FILLER_39_130 ();
 sg13g2_fill_1 FILLER_39_132 ();
 sg13g2_fill_1 FILLER_39_221 ();
 sg13g2_fill_1 FILLER_39_233 ();
 sg13g2_fill_1 FILLER_39_244 ();
 sg13g2_fill_2 FILLER_39_306 ();
 sg13g2_fill_2 FILLER_39_327 ();
 sg13g2_fill_2 FILLER_39_368 ();
 sg13g2_fill_1 FILLER_39_370 ();
 sg13g2_decap_8 FILLER_39_384 ();
 sg13g2_decap_8 FILLER_39_391 ();
 sg13g2_decap_8 FILLER_39_398 ();
 sg13g2_decap_4 FILLER_39_405 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_52 ();
 sg13g2_fill_1 FILLER_40_54 ();
 sg13g2_fill_1 FILLER_40_63 ();
 sg13g2_fill_1 FILLER_40_213 ();
 sg13g2_fill_2 FILLER_40_236 ();
 sg13g2_fill_1 FILLER_40_238 ();
 sg13g2_fill_1 FILLER_40_253 ();
 sg13g2_fill_2 FILLER_40_278 ();
 sg13g2_decap_8 FILLER_40_292 ();
 sg13g2_fill_2 FILLER_40_299 ();
 sg13g2_fill_2 FILLER_40_356 ();
 sg13g2_fill_1 FILLER_40_358 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_50 ();
 sg13g2_fill_1 FILLER_41_74 ();
 sg13g2_fill_2 FILLER_41_85 ();
 sg13g2_fill_1 FILLER_41_87 ();
 sg13g2_fill_2 FILLER_41_106 ();
 sg13g2_fill_1 FILLER_41_108 ();
 sg13g2_fill_2 FILLER_41_182 ();
 sg13g2_fill_1 FILLER_41_184 ();
 sg13g2_fill_1 FILLER_41_200 ();
 sg13g2_fill_2 FILLER_41_210 ();
 sg13g2_fill_1 FILLER_41_212 ();
 sg13g2_fill_2 FILLER_41_233 ();
 sg13g2_fill_1 FILLER_41_235 ();
 sg13g2_fill_1 FILLER_41_254 ();
 sg13g2_decap_4 FILLER_41_290 ();
 sg13g2_decap_4 FILLER_41_312 ();
 sg13g2_fill_1 FILLER_41_338 ();
 sg13g2_fill_2 FILLER_41_356 ();
 sg13g2_decap_8 FILLER_41_375 ();
 sg13g2_decap_8 FILLER_41_382 ();
 sg13g2_decap_8 FILLER_41_389 ();
 sg13g2_decap_8 FILLER_41_396 ();
 sg13g2_decap_4 FILLER_41_403 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_28 ();
 sg13g2_fill_1 FILLER_42_48 ();
 sg13g2_fill_2 FILLER_42_93 ();
 sg13g2_fill_1 FILLER_42_128 ();
 sg13g2_fill_2 FILLER_42_134 ();
 sg13g2_fill_2 FILLER_42_202 ();
 sg13g2_fill_2 FILLER_42_209 ();
 sg13g2_fill_1 FILLER_42_211 ();
 sg13g2_fill_2 FILLER_42_216 ();
 sg13g2_fill_2 FILLER_42_270 ();
 sg13g2_fill_2 FILLER_42_347 ();
 sg13g2_fill_1 FILLER_42_349 ();
 sg13g2_decap_8 FILLER_42_369 ();
 sg13g2_decap_8 FILLER_42_376 ();
 sg13g2_decap_8 FILLER_42_383 ();
 sg13g2_decap_8 FILLER_42_390 ();
 sg13g2_decap_8 FILLER_42_397 ();
 sg13g2_decap_4 FILLER_42_404 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_2 ();
 sg13g2_fill_2 FILLER_43_72 ();
 sg13g2_fill_2 FILLER_43_83 ();
 sg13g2_fill_1 FILLER_43_85 ();
 sg13g2_fill_2 FILLER_43_131 ();
 sg13g2_fill_1 FILLER_43_133 ();
 sg13g2_fill_1 FILLER_43_143 ();
 sg13g2_fill_2 FILLER_43_157 ();
 sg13g2_fill_2 FILLER_43_194 ();
 sg13g2_fill_1 FILLER_43_231 ();
 sg13g2_fill_1 FILLER_43_255 ();
 sg13g2_fill_2 FILLER_43_270 ();
 sg13g2_fill_1 FILLER_43_272 ();
 sg13g2_decap_8 FILLER_43_376 ();
 sg13g2_decap_8 FILLER_43_383 ();
 sg13g2_decap_8 FILLER_43_390 ();
 sg13g2_decap_8 FILLER_43_397 ();
 sg13g2_decap_4 FILLER_43_404 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_27 ();
 sg13g2_fill_1 FILLER_44_69 ();
 sg13g2_fill_2 FILLER_44_82 ();
 sg13g2_fill_2 FILLER_44_115 ();
 sg13g2_fill_1 FILLER_44_133 ();
 sg13g2_fill_2 FILLER_44_160 ();
 sg13g2_fill_1 FILLER_44_162 ();
 sg13g2_fill_2 FILLER_44_172 ();
 sg13g2_fill_2 FILLER_44_183 ();
 sg13g2_fill_1 FILLER_44_203 ();
 sg13g2_decap_4 FILLER_44_291 ();
 sg13g2_fill_1 FILLER_44_322 ();
 sg13g2_decap_8 FILLER_44_386 ();
 sg13g2_decap_8 FILLER_44_393 ();
 sg13g2_decap_8 FILLER_44_400 ();
 sg13g2_fill_2 FILLER_44_407 ();
 sg13g2_fill_2 FILLER_45_88 ();
 sg13g2_fill_2 FILLER_45_162 ();
 sg13g2_fill_1 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_271 ();
 sg13g2_decap_8 FILLER_45_278 ();
 sg13g2_decap_8 FILLER_45_285 ();
 sg13g2_fill_1 FILLER_45_292 ();
 sg13g2_fill_2 FILLER_45_344 ();
 sg13g2_fill_1 FILLER_45_346 ();
 sg13g2_decap_8 FILLER_45_370 ();
 sg13g2_decap_8 FILLER_45_377 ();
 sg13g2_decap_8 FILLER_45_384 ();
 sg13g2_decap_8 FILLER_45_391 ();
 sg13g2_decap_8 FILLER_45_398 ();
 sg13g2_decap_4 FILLER_45_405 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_2 ();
 sg13g2_fill_2 FILLER_46_20 ();
 sg13g2_fill_1 FILLER_46_22 ();
 sg13g2_fill_1 FILLER_46_56 ();
 sg13g2_fill_2 FILLER_46_66 ();
 sg13g2_fill_1 FILLER_46_68 ();
 sg13g2_fill_2 FILLER_46_126 ();
 sg13g2_fill_1 FILLER_46_235 ();
 sg13g2_decap_8 FILLER_46_270 ();
 sg13g2_decap_8 FILLER_46_277 ();
 sg13g2_fill_2 FILLER_46_313 ();
 sg13g2_decap_8 FILLER_46_334 ();
 sg13g2_fill_2 FILLER_46_341 ();
 sg13g2_fill_1 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_361 ();
 sg13g2_decap_8 FILLER_46_368 ();
 sg13g2_decap_8 FILLER_46_375 ();
 sg13g2_decap_8 FILLER_46_382 ();
 sg13g2_decap_8 FILLER_46_389 ();
 sg13g2_decap_8 FILLER_46_396 ();
 sg13g2_decap_4 FILLER_46_403 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_fill_2 FILLER_47_26 ();
 sg13g2_fill_1 FILLER_47_28 ();
 sg13g2_fill_2 FILLER_47_38 ();
 sg13g2_fill_1 FILLER_47_40 ();
 sg13g2_fill_1 FILLER_47_50 ();
 sg13g2_fill_2 FILLER_47_102 ();
 sg13g2_fill_2 FILLER_47_167 ();
 sg13g2_fill_1 FILLER_47_169 ();
 sg13g2_fill_1 FILLER_47_205 ();
 sg13g2_fill_1 FILLER_47_214 ();
 sg13g2_fill_1 FILLER_47_254 ();
 sg13g2_fill_1 FILLER_47_327 ();
 sg13g2_decap_8 FILLER_47_333 ();
 sg13g2_decap_4 FILLER_47_340 ();
 sg13g2_fill_1 FILLER_47_344 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_fill_2 FILLER_47_406 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_49 ();
 sg13g2_fill_2 FILLER_48_72 ();
 sg13g2_fill_1 FILLER_48_74 ();
 sg13g2_fill_1 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_173 ();
 sg13g2_fill_2 FILLER_48_180 ();
 sg13g2_fill_1 FILLER_48_190 ();
 sg13g2_fill_2 FILLER_48_204 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_4 FILLER_48_217 ();
 sg13g2_fill_1 FILLER_48_221 ();
 sg13g2_fill_2 FILLER_48_242 ();
 sg13g2_fill_1 FILLER_48_244 ();
 sg13g2_fill_1 FILLER_48_276 ();
 sg13g2_fill_2 FILLER_48_331 ();
 sg13g2_fill_1 FILLER_48_333 ();
 sg13g2_decap_8 FILLER_48_391 ();
 sg13g2_decap_8 FILLER_48_398 ();
 sg13g2_decap_4 FILLER_48_405 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_27 ();
 sg13g2_fill_1 FILLER_49_85 ();
 sg13g2_fill_2 FILLER_49_128 ();
 sg13g2_fill_1 FILLER_49_136 ();
 sg13g2_decap_8 FILLER_49_172 ();
 sg13g2_decap_4 FILLER_49_179 ();
 sg13g2_fill_2 FILLER_49_183 ();
 sg13g2_fill_1 FILLER_49_190 ();
 sg13g2_fill_2 FILLER_49_210 ();
 sg13g2_decap_8 FILLER_49_221 ();
 sg13g2_fill_2 FILLER_49_228 ();
 sg13g2_fill_2 FILLER_49_234 ();
 sg13g2_fill_1 FILLER_49_236 ();
 sg13g2_fill_1 FILLER_49_304 ();
 sg13g2_fill_1 FILLER_49_314 ();
 sg13g2_fill_2 FILLER_49_325 ();
 sg13g2_fill_1 FILLER_49_327 ();
 sg13g2_fill_2 FILLER_49_354 ();
 sg13g2_fill_1 FILLER_49_356 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_decap_4 FILLER_49_403 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_fill_2 FILLER_50_28 ();
 sg13g2_fill_2 FILLER_50_71 ();
 sg13g2_fill_1 FILLER_50_73 ();
 sg13g2_fill_2 FILLER_50_100 ();
 sg13g2_fill_2 FILLER_50_154 ();
 sg13g2_fill_1 FILLER_50_156 ();
 sg13g2_fill_2 FILLER_50_166 ();
 sg13g2_fill_1 FILLER_50_168 ();
 sg13g2_decap_4 FILLER_50_181 ();
 sg13g2_fill_1 FILLER_50_185 ();
 sg13g2_fill_1 FILLER_50_192 ();
 sg13g2_fill_2 FILLER_50_254 ();
 sg13g2_fill_2 FILLER_50_261 ();
 sg13g2_fill_2 FILLER_50_271 ();
 sg13g2_fill_1 FILLER_50_273 ();
 sg13g2_decap_4 FILLER_50_279 ();
 sg13g2_fill_1 FILLER_50_313 ();
 sg13g2_decap_4 FILLER_50_327 ();
 sg13g2_fill_1 FILLER_50_331 ();
 sg13g2_fill_1 FILLER_50_337 ();
 sg13g2_fill_2 FILLER_50_342 ();
 sg13g2_fill_1 FILLER_50_344 ();
 sg13g2_fill_2 FILLER_50_353 ();
 sg13g2_fill_2 FILLER_50_359 ();
 sg13g2_fill_2 FILLER_50_366 ();
 sg13g2_fill_2 FILLER_50_376 ();
 sg13g2_decap_8 FILLER_50_388 ();
 sg13g2_decap_8 FILLER_50_395 ();
 sg13g2_decap_8 FILLER_50_402 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_27 ();
 sg13g2_fill_2 FILLER_51_131 ();
 sg13g2_decap_4 FILLER_51_174 ();
 sg13g2_fill_1 FILLER_51_178 ();
 sg13g2_fill_2 FILLER_51_199 ();
 sg13g2_decap_4 FILLER_51_229 ();
 sg13g2_fill_1 FILLER_51_233 ();
 sg13g2_fill_1 FILLER_51_238 ();
 sg13g2_decap_4 FILLER_51_243 ();
 sg13g2_fill_1 FILLER_51_247 ();
 sg13g2_fill_1 FILLER_51_256 ();
 sg13g2_fill_2 FILLER_51_279 ();
 sg13g2_fill_2 FILLER_51_336 ();
 sg13g2_fill_1 FILLER_51_338 ();
 sg13g2_decap_8 FILLER_51_343 ();
 sg13g2_decap_8 FILLER_51_350 ();
 sg13g2_decap_8 FILLER_51_357 ();
 sg13g2_decap_8 FILLER_51_364 ();
 sg13g2_decap_8 FILLER_51_371 ();
 sg13g2_decap_8 FILLER_51_378 ();
 sg13g2_decap_8 FILLER_51_385 ();
 sg13g2_decap_8 FILLER_51_392 ();
 sg13g2_decap_8 FILLER_51_399 ();
 sg13g2_fill_2 FILLER_51_406 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_fill_1 FILLER_52_31 ();
 sg13g2_fill_1 FILLER_52_106 ();
 sg13g2_fill_2 FILLER_52_201 ();
 sg13g2_fill_1 FILLER_52_203 ();
 sg13g2_fill_2 FILLER_52_213 ();
 sg13g2_fill_2 FILLER_52_221 ();
 sg13g2_fill_2 FILLER_52_277 ();
 sg13g2_fill_1 FILLER_52_279 ();
 sg13g2_fill_1 FILLER_52_306 ();
 sg13g2_fill_1 FILLER_52_362 ();
 sg13g2_decap_8 FILLER_52_368 ();
 sg13g2_decap_4 FILLER_52_375 ();
 sg13g2_decap_8 FILLER_52_384 ();
 sg13g2_decap_8 FILLER_52_391 ();
 sg13g2_decap_8 FILLER_52_398 ();
 sg13g2_decap_4 FILLER_52_405 ();
 sg13g2_fill_1 FILLER_53_45 ();
 sg13g2_fill_2 FILLER_53_92 ();
 sg13g2_fill_1 FILLER_53_107 ();
 sg13g2_fill_2 FILLER_53_128 ();
 sg13g2_fill_1 FILLER_53_158 ();
 sg13g2_decap_4 FILLER_53_177 ();
 sg13g2_fill_2 FILLER_53_181 ();
 sg13g2_fill_2 FILLER_53_189 ();
 sg13g2_fill_1 FILLER_53_191 ();
 sg13g2_decap_8 FILLER_53_239 ();
 sg13g2_decap_4 FILLER_53_246 ();
 sg13g2_fill_2 FILLER_53_250 ();
 sg13g2_fill_2 FILLER_53_257 ();
 sg13g2_fill_1 FILLER_53_259 ();
 sg13g2_fill_2 FILLER_53_273 ();
 sg13g2_fill_2 FILLER_53_284 ();
 sg13g2_decap_4 FILLER_53_324 ();
 sg13g2_fill_2 FILLER_53_373 ();
 sg13g2_fill_1 FILLER_53_375 ();
 sg13g2_fill_1 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_49 ();
 sg13g2_fill_1 FILLER_54_132 ();
 sg13g2_fill_2 FILLER_54_147 ();
 sg13g2_fill_1 FILLER_54_149 ();
 sg13g2_decap_8 FILLER_54_176 ();
 sg13g2_decap_8 FILLER_54_183 ();
 sg13g2_decap_8 FILLER_54_199 ();
 sg13g2_fill_2 FILLER_54_206 ();
 sg13g2_fill_1 FILLER_54_217 ();
 sg13g2_fill_2 FILLER_54_222 ();
 sg13g2_fill_1 FILLER_54_224 ();
 sg13g2_fill_2 FILLER_54_251 ();
 sg13g2_fill_2 FILLER_54_258 ();
 sg13g2_fill_1 FILLER_54_352 ();
 sg13g2_fill_2 FILLER_55_42 ();
 sg13g2_fill_2 FILLER_55_53 ();
 sg13g2_fill_1 FILLER_55_55 ();
 sg13g2_fill_2 FILLER_55_91 ();
 sg13g2_fill_1 FILLER_55_93 ();
 sg13g2_fill_2 FILLER_55_120 ();
 sg13g2_fill_2 FILLER_55_173 ();
 sg13g2_fill_1 FILLER_55_175 ();
 sg13g2_decap_8 FILLER_55_181 ();
 sg13g2_fill_1 FILLER_55_188 ();
 sg13g2_fill_1 FILLER_55_199 ();
 sg13g2_decap_4 FILLER_55_206 ();
 sg13g2_fill_1 FILLER_55_210 ();
 sg13g2_fill_1 FILLER_55_219 ();
 sg13g2_fill_2 FILLER_55_226 ();
 sg13g2_decap_8 FILLER_55_240 ();
 sg13g2_decap_8 FILLER_55_247 ();
 sg13g2_fill_1 FILLER_55_284 ();
 sg13g2_decap_8 FILLER_55_331 ();
 sg13g2_decap_4 FILLER_55_338 ();
 sg13g2_fill_1 FILLER_55_350 ();
 sg13g2_fill_2 FILLER_55_371 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_2 ();
 sg13g2_fill_2 FILLER_56_34 ();
 sg13g2_fill_2 FILLER_56_106 ();
 sg13g2_fill_1 FILLER_56_108 ();
 sg13g2_fill_2 FILLER_56_134 ();
 sg13g2_fill_1 FILLER_56_136 ();
 sg13g2_fill_2 FILLER_56_142 ();
 sg13g2_fill_2 FILLER_56_153 ();
 sg13g2_fill_1 FILLER_56_155 ();
 sg13g2_fill_2 FILLER_56_165 ();
 sg13g2_fill_1 FILLER_56_167 ();
 sg13g2_fill_1 FILLER_56_179 ();
 sg13g2_decap_8 FILLER_56_192 ();
 sg13g2_decap_4 FILLER_56_199 ();
 sg13g2_fill_1 FILLER_56_240 ();
 sg13g2_fill_2 FILLER_56_248 ();
 sg13g2_fill_1 FILLER_56_250 ();
 sg13g2_fill_2 FILLER_56_259 ();
 sg13g2_decap_4 FILLER_56_326 ();
 sg13g2_fill_2 FILLER_56_356 ();
 sg13g2_fill_1 FILLER_56_358 ();
 sg13g2_fill_1 FILLER_56_372 ();
 sg13g2_fill_2 FILLER_56_378 ();
 sg13g2_decap_8 FILLER_56_398 ();
 sg13g2_decap_4 FILLER_56_405 ();
 sg13g2_fill_1 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_31 ();
 sg13g2_fill_1 FILLER_57_33 ();
 sg13g2_fill_1 FILLER_57_138 ();
 sg13g2_fill_2 FILLER_57_172 ();
 sg13g2_fill_1 FILLER_57_174 ();
 sg13g2_fill_2 FILLER_57_205 ();
 sg13g2_fill_2 FILLER_57_227 ();
 sg13g2_fill_1 FILLER_57_229 ();
 sg13g2_fill_2 FILLER_57_328 ();
 sg13g2_decap_8 FILLER_57_361 ();
 sg13g2_decap_8 FILLER_57_368 ();
 sg13g2_fill_2 FILLER_57_375 ();
 sg13g2_fill_1 FILLER_57_377 ();
 sg13g2_fill_2 FILLER_57_385 ();
 sg13g2_fill_1 FILLER_57_387 ();
 sg13g2_decap_8 FILLER_57_391 ();
 sg13g2_decap_8 FILLER_57_398 ();
 sg13g2_decap_4 FILLER_57_405 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_56 ();
 sg13g2_fill_2 FILLER_58_79 ();
 sg13g2_fill_1 FILLER_58_90 ();
 sg13g2_fill_1 FILLER_58_100 ();
 sg13g2_fill_1 FILLER_58_123 ();
 sg13g2_fill_1 FILLER_58_138 ();
 sg13g2_fill_2 FILLER_58_149 ();
 sg13g2_fill_1 FILLER_58_151 ();
 sg13g2_fill_2 FILLER_58_178 ();
 sg13g2_fill_1 FILLER_58_180 ();
 sg13g2_fill_1 FILLER_58_210 ();
 sg13g2_fill_2 FILLER_58_275 ();
 sg13g2_fill_1 FILLER_58_277 ();
 sg13g2_decap_8 FILLER_58_355 ();
 sg13g2_fill_2 FILLER_58_362 ();
 sg13g2_decap_4 FILLER_58_371 ();
 sg13g2_fill_1 FILLER_59_54 ();
 sg13g2_fill_2 FILLER_59_66 ();
 sg13g2_fill_1 FILLER_59_82 ();
 sg13g2_fill_1 FILLER_59_96 ();
 sg13g2_decap_8 FILLER_59_109 ();
 sg13g2_decap_4 FILLER_59_161 ();
 sg13g2_decap_8 FILLER_59_173 ();
 sg13g2_fill_1 FILLER_59_180 ();
 sg13g2_decap_4 FILLER_59_195 ();
 sg13g2_decap_8 FILLER_59_230 ();
 sg13g2_fill_1 FILLER_59_240 ();
 sg13g2_fill_1 FILLER_59_308 ();
 sg13g2_fill_2 FILLER_59_321 ();
 sg13g2_fill_2 FILLER_59_328 ();
 sg13g2_decap_8 FILLER_59_387 ();
 sg13g2_decap_8 FILLER_59_398 ();
 sg13g2_decap_4 FILLER_59_405 ();
 sg13g2_fill_1 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_32 ();
 sg13g2_fill_1 FILLER_60_52 ();
 sg13g2_fill_1 FILLER_60_74 ();
 sg13g2_fill_1 FILLER_60_87 ();
 sg13g2_fill_1 FILLER_60_134 ();
 sg13g2_fill_2 FILLER_60_140 ();
 sg13g2_decap_8 FILLER_60_174 ();
 sg13g2_decap_8 FILLER_60_181 ();
 sg13g2_decap_8 FILLER_60_188 ();
 sg13g2_decap_4 FILLER_60_195 ();
 sg13g2_fill_2 FILLER_60_199 ();
 sg13g2_decap_8 FILLER_60_206 ();
 sg13g2_fill_1 FILLER_60_213 ();
 sg13g2_decap_4 FILLER_60_234 ();
 sg13g2_fill_2 FILLER_60_238 ();
 sg13g2_decap_4 FILLER_60_244 ();
 sg13g2_fill_1 FILLER_60_302 ();
 sg13g2_fill_1 FILLER_60_320 ();
 sg13g2_decap_8 FILLER_60_333 ();
 sg13g2_decap_4 FILLER_60_348 ();
 sg13g2_fill_2 FILLER_60_352 ();
 sg13g2_fill_2 FILLER_60_359 ();
 sg13g2_fill_1 FILLER_60_361 ();
 sg13g2_fill_2 FILLER_60_367 ();
 sg13g2_fill_2 FILLER_60_374 ();
 sg13g2_fill_1 FILLER_60_376 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_fill_1 FILLER_61_16 ();
 sg13g2_fill_2 FILLER_61_122 ();
 sg13g2_fill_2 FILLER_61_157 ();
 sg13g2_decap_8 FILLER_61_180 ();
 sg13g2_fill_2 FILLER_61_187 ();
 sg13g2_decap_4 FILLER_61_202 ();
 sg13g2_fill_2 FILLER_61_206 ();
 sg13g2_fill_2 FILLER_61_236 ();
 sg13g2_fill_1 FILLER_61_238 ();
 sg13g2_fill_1 FILLER_61_288 ();
 sg13g2_fill_1 FILLER_61_303 ();
 sg13g2_decap_8 FILLER_61_336 ();
 sg13g2_decap_8 FILLER_61_343 ();
 sg13g2_decap_8 FILLER_61_350 ();
 sg13g2_decap_8 FILLER_61_357 ();
 sg13g2_fill_1 FILLER_61_364 ();
 sg13g2_decap_4 FILLER_61_379 ();
 sg13g2_fill_1 FILLER_62_48 ();
 sg13g2_fill_1 FILLER_62_100 ();
 sg13g2_decap_4 FILLER_62_181 ();
 sg13g2_fill_1 FILLER_62_185 ();
 sg13g2_fill_2 FILLER_62_214 ();
 sg13g2_fill_2 FILLER_62_227 ();
 sg13g2_fill_1 FILLER_62_229 ();
 sg13g2_decap_8 FILLER_62_338 ();
 sg13g2_decap_8 FILLER_62_345 ();
 sg13g2_decap_8 FILLER_62_352 ();
 sg13g2_decap_8 FILLER_62_359 ();
 sg13g2_decap_8 FILLER_62_366 ();
 sg13g2_decap_8 FILLER_62_373 ();
 sg13g2_decap_8 FILLER_62_380 ();
 sg13g2_fill_2 FILLER_62_391 ();
 sg13g2_fill_1 FILLER_62_393 ();
 sg13g2_decap_4 FILLER_62_403 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_2 ();
 sg13g2_fill_1 FILLER_63_52 ();
 sg13g2_fill_1 FILLER_63_58 ();
 sg13g2_fill_1 FILLER_63_78 ();
 sg13g2_fill_2 FILLER_63_135 ();
 sg13g2_fill_2 FILLER_63_155 ();
 sg13g2_fill_1 FILLER_63_175 ();
 sg13g2_fill_2 FILLER_63_181 ();
 sg13g2_fill_1 FILLER_63_187 ();
 sg13g2_fill_2 FILLER_63_193 ();
 sg13g2_fill_1 FILLER_63_195 ();
 sg13g2_fill_2 FILLER_63_219 ();
 sg13g2_fill_1 FILLER_63_221 ();
 sg13g2_fill_2 FILLER_63_228 ();
 sg13g2_fill_1 FILLER_63_230 ();
 sg13g2_fill_2 FILLER_63_253 ();
 sg13g2_decap_4 FILLER_63_340 ();
 sg13g2_fill_2 FILLER_63_344 ();
 sg13g2_fill_2 FILLER_63_351 ();
 sg13g2_fill_1 FILLER_63_353 ();
 sg13g2_fill_2 FILLER_63_358 ();
 sg13g2_fill_1 FILLER_63_360 ();
 sg13g2_decap_8 FILLER_63_365 ();
 sg13g2_fill_2 FILLER_63_372 ();
 sg13g2_fill_1 FILLER_63_374 ();
 sg13g2_decap_8 FILLER_63_380 ();
 sg13g2_fill_1 FILLER_63_387 ();
 sg13g2_decap_8 FILLER_63_392 ();
 sg13g2_decap_8 FILLER_63_399 ();
 sg13g2_fill_2 FILLER_63_406 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_fill_1 FILLER_64_126 ();
 sg13g2_fill_1 FILLER_64_141 ();
 sg13g2_fill_1 FILLER_64_156 ();
 sg13g2_fill_2 FILLER_64_186 ();
 sg13g2_fill_2 FILLER_64_202 ();
 sg13g2_fill_1 FILLER_64_204 ();
 sg13g2_fill_2 FILLER_64_210 ();
 sg13g2_fill_1 FILLER_64_212 ();
 sg13g2_fill_2 FILLER_64_227 ();
 sg13g2_fill_1 FILLER_64_240 ();
 sg13g2_fill_2 FILLER_64_246 ();
 sg13g2_fill_1 FILLER_64_248 ();
 sg13g2_fill_1 FILLER_64_267 ();
 sg13g2_decap_8 FILLER_64_333 ();
 sg13g2_fill_2 FILLER_64_340 ();
 sg13g2_fill_1 FILLER_64_342 ();
 sg13g2_decap_4 FILLER_64_403 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_fill_1 FILLER_65_49 ();
 sg13g2_fill_1 FILLER_65_89 ();
 sg13g2_fill_2 FILLER_65_134 ();
 sg13g2_fill_2 FILLER_65_193 ();
 sg13g2_fill_1 FILLER_65_195 ();
 sg13g2_fill_2 FILLER_65_203 ();
 sg13g2_fill_2 FILLER_65_211 ();
 sg13g2_fill_1 FILLER_65_213 ();
 sg13g2_fill_2 FILLER_65_224 ();
 sg13g2_fill_1 FILLER_65_240 ();
 sg13g2_fill_2 FILLER_65_252 ();
 sg13g2_fill_1 FILLER_65_272 ();
 sg13g2_fill_1 FILLER_65_290 ();
 sg13g2_fill_2 FILLER_65_318 ();
 sg13g2_decap_8 FILLER_65_324 ();
 sg13g2_decap_4 FILLER_65_331 ();
 sg13g2_fill_1 FILLER_65_335 ();
 sg13g2_fill_1 FILLER_65_357 ();
 sg13g2_fill_2 FILLER_65_363 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_28 ();
 sg13g2_fill_2 FILLER_66_53 ();
 sg13g2_fill_2 FILLER_66_73 ();
 sg13g2_fill_1 FILLER_66_106 ();
 sg13g2_fill_2 FILLER_66_112 ();
 sg13g2_fill_1 FILLER_66_161 ();
 sg13g2_fill_2 FILLER_66_173 ();
 sg13g2_fill_1 FILLER_66_235 ();
 sg13g2_fill_2 FILLER_66_288 ();
 sg13g2_fill_1 FILLER_66_290 ();
 sg13g2_decap_4 FILLER_66_295 ();
 sg13g2_decap_8 FILLER_66_303 ();
 sg13g2_decap_8 FILLER_66_310 ();
 sg13g2_decap_8 FILLER_66_317 ();
 sg13g2_decap_8 FILLER_66_324 ();
 sg13g2_fill_1 FILLER_66_331 ();
 sg13g2_fill_2 FILLER_66_337 ();
 sg13g2_fill_1 FILLER_66_366 ();
 sg13g2_fill_1 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_83 ();
 sg13g2_fill_1 FILLER_67_85 ();
 sg13g2_fill_2 FILLER_67_111 ();
 sg13g2_fill_1 FILLER_67_113 ();
 sg13g2_fill_1 FILLER_67_127 ();
 sg13g2_fill_1 FILLER_67_223 ();
 sg13g2_fill_2 FILLER_67_259 ();
 sg13g2_fill_2 FILLER_67_270 ();
 sg13g2_fill_1 FILLER_67_272 ();
 sg13g2_fill_2 FILLER_67_277 ();
 sg13g2_fill_1 FILLER_67_284 ();
 sg13g2_fill_1 FILLER_67_324 ();
 sg13g2_decap_8 FILLER_67_349 ();
 sg13g2_fill_2 FILLER_67_356 ();
 sg13g2_fill_1 FILLER_67_358 ();
 sg13g2_fill_2 FILLER_67_363 ();
 sg13g2_fill_1 FILLER_67_365 ();
 sg13g2_fill_2 FILLER_67_376 ();
 sg13g2_decap_4 FILLER_67_382 ();
 sg13g2_fill_1 FILLER_67_386 ();
 sg13g2_fill_2 FILLER_67_395 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_83 ();
 sg13g2_fill_1 FILLER_68_121 ();
 sg13g2_fill_1 FILLER_68_127 ();
 sg13g2_fill_1 FILLER_68_133 ();
 sg13g2_fill_2 FILLER_68_186 ();
 sg13g2_fill_1 FILLER_68_188 ();
 sg13g2_fill_2 FILLER_68_198 ();
 sg13g2_fill_1 FILLER_68_200 ();
 sg13g2_decap_8 FILLER_68_220 ();
 sg13g2_fill_2 FILLER_68_236 ();
 sg13g2_fill_2 FILLER_68_247 ();
 sg13g2_fill_1 FILLER_68_249 ();
 sg13g2_decap_8 FILLER_68_325 ();
 sg13g2_decap_8 FILLER_68_332 ();
 sg13g2_decap_4 FILLER_68_339 ();
 sg13g2_fill_2 FILLER_68_343 ();
 sg13g2_fill_2 FILLER_68_350 ();
 sg13g2_fill_1 FILLER_68_352 ();
 sg13g2_fill_2 FILLER_68_358 ();
 sg13g2_fill_1 FILLER_68_360 ();
 sg13g2_decap_8 FILLER_68_375 ();
 sg13g2_decap_8 FILLER_68_382 ();
 sg13g2_decap_8 FILLER_68_389 ();
 sg13g2_decap_8 FILLER_68_396 ();
 sg13g2_decap_4 FILLER_68_403 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_fill_1 FILLER_69_26 ();
 sg13g2_fill_2 FILLER_69_93 ();
 sg13g2_fill_1 FILLER_69_164 ();
 sg13g2_fill_1 FILLER_69_195 ();
 sg13g2_fill_2 FILLER_69_205 ();
 sg13g2_fill_1 FILLER_69_207 ();
 sg13g2_fill_1 FILLER_69_217 ();
 sg13g2_decap_8 FILLER_69_223 ();
 sg13g2_decap_8 FILLER_69_230 ();
 sg13g2_decap_8 FILLER_69_237 ();
 sg13g2_decap_4 FILLER_69_244 ();
 sg13g2_fill_1 FILLER_69_248 ();
 sg13g2_fill_2 FILLER_69_298 ();
 sg13g2_fill_1 FILLER_69_300 ();
 sg13g2_fill_2 FILLER_69_305 ();
 sg13g2_fill_2 FILLER_69_323 ();
 sg13g2_fill_1 FILLER_69_325 ();
 sg13g2_fill_1 FILLER_69_368 ();
 sg13g2_fill_1 FILLER_69_381 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_fill_2 FILLER_70_60 ();
 sg13g2_fill_1 FILLER_70_62 ();
 sg13g2_fill_1 FILLER_70_107 ();
 sg13g2_fill_2 FILLER_70_117 ();
 sg13g2_fill_2 FILLER_70_132 ();
 sg13g2_fill_2 FILLER_70_151 ();
 sg13g2_fill_1 FILLER_70_165 ();
 sg13g2_fill_2 FILLER_70_196 ();
 sg13g2_fill_1 FILLER_70_198 ();
 sg13g2_fill_2 FILLER_70_223 ();
 sg13g2_decap_8 FILLER_70_244 ();
 sg13g2_decap_4 FILLER_70_251 ();
 sg13g2_fill_1 FILLER_70_255 ();
 sg13g2_decap_8 FILLER_70_284 ();
 sg13g2_decap_8 FILLER_70_291 ();
 sg13g2_fill_2 FILLER_70_298 ();
 sg13g2_fill_1 FILLER_70_300 ();
 sg13g2_decap_8 FILLER_70_305 ();
 sg13g2_decap_8 FILLER_70_312 ();
 sg13g2_decap_8 FILLER_70_319 ();
 sg13g2_decap_8 FILLER_70_326 ();
 sg13g2_fill_2 FILLER_70_341 ();
 sg13g2_fill_1 FILLER_70_343 ();
 sg13g2_fill_2 FILLER_70_358 ();
 sg13g2_fill_1 FILLER_70_360 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_fill_2 FILLER_71_25 ();
 sg13g2_fill_1 FILLER_71_27 ();
 sg13g2_fill_1 FILLER_71_43 ();
 sg13g2_fill_1 FILLER_71_65 ();
 sg13g2_fill_2 FILLER_71_98 ();
 sg13g2_fill_1 FILLER_71_106 ();
 sg13g2_fill_1 FILLER_71_113 ();
 sg13g2_fill_2 FILLER_71_167 ();
 sg13g2_fill_1 FILLER_71_169 ();
 sg13g2_fill_2 FILLER_71_188 ();
 sg13g2_fill_2 FILLER_71_200 ();
 sg13g2_decap_4 FILLER_71_261 ();
 sg13g2_decap_4 FILLER_71_270 ();
 sg13g2_fill_2 FILLER_71_274 ();
 sg13g2_decap_8 FILLER_71_281 ();
 sg13g2_decap_8 FILLER_71_288 ();
 sg13g2_decap_8 FILLER_71_295 ();
 sg13g2_decap_8 FILLER_71_309 ();
 sg13g2_decap_8 FILLER_71_316 ();
 sg13g2_decap_8 FILLER_71_323 ();
 sg13g2_decap_8 FILLER_71_333 ();
 sg13g2_decap_4 FILLER_71_340 ();
 sg13g2_decap_8 FILLER_71_348 ();
 sg13g2_fill_2 FILLER_71_355 ();
 sg13g2_fill_2 FILLER_71_361 ();
 sg13g2_fill_1 FILLER_71_363 ();
 sg13g2_decap_8 FILLER_71_379 ();
 sg13g2_decap_4 FILLER_71_386 ();
 sg13g2_fill_2 FILLER_71_390 ();
 sg13g2_decap_8 FILLER_71_400 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_fill_1 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_63 ();
 sg13g2_fill_2 FILLER_72_80 ();
 sg13g2_fill_1 FILLER_72_82 ();
 sg13g2_fill_1 FILLER_72_105 ();
 sg13g2_fill_2 FILLER_72_115 ();
 sg13g2_fill_2 FILLER_72_194 ();
 sg13g2_fill_1 FILLER_72_205 ();
 sg13g2_fill_1 FILLER_72_215 ();
 sg13g2_fill_2 FILLER_72_271 ();
 sg13g2_fill_1 FILLER_72_273 ();
 sg13g2_fill_2 FILLER_72_284 ();
 sg13g2_fill_1 FILLER_72_286 ();
 sg13g2_fill_2 FILLER_72_321 ();
 sg13g2_fill_1 FILLER_72_333 ();
 sg13g2_fill_1 FILLER_72_338 ();
 sg13g2_fill_2 FILLER_72_344 ();
 sg13g2_fill_1 FILLER_72_346 ();
 sg13g2_decap_8 FILLER_72_357 ();
 sg13g2_decap_8 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_371 ();
 sg13g2_decap_4 FILLER_72_378 ();
 sg13g2_fill_1 FILLER_72_382 ();
 sg13g2_fill_2 FILLER_73_38 ();
 sg13g2_fill_1 FILLER_73_40 ();
 sg13g2_fill_2 FILLER_73_189 ();
 sg13g2_fill_1 FILLER_73_191 ();
 sg13g2_fill_2 FILLER_73_224 ();
 sg13g2_decap_8 FILLER_73_257 ();
 sg13g2_decap_8 FILLER_73_264 ();
 sg13g2_decap_8 FILLER_73_271 ();
 sg13g2_decap_4 FILLER_73_282 ();
 sg13g2_fill_2 FILLER_73_286 ();
 sg13g2_fill_1 FILLER_73_314 ();
 sg13g2_fill_2 FILLER_73_362 ();
 sg13g2_fill_1 FILLER_73_364 ();
 sg13g2_fill_2 FILLER_73_391 ();
 sg13g2_fill_1 FILLER_73_393 ();
 sg13g2_decap_8 FILLER_73_398 ();
 sg13g2_decap_4 FILLER_73_405 ();
 sg13g2_fill_1 FILLER_74_26 ();
 sg13g2_fill_2 FILLER_74_42 ();
 sg13g2_fill_1 FILLER_74_164 ();
 sg13g2_decap_4 FILLER_74_243 ();
 sg13g2_decap_8 FILLER_74_251 ();
 sg13g2_decap_4 FILLER_74_258 ();
 sg13g2_decap_4 FILLER_74_266 ();
 sg13g2_fill_1 FILLER_74_270 ();
 sg13g2_decap_8 FILLER_74_286 ();
 sg13g2_decap_8 FILLER_74_308 ();
 sg13g2_decap_8 FILLER_74_320 ();
 sg13g2_fill_2 FILLER_74_327 ();
 sg13g2_fill_1 FILLER_74_329 ();
 sg13g2_decap_8 FILLER_74_350 ();
 sg13g2_decap_8 FILLER_74_363 ();
 sg13g2_decap_4 FILLER_74_370 ();
 sg13g2_decap_8 FILLER_74_383 ();
 sg13g2_decap_8 FILLER_74_390 ();
 sg13g2_decap_8 FILLER_74_397 ();
 sg13g2_decap_4 FILLER_74_404 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_fill_1 FILLER_75_38 ();
 sg13g2_fill_2 FILLER_75_48 ();
 sg13g2_fill_2 FILLER_75_135 ();
 sg13g2_fill_1 FILLER_75_154 ();
 sg13g2_fill_2 FILLER_75_168 ();
 sg13g2_fill_1 FILLER_75_170 ();
 sg13g2_fill_1 FILLER_75_184 ();
 sg13g2_fill_1 FILLER_75_198 ();
 sg13g2_decap_8 FILLER_75_234 ();
 sg13g2_fill_2 FILLER_75_241 ();
 sg13g2_fill_1 FILLER_75_243 ();
 sg13g2_decap_8 FILLER_75_249 ();
 sg13g2_fill_2 FILLER_75_256 ();
 sg13g2_decap_8 FILLER_75_288 ();
 sg13g2_decap_8 FILLER_75_295 ();
 sg13g2_decap_8 FILLER_75_302 ();
 sg13g2_decap_4 FILLER_75_309 ();
 sg13g2_fill_1 FILLER_75_327 ();
 sg13g2_fill_1 FILLER_75_341 ();
 sg13g2_fill_1 FILLER_75_351 ();
 sg13g2_fill_1 FILLER_75_364 ();
 sg13g2_fill_2 FILLER_76_72 ();
 sg13g2_fill_1 FILLER_76_74 ();
 sg13g2_fill_2 FILLER_76_130 ();
 sg13g2_fill_1 FILLER_76_220 ();
 sg13g2_decap_8 FILLER_76_229 ();
 sg13g2_decap_4 FILLER_76_236 ();
 sg13g2_fill_1 FILLER_76_240 ();
 sg13g2_fill_2 FILLER_76_272 ();
 sg13g2_decap_8 FILLER_76_284 ();
 sg13g2_decap_8 FILLER_76_291 ();
 sg13g2_fill_2 FILLER_76_298 ();
 sg13g2_decap_8 FILLER_76_307 ();
 sg13g2_fill_2 FILLER_76_347 ();
 sg13g2_fill_1 FILLER_76_349 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_fill_2 FILLER_76_392 ();
 sg13g2_decap_8 FILLER_76_398 ();
 sg13g2_decap_4 FILLER_76_405 ();
 sg13g2_fill_2 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_71 ();
 sg13g2_fill_2 FILLER_77_139 ();
 sg13g2_fill_1 FILLER_77_141 ();
 sg13g2_fill_2 FILLER_77_207 ();
 sg13g2_fill_1 FILLER_77_209 ();
 sg13g2_fill_2 FILLER_77_214 ();
 sg13g2_fill_1 FILLER_77_216 ();
 sg13g2_fill_2 FILLER_77_225 ();
 sg13g2_fill_2 FILLER_77_330 ();
 sg13g2_fill_1 FILLER_77_332 ();
 sg13g2_fill_2 FILLER_77_341 ();
 sg13g2_fill_1 FILLER_77_343 ();
 sg13g2_fill_2 FILLER_77_357 ();
 sg13g2_fill_1 FILLER_77_359 ();
 sg13g2_fill_2 FILLER_77_366 ();
 sg13g2_fill_1 FILLER_77_368 ();
 sg13g2_fill_2 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_152 ();
 sg13g2_fill_1 FILLER_78_225 ();
 sg13g2_decap_4 FILLER_78_268 ();
 sg13g2_fill_2 FILLER_78_272 ();
 sg13g2_decap_4 FILLER_78_279 ();
 sg13g2_decap_4 FILLER_78_313 ();
 sg13g2_fill_1 FILLER_78_317 ();
 sg13g2_fill_2 FILLER_78_333 ();
 sg13g2_fill_2 FILLER_78_343 ();
 sg13g2_fill_1 FILLER_78_345 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_2 ();
 sg13g2_fill_2 FILLER_79_45 ();
 sg13g2_fill_1 FILLER_79_79 ();
 sg13g2_fill_1 FILLER_79_89 ();
 sg13g2_fill_1 FILLER_79_95 ();
 sg13g2_fill_1 FILLER_79_171 ();
 sg13g2_fill_1 FILLER_79_194 ();
 sg13g2_fill_1 FILLER_79_251 ();
 sg13g2_decap_8 FILLER_79_278 ();
 sg13g2_fill_1 FILLER_79_285 ();
 sg13g2_decap_8 FILLER_79_312 ();
 sg13g2_fill_2 FILLER_79_319 ();
 sg13g2_fill_1 FILLER_79_321 ();
 sg13g2_decap_4 FILLER_79_346 ();
 sg13g2_fill_2 FILLER_79_358 ();
 sg13g2_fill_1 FILLER_79_360 ();
 sg13g2_decap_8 FILLER_79_370 ();
 sg13g2_decap_8 FILLER_79_377 ();
 sg13g2_fill_2 FILLER_79_384 ();
 sg13g2_fill_1 FILLER_79_386 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_2 ();
 sg13g2_fill_1 FILLER_80_32 ();
 sg13g2_fill_2 FILLER_80_57 ();
 sg13g2_fill_1 FILLER_80_73 ();
 sg13g2_fill_1 FILLER_80_106 ();
 sg13g2_fill_1 FILLER_80_134 ();
 sg13g2_fill_2 FILLER_80_153 ();
 sg13g2_fill_1 FILLER_80_155 ();
 sg13g2_fill_2 FILLER_80_197 ();
 sg13g2_decap_8 FILLER_80_245 ();
 sg13g2_decap_8 FILLER_80_252 ();
 sg13g2_decap_4 FILLER_80_259 ();
 sg13g2_decap_8 FILLER_80_267 ();
 sg13g2_decap_4 FILLER_80_274 ();
 sg13g2_fill_2 FILLER_80_278 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_fill_2 FILLER_80_292 ();
 sg13g2_fill_2 FILLER_80_302 ();
 sg13g2_decap_8 FILLER_80_309 ();
 sg13g2_decap_8 FILLER_80_316 ();
 sg13g2_decap_8 FILLER_80_323 ();
 sg13g2_decap_8 FILLER_80_330 ();
 sg13g2_decap_8 FILLER_80_337 ();
 sg13g2_decap_8 FILLER_80_344 ();
 sg13g2_fill_1 FILLER_80_351 ();
 sg13g2_fill_2 FILLER_80_357 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_decap_8 FILLER_80_373 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[1] = net311;
 assign uio_oe[6] = net312;
 assign uio_oe[7] = net313;
endmodule

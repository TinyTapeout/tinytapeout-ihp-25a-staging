VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_torurstrom_async_lock
  CLASS BLOCK ;
  FOREIGN tt_um_torurstrom_async_lock ;
  ORIGIN 0.000 0.000 ;
  SIZE 202.080 BY 154.980 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 21.580 3.560 23.780 151.420 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 60.450 3.560 62.650 151.420 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 99.320 3.560 101.520 151.420 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 138.190 3.560 140.390 151.420 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 177.060 3.560 179.260 151.420 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 15.380 3.560 17.580 151.420 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 54.250 3.560 56.450 151.420 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 93.120 3.560 95.320 151.420 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 131.990 3.560 134.190 151.420 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 170.860 3.560 173.060 151.420 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 187.050 153.980 187.350 154.980 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 190.890 153.980 191.190 154.980 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 183.210 153.980 183.510 154.980 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal5 ;
        RECT 179.370 153.980 179.670 154.980 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal5 ;
        RECT 175.530 153.980 175.830 154.980 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal5 ;
        RECT 171.690 153.980 171.990 154.980 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal5 ;
        RECT 167.850 153.980 168.150 154.980 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal5 ;
        RECT 164.010 153.980 164.310 154.980 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal5 ;
        RECT 160.170 153.980 160.470 154.980 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal5 ;
        RECT 156.330 153.980 156.630 154.980 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal5 ;
        RECT 152.490 153.980 152.790 154.980 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 148.650 153.980 148.950 154.980 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 144.810 153.980 145.110 154.980 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 140.970 153.980 141.270 154.980 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 137.130 153.980 137.430 154.980 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 133.290 153.980 133.590 154.980 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 129.450 153.980 129.750 154.980 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 125.610 153.980 125.910 154.980 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 121.770 153.980 122.070 154.980 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 56.490 153.980 56.790 154.980 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 52.650 153.980 52.950 154.980 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 48.810 153.980 49.110 154.980 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 44.970 153.980 45.270 154.980 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 41.130 153.980 41.430 154.980 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 37.290 153.980 37.590 154.980 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 33.450 153.980 33.750 154.980 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 29.610 153.980 29.910 154.980 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 87.210 153.980 87.510 154.980 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 83.370 153.980 83.670 154.980 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 79.530 153.980 79.830 154.980 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 75.690 153.980 75.990 154.980 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 71.850 153.980 72.150 154.980 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 68.010 153.980 68.310 154.980 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 64.170 153.980 64.470 154.980 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 60.330 153.980 60.630 154.980 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434200 ;
    ANTENNADIFFAREA 0.706800 ;
    PORT
      LAYER Metal5 ;
        RECT 117.930 153.980 118.230 154.980 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434200 ;
    ANTENNADIFFAREA 0.706800 ;
    PORT
      LAYER Metal5 ;
        RECT 114.090 153.980 114.390 154.980 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434200 ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal5 ;
        RECT 110.250 153.980 110.550 154.980 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434200 ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal5 ;
        RECT 106.410 153.980 106.710 154.980 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434200 ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal5 ;
        RECT 102.570 153.980 102.870 154.980 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434200 ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal5 ;
        RECT 98.730 153.980 99.030 154.980 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434200 ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal5 ;
        RECT 94.890 153.980 95.190 154.980 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434200 ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal5 ;
        RECT 91.050 153.980 91.350 154.980 ;
    END
  END uo_out[7]
  OBS
      LAYER GatPoly ;
        RECT 2.880 3.630 199.200 151.350 ;
      LAYER Metal1 ;
        RECT 2.880 3.560 199.200 151.420 ;
      LAYER Metal2 ;
        RECT 15.515 3.680 181.105 152.140 ;
      LAYER Metal3 ;
        RECT 15.560 3.635 181.060 152.185 ;
      LAYER Metal4 ;
        RECT 15.515 3.680 181.105 152.140 ;
      LAYER Metal5 ;
        RECT 30.120 153.770 33.240 153.980 ;
        RECT 33.960 153.770 37.080 153.980 ;
        RECT 37.800 153.770 40.920 153.980 ;
        RECT 41.640 153.770 44.760 153.980 ;
        RECT 45.480 153.770 48.600 153.980 ;
        RECT 49.320 153.770 52.440 153.980 ;
        RECT 53.160 153.770 56.280 153.980 ;
        RECT 57.000 153.770 60.120 153.980 ;
        RECT 60.840 153.770 63.960 153.980 ;
        RECT 64.680 153.770 67.800 153.980 ;
        RECT 68.520 153.770 71.640 153.980 ;
        RECT 72.360 153.770 75.480 153.980 ;
        RECT 76.200 153.770 79.320 153.980 ;
        RECT 80.040 153.770 83.160 153.980 ;
        RECT 83.880 153.770 87.000 153.980 ;
        RECT 87.720 153.770 90.840 153.980 ;
        RECT 91.560 153.770 94.680 153.980 ;
        RECT 95.400 153.770 98.520 153.980 ;
        RECT 99.240 153.770 102.360 153.980 ;
        RECT 103.080 153.770 106.200 153.980 ;
        RECT 106.920 153.770 110.040 153.980 ;
        RECT 110.760 153.770 113.880 153.980 ;
        RECT 114.600 153.770 117.720 153.980 ;
        RECT 118.440 153.770 121.560 153.980 ;
        RECT 122.280 153.770 125.400 153.980 ;
        RECT 126.120 153.770 129.240 153.980 ;
        RECT 129.960 153.770 133.080 153.980 ;
        RECT 133.800 153.770 136.920 153.980 ;
        RECT 137.640 153.770 140.760 153.980 ;
        RECT 141.480 153.770 144.600 153.980 ;
        RECT 145.320 153.770 148.440 153.980 ;
        RECT 149.160 153.770 152.280 153.980 ;
        RECT 153.000 153.770 156.120 153.980 ;
        RECT 156.840 153.770 159.960 153.980 ;
        RECT 160.680 153.770 163.800 153.980 ;
        RECT 164.520 153.770 167.640 153.980 ;
        RECT 168.360 153.770 171.480 153.980 ;
        RECT 172.200 153.770 175.320 153.980 ;
        RECT 176.040 153.770 179.160 153.980 ;
        RECT 29.660 151.630 179.620 153.770 ;
        RECT 29.660 126.275 54.040 151.630 ;
        RECT 56.660 126.275 60.240 151.630 ;
        RECT 62.860 126.275 92.910 151.630 ;
        RECT 95.530 126.275 99.110 151.630 ;
        RECT 101.730 126.275 131.780 151.630 ;
        RECT 134.400 126.275 137.980 151.630 ;
        RECT 140.600 126.275 170.650 151.630 ;
        RECT 173.270 126.275 176.850 151.630 ;
        RECT 179.470 126.275 179.620 151.630 ;
  END
END tt_um_torurstrom_async_lock
END LIBRARY


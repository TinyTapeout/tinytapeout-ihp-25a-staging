module tt_um_rejunity_sn76489 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net252;
 wire \chan[0].attenuation.control[0] ;
 wire \chan[0].attenuation.control[1] ;
 wire \chan[0].attenuation.control[2] ;
 wire \chan[0].attenuation.control[3] ;
 wire \chan[0].attenuation.in ;
 wire \chan[1].attenuation.control[0] ;
 wire \chan[1].attenuation.control[1] ;
 wire \chan[1].attenuation.control[2] ;
 wire \chan[1].attenuation.control[3] ;
 wire \chan[1].attenuation.in ;
 wire \chan[2].attenuation.control[0] ;
 wire \chan[2].attenuation.control[1] ;
 wire \chan[2].attenuation.control[2] ;
 wire \chan[2].attenuation.control[3] ;
 wire \chan[2].attenuation.in ;
 wire \chan[3].attenuation.control[0] ;
 wire \chan[3].attenuation.control[1] ;
 wire \chan[3].attenuation.control[2] ;
 wire \chan[3].attenuation.control[3] ;
 wire \chan[3].attenuation.in ;
 wire \clk_counter[0] ;
 wire \clk_counter[1] ;
 wire \clk_counter[2] ;
 wire \clk_counter[3] ;
 wire \clk_counter[4] ;
 wire \clk_counter[5] ;
 wire \clk_counter[6] ;
 wire \control_noise[0][0] ;
 wire \control_noise[0][1] ;
 wire \control_noise[0][2] ;
 wire \control_tone_freq[0][0] ;
 wire \control_tone_freq[0][1] ;
 wire \control_tone_freq[0][2] ;
 wire \control_tone_freq[0][3] ;
 wire \control_tone_freq[0][4] ;
 wire \control_tone_freq[0][5] ;
 wire \control_tone_freq[0][6] ;
 wire \control_tone_freq[0][7] ;
 wire \control_tone_freq[0][8] ;
 wire \control_tone_freq[0][9] ;
 wire \control_tone_freq[1][0] ;
 wire \control_tone_freq[1][1] ;
 wire \control_tone_freq[1][2] ;
 wire \control_tone_freq[1][3] ;
 wire \control_tone_freq[1][4] ;
 wire \control_tone_freq[1][5] ;
 wire \control_tone_freq[1][6] ;
 wire \control_tone_freq[1][7] ;
 wire \control_tone_freq[1][8] ;
 wire \control_tone_freq[1][9] ;
 wire \control_tone_freq[2][0] ;
 wire \control_tone_freq[2][1] ;
 wire \control_tone_freq[2][2] ;
 wire \control_tone_freq[2][3] ;
 wire \control_tone_freq[2][4] ;
 wire \control_tone_freq[2][5] ;
 wire \control_tone_freq[2][6] ;
 wire \control_tone_freq[2][7] ;
 wire \control_tone_freq[2][8] ;
 wire \control_tone_freq[2][9] ;
 wire \genblk4[0].pwm.accumulator[0] ;
 wire \genblk4[0].pwm.accumulator[10] ;
 wire \genblk4[0].pwm.accumulator[1] ;
 wire \genblk4[0].pwm.accumulator[2] ;
 wire \genblk4[0].pwm.accumulator[3] ;
 wire \genblk4[0].pwm.accumulator[4] ;
 wire \genblk4[0].pwm.accumulator[5] ;
 wire \genblk4[0].pwm.accumulator[6] ;
 wire \genblk4[0].pwm.accumulator[7] ;
 wire \genblk4[0].pwm.accumulator[8] ;
 wire \genblk4[0].pwm.accumulator[9] ;
 wire \genblk4[1].pwm.accumulator[0] ;
 wire \genblk4[1].pwm.accumulator[10] ;
 wire \genblk4[1].pwm.accumulator[1] ;
 wire \genblk4[1].pwm.accumulator[2] ;
 wire \genblk4[1].pwm.accumulator[3] ;
 wire \genblk4[1].pwm.accumulator[4] ;
 wire \genblk4[1].pwm.accumulator[5] ;
 wire \genblk4[1].pwm.accumulator[6] ;
 wire \genblk4[1].pwm.accumulator[7] ;
 wire \genblk4[1].pwm.accumulator[8] ;
 wire \genblk4[1].pwm.accumulator[9] ;
 wire \genblk4[2].pwm.accumulator[0] ;
 wire \genblk4[2].pwm.accumulator[10] ;
 wire \genblk4[2].pwm.accumulator[1] ;
 wire \genblk4[2].pwm.accumulator[2] ;
 wire \genblk4[2].pwm.accumulator[3] ;
 wire \genblk4[2].pwm.accumulator[4] ;
 wire \genblk4[2].pwm.accumulator[5] ;
 wire \genblk4[2].pwm.accumulator[6] ;
 wire \genblk4[2].pwm.accumulator[7] ;
 wire \genblk4[2].pwm.accumulator[8] ;
 wire \genblk4[2].pwm.accumulator[9] ;
 wire \genblk4[3].pwm.accumulator[0] ;
 wire \genblk4[3].pwm.accumulator[10] ;
 wire \genblk4[3].pwm.accumulator[1] ;
 wire \genblk4[3].pwm.accumulator[2] ;
 wire \genblk4[3].pwm.accumulator[3] ;
 wire \genblk4[3].pwm.accumulator[4] ;
 wire \genblk4[3].pwm.accumulator[5] ;
 wire \genblk4[3].pwm.accumulator[6] ;
 wire \genblk4[3].pwm.accumulator[7] ;
 wire \genblk4[3].pwm.accumulator[8] ;
 wire \genblk4[3].pwm.accumulator[9] ;
 wire \latch_control_reg[0] ;
 wire \latch_control_reg[1] ;
 wire \latch_control_reg[2] ;
 wire \noise[0].gen.counter[0] ;
 wire \noise[0].gen.counter[1] ;
 wire \noise[0].gen.counter[2] ;
 wire \noise[0].gen.counter[3] ;
 wire \noise[0].gen.counter[4] ;
 wire \noise[0].gen.counter[5] ;
 wire \noise[0].gen.counter[6] ;
 wire \noise[0].gen.lfsr[10] ;
 wire \noise[0].gen.lfsr[11] ;
 wire \noise[0].gen.lfsr[12] ;
 wire \noise[0].gen.lfsr[13] ;
 wire \noise[0].gen.lfsr[14] ;
 wire \noise[0].gen.lfsr[1] ;
 wire \noise[0].gen.lfsr[2] ;
 wire \noise[0].gen.lfsr[3] ;
 wire \noise[0].gen.lfsr[4] ;
 wire \noise[0].gen.lfsr[5] ;
 wire \noise[0].gen.lfsr[6] ;
 wire \noise[0].gen.lfsr[7] ;
 wire \noise[0].gen.lfsr[8] ;
 wire \noise[0].gen.lfsr[9] ;
 wire \noise[0].gen.restart_noise ;
 wire \noise[0].gen.signal_edge.previous_signal_state_0 ;
 wire \pwm.accumulator[0] ;
 wire \pwm.accumulator[10] ;
 wire \pwm.accumulator[11] ;
 wire \pwm.accumulator[12] ;
 wire \pwm.accumulator[1] ;
 wire \pwm.accumulator[2] ;
 wire \pwm.accumulator[3] ;
 wire \pwm.accumulator[4] ;
 wire \pwm.accumulator[5] ;
 wire \pwm.accumulator[6] ;
 wire \pwm.accumulator[7] ;
 wire \pwm.accumulator[8] ;
 wire \pwm.accumulator[9] ;
 wire \tone[0].gen.counter[0] ;
 wire \tone[0].gen.counter[1] ;
 wire \tone[0].gen.counter[2] ;
 wire \tone[0].gen.counter[3] ;
 wire \tone[0].gen.counter[4] ;
 wire \tone[0].gen.counter[5] ;
 wire \tone[0].gen.counter[6] ;
 wire \tone[0].gen.counter[7] ;
 wire \tone[0].gen.counter[8] ;
 wire \tone[0].gen.counter[9] ;
 wire \tone[1].gen.counter[0] ;
 wire \tone[1].gen.counter[1] ;
 wire \tone[1].gen.counter[2] ;
 wire \tone[1].gen.counter[3] ;
 wire \tone[1].gen.counter[4] ;
 wire \tone[1].gen.counter[5] ;
 wire \tone[1].gen.counter[6] ;
 wire \tone[1].gen.counter[7] ;
 wire \tone[1].gen.counter[8] ;
 wire \tone[1].gen.counter[9] ;
 wire \tone[2].gen.counter[0] ;
 wire \tone[2].gen.counter[1] ;
 wire \tone[2].gen.counter[2] ;
 wire \tone[2].gen.counter[3] ;
 wire \tone[2].gen.counter[4] ;
 wire \tone[2].gen.counter[5] ;
 wire \tone[2].gen.counter[6] ;
 wire \tone[2].gen.counter[7] ;
 wire \tone[2].gen.counter[8] ;
 wire \tone[2].gen.counter[9] ;
 wire net13;
 wire net14;
 wire net15;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire clknet_0_clk;
 wire net16;
 wire net17;
 wire net18;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;

 sg13g2_inv_1 _1362_ (.Y(_0478_),
    .A(net297));
 sg13g2_inv_4 _1363_ (.A(net4),
    .Y(_0479_));
 sg13g2_inv_1 _1364_ (.Y(_0480_),
    .A(net271));
 sg13g2_inv_4 _1365_ (.A(net3),
    .Y(_0481_));
 sg13g2_inv_1 _1366_ (.Y(_0482_),
    .A(net268));
 sg13g2_inv_2 _1367_ (.Y(_0483_),
    .A(net2));
 sg13g2_inv_2 _1368_ (.Y(_0484_),
    .A(net1));
 sg13g2_inv_1 _1369_ (.Y(_0485_),
    .A(net344));
 sg13g2_inv_1 _1370_ (.Y(_0486_),
    .A(net332));
 sg13g2_inv_1 _1371_ (.Y(_0487_),
    .A(net422));
 sg13g2_inv_1 _1372_ (.Y(_0488_),
    .A(net258));
 sg13g2_inv_1 _1373_ (.Y(_0489_),
    .A(net343));
 sg13g2_inv_1 _1374_ (.Y(_0490_),
    .A(net345));
 sg13g2_inv_1 _1375_ (.Y(_0491_),
    .A(net260));
 sg13g2_inv_1 _1376_ (.Y(_0492_),
    .A(net336));
 sg13g2_inv_1 _1377_ (.Y(_0493_),
    .A(net262));
 sg13g2_inv_1 _1378_ (.Y(_0494_),
    .A(net306));
 sg13g2_inv_1 _1379_ (.Y(_0495_),
    .A(net264));
 sg13g2_inv_1 _1380_ (.Y(_0496_),
    .A(net310));
 sg13g2_inv_1 _1381_ (.Y(_0497_),
    .A(net362));
 sg13g2_inv_1 _1382_ (.Y(_0498_),
    .A(net269));
 sg13g2_inv_1 _1383_ (.Y(_0499_),
    .A(net6));
 sg13g2_inv_1 _1384_ (.Y(_0500_),
    .A(net292));
 sg13g2_inv_1 _1385_ (.Y(_0501_),
    .A(net5));
 sg13g2_inv_1 _1386_ (.Y(_0502_),
    .A(net295));
 sg13g2_inv_1 _1387_ (.Y(_0503_),
    .A(net284));
 sg13g2_inv_1 _1388_ (.Y(_0504_),
    .A(net290));
 sg13g2_inv_1 _1389_ (.Y(_0505_),
    .A(net330));
 sg13g2_inv_1 _1390_ (.Y(_0506_),
    .A(net294));
 sg13g2_inv_1 _1391_ (.Y(_0507_),
    .A(net334));
 sg13g2_inv_1 _1392_ (.Y(_0508_),
    .A(net320));
 sg13g2_inv_1 _1393_ (.Y(_0509_),
    .A(net276));
 sg13g2_inv_1 _1394_ (.Y(_0510_),
    .A(net281));
 sg13g2_inv_1 _1395_ (.Y(_0511_),
    .A(net279));
 sg13g2_inv_1 _1396_ (.Y(_0512_),
    .A(net298));
 sg13g2_inv_1 _1397_ (.Y(_0513_),
    .A(net266));
 sg13g2_inv_1 _1398_ (.Y(_0514_),
    .A(net277));
 sg13g2_inv_1 _1399_ (.Y(_0515_),
    .A(net286));
 sg13g2_inv_1 _1400_ (.Y(_0516_),
    .A(net272));
 sg13g2_inv_1 _1401_ (.Y(_0517_),
    .A(net283));
 sg13g2_inv_1 _1402_ (.Y(_0518_),
    .A(\chan[3].attenuation.control[2] ));
 sg13g2_inv_1 _1403_ (.Y(_0519_),
    .A(\chan[2].attenuation.control[1] ));
 sg13g2_inv_1 _1404_ (.Y(_0520_),
    .A(\chan[1].attenuation.control[3] ));
 sg13g2_inv_1 _1405_ (.Y(_0521_),
    .A(\chan[1].attenuation.control[2] ));
 sg13g2_inv_1 _1406_ (.Y(_0522_),
    .A(\chan[1].attenuation.control[0] ));
 sg13g2_inv_1 _1407_ (.Y(_0523_),
    .A(\chan[0].attenuation.control[2] ));
 sg13g2_inv_1 _1408_ (.Y(_0524_),
    .A(net443));
 sg13g2_inv_1 _1409_ (.Y(_0525_),
    .A(net11));
 sg13g2_inv_1 _1410_ (.Y(_0526_),
    .A(net352));
 sg13g2_inv_1 _1411_ (.Y(_0527_),
    .A(net244));
 sg13g2_inv_1 _1412_ (.Y(_0528_),
    .A(_0004_));
 sg13g2_inv_1 _1413_ (.Y(_0529_),
    .A(net267));
 sg13g2_inv_1 _1414_ (.Y(_0530_),
    .A(net505));
 sg13g2_inv_1 _1415_ (.Y(_0531_),
    .A(\genblk4[2].pwm.accumulator[4] ));
 sg13g2_inv_1 _1416_ (.Y(_0532_),
    .A(net450));
 sg13g2_inv_1 _1417_ (.Y(_0533_),
    .A(net278));
 sg13g2_nor2b_2 _1418_ (.A(\chan[0].attenuation.control[3] ),
    .B_N(net221),
    .Y(_0534_));
 sg13g2_nand2b_2 _1419_ (.Y(_0535_),
    .B(\chan[0].attenuation.in ),
    .A_N(\chan[0].attenuation.control[3] ));
 sg13g2_nor2b_2 _1420_ (.A(\chan[0].attenuation.control[2] ),
    .B_N(net221),
    .Y(_0536_));
 sg13g2_nor2b_1 _1421_ (.A(\chan[0].attenuation.control[1] ),
    .B_N(net221),
    .Y(_0537_));
 sg13g2_nand2b_1 _1422_ (.Y(_0538_),
    .B(net221),
    .A_N(\chan[0].attenuation.control[1] ));
 sg13g2_a221oi_1 _1423_ (.B2(_0537_),
    .C1(_0534_),
    .B1(net223),
    .A1(net221),
    .Y(_0539_),
    .A2(_0523_));
 sg13g2_nand2_1 _1424_ (.Y(_0540_),
    .A(net223),
    .B(_0536_));
 sg13g2_a221oi_1 _1425_ (.B2(net223),
    .C1(_0539_),
    .B1(_0536_),
    .A1(\chan[0].attenuation.control[1] ),
    .Y(_0541_),
    .A2(_0534_));
 sg13g2_nor2b_2 _1426_ (.A(\chan[1].attenuation.control[2] ),
    .B_N(\chan[1].attenuation.in ),
    .Y(_0542_));
 sg13g2_nand3b_1 _1427_ (.B(\chan[1].attenuation.control[0] ),
    .C(net220),
    .Y(_0543_),
    .A_N(\chan[1].attenuation.control[2] ));
 sg13g2_xnor2_1 _1428_ (.Y(_0544_),
    .A(\chan[1].attenuation.control[0] ),
    .B(_0542_));
 sg13g2_nor2b_1 _1429_ (.A(\chan[1].attenuation.control[1] ),
    .B_N(net220),
    .Y(_0545_));
 sg13g2_or2_1 _1430_ (.X(_0546_),
    .B(_0545_),
    .A(_0542_));
 sg13g2_nor2b_1 _1431_ (.A(\chan[1].attenuation.control[3] ),
    .B_N(net220),
    .Y(_0547_));
 sg13g2_nand2b_2 _1432_ (.Y(_0548_),
    .B(net220),
    .A_N(\chan[1].attenuation.control[3] ));
 sg13g2_o21ai_1 _1433_ (.B1(\chan[1].attenuation.control[3] ),
    .Y(_0549_),
    .A1(_0542_),
    .A2(net216));
 sg13g2_and2_1 _1434_ (.A(_0543_),
    .B(_0547_),
    .X(_0550_));
 sg13g2_nand3b_1 _1435_ (.B(_0543_),
    .C(_0547_),
    .Y(_0551_),
    .A_N(\chan[1].attenuation.control[1] ));
 sg13g2_o21ai_1 _1436_ (.B1(_0551_),
    .Y(_0552_),
    .A1(_0544_),
    .A2(_0549_));
 sg13g2_nand2_1 _1437_ (.Y(_0553_),
    .A(_0541_),
    .B(_0552_));
 sg13g2_nor2b_2 _1438_ (.A(net222),
    .B_N(net219),
    .Y(_0554_));
 sg13g2_nand2b_1 _1439_ (.Y(_0555_),
    .B(net218),
    .A_N(net222));
 sg13g2_nand2b_2 _1440_ (.Y(_0556_),
    .B(net218),
    .A_N(\chan[2].attenuation.control[1] ));
 sg13g2_nand2_2 _1441_ (.Y(_0557_),
    .A(_0555_),
    .B(_0556_));
 sg13g2_nor2b_2 _1442_ (.A(\chan[2].attenuation.control[3] ),
    .B_N(net218),
    .Y(_0558_));
 sg13g2_nand2b_2 _1443_ (.Y(_0559_),
    .B(net219),
    .A_N(\chan[2].attenuation.control[3] ));
 sg13g2_nor2b_2 _1444_ (.A(\chan[2].attenuation.control[0] ),
    .B_N(net218),
    .Y(_0560_));
 sg13g2_and2_1 _1445_ (.A(net222),
    .B(_0560_),
    .X(_0561_));
 sg13g2_nand3b_1 _1446_ (.B(net222),
    .C(net218),
    .Y(_0562_),
    .A_N(\chan[2].attenuation.control[0] ));
 sg13g2_nand3b_1 _1447_ (.B(\chan[2].attenuation.control[0] ),
    .C(net218),
    .Y(_0563_),
    .A_N(net222));
 sg13g2_nand3_1 _1448_ (.B(_0562_),
    .C(_0563_),
    .A(_0559_),
    .Y(_0564_));
 sg13g2_nor2_2 _1449_ (.A(\chan[2].attenuation.control[0] ),
    .B(_0556_),
    .Y(_0565_));
 sg13g2_nand3_1 _1450_ (.B(_0558_),
    .C(_0560_),
    .A(_0519_),
    .Y(_0566_));
 sg13g2_nand3b_1 _1451_ (.B(net222),
    .C(net218),
    .Y(_0567_),
    .A_N(\chan[2].attenuation.control[3] ));
 sg13g2_and2_1 _1452_ (.A(_0566_),
    .B(_0567_),
    .X(_0568_));
 sg13g2_nand3_1 _1453_ (.B(_0566_),
    .C(_0567_),
    .A(_0564_),
    .Y(_0569_));
 sg13g2_nand2_2 _1454_ (.Y(_0570_),
    .A(_0557_),
    .B(_0569_));
 sg13g2_xnor2_1 _1455_ (.Y(_0571_),
    .A(_0541_),
    .B(_0552_));
 sg13g2_o21ai_1 _1456_ (.B1(_0553_),
    .Y(_0572_),
    .A1(_0570_),
    .A2(_0571_));
 sg13g2_a21oi_2 _1457_ (.B1(_0560_),
    .Y(_0573_),
    .A2(_0519_),
    .A1(net218));
 sg13g2_nor3_1 _1458_ (.A(_0554_),
    .B(_0565_),
    .C(_0573_),
    .Y(_0574_));
 sg13g2_o21ai_1 _1459_ (.B1(_0567_),
    .Y(_0575_),
    .A1(\chan[2].attenuation.control[1] ),
    .A2(_0559_));
 sg13g2_a21oi_1 _1460_ (.A1(\chan[2].attenuation.control[1] ),
    .A2(_0560_),
    .Y(_0576_),
    .B1(_0575_));
 sg13g2_nor2_2 _1461_ (.A(_0574_),
    .B(_0576_),
    .Y(_0577_));
 sg13g2_nand2_2 _1462_ (.Y(_0578_),
    .A(\chan[0].attenuation.control[1] ),
    .B(\chan[0].attenuation.control[0] ));
 sg13g2_and3_1 _1463_ (.X(_0579_),
    .A(net221),
    .B(\chan[0].attenuation.control[2] ),
    .C(_0578_));
 sg13g2_nand3_1 _1464_ (.B(\chan[0].attenuation.control[2] ),
    .C(_0578_),
    .A(net221),
    .Y(_0580_));
 sg13g2_nor2_1 _1465_ (.A(net223),
    .B(_0538_),
    .Y(_0581_));
 sg13g2_nand2b_1 _1466_ (.Y(_0582_),
    .B(_0537_),
    .A_N(net223));
 sg13g2_a21oi_2 _1467_ (.B1(_0535_),
    .Y(_0583_),
    .A2(_0536_),
    .A1(\chan[0].attenuation.control[1] ));
 sg13g2_a21o_1 _1468_ (.A2(_0536_),
    .A1(\chan[0].attenuation.control[1] ),
    .B1(_0535_),
    .X(_0584_));
 sg13g2_nand3b_1 _1469_ (.B(_0536_),
    .C(\chan[0].attenuation.control[1] ),
    .Y(_0585_),
    .A_N(net223));
 sg13g2_a22oi_1 _1470_ (.Y(_0586_),
    .B1(_0584_),
    .B2(_0585_),
    .A2(_0582_),
    .A1(_0579_));
 sg13g2_a21o_1 _1471_ (.A2(_0522_),
    .A1(net220),
    .B1(net216),
    .X(_0587_));
 sg13g2_and2_1 _1472_ (.A(_0522_),
    .B(net216),
    .X(_0588_));
 sg13g2_a21oi_1 _1473_ (.A1(_0522_),
    .A2(net216),
    .Y(_0589_),
    .B1(_0542_));
 sg13g2_nand3_1 _1474_ (.B(\chan[1].attenuation.control[1] ),
    .C(_0522_),
    .A(net220),
    .Y(_0590_));
 sg13g2_a21o_1 _1475_ (.A2(_0542_),
    .A1(\chan[1].attenuation.control[1] ),
    .B1(_0548_),
    .X(_0591_));
 sg13g2_a22oi_1 _1476_ (.Y(_0592_),
    .B1(_0590_),
    .B2(_0591_),
    .A2(_0589_),
    .A1(_0587_));
 sg13g2_and2_1 _1477_ (.A(_0586_),
    .B(_0592_),
    .X(_0593_));
 sg13g2_or2_1 _1478_ (.X(_0594_),
    .B(_0592_),
    .A(_0586_));
 sg13g2_xor2_1 _1479_ (.B(_0592_),
    .A(_0586_),
    .X(_0595_));
 sg13g2_xnor2_1 _1480_ (.Y(_0596_),
    .A(_0577_),
    .B(_0595_));
 sg13g2_nand2b_1 _1481_ (.Y(_0597_),
    .B(_0572_),
    .A_N(_0596_));
 sg13g2_nor2b_1 _1482_ (.A(\chan[3].attenuation.control[1] ),
    .B_N(\chan[3].attenuation.in ),
    .Y(_0598_));
 sg13g2_nand2b_1 _1483_ (.Y(_0599_),
    .B(net217),
    .A_N(\chan[3].attenuation.control[1] ));
 sg13g2_nand2b_1 _1484_ (.Y(_0600_),
    .B(net217),
    .A_N(\chan[3].attenuation.control[0] ));
 sg13g2_nand2_1 _1485_ (.Y(_0601_),
    .A(_0599_),
    .B(_0600_));
 sg13g2_nor2b_2 _1486_ (.A(\chan[3].attenuation.control[2] ),
    .B_N(net217),
    .Y(_0602_));
 sg13g2_a21oi_2 _1487_ (.B1(_0518_),
    .Y(_0603_),
    .A2(_0600_),
    .A1(_0599_));
 sg13g2_nand2b_2 _1488_ (.Y(_0604_),
    .B(_0598_),
    .A_N(\chan[3].attenuation.control[0] ));
 sg13g2_nand2_1 _1489_ (.Y(_0605_),
    .A(_0603_),
    .B(_0604_));
 sg13g2_nor2b_2 _1490_ (.A(\chan[3].attenuation.control[3] ),
    .B_N(net217),
    .Y(_0606_));
 sg13g2_nand2b_2 _1491_ (.Y(_0607_),
    .B(net217),
    .A_N(\chan[3].attenuation.control[3] ));
 sg13g2_a21oi_1 _1492_ (.A1(\chan[3].attenuation.control[1] ),
    .A2(_0602_),
    .Y(_0608_),
    .B1(_0607_));
 sg13g2_inv_1 _1493_ (.Y(_0609_),
    .A(_0608_));
 sg13g2_nand3b_1 _1494_ (.B(_0602_),
    .C(\chan[3].attenuation.control[1] ),
    .Y(_0610_),
    .A_N(\chan[3].attenuation.control[0] ));
 sg13g2_a22oi_1 _1495_ (.Y(_0611_),
    .B1(_0609_),
    .B2(_0610_),
    .A2(_0604_),
    .A1(_0603_));
 sg13g2_inv_1 _1496_ (.Y(_0612_),
    .A(_0611_));
 sg13g2_xor2_1 _1497_ (.B(_0596_),
    .A(_0572_),
    .X(_0613_));
 sg13g2_o21ai_1 _1498_ (.B1(_0597_),
    .Y(_0614_),
    .A1(_0612_),
    .A2(_0613_));
 sg13g2_a21oi_2 _1499_ (.B1(_0593_),
    .Y(_0615_),
    .A2(_0594_),
    .A1(_0577_));
 sg13g2_nor2_1 _1500_ (.A(\chan[2].attenuation.control[1] ),
    .B(_0555_),
    .Y(_0616_));
 sg13g2_mux2_1 _1501_ (.A0(net222),
    .A1(_0554_),
    .S(_0556_),
    .X(_0617_));
 sg13g2_a21oi_1 _1502_ (.A1(_0559_),
    .A2(_0562_),
    .Y(_0618_),
    .B1(_0617_));
 sg13g2_o21ai_1 _1503_ (.B1(_0618_),
    .Y(_0619_),
    .A1(\chan[2].attenuation.control[0] ),
    .A2(_0567_));
 sg13g2_inv_1 _1504_ (.Y(_0620_),
    .A(_0619_));
 sg13g2_a22oi_1 _1505_ (.Y(_0621_),
    .B1(net216),
    .B2(\chan[1].attenuation.control[2] ),
    .A2(_0542_),
    .A1(\chan[1].attenuation.control[1] ));
 sg13g2_o21ai_1 _1506_ (.B1(_0621_),
    .Y(_0622_),
    .A1(\chan[1].attenuation.control[3] ),
    .A2(_0590_));
 sg13g2_a21oi_2 _1507_ (.B1(_0622_),
    .Y(_0623_),
    .A2(_0590_),
    .A1(_0548_));
 sg13g2_and3_1 _1508_ (.X(_0624_),
    .A(net221),
    .B(\chan[0].attenuation.control[3] ),
    .C(_0578_));
 sg13g2_nor2_1 _1509_ (.A(_0523_),
    .B(_0537_),
    .Y(_0625_));
 sg13g2_a22oi_1 _1510_ (.Y(_0626_),
    .B1(_0624_),
    .B2(_0625_),
    .A2(_0583_),
    .A1(_0580_));
 sg13g2_inv_1 _1511_ (.Y(_0627_),
    .A(_0626_));
 sg13g2_and2_1 _1512_ (.A(_0623_),
    .B(_0627_),
    .X(_0628_));
 sg13g2_xnor2_1 _1513_ (.Y(_0629_),
    .A(_0623_),
    .B(_0626_));
 sg13g2_xnor2_1 _1514_ (.Y(_0630_),
    .A(_0619_),
    .B(_0629_));
 sg13g2_nor2b_1 _1515_ (.A(_0615_),
    .B_N(_0630_),
    .Y(_0631_));
 sg13g2_xnor2_1 _1516_ (.Y(_0632_),
    .A(_0615_),
    .B(_0630_));
 sg13g2_nor2_1 _1517_ (.A(_0603_),
    .B(_0609_),
    .Y(_0633_));
 sg13g2_or2_1 _1518_ (.X(_0634_),
    .B(_0602_),
    .A(_0598_));
 sg13g2_nor2_1 _1519_ (.A(_0606_),
    .B(_0634_),
    .Y(_0635_));
 sg13g2_a21oi_2 _1520_ (.B1(_0633_),
    .Y(_0636_),
    .A2(_0635_),
    .A1(_0603_));
 sg13g2_inv_1 _1521_ (.Y(_0637_),
    .A(_0636_));
 sg13g2_xnor2_1 _1522_ (.Y(_0638_),
    .A(_0632_),
    .B(_0636_));
 sg13g2_nand2_1 _1523_ (.Y(_0639_),
    .A(_0614_),
    .B(_0638_));
 sg13g2_a21oi_1 _1524_ (.A1(_0523_),
    .A2(_0624_),
    .Y(_0640_),
    .B1(_0539_));
 sg13g2_mux2_1 _1525_ (.A0(_0538_),
    .A1(net223),
    .S(_0536_),
    .X(_0641_));
 sg13g2_a221oi_1 _1526_ (.B2(_0534_),
    .C1(_0539_),
    .B1(_0641_),
    .A1(_0523_),
    .Y(_0642_),
    .A2(_0624_));
 sg13g2_and2_1 _1527_ (.A(_0521_),
    .B(net216),
    .X(_0643_));
 sg13g2_a221oi_1 _1528_ (.B2(net216),
    .C1(_0522_),
    .B1(_0521_),
    .A1(net220),
    .Y(_0644_),
    .A2(_0520_));
 sg13g2_or2_1 _1529_ (.X(_0645_),
    .B(_0644_),
    .A(_0550_));
 sg13g2_o21ai_1 _1530_ (.B1(\chan[1].attenuation.control[0] ),
    .Y(_0646_),
    .A1(_0542_),
    .A2(net216));
 sg13g2_o21ai_1 _1531_ (.B1(_0548_),
    .Y(_0647_),
    .A1(_0643_),
    .A2(_0646_));
 sg13g2_o21ai_1 _1532_ (.B1(_0546_),
    .Y(_0648_),
    .A1(_0550_),
    .A2(_0644_));
 sg13g2_and3_1 _1533_ (.X(_0649_),
    .A(_0546_),
    .B(_0642_),
    .C(_0645_));
 sg13g2_nor2_1 _1534_ (.A(_0558_),
    .B(_0616_),
    .Y(_0650_));
 sg13g2_and2_1 _1535_ (.A(\chan[2].attenuation.control[0] ),
    .B(_0559_),
    .X(_0651_));
 sg13g2_a22oi_1 _1536_ (.Y(_0652_),
    .B1(_0617_),
    .B2(_0651_),
    .A2(_0565_),
    .A1(_0558_));
 sg13g2_nor2_2 _1537_ (.A(net428),
    .B(_0559_),
    .Y(_0653_));
 sg13g2_nand3b_1 _1538_ (.B(_0557_),
    .C(_0563_),
    .Y(_0654_),
    .A_N(\chan[2].attenuation.control[3] ));
 sg13g2_nand2_2 _1539_ (.Y(_0655_),
    .A(_0652_),
    .B(_0654_));
 sg13g2_xnor2_1 _1540_ (.Y(_0656_),
    .A(_0642_),
    .B(_0648_));
 sg13g2_a21oi_1 _1541_ (.A1(_0655_),
    .A2(_0656_),
    .Y(_0657_),
    .B1(_0649_));
 sg13g2_xnor2_1 _1542_ (.Y(_0658_),
    .A(_0570_),
    .B(_0571_));
 sg13g2_nor2_1 _1543_ (.A(_0657_),
    .B(_0658_),
    .Y(_0659_));
 sg13g2_a221oi_1 _1544_ (.B2(_0598_),
    .C1(_0606_),
    .B1(\chan[3].attenuation.control[0] ),
    .A1(net217),
    .Y(_0660_),
    .A2(_0518_));
 sg13g2_inv_1 _1545_ (.Y(_0661_),
    .A(_0660_));
 sg13g2_nand2_1 _1546_ (.Y(_0662_),
    .A(\chan[3].attenuation.control[0] ),
    .B(_0602_));
 sg13g2_a221oi_1 _1547_ (.B2(\chan[3].attenuation.control[1] ),
    .C1(_0660_),
    .B1(_0606_),
    .A1(\chan[3].attenuation.control[0] ),
    .Y(_0663_),
    .A2(_0602_));
 sg13g2_xor2_1 _1548_ (.B(_0658_),
    .A(_0657_),
    .X(_0664_));
 sg13g2_a21oi_1 _1549_ (.A1(_0663_),
    .A2(_0664_),
    .Y(_0665_),
    .B1(_0659_));
 sg13g2_xnor2_1 _1550_ (.Y(_0666_),
    .A(_0612_),
    .B(_0613_));
 sg13g2_nor2_1 _1551_ (.A(_0665_),
    .B(_0666_),
    .Y(_0667_));
 sg13g2_nand3_1 _1552_ (.B(_0518_),
    .C(_0601_),
    .A(\chan[3].attenuation.control[3] ),
    .Y(_0668_));
 sg13g2_a21o_1 _1553_ (.A2(_0662_),
    .A1(_0634_),
    .B1(_0607_),
    .X(_0669_));
 sg13g2_nand3_1 _1554_ (.B(_0668_),
    .C(_0669_),
    .A(_0661_),
    .Y(_0670_));
 sg13g2_xnor2_1 _1555_ (.Y(_0671_),
    .A(_0655_),
    .B(_0656_));
 sg13g2_nor2_1 _1556_ (.A(_0670_),
    .B(_0671_),
    .Y(_0672_));
 sg13g2_xor2_1 _1557_ (.B(_0664_),
    .A(_0663_),
    .X(_0673_));
 sg13g2_and2_1 _1558_ (.A(_0672_),
    .B(_0673_),
    .X(_0674_));
 sg13g2_xor2_1 _1559_ (.B(_0666_),
    .A(_0665_),
    .X(_0675_));
 sg13g2_a21oi_1 _1560_ (.A1(_0674_),
    .A2(_0675_),
    .Y(_0676_),
    .B1(_0667_));
 sg13g2_nor2_1 _1561_ (.A(_0614_),
    .B(_0638_),
    .Y(_0677_));
 sg13g2_xor2_1 _1562_ (.B(_0638_),
    .A(_0614_),
    .X(_0678_));
 sg13g2_o21ai_1 _1563_ (.B1(_0639_),
    .Y(_0679_),
    .A1(_0676_),
    .A2(_0677_));
 sg13g2_nand2_1 _1564_ (.Y(_0680_),
    .A(_0604_),
    .B(_0606_));
 sg13g2_nand3_1 _1565_ (.B(_0668_),
    .C(_0680_),
    .A(_0661_),
    .Y(_0681_));
 sg13g2_inv_1 _1566_ (.Y(_0682_),
    .A(_0681_));
 sg13g2_a21oi_2 _1567_ (.B1(_0628_),
    .Y(_0683_),
    .A2(_0629_),
    .A1(_0620_));
 sg13g2_o21ai_1 _1568_ (.B1(_0640_),
    .Y(_0684_),
    .A1(_0535_),
    .A2(_0581_));
 sg13g2_inv_1 _1569_ (.Y(_0685_),
    .A(_0684_));
 sg13g2_o21ai_1 _1570_ (.B1(_0647_),
    .Y(_0686_),
    .A1(_0548_),
    .A2(_0588_));
 sg13g2_or2_1 _1571_ (.X(_0687_),
    .B(_0686_),
    .A(_0684_));
 sg13g2_xnor2_1 _1572_ (.Y(_0688_),
    .A(_0684_),
    .B(_0686_));
 sg13g2_xnor2_1 _1573_ (.Y(_0689_),
    .A(_0652_),
    .B(_0688_));
 sg13g2_or2_1 _1574_ (.X(_0690_),
    .B(_0689_),
    .A(_0683_));
 sg13g2_xnor2_1 _1575_ (.Y(_0691_),
    .A(_0683_),
    .B(_0689_));
 sg13g2_xnor2_1 _1576_ (.Y(_0692_),
    .A(_0682_),
    .B(_0691_));
 sg13g2_a21oi_2 _1577_ (.B1(_0631_),
    .Y(_0693_),
    .A2(_0637_),
    .A1(_0632_));
 sg13g2_nor2b_1 _1578_ (.A(_0693_),
    .B_N(_0692_),
    .Y(_0694_));
 sg13g2_xnor2_1 _1579_ (.Y(_0695_),
    .A(_0692_),
    .B(_0693_));
 sg13g2_xor2_1 _1580_ (.B(_0695_),
    .A(_0679_),
    .X(uo_out[0]));
 sg13g2_a21oi_1 _1581_ (.A1(_0679_),
    .A2(_0695_),
    .Y(_0696_),
    .B1(_0694_));
 sg13g2_o21ai_1 _1582_ (.B1(_0690_),
    .Y(_0697_),
    .A1(_0681_),
    .A2(_0691_));
 sg13g2_o21ai_1 _1583_ (.B1(_0687_),
    .Y(_0698_),
    .A1(_0652_),
    .A2(_0688_));
 sg13g2_nor2_1 _1584_ (.A(\chan[0].attenuation.control[2] ),
    .B(_0538_),
    .Y(_0699_));
 sg13g2_nand2_1 _1585_ (.Y(_0700_),
    .A(_0582_),
    .B(_0624_));
 sg13g2_xnor2_1 _1586_ (.Y(_0701_),
    .A(_0699_),
    .B(_0700_));
 sg13g2_nand3b_1 _1587_ (.B(\chan[1].attenuation.control[3] ),
    .C(_0587_),
    .Y(_0702_),
    .A_N(_0588_));
 sg13g2_xnor2_1 _1588_ (.Y(_0703_),
    .A(_0643_),
    .B(_0702_));
 sg13g2_and2_1 _1589_ (.A(_0701_),
    .B(_0703_),
    .X(_0704_));
 sg13g2_xor2_1 _1590_ (.B(_0703_),
    .A(_0701_),
    .X(_0705_));
 sg13g2_nor3_1 _1591_ (.A(_0558_),
    .B(_0565_),
    .C(_0573_),
    .Y(_0706_));
 sg13g2_xnor2_1 _1592_ (.Y(_0707_),
    .A(_0616_),
    .B(_0706_));
 sg13g2_inv_1 _1593_ (.Y(_0708_),
    .A(_0707_));
 sg13g2_xnor2_1 _1594_ (.Y(_0709_),
    .A(_0705_),
    .B(_0707_));
 sg13g2_and2_1 _1595_ (.A(_0698_),
    .B(_0709_),
    .X(_0710_));
 sg13g2_xnor2_1 _1596_ (.Y(_0711_),
    .A(_0698_),
    .B(_0709_));
 sg13g2_nor2_1 _1597_ (.A(\chan[3].attenuation.control[2] ),
    .B(_0599_),
    .Y(_0712_));
 sg13g2_nand3_1 _1598_ (.B(_0601_),
    .C(_0604_),
    .A(\chan[3].attenuation.control[3] ),
    .Y(_0713_));
 sg13g2_xnor2_1 _1599_ (.Y(_0714_),
    .A(_0712_),
    .B(_0713_));
 sg13g2_nor2b_1 _1600_ (.A(_0711_),
    .B_N(_0714_),
    .Y(_0715_));
 sg13g2_xnor2_1 _1601_ (.Y(_0716_),
    .A(_0711_),
    .B(_0714_));
 sg13g2_nand2_1 _1602_ (.Y(_0717_),
    .A(_0697_),
    .B(_0716_));
 sg13g2_xor2_1 _1603_ (.B(_0716_),
    .A(_0697_),
    .X(_0718_));
 sg13g2_xnor2_1 _1604_ (.Y(uo_out[1]),
    .A(_0696_),
    .B(_0718_));
 sg13g2_nor2_1 _1605_ (.A(_0606_),
    .B(_0712_),
    .Y(_0719_));
 sg13g2_nand2b_1 _1606_ (.Y(_0720_),
    .B(_0604_),
    .A_N(_0602_));
 sg13g2_xor2_1 _1607_ (.B(_0602_),
    .A(\chan[3].attenuation.control[0] ),
    .X(_0721_));
 sg13g2_a22oi_1 _1608_ (.Y(_0722_),
    .B1(_0721_),
    .B2(_0608_),
    .A2(_0720_),
    .A1(_0719_));
 sg13g2_a21o_1 _1609_ (.A2(_0708_),
    .A1(_0705_),
    .B1(_0704_),
    .X(_0723_));
 sg13g2_o21ai_1 _1610_ (.B1(_0650_),
    .Y(_0724_),
    .A1(_0554_),
    .A2(_0565_));
 sg13g2_o21ai_1 _1611_ (.B1(_0724_),
    .Y(_0725_),
    .A1(_0561_),
    .A2(_0568_));
 sg13g2_nor2_1 _1612_ (.A(_0534_),
    .B(_0699_),
    .Y(_0726_));
 sg13g2_nand2b_1 _1613_ (.Y(_0727_),
    .B(_0582_),
    .A_N(_0536_));
 sg13g2_xor2_1 _1614_ (.B(_0536_),
    .A(net223),
    .X(_0728_));
 sg13g2_a22oi_1 _1615_ (.Y(_0729_),
    .B1(_0728_),
    .B2(_0583_),
    .A2(_0727_),
    .A1(_0726_));
 sg13g2_nor2_1 _1616_ (.A(_0544_),
    .B(_0591_),
    .Y(_0730_));
 sg13g2_nor3_1 _1617_ (.A(_0547_),
    .B(_0589_),
    .C(_0643_),
    .Y(_0731_));
 sg13g2_nor2_2 _1618_ (.A(_0730_),
    .B(_0731_),
    .Y(_0732_));
 sg13g2_nor2_1 _1619_ (.A(_0729_),
    .B(_0732_),
    .Y(_0733_));
 sg13g2_xor2_1 _1620_ (.B(_0732_),
    .A(_0729_),
    .X(_0734_));
 sg13g2_xnor2_1 _1621_ (.Y(_0735_),
    .A(_0725_),
    .B(_0734_));
 sg13g2_nor2b_1 _1622_ (.A(_0735_),
    .B_N(_0723_),
    .Y(_0736_));
 sg13g2_xor2_1 _1623_ (.B(_0735_),
    .A(_0723_),
    .X(_0737_));
 sg13g2_nor2_1 _1624_ (.A(_0722_),
    .B(_0737_),
    .Y(_0738_));
 sg13g2_xor2_1 _1625_ (.B(_0737_),
    .A(_0722_),
    .X(_0739_));
 sg13g2_o21ai_1 _1626_ (.B1(_0739_),
    .Y(_0740_),
    .A1(_0710_),
    .A2(_0715_));
 sg13g2_or3_1 _1627_ (.A(_0710_),
    .B(_0715_),
    .C(_0739_),
    .X(_0741_));
 sg13g2_and2_1 _1628_ (.A(_0740_),
    .B(_0741_),
    .X(_0742_));
 sg13g2_and3_1 _1629_ (.X(_0743_),
    .A(_0679_),
    .B(_0695_),
    .C(_0718_));
 sg13g2_o21ai_1 _1630_ (.B1(_0694_),
    .Y(_0744_),
    .A1(_0697_),
    .A2(_0716_));
 sg13g2_nand2_1 _1631_ (.Y(_0745_),
    .A(_0717_),
    .B(_0744_));
 sg13g2_nor2_1 _1632_ (.A(_0743_),
    .B(_0745_),
    .Y(_0746_));
 sg13g2_o21ai_1 _1633_ (.B1(_0742_),
    .Y(_0747_),
    .A1(_0743_),
    .A2(_0745_));
 sg13g2_xnor2_1 _1634_ (.Y(uo_out[2]),
    .A(_0742_),
    .B(_0746_));
 sg13g2_a21oi_1 _1635_ (.A1(_0605_),
    .A2(_0662_),
    .Y(_0748_),
    .B1(_0607_));
 sg13g2_nor2_2 _1636_ (.A(_0719_),
    .B(_0748_),
    .Y(_0749_));
 sg13g2_a21oi_1 _1637_ (.A1(_0725_),
    .A2(_0734_),
    .Y(_0750_),
    .B1(_0733_));
 sg13g2_a21oi_1 _1638_ (.A1(\chan[2].attenuation.control[0] ),
    .A2(_0554_),
    .Y(_0751_),
    .B1(_0574_));
 sg13g2_nor2_1 _1639_ (.A(_0559_),
    .B(_0751_),
    .Y(_0752_));
 sg13g2_or2_2 _1640_ (.X(_0753_),
    .B(_0752_),
    .A(_0650_));
 sg13g2_inv_1 _1641_ (.Y(_0754_),
    .A(_0753_));
 sg13g2_o21ai_1 _1642_ (.B1(_0540_),
    .Y(_0755_),
    .A1(_0580_),
    .A2(_0581_));
 sg13g2_a21oi_2 _1643_ (.B1(_0726_),
    .Y(_0756_),
    .A2(_0755_),
    .A1(_0534_));
 sg13g2_a221oi_1 _1644_ (.B2(_0589_),
    .C1(_0548_),
    .B1(_0587_),
    .A1(\chan[1].attenuation.control[0] ),
    .Y(_0757_),
    .A2(_0542_));
 sg13g2_a21o_2 _1645_ (.A2(_0643_),
    .A1(\chan[1].attenuation.control[3] ),
    .B1(_0757_),
    .X(_0758_));
 sg13g2_nand2_1 _1646_ (.Y(_0759_),
    .A(_0756_),
    .B(_0758_));
 sg13g2_xnor2_1 _1647_ (.Y(_0760_),
    .A(_0756_),
    .B(_0758_));
 sg13g2_xor2_1 _1648_ (.B(_0760_),
    .A(_0753_),
    .X(_0761_));
 sg13g2_nor2b_1 _1649_ (.A(_0750_),
    .B_N(_0761_),
    .Y(_0762_));
 sg13g2_xnor2_1 _1650_ (.Y(_0763_),
    .A(_0750_),
    .B(_0761_));
 sg13g2_xor2_1 _1651_ (.B(_0763_),
    .A(_0749_),
    .X(_0764_));
 sg13g2_nor3_1 _1652_ (.A(_0736_),
    .B(_0738_),
    .C(_0764_),
    .Y(_0765_));
 sg13g2_o21ai_1 _1653_ (.B1(_0764_),
    .Y(_0766_),
    .A1(_0736_),
    .A2(_0738_));
 sg13g2_nand2b_1 _1654_ (.Y(_0767_),
    .B(_0766_),
    .A_N(_0765_));
 sg13g2_nand2_1 _1655_ (.Y(_0768_),
    .A(_0740_),
    .B(_0747_));
 sg13g2_xnor2_1 _1656_ (.Y(uo_out[3]),
    .A(_0767_),
    .B(_0768_));
 sg13g2_a21oi_1 _1657_ (.A1(_0749_),
    .A2(_0763_),
    .Y(_0769_),
    .B1(_0762_));
 sg13g2_and2_2 _1658_ (.A(_0601_),
    .B(_0608_),
    .X(_0770_));
 sg13g2_inv_1 _1659_ (.Y(_0771_),
    .A(_0770_));
 sg13g2_o21ai_1 _1660_ (.B1(_0759_),
    .Y(_0772_),
    .A1(_0753_),
    .A2(_0760_));
 sg13g2_nor2b_2 _1661_ (.A(_0573_),
    .B_N(_0575_),
    .Y(_0773_));
 sg13g2_nand2_2 _1662_ (.Y(_0774_),
    .A(_0578_),
    .B(_0583_));
 sg13g2_inv_1 _1663_ (.Y(_0775_),
    .A(_0774_));
 sg13g2_nand2b_2 _1664_ (.Y(_0776_),
    .B(_0587_),
    .A_N(_0591_));
 sg13g2_inv_1 _1665_ (.Y(_0777_),
    .A(_0776_));
 sg13g2_xor2_1 _1666_ (.B(_0776_),
    .A(_0774_),
    .X(_0778_));
 sg13g2_nand2_1 _1667_ (.Y(_0779_),
    .A(_0773_),
    .B(_0778_));
 sg13g2_xor2_1 _1668_ (.B(_0778_),
    .A(_0773_),
    .X(_0780_));
 sg13g2_nand2_1 _1669_ (.Y(_0781_),
    .A(_0772_),
    .B(_0780_));
 sg13g2_xnor2_1 _1670_ (.Y(_0782_),
    .A(_0772_),
    .B(_0780_));
 sg13g2_xnor2_1 _1671_ (.Y(_0783_),
    .A(_0771_),
    .B(_0782_));
 sg13g2_nor2_1 _1672_ (.A(_0769_),
    .B(_0783_),
    .Y(_0784_));
 sg13g2_nand2_1 _1673_ (.Y(_0785_),
    .A(_0769_),
    .B(_0783_));
 sg13g2_nand2b_1 _1674_ (.Y(_0786_),
    .B(_0785_),
    .A_N(_0784_));
 sg13g2_and2_1 _1675_ (.A(_0740_),
    .B(_0766_),
    .X(_0787_));
 sg13g2_a21oi_1 _1676_ (.A1(_0747_),
    .A2(_0787_),
    .Y(_0788_),
    .B1(_0765_));
 sg13g2_xnor2_1 _1677_ (.Y(uo_out[4]),
    .A(_0786_),
    .B(_0788_));
 sg13g2_a21oi_1 _1678_ (.A1(_0785_),
    .A2(_0788_),
    .Y(_0789_),
    .B1(_0784_));
 sg13g2_o21ai_1 _1679_ (.B1(_0781_),
    .Y(_0790_),
    .A1(_0771_),
    .A2(_0782_));
 sg13g2_nor2_2 _1680_ (.A(\chan[3].attenuation.control[2] ),
    .B(_0607_),
    .Y(_0791_));
 sg13g2_o21ai_1 _1681_ (.B1(_0779_),
    .Y(_0792_),
    .A1(_0774_),
    .A2(_0776_));
 sg13g2_nor2_2 _1682_ (.A(\chan[0].attenuation.control[2] ),
    .B(_0535_),
    .Y(_0793_));
 sg13g2_nor2_2 _1683_ (.A(\chan[1].attenuation.control[2] ),
    .B(_0548_),
    .Y(_0794_));
 sg13g2_xnor2_1 _1684_ (.Y(_0795_),
    .A(_0793_),
    .B(_0794_));
 sg13g2_nor3_1 _1685_ (.A(net222),
    .B(_0559_),
    .C(_0795_),
    .Y(_0796_));
 sg13g2_xor2_1 _1686_ (.B(_0795_),
    .A(_0653_),
    .X(_0797_));
 sg13g2_inv_1 _1687_ (.Y(_0798_),
    .A(_0797_));
 sg13g2_xnor2_1 _1688_ (.Y(_0799_),
    .A(_0792_),
    .B(_0798_));
 sg13g2_nor3_1 _1689_ (.A(\chan[3].attenuation.control[2] ),
    .B(_0607_),
    .C(_0799_),
    .Y(_0800_));
 sg13g2_xor2_1 _1690_ (.B(_0799_),
    .A(_0791_),
    .X(_0801_));
 sg13g2_nand2b_1 _1691_ (.Y(_0802_),
    .B(_0790_),
    .A_N(_0801_));
 sg13g2_xnor2_1 _1692_ (.Y(_0803_),
    .A(_0790_),
    .B(_0801_));
 sg13g2_inv_1 _1693_ (.Y(_0804_),
    .A(_0803_));
 sg13g2_xnor2_1 _1694_ (.Y(uo_out[5]),
    .A(_0789_),
    .B(_0803_));
 sg13g2_o21ai_1 _1695_ (.B1(_0802_),
    .Y(_0805_),
    .A1(_0789_),
    .A2(_0804_));
 sg13g2_a21oi_2 _1696_ (.B1(_0796_),
    .Y(_0806_),
    .A2(_0794_),
    .A1(_0793_));
 sg13g2_a21o_1 _1697_ (.A2(_0798_),
    .A1(_0792_),
    .B1(_0800_),
    .X(_0807_));
 sg13g2_nor2b_1 _1698_ (.A(_0806_),
    .B_N(_0807_),
    .Y(_0808_));
 sg13g2_xor2_1 _1699_ (.B(_0807_),
    .A(_0806_),
    .X(_0809_));
 sg13g2_nor2b_1 _1700_ (.A(_0809_),
    .B_N(_0805_),
    .Y(_0810_));
 sg13g2_xnor2_1 _1701_ (.Y(uo_out[6]),
    .A(_0805_),
    .B(_0809_));
 sg13g2_nor2_1 _1702_ (.A(_0808_),
    .B(_0810_),
    .Y(_0811_));
 sg13g2_inv_1 _1703_ (.Y(uo_out[7]),
    .A(_0811_));
 sg13g2_xor2_1 _1704_ (.B(_0671_),
    .A(_0670_),
    .X(_0812_));
 sg13g2_or2_1 _1705_ (.X(_0813_),
    .B(_0812_),
    .A(net415));
 sg13g2_nand2_1 _1706_ (.Y(_0814_),
    .A(net415),
    .B(_0812_));
 sg13g2_and3_1 _1707_ (.X(_0007_),
    .A(net233),
    .B(_0813_),
    .C(_0814_));
 sg13g2_xor2_1 _1708_ (.B(_0673_),
    .A(_0672_),
    .X(_0815_));
 sg13g2_nand2_1 _1709_ (.Y(_0816_),
    .A(net482),
    .B(_0815_));
 sg13g2_xnor2_1 _1710_ (.Y(_0817_),
    .A(\pwm.accumulator[1] ),
    .B(_0815_));
 sg13g2_o21ai_1 _1711_ (.B1(net245),
    .Y(_0818_),
    .A1(_0814_),
    .A2(_0817_));
 sg13g2_a21oi_1 _1712_ (.A1(_0814_),
    .A2(_0817_),
    .Y(_0008_),
    .B1(_0818_));
 sg13g2_o21ai_1 _1713_ (.B1(_0816_),
    .Y(_0819_),
    .A1(_0814_),
    .A2(_0817_));
 sg13g2_xor2_1 _1714_ (.B(_0675_),
    .A(_0674_),
    .X(_0820_));
 sg13g2_and2_1 _1715_ (.A(\pwm.accumulator[2] ),
    .B(_0820_),
    .X(_0821_));
 sg13g2_or2_1 _1716_ (.X(_0822_),
    .B(_0820_),
    .A(\pwm.accumulator[2] ));
 sg13g2_nor2b_1 _1717_ (.A(_0821_),
    .B_N(_0822_),
    .Y(_0823_));
 sg13g2_o21ai_1 _1718_ (.B1(net245),
    .Y(_0824_),
    .A1(_0819_),
    .A2(_0823_));
 sg13g2_a21oi_1 _1719_ (.A1(_0819_),
    .A2(_0823_),
    .Y(_0009_),
    .B1(_0824_));
 sg13g2_a21oi_1 _1720_ (.A1(_0819_),
    .A2(_0822_),
    .Y(_0825_),
    .B1(_0821_));
 sg13g2_xnor2_1 _1721_ (.Y(_0826_),
    .A(_0676_),
    .B(_0678_));
 sg13g2_nand2_1 _1722_ (.Y(_0827_),
    .A(net469),
    .B(_0826_));
 sg13g2_xnor2_1 _1723_ (.Y(_0828_),
    .A(net469),
    .B(_0826_));
 sg13g2_o21ai_1 _1724_ (.B1(net245),
    .Y(_0829_),
    .A1(_0825_),
    .A2(_0828_));
 sg13g2_a21oi_1 _1725_ (.A1(_0825_),
    .A2(_0828_),
    .Y(_0010_),
    .B1(_0829_));
 sg13g2_and2_1 _1726_ (.A(\pwm.accumulator[4] ),
    .B(uo_out[0]),
    .X(_0830_));
 sg13g2_xor2_1 _1727_ (.B(uo_out[0]),
    .A(net503),
    .X(_0831_));
 sg13g2_o21ai_1 _1728_ (.B1(_0827_),
    .Y(_0832_),
    .A1(_0825_),
    .A2(_0828_));
 sg13g2_nor2_1 _1729_ (.A(_0831_),
    .B(_0832_),
    .Y(_0833_));
 sg13g2_a21oi_1 _1730_ (.A1(_0831_),
    .A2(_0832_),
    .Y(_0834_),
    .B1(net228));
 sg13g2_nor2b_1 _1731_ (.A(_0833_),
    .B_N(_0834_),
    .Y(_0011_));
 sg13g2_nand2_1 _1732_ (.Y(_0835_),
    .A(net511),
    .B(uo_out[1]));
 sg13g2_xnor2_1 _1733_ (.Y(_0836_),
    .A(net465),
    .B(uo_out[1]));
 sg13g2_a21oi_2 _1734_ (.B1(_0830_),
    .Y(_0837_),
    .A2(_0832_),
    .A1(_0831_));
 sg13g2_o21ai_1 _1735_ (.B1(net244),
    .Y(_0838_),
    .A1(_0836_),
    .A2(_0837_));
 sg13g2_a21oi_1 _1736_ (.A1(_0836_),
    .A2(_0837_),
    .Y(_0012_),
    .B1(_0838_));
 sg13g2_o21ai_1 _1737_ (.B1(_0835_),
    .Y(_0839_),
    .A1(_0836_),
    .A2(_0837_));
 sg13g2_and2_1 _1738_ (.A(\pwm.accumulator[6] ),
    .B(uo_out[2]),
    .X(_0840_));
 sg13g2_xor2_1 _1739_ (.B(uo_out[2]),
    .A(\pwm.accumulator[6] ),
    .X(_0841_));
 sg13g2_or2_1 _1740_ (.X(_0842_),
    .B(_0841_),
    .A(_0839_));
 sg13g2_nand2_1 _1741_ (.Y(_0843_),
    .A(_0839_),
    .B(_0841_));
 sg13g2_and3_1 _1742_ (.X(_0013_),
    .A(net244),
    .B(_0842_),
    .C(_0843_));
 sg13g2_nor2_1 _1743_ (.A(net458),
    .B(uo_out[3]),
    .Y(_0844_));
 sg13g2_xor2_1 _1744_ (.B(uo_out[3]),
    .A(net458),
    .X(_0845_));
 sg13g2_nand2b_1 _1745_ (.Y(_0846_),
    .B(_0843_),
    .A_N(_0840_));
 sg13g2_o21ai_1 _1746_ (.B1(net244),
    .Y(_0847_),
    .A1(_0845_),
    .A2(_0846_));
 sg13g2_a21oi_1 _1747_ (.A1(_0845_),
    .A2(_0846_),
    .Y(_0014_),
    .B1(_0847_));
 sg13g2_and2_1 _1748_ (.A(\pwm.accumulator[8] ),
    .B(uo_out[4]),
    .X(_0848_));
 sg13g2_xnor2_1 _1749_ (.Y(_0849_),
    .A(net499),
    .B(uo_out[4]));
 sg13g2_a221oi_1 _1750_ (.B2(_0841_),
    .C1(_0840_),
    .B1(_0839_),
    .A1(\pwm.accumulator[7] ),
    .Y(_0850_),
    .A2(uo_out[3]));
 sg13g2_o21ai_1 _1751_ (.B1(_0849_),
    .Y(_0851_),
    .A1(_0844_),
    .A2(_0850_));
 sg13g2_or3_1 _1752_ (.A(_0844_),
    .B(_0849_),
    .C(_0850_),
    .X(_0852_));
 sg13g2_and3_1 _1753_ (.X(_0015_),
    .A(net236),
    .B(_0851_),
    .C(_0852_));
 sg13g2_nor2_1 _1754_ (.A(net452),
    .B(uo_out[5]),
    .Y(_0853_));
 sg13g2_xnor2_1 _1755_ (.Y(_0854_),
    .A(net452),
    .B(uo_out[5]));
 sg13g2_nor2b_1 _1756_ (.A(_0848_),
    .B_N(_0852_),
    .Y(_0855_));
 sg13g2_o21ai_1 _1757_ (.B1(net236),
    .Y(_0856_),
    .A1(_0854_),
    .A2(_0855_));
 sg13g2_a21oi_1 _1758_ (.A1(_0854_),
    .A2(_0855_),
    .Y(_0016_),
    .B1(_0856_));
 sg13g2_nand2_1 _1759_ (.Y(_0857_),
    .A(net467),
    .B(uo_out[6]));
 sg13g2_xnor2_1 _1760_ (.Y(_0858_),
    .A(net467),
    .B(uo_out[6]));
 sg13g2_a21oi_1 _1761_ (.A1(\pwm.accumulator[9] ),
    .A2(uo_out[5]),
    .Y(_0859_),
    .B1(_0848_));
 sg13g2_a21o_1 _1762_ (.A2(_0859_),
    .A1(_0852_),
    .B1(_0853_),
    .X(_0860_));
 sg13g2_o21ai_1 _1763_ (.B1(net236),
    .Y(_0861_),
    .A1(_0858_),
    .A2(_0860_));
 sg13g2_a21oi_1 _1764_ (.A1(_0858_),
    .A2(_0860_),
    .Y(_0017_),
    .B1(_0861_));
 sg13g2_nand2_1 _1765_ (.Y(_0862_),
    .A(net347),
    .B(uo_out[7]));
 sg13g2_xnor2_1 _1766_ (.Y(_0863_),
    .A(net347),
    .B(_0811_));
 sg13g2_o21ai_1 _1767_ (.B1(_0857_),
    .Y(_0864_),
    .A1(_0858_),
    .A2(_0860_));
 sg13g2_nand2_1 _1768_ (.Y(_0865_),
    .A(_0863_),
    .B(_0864_));
 sg13g2_o21ai_1 _1769_ (.B1(net236),
    .Y(_0866_),
    .A1(_0863_),
    .A2(_0864_));
 sg13g2_nor2b_1 _1770_ (.A(_0866_),
    .B_N(_0865_),
    .Y(_0018_));
 sg13g2_a21oi_1 _1771_ (.A1(_0862_),
    .A2(_0865_),
    .Y(_0019_),
    .B1(net224));
 sg13g2_nor2b_2 _1772_ (.A(net9),
    .B_N(net8),
    .Y(_0867_));
 sg13g2_o21ai_1 _1773_ (.B1(net243),
    .Y(_0868_),
    .A1(net427),
    .A2(_0867_));
 sg13g2_a21oi_1 _1774_ (.A1(_0501_),
    .A2(_0867_),
    .Y(_0020_),
    .B1(_0868_));
 sg13g2_o21ai_1 _1775_ (.B1(net237),
    .Y(_0869_),
    .A1(net429),
    .A2(_0867_));
 sg13g2_a21oi_1 _1776_ (.A1(_0499_),
    .A2(_0867_),
    .Y(_0021_),
    .B1(_0869_));
 sg13g2_nor2_1 _1777_ (.A(net361),
    .B(_0867_),
    .Y(_0870_));
 sg13g2_nor2b_2 _1778_ (.A(net7),
    .B_N(_0867_),
    .Y(_0871_));
 sg13g2_nor3_1 _1779_ (.A(net227),
    .B(_0870_),
    .C(_0871_),
    .Y(_0022_));
 sg13g2_and2_1 _1780_ (.A(net244),
    .B(net257),
    .X(_0023_));
 sg13g2_o21ai_1 _1781_ (.B1(net244),
    .Y(_0872_),
    .A1(net350),
    .A2(\clk_counter[0] ));
 sg13g2_a21oi_1 _1782_ (.A1(net350),
    .A2(\clk_counter[0] ),
    .Y(_0024_),
    .B1(_0872_));
 sg13g2_a21oi_1 _1783_ (.A1(\clk_counter[1] ),
    .A2(\clk_counter[0] ),
    .Y(_0873_),
    .B1(net287));
 sg13g2_nand3_1 _1784_ (.B(\clk_counter[0] ),
    .C(net287),
    .A(net350),
    .Y(_0874_));
 sg13g2_nand2_1 _1785_ (.Y(_0875_),
    .A(net244),
    .B(_0874_));
 sg13g2_nor2_1 _1786_ (.A(net288),
    .B(_0875_),
    .Y(_0025_));
 sg13g2_and2_1 _1787_ (.A(_0524_),
    .B(_0874_),
    .X(_0876_));
 sg13g2_nor2_1 _1788_ (.A(_0524_),
    .B(_0874_),
    .Y(_0877_));
 sg13g2_nor3_1 _1789_ (.A(net228),
    .B(net444),
    .C(_0877_),
    .Y(_0026_));
 sg13g2_and2_1 _1790_ (.A(net405),
    .B(_0877_),
    .X(_0878_));
 sg13g2_o21ai_1 _1791_ (.B1(net245),
    .Y(_0879_),
    .A1(net405),
    .A2(_0877_));
 sg13g2_nor2_1 _1792_ (.A(_0878_),
    .B(net406),
    .Y(_0027_));
 sg13g2_or2_1 _1793_ (.X(_0880_),
    .B(_0878_),
    .A(net455));
 sg13g2_nand2_1 _1794_ (.Y(_0881_),
    .A(net455),
    .B(_0878_));
 sg13g2_and3_1 _1795_ (.X(_0028_),
    .A(net244),
    .B(_0880_),
    .C(_0881_));
 sg13g2_o21ai_1 _1796_ (.B1(net245),
    .Y(_0882_),
    .A1(_0526_),
    .A2(_0881_));
 sg13g2_a21oi_1 _1797_ (.A1(_0526_),
    .A2(_0881_),
    .Y(_0029_),
    .B1(_0882_));
 sg13g2_nor2b_1 _1798_ (.A(\latch_control_reg[1] ),
    .B_N(\latch_control_reg[0] ),
    .Y(_0883_));
 sg13g2_nor3_2 _1799_ (.A(\latch_control_reg[2] ),
    .B(net8),
    .C(net9),
    .Y(_0884_));
 sg13g2_nor2_1 _1800_ (.A(net6),
    .B(_0501_),
    .Y(_0885_));
 sg13g2_a22oi_1 _1801_ (.Y(_0886_),
    .B1(_0885_),
    .B2(_0871_),
    .A2(_0884_),
    .A1(_0883_));
 sg13g2_a21oi_1 _1802_ (.A1(net419),
    .A2(_0886_),
    .Y(_0887_),
    .B1(net226));
 sg13g2_o21ai_1 _1803_ (.B1(_0887_),
    .Y(_0030_),
    .A1(_0484_),
    .A2(_0886_));
 sg13g2_a21oi_1 _1804_ (.A1(net479),
    .A2(_0886_),
    .Y(_0888_),
    .B1(net226));
 sg13g2_o21ai_1 _1805_ (.B1(_0888_),
    .Y(_0031_),
    .A1(_0483_),
    .A2(_0886_));
 sg13g2_a21oi_1 _1806_ (.A1(net480),
    .A2(_0886_),
    .Y(_0889_),
    .B1(net226));
 sg13g2_o21ai_1 _1807_ (.B1(_0889_),
    .Y(_0032_),
    .A1(_0481_),
    .A2(_0886_));
 sg13g2_a21oi_1 _1808_ (.A1(net439),
    .A2(_0886_),
    .Y(_0890_),
    .B1(net226));
 sg13g2_o21ai_1 _1809_ (.B1(_0890_),
    .Y(_0033_),
    .A1(_0479_),
    .A2(_0886_));
 sg13g2_nor2_1 _1810_ (.A(_0499_),
    .B(_0501_),
    .Y(_0891_));
 sg13g2_and2_1 _1811_ (.A(\latch_control_reg[1] ),
    .B(\latch_control_reg[0] ),
    .X(_0892_));
 sg13g2_a22oi_1 _1812_ (.Y(_0893_),
    .B1(_0892_),
    .B2(_0884_),
    .A2(_0891_),
    .A1(_0871_));
 sg13g2_a21oi_1 _1813_ (.A1(net460),
    .A2(_0893_),
    .Y(_0894_),
    .B1(net225));
 sg13g2_o21ai_1 _1814_ (.B1(_0894_),
    .Y(_0034_),
    .A1(_0484_),
    .A2(_0893_));
 sg13g2_a21oi_1 _1815_ (.A1(net430),
    .A2(_0893_),
    .Y(_0895_),
    .B1(net225));
 sg13g2_o21ai_1 _1816_ (.B1(_0895_),
    .Y(_0035_),
    .A1(_0483_),
    .A2(_0893_));
 sg13g2_a21oi_1 _1817_ (.A1(net474),
    .A2(_0893_),
    .Y(_0896_),
    .B1(net225));
 sg13g2_o21ai_1 _1818_ (.B1(_0896_),
    .Y(_0036_),
    .A1(_0481_),
    .A2(_0893_));
 sg13g2_a21oi_1 _1819_ (.A1(net481),
    .A2(_0893_),
    .Y(_0897_),
    .B1(net225));
 sg13g2_o21ai_1 _1820_ (.B1(_0897_),
    .Y(_0037_),
    .A1(_0479_),
    .A2(_0893_));
 sg13g2_nor3_2 _1821_ (.A(net8),
    .B(net9),
    .C(_0003_),
    .Y(_0898_));
 sg13g2_and2_2 _1822_ (.A(net7),
    .B(_0867_),
    .X(_0899_));
 sg13g2_a22oi_1 _1823_ (.Y(_0900_),
    .B1(_0899_),
    .B2(_0885_),
    .A2(_0898_),
    .A1(_0883_));
 sg13g2_a21oi_1 _1824_ (.A1(net492),
    .A2(_0900_),
    .Y(_0901_),
    .B1(net229));
 sg13g2_o21ai_1 _1825_ (.B1(_0901_),
    .Y(_0038_),
    .A1(_0484_),
    .A2(_0900_));
 sg13g2_a21oi_1 _1826_ (.A1(net471),
    .A2(_0900_),
    .Y(_0902_),
    .B1(net225));
 sg13g2_o21ai_1 _1827_ (.B1(_0902_),
    .Y(_0039_),
    .A1(_0483_),
    .A2(_0900_));
 sg13g2_a21oi_1 _1828_ (.A1(net428),
    .A2(_0900_),
    .Y(_0903_),
    .B1(net228));
 sg13g2_o21ai_1 _1829_ (.B1(_0903_),
    .Y(_0040_),
    .A1(_0481_),
    .A2(_0900_));
 sg13g2_a21oi_1 _1830_ (.A1(net454),
    .A2(_0900_),
    .Y(_0904_),
    .B1(net227));
 sg13g2_o21ai_1 _1831_ (.B1(_0904_),
    .Y(_0041_),
    .A1(_0479_),
    .A2(_0900_));
 sg13g2_a22oi_1 _1832_ (.Y(_0905_),
    .B1(_0899_),
    .B2(_0891_),
    .A2(_0898_),
    .A1(_0892_));
 sg13g2_a21oi_1 _1833_ (.A1(net472),
    .A2(_0905_),
    .Y(_0906_),
    .B1(net229));
 sg13g2_o21ai_1 _1834_ (.B1(_0906_),
    .Y(_0042_),
    .A1(_0484_),
    .A2(_0905_));
 sg13g2_a21oi_1 _1835_ (.A1(net449),
    .A2(_0905_),
    .Y(_0907_),
    .B1(net228));
 sg13g2_o21ai_1 _1836_ (.B1(_0907_),
    .Y(_0043_),
    .A1(_0483_),
    .A2(_0905_));
 sg13g2_a21oi_1 _1837_ (.A1(net473),
    .A2(_0905_),
    .Y(_0908_),
    .B1(net228));
 sg13g2_o21ai_1 _1838_ (.B1(_0908_),
    .Y(_0044_),
    .A1(_0481_),
    .A2(_0905_));
 sg13g2_a21oi_1 _1839_ (.A1(net438),
    .A2(_0905_),
    .Y(_0909_),
    .B1(net228));
 sg13g2_o21ai_1 _1840_ (.B1(_0909_),
    .Y(_0045_),
    .A1(_0479_),
    .A2(_0905_));
 sg13g2_nor2_1 _1841_ (.A(\latch_control_reg[1] ),
    .B(\latch_control_reg[0] ),
    .Y(_0910_));
 sg13g2_nand2_1 _1842_ (.Y(_0911_),
    .A(_0884_),
    .B(_0910_));
 sg13g2_o21ai_1 _1843_ (.B1(net246),
    .Y(_0912_),
    .A1(net1),
    .A2(net212));
 sg13g2_a21oi_1 _1844_ (.A1(_0517_),
    .A2(net213),
    .Y(_0046_),
    .B1(_0912_));
 sg13g2_o21ai_1 _1845_ (.B1(net246),
    .Y(_0913_),
    .A1(net2),
    .A2(net212));
 sg13g2_a21oi_1 _1846_ (.A1(_0516_),
    .A2(net213),
    .Y(_0047_),
    .B1(_0913_));
 sg13g2_o21ai_1 _1847_ (.B1(net246),
    .Y(_0914_),
    .A1(net3),
    .A2(net212));
 sg13g2_a21oi_1 _1848_ (.A1(_0515_),
    .A2(net213),
    .Y(_0048_),
    .B1(_0914_));
 sg13g2_o21ai_1 _1849_ (.B1(net246),
    .Y(_0915_),
    .A1(net4),
    .A2(net212));
 sg13g2_a21oi_1 _1850_ (.A1(_0514_),
    .A2(net213),
    .Y(_0049_),
    .B1(_0915_));
 sg13g2_o21ai_1 _1851_ (.B1(net247),
    .Y(_0916_),
    .A1(net5),
    .A2(net212));
 sg13g2_a21oi_1 _1852_ (.A1(_0513_),
    .A2(net212),
    .Y(_0050_),
    .B1(_0916_));
 sg13g2_o21ai_1 _1853_ (.B1(net247),
    .Y(_0917_),
    .A1(net6),
    .A2(net212));
 sg13g2_a21oi_1 _1854_ (.A1(_0512_),
    .A2(net212),
    .Y(_0051_),
    .B1(_0917_));
 sg13g2_nand3b_1 _1855_ (.B(_0884_),
    .C(net508),
    .Y(_0918_),
    .A_N(\latch_control_reg[0] ));
 sg13g2_o21ai_1 _1856_ (.B1(net238),
    .Y(_0919_),
    .A1(net1),
    .A2(net211));
 sg13g2_a21oi_1 _1857_ (.A1(_0511_),
    .A2(net211),
    .Y(_0052_),
    .B1(_0919_));
 sg13g2_o21ai_1 _1858_ (.B1(net239),
    .Y(_0920_),
    .A1(net2),
    .A2(net211));
 sg13g2_a21oi_1 _1859_ (.A1(_0510_),
    .A2(net211),
    .Y(_0053_),
    .B1(_0920_));
 sg13g2_o21ai_1 _1860_ (.B1(net241),
    .Y(_0921_),
    .A1(net3),
    .A2(net210));
 sg13g2_a21oi_1 _1861_ (.A1(_0509_),
    .A2(net210),
    .Y(_0054_),
    .B1(_0921_));
 sg13g2_o21ai_1 _1862_ (.B1(net241),
    .Y(_0922_),
    .A1(net4),
    .A2(net210));
 sg13g2_a21oi_1 _1863_ (.A1(_0508_),
    .A2(net210),
    .Y(_0055_),
    .B1(_0922_));
 sg13g2_o21ai_1 _1864_ (.B1(net240),
    .Y(_0923_),
    .A1(net5),
    .A2(net210));
 sg13g2_a21oi_1 _1865_ (.A1(_0507_),
    .A2(net210),
    .Y(_0056_),
    .B1(_0923_));
 sg13g2_o21ai_1 _1866_ (.B1(net240),
    .Y(_0924_),
    .A1(net6),
    .A2(net210));
 sg13g2_a21oi_1 _1867_ (.A1(_0506_),
    .A2(net210),
    .Y(_0057_),
    .B1(_0924_));
 sg13g2_nand2_1 _1868_ (.Y(_0925_),
    .A(_0898_),
    .B(_0910_));
 sg13g2_o21ai_1 _1869_ (.B1(net249),
    .Y(_0926_),
    .A1(net1),
    .A2(net209));
 sg13g2_a21oi_1 _1870_ (.A1(_0505_),
    .A2(net209),
    .Y(_0058_),
    .B1(_0926_));
 sg13g2_o21ai_1 _1871_ (.B1(net248),
    .Y(_0927_),
    .A1(net2),
    .A2(net209));
 sg13g2_a21oi_1 _1872_ (.A1(_0504_),
    .A2(net209),
    .Y(_0059_),
    .B1(_0927_));
 sg13g2_o21ai_1 _1873_ (.B1(net250),
    .Y(_0928_),
    .A1(net3),
    .A2(net208));
 sg13g2_a21oi_1 _1874_ (.A1(_0503_),
    .A2(net208),
    .Y(_0060_),
    .B1(_0928_));
 sg13g2_o21ai_1 _1875_ (.B1(net249),
    .Y(_0929_),
    .A1(net4),
    .A2(net208));
 sg13g2_a21oi_1 _1876_ (.A1(_0502_),
    .A2(net208),
    .Y(_0061_),
    .B1(_0929_));
 sg13g2_o21ai_1 _1877_ (.B1(net249),
    .Y(_0930_),
    .A1(net5),
    .A2(net208));
 sg13g2_a21oi_1 _1878_ (.A1(_0500_),
    .A2(net208),
    .Y(_0062_),
    .B1(_0930_));
 sg13g2_o21ai_1 _1879_ (.B1(net249),
    .Y(_0931_),
    .A1(net6),
    .A2(net208));
 sg13g2_a21oi_1 _1880_ (.A1(_0498_),
    .A2(net208),
    .Y(_0063_),
    .B1(_0931_));
 sg13g2_nor2_1 _1881_ (.A(_0499_),
    .B(net5),
    .Y(_0932_));
 sg13g2_nand2_2 _1882_ (.Y(_0933_),
    .A(_0899_),
    .B(_0932_));
 sg13g2_o21ai_1 _1883_ (.B1(net237),
    .Y(_0934_),
    .A1(net1),
    .A2(_0933_));
 sg13g2_a21oi_1 _1884_ (.A1(_0497_),
    .A2(_0933_),
    .Y(_0064_),
    .B1(_0934_));
 sg13g2_o21ai_1 _1885_ (.B1(net243),
    .Y(_0935_),
    .A1(net2),
    .A2(_0933_));
 sg13g2_a21oi_1 _1886_ (.A1(_0496_),
    .A2(_0933_),
    .Y(_0065_),
    .B1(_0935_));
 sg13g2_a21oi_1 _1887_ (.A1(net376),
    .A2(_0933_),
    .Y(_0936_),
    .B1(net225));
 sg13g2_o21ai_1 _1888_ (.B1(_0936_),
    .Y(_0066_),
    .A1(_0481_),
    .A2(_0933_));
 sg13g2_mux4_1 _1889_ (.S0(_0497_),
    .A0(net500),
    .A1(_0528_),
    .A2(net219),
    .A3(\noise[0].gen.counter[6] ),
    .S1(net310),
    .X(_0937_));
 sg13g2_and2_1 _1890_ (.A(net237),
    .B(_0937_),
    .X(_0067_));
 sg13g2_nor3_1 _1891_ (.A(\tone[0].gen.counter[3] ),
    .B(\tone[0].gen.counter[2] ),
    .C(\tone[0].gen.counter[1] ),
    .Y(_0938_));
 sg13g2_nor4_1 _1892_ (.A(\tone[0].gen.counter[9] ),
    .B(\tone[0].gen.counter[8] ),
    .C(\tone[0].gen.counter[7] ),
    .D(\tone[0].gen.counter[4] ),
    .Y(_0939_));
 sg13g2_nand3_1 _1893_ (.B(_0938_),
    .C(_0939_),
    .A(_0494_),
    .Y(_0940_));
 sg13g2_nor3_1 _1894_ (.A(\tone[0].gen.counter[6] ),
    .B(\tone[0].gen.counter[5] ),
    .C(_0940_),
    .Y(_0941_));
 sg13g2_nor4_1 _1895_ (.A(\clk_counter[1] ),
    .B(\clk_counter[0] ),
    .C(\clk_counter[3] ),
    .D(\clk_counter[2] ),
    .Y(_0942_));
 sg13g2_a21oi_1 _1896_ (.A1(_0525_),
    .A2(net10),
    .Y(_0943_),
    .B1(_0942_));
 sg13g2_nor3_1 _1897_ (.A(\clk_counter[5] ),
    .B(\clk_counter[4] ),
    .C(\clk_counter[6] ),
    .Y(_0944_));
 sg13g2_or3_1 _1898_ (.A(_0525_),
    .B(net10),
    .C(_0944_),
    .X(_0945_));
 sg13g2_nor2b_1 _1899_ (.A(_0943_),
    .B_N(_0945_),
    .Y(_0946_));
 sg13g2_nand2b_1 _1900_ (.Y(_0947_),
    .B(_0945_),
    .A_N(_0943_));
 sg13g2_and2_1 _1901_ (.A(net207),
    .B(net202),
    .X(_0948_));
 sg13g2_o21ai_1 _1902_ (.B1(net233),
    .Y(_0949_),
    .A1(\chan[0].attenuation.in ),
    .A2(_0948_));
 sg13g2_a21oi_1 _1903_ (.A1(_0495_),
    .A2(_0948_),
    .Y(_0068_),
    .B1(_0949_));
 sg13g2_a21oi_1 _1904_ (.A1(net343),
    .A2(net207),
    .Y(_0950_),
    .B1(net306));
 sg13g2_o21ai_1 _1905_ (.B1(net240),
    .Y(_0951_),
    .A1(net197),
    .A2(_0950_));
 sg13g2_a21oi_1 _1906_ (.A1(_0494_),
    .A2(net197),
    .Y(_0069_),
    .B1(_0951_));
 sg13g2_a21oi_1 _1907_ (.A1(net375),
    .A2(net207),
    .Y(_0952_),
    .B1(net399));
 sg13g2_nand2_1 _1908_ (.Y(_0953_),
    .A(_0950_),
    .B(_0952_));
 sg13g2_o21ai_1 _1909_ (.B1(net202),
    .Y(_0954_),
    .A1(_0950_),
    .A2(_0952_));
 sg13g2_inv_1 _1910_ (.Y(_0955_),
    .A(_0954_));
 sg13g2_o21ai_1 _1911_ (.B1(net241),
    .Y(_0956_),
    .A1(net399),
    .A2(net202));
 sg13g2_a21oi_1 _1912_ (.A1(_0953_),
    .A2(_0955_),
    .Y(_0070_),
    .B1(_0956_));
 sg13g2_a21o_1 _1913_ (.A2(net207),
    .A1(net363),
    .B1(net381),
    .X(_0957_));
 sg13g2_nand2_1 _1914_ (.Y(_0958_),
    .A(_0953_),
    .B(_0957_));
 sg13g2_nor2_1 _1915_ (.A(_0953_),
    .B(_0957_),
    .Y(_0959_));
 sg13g2_nor2_1 _1916_ (.A(net197),
    .B(_0959_),
    .Y(_0960_));
 sg13g2_o21ai_1 _1917_ (.B1(net241),
    .Y(_0961_),
    .A1(net381),
    .A2(net202));
 sg13g2_a21oi_1 _1918_ (.A1(_0958_),
    .A2(_0960_),
    .Y(_0071_),
    .B1(_0961_));
 sg13g2_a21oi_1 _1919_ (.A1(net372),
    .A2(net207),
    .Y(_0962_),
    .B1(net414));
 sg13g2_and2_1 _1920_ (.A(_0959_),
    .B(_0962_),
    .X(_0963_));
 sg13g2_o21ai_1 _1921_ (.B1(net202),
    .Y(_0964_),
    .A1(_0959_),
    .A2(_0962_));
 sg13g2_nor2_1 _1922_ (.A(_0963_),
    .B(_0964_),
    .Y(_0965_));
 sg13g2_o21ai_1 _1923_ (.B1(net240),
    .Y(_0966_),
    .A1(net414),
    .A2(net206));
 sg13g2_nor2_1 _1924_ (.A(_0965_),
    .B(_0966_),
    .Y(_0072_));
 sg13g2_a21oi_1 _1925_ (.A1(net283),
    .A2(_0941_),
    .Y(_0967_),
    .B1(net392));
 sg13g2_and2_1 _1926_ (.A(_0963_),
    .B(_0967_),
    .X(_0968_));
 sg13g2_o21ai_1 _1927_ (.B1(net202),
    .Y(_0969_),
    .A1(_0963_),
    .A2(_0967_));
 sg13g2_nor2_1 _1928_ (.A(_0968_),
    .B(_0969_),
    .Y(_0970_));
 sg13g2_o21ai_1 _1929_ (.B1(net241),
    .Y(_0971_),
    .A1(net392),
    .A2(net202));
 sg13g2_nor2_1 _1930_ (.A(_0970_),
    .B(_0971_),
    .Y(_0073_));
 sg13g2_a21oi_1 _1931_ (.A1(net272),
    .A2(_0941_),
    .Y(_0972_),
    .B1(net402));
 sg13g2_nand2_1 _1932_ (.Y(_0973_),
    .A(_0968_),
    .B(_0972_));
 sg13g2_o21ai_1 _1933_ (.B1(net205),
    .Y(_0974_),
    .A1(_0968_),
    .A2(_0972_));
 sg13g2_inv_1 _1934_ (.Y(_0975_),
    .A(_0974_));
 sg13g2_o21ai_1 _1935_ (.B1(net241),
    .Y(_0976_),
    .A1(net402),
    .A2(net205));
 sg13g2_a21oi_1 _1936_ (.A1(_0973_),
    .A2(_0975_),
    .Y(_0074_),
    .B1(_0976_));
 sg13g2_a21o_1 _1937_ (.A2(net207),
    .A1(net286),
    .B1(net394),
    .X(_0977_));
 sg13g2_nand2_1 _1938_ (.Y(_0978_),
    .A(_0973_),
    .B(_0977_));
 sg13g2_nor2_1 _1939_ (.A(_0973_),
    .B(_0977_),
    .Y(_0979_));
 sg13g2_nor2_1 _1940_ (.A(net198),
    .B(_0979_),
    .Y(_0980_));
 sg13g2_o21ai_1 _1941_ (.B1(net246),
    .Y(_0981_),
    .A1(net394),
    .A2(net205));
 sg13g2_a21oi_1 _1942_ (.A1(_0978_),
    .A2(_0980_),
    .Y(_0075_),
    .B1(_0981_));
 sg13g2_a21oi_1 _1943_ (.A1(net277),
    .A2(net207),
    .Y(_0982_),
    .B1(net384));
 sg13g2_and2_1 _1944_ (.A(_0979_),
    .B(_0982_),
    .X(_0983_));
 sg13g2_o21ai_1 _1945_ (.B1(net205),
    .Y(_0984_),
    .A1(_0979_),
    .A2(_0982_));
 sg13g2_nor2_1 _1946_ (.A(_0983_),
    .B(_0984_),
    .Y(_0985_));
 sg13g2_o21ai_1 _1947_ (.B1(net246),
    .Y(_0986_),
    .A1(net384),
    .A2(net205));
 sg13g2_nor2_1 _1948_ (.A(_0985_),
    .B(_0986_),
    .Y(_0076_));
 sg13g2_a21oi_1 _1949_ (.A1(net266),
    .A2(net207),
    .Y(_0987_),
    .B1(net411));
 sg13g2_and2_1 _1950_ (.A(_0983_),
    .B(_0987_),
    .X(_0988_));
 sg13g2_o21ai_1 _1951_ (.B1(net205),
    .Y(_0989_),
    .A1(_0983_),
    .A2(_0987_));
 sg13g2_nor2_1 _1952_ (.A(_0988_),
    .B(_0989_),
    .Y(_0990_));
 sg13g2_o21ai_1 _1953_ (.B1(net246),
    .Y(_0991_),
    .A1(net411),
    .A2(net205));
 sg13g2_nor2_1 _1954_ (.A(_0990_),
    .B(_0991_),
    .Y(_0077_));
 sg13g2_nand2_1 _1955_ (.Y(_0992_),
    .A(net205),
    .B(_0988_));
 sg13g2_a21oi_1 _1956_ (.A1(net298),
    .A2(_0948_),
    .Y(_0993_),
    .B1(net386));
 sg13g2_o21ai_1 _1957_ (.B1(net240),
    .Y(_0994_),
    .A1(_0992_),
    .A2(_0993_));
 sg13g2_a21oi_1 _1958_ (.A1(_0992_),
    .A2(_0993_),
    .Y(_0078_),
    .B1(_0994_));
 sg13g2_nor3_1 _1959_ (.A(\tone[1].gen.counter[3] ),
    .B(\tone[1].gen.counter[2] ),
    .C(\tone[1].gen.counter[1] ),
    .Y(_0995_));
 sg13g2_nor4_1 _1960_ (.A(\tone[1].gen.counter[9] ),
    .B(\tone[1].gen.counter[8] ),
    .C(\tone[1].gen.counter[7] ),
    .D(\tone[1].gen.counter[4] ),
    .Y(_0996_));
 sg13g2_nand3_1 _1961_ (.B(_0995_),
    .C(_0996_),
    .A(_0492_),
    .Y(_0997_));
 sg13g2_nor3_1 _1962_ (.A(\tone[1].gen.counter[6] ),
    .B(\tone[1].gen.counter[5] ),
    .C(_0997_),
    .Y(_0998_));
 sg13g2_and2_1 _1963_ (.A(net201),
    .B(net196),
    .X(_0999_));
 sg13g2_o21ai_1 _1964_ (.B1(net233),
    .Y(_1000_),
    .A1(net220),
    .A2(_0999_));
 sg13g2_a21oi_1 _1965_ (.A1(_0493_),
    .A2(_0999_),
    .Y(_0079_),
    .B1(_1000_));
 sg13g2_a21oi_1 _1966_ (.A1(net344),
    .A2(net196),
    .Y(_1001_),
    .B1(net336));
 sg13g2_o21ai_1 _1967_ (.B1(net238),
    .Y(_1002_),
    .A1(net197),
    .A2(_1001_));
 sg13g2_a21oi_1 _1968_ (.A1(_0492_),
    .A2(net197),
    .Y(_0080_),
    .B1(_1002_));
 sg13g2_a21oi_1 _1969_ (.A1(net391),
    .A2(net196),
    .Y(_1003_),
    .B1(net413));
 sg13g2_nand2_1 _1970_ (.Y(_1004_),
    .A(_1001_),
    .B(_1003_));
 sg13g2_o21ai_1 _1971_ (.B1(net201),
    .Y(_1005_),
    .A1(_1001_),
    .A2(_1003_));
 sg13g2_inv_1 _1972_ (.Y(_1006_),
    .A(_1005_));
 sg13g2_o21ai_1 _1973_ (.B1(net238),
    .Y(_1007_),
    .A1(net413),
    .A2(net199));
 sg13g2_a21oi_1 _1974_ (.A1(_1004_),
    .A2(_1006_),
    .Y(_0081_),
    .B1(_1007_));
 sg13g2_a21o_1 _1975_ (.A2(net196),
    .A1(net383),
    .B1(net397),
    .X(_1008_));
 sg13g2_nand2_1 _1976_ (.Y(_1009_),
    .A(_1004_),
    .B(_1008_));
 sg13g2_nor2_1 _1977_ (.A(_1004_),
    .B(_1008_),
    .Y(_1010_));
 sg13g2_nor2_1 _1978_ (.A(net197),
    .B(_1010_),
    .Y(_1011_));
 sg13g2_o21ai_1 _1979_ (.B1(net238),
    .Y(_1012_),
    .A1(net397),
    .A2(net199));
 sg13g2_a21oi_1 _1980_ (.A1(_1009_),
    .A2(_1011_),
    .Y(_0082_),
    .B1(_1012_));
 sg13g2_a21oi_1 _1981_ (.A1(\control_tone_freq[1][3] ),
    .A2(net196),
    .Y(_1013_),
    .B1(net400));
 sg13g2_and2_1 _1982_ (.A(_1010_),
    .B(_1013_),
    .X(_1014_));
 sg13g2_o21ai_1 _1983_ (.B1(net199),
    .Y(_1015_),
    .A1(_1010_),
    .A2(_1013_));
 sg13g2_nor2_1 _1984_ (.A(_1014_),
    .B(_1015_),
    .Y(_1016_));
 sg13g2_o21ai_1 _1985_ (.B1(net238),
    .Y(_1017_),
    .A1(net400),
    .A2(net199));
 sg13g2_nor2_1 _1986_ (.A(_1016_),
    .B(_1017_),
    .Y(_0083_));
 sg13g2_a21oi_1 _1987_ (.A1(net279),
    .A2(_0998_),
    .Y(_1018_),
    .B1(net417));
 sg13g2_and2_1 _1988_ (.A(_1014_),
    .B(_1018_),
    .X(_1019_));
 sg13g2_o21ai_1 _1989_ (.B1(net200),
    .Y(_1020_),
    .A1(_1014_),
    .A2(_1018_));
 sg13g2_nor2_1 _1990_ (.A(_1019_),
    .B(_1020_),
    .Y(_1021_));
 sg13g2_o21ai_1 _1991_ (.B1(net239),
    .Y(_1022_),
    .A1(net417),
    .A2(net200));
 sg13g2_nor2_1 _1992_ (.A(_1021_),
    .B(_1022_),
    .Y(_0084_));
 sg13g2_a21oi_1 _1993_ (.A1(net281),
    .A2(_0998_),
    .Y(_0180_),
    .B1(net385));
 sg13g2_nand2_1 _1994_ (.Y(_0181_),
    .A(_1019_),
    .B(_0180_));
 sg13g2_o21ai_1 _1995_ (.B1(net200),
    .Y(_0182_),
    .A1(_1019_),
    .A2(_0180_));
 sg13g2_inv_1 _1996_ (.Y(_0183_),
    .A(_0182_));
 sg13g2_o21ai_1 _1997_ (.B1(net239),
    .Y(_0184_),
    .A1(net385),
    .A2(net200));
 sg13g2_a21oi_1 _1998_ (.A1(_0181_),
    .A2(_0183_),
    .Y(_0085_),
    .B1(_0184_));
 sg13g2_a21o_1 _1999_ (.A2(net196),
    .A1(net276),
    .B1(net388),
    .X(_0185_));
 sg13g2_nand2_1 _2000_ (.Y(_0186_),
    .A(_0181_),
    .B(_0185_));
 sg13g2_nor2_1 _2001_ (.A(_0181_),
    .B(_0185_),
    .Y(_0187_));
 sg13g2_nor2_1 _2002_ (.A(net197),
    .B(_0187_),
    .Y(_0188_));
 sg13g2_o21ai_1 _2003_ (.B1(net239),
    .Y(_0189_),
    .A1(net388),
    .A2(net201));
 sg13g2_a21oi_1 _2004_ (.A1(_0186_),
    .A2(_0188_),
    .Y(_0086_),
    .B1(_0189_));
 sg13g2_a21oi_1 _2005_ (.A1(net320),
    .A2(net196),
    .Y(_0190_),
    .B1(net418));
 sg13g2_and2_1 _2006_ (.A(_0187_),
    .B(_0190_),
    .X(_0191_));
 sg13g2_o21ai_1 _2007_ (.B1(net200),
    .Y(_0192_),
    .A1(_0187_),
    .A2(_0190_));
 sg13g2_nor2_1 _2008_ (.A(_0191_),
    .B(_0192_),
    .Y(_0193_));
 sg13g2_o21ai_1 _2009_ (.B1(net239),
    .Y(_0194_),
    .A1(net418),
    .A2(net201));
 sg13g2_nor2_1 _2010_ (.A(_0193_),
    .B(_0194_),
    .Y(_0087_));
 sg13g2_a21oi_1 _2011_ (.A1(net334),
    .A2(net196),
    .Y(_0195_),
    .B1(net408));
 sg13g2_and2_1 _2012_ (.A(_0191_),
    .B(_0195_),
    .X(_0196_));
 sg13g2_o21ai_1 _2013_ (.B1(net200),
    .Y(_0197_),
    .A1(_0191_),
    .A2(_0195_));
 sg13g2_nor2_1 _2014_ (.A(_0196_),
    .B(_0197_),
    .Y(_0198_));
 sg13g2_o21ai_1 _2015_ (.B1(net239),
    .Y(_0199_),
    .A1(net408),
    .A2(net200));
 sg13g2_nor2_1 _2016_ (.A(_0198_),
    .B(_0199_),
    .Y(_0088_));
 sg13g2_nand2_1 _2017_ (.Y(_0200_),
    .A(net200),
    .B(_0196_));
 sg13g2_a21oi_1 _2018_ (.A1(net294),
    .A2(_0999_),
    .Y(_0201_),
    .B1(net389));
 sg13g2_o21ai_1 _2019_ (.B1(net239),
    .Y(_0202_),
    .A1(_0200_),
    .A2(_0201_));
 sg13g2_a21oi_1 _2020_ (.A1(_0200_),
    .A2(_0201_),
    .Y(_0089_),
    .B1(_0202_));
 sg13g2_nor3_1 _2021_ (.A(\tone[2].gen.counter[3] ),
    .B(\tone[2].gen.counter[2] ),
    .C(\tone[2].gen.counter[1] ),
    .Y(_0203_));
 sg13g2_nor4_1 _2022_ (.A(\tone[2].gen.counter[9] ),
    .B(\tone[2].gen.counter[8] ),
    .C(\tone[2].gen.counter[7] ),
    .D(\tone[2].gen.counter[4] ),
    .Y(_0204_));
 sg13g2_nand3_1 _2023_ (.B(_0203_),
    .C(_0204_),
    .A(_0490_),
    .Y(_0205_));
 sg13g2_nor3_2 _2024_ (.A(\tone[2].gen.counter[6] ),
    .B(net509),
    .C(_0205_),
    .Y(_0206_));
 sg13g2_and2_1 _2025_ (.A(net206),
    .B(net195),
    .X(_0207_));
 sg13g2_o21ai_1 _2026_ (.B1(net247),
    .Y(_0208_),
    .A1(net219),
    .A2(_0207_));
 sg13g2_a21oi_1 _2027_ (.A1(_0491_),
    .A2(_0207_),
    .Y(_0090_),
    .B1(_0208_));
 sg13g2_a21oi_1 _2028_ (.A1(\control_tone_freq[2][0] ),
    .A2(net195),
    .Y(_0209_),
    .B1(net345));
 sg13g2_o21ai_1 _2029_ (.B1(net248),
    .Y(_0210_),
    .A1(net198),
    .A2(_0209_));
 sg13g2_a21oi_1 _2030_ (.A1(_0490_),
    .A2(net198),
    .Y(_0091_),
    .B1(_0210_));
 sg13g2_a21oi_1 _2031_ (.A1(net268),
    .A2(_0206_),
    .Y(_0211_),
    .B1(net377));
 sg13g2_nand2_1 _2032_ (.Y(_0212_),
    .A(_0209_),
    .B(_0211_));
 sg13g2_o21ai_1 _2033_ (.B1(net204),
    .Y(_0213_),
    .A1(_0209_),
    .A2(_0211_));
 sg13g2_inv_1 _2034_ (.Y(_0214_),
    .A(_0213_));
 sg13g2_o21ai_1 _2035_ (.B1(net248),
    .Y(_0215_),
    .A1(net377),
    .A2(net204));
 sg13g2_a21oi_1 _2036_ (.A1(_0212_),
    .A2(_0214_),
    .Y(_0092_),
    .B1(_0215_));
 sg13g2_a21o_1 _2037_ (.A2(net510),
    .A1(net271),
    .B1(net380),
    .X(_0216_));
 sg13g2_nand2_1 _2038_ (.Y(_0217_),
    .A(_0212_),
    .B(_0216_));
 sg13g2_nor2_1 _2039_ (.A(_0212_),
    .B(_0216_),
    .Y(_0218_));
 sg13g2_nor2_1 _2040_ (.A(net198),
    .B(_0218_),
    .Y(_0219_));
 sg13g2_o21ai_1 _2041_ (.B1(net248),
    .Y(_0220_),
    .A1(net380),
    .A2(net204));
 sg13g2_a21oi_1 _2042_ (.A1(_0217_),
    .A2(_0219_),
    .Y(_0093_),
    .B1(_0220_));
 sg13g2_a21oi_1 _2043_ (.A1(net297),
    .A2(net195),
    .Y(_0221_),
    .B1(net412));
 sg13g2_and2_1 _2044_ (.A(_0218_),
    .B(_0221_),
    .X(_0222_));
 sg13g2_o21ai_1 _2045_ (.B1(net204),
    .Y(_0223_),
    .A1(_0218_),
    .A2(_0221_));
 sg13g2_nor2_1 _2046_ (.A(_0222_),
    .B(_0223_),
    .Y(_0224_));
 sg13g2_o21ai_1 _2047_ (.B1(net248),
    .Y(_0225_),
    .A1(net412),
    .A2(net204));
 sg13g2_nor2_1 _2048_ (.A(_0224_),
    .B(_0225_),
    .Y(_0094_));
 sg13g2_a21oi_1 _2049_ (.A1(\control_tone_freq[2][4] ),
    .A2(net195),
    .Y(_0226_),
    .B1(net425));
 sg13g2_and2_1 _2050_ (.A(_0222_),
    .B(_0226_),
    .X(_0227_));
 sg13g2_o21ai_1 _2051_ (.B1(net203),
    .Y(_0228_),
    .A1(_0222_),
    .A2(_0226_));
 sg13g2_nor2_1 _2052_ (.A(_0227_),
    .B(_0228_),
    .Y(_0229_));
 sg13g2_o21ai_1 _2053_ (.B1(net248),
    .Y(_0230_),
    .A1(net425),
    .A2(net204));
 sg13g2_nor2_1 _2054_ (.A(_0229_),
    .B(_0230_),
    .Y(_0095_));
 sg13g2_a21oi_1 _2055_ (.A1(net290),
    .A2(net195),
    .Y(_0231_),
    .B1(net421));
 sg13g2_nand2_1 _2056_ (.Y(_0232_),
    .A(_0227_),
    .B(_0231_));
 sg13g2_o21ai_1 _2057_ (.B1(net203),
    .Y(_0233_),
    .A1(_0227_),
    .A2(_0231_));
 sg13g2_inv_1 _2058_ (.Y(_0234_),
    .A(_0233_));
 sg13g2_o21ai_1 _2059_ (.B1(net248),
    .Y(_0235_),
    .A1(net421),
    .A2(net203));
 sg13g2_a21oi_1 _2060_ (.A1(_0232_),
    .A2(_0234_),
    .Y(_0096_),
    .B1(_0235_));
 sg13g2_a21o_1 _2061_ (.A2(net195),
    .A1(net284),
    .B1(net420),
    .X(_0236_));
 sg13g2_nand2_1 _2062_ (.Y(_0237_),
    .A(_0232_),
    .B(_0236_));
 sg13g2_nor2_1 _2063_ (.A(_0232_),
    .B(_0236_),
    .Y(_0238_));
 sg13g2_nor2_1 _2064_ (.A(net197),
    .B(_0238_),
    .Y(_0239_));
 sg13g2_o21ai_1 _2065_ (.B1(net248),
    .Y(_0240_),
    .A1(net420),
    .A2(net203));
 sg13g2_a21oi_1 _2066_ (.A1(_0237_),
    .A2(_0239_),
    .Y(_0097_),
    .B1(_0240_));
 sg13g2_a21oi_1 _2067_ (.A1(net295),
    .A2(net195),
    .Y(_0241_),
    .B1(net407));
 sg13g2_and2_1 _2068_ (.A(_0238_),
    .B(_0241_),
    .X(_0242_));
 sg13g2_o21ai_1 _2069_ (.B1(net203),
    .Y(_0243_),
    .A1(_0238_),
    .A2(_0241_));
 sg13g2_nor2_1 _2070_ (.A(_0242_),
    .B(_0243_),
    .Y(_0244_));
 sg13g2_o21ai_1 _2071_ (.B1(net249),
    .Y(_0245_),
    .A1(net407),
    .A2(net203));
 sg13g2_nor2_1 _2072_ (.A(_0244_),
    .B(_0245_),
    .Y(_0098_));
 sg13g2_a21oi_1 _2073_ (.A1(net292),
    .A2(net195),
    .Y(_0246_),
    .B1(net409));
 sg13g2_and2_1 _2074_ (.A(_0242_),
    .B(_0246_),
    .X(_0247_));
 sg13g2_o21ai_1 _2075_ (.B1(net203),
    .Y(_0248_),
    .A1(_0242_),
    .A2(_0246_));
 sg13g2_nor2_1 _2076_ (.A(_0247_),
    .B(_0248_),
    .Y(_0249_));
 sg13g2_o21ai_1 _2077_ (.B1(net249),
    .Y(_0250_),
    .A1(net409),
    .A2(net203));
 sg13g2_nor2_1 _2078_ (.A(_0249_),
    .B(_0250_),
    .Y(_0099_));
 sg13g2_nand2_1 _2079_ (.Y(_0251_),
    .A(net206),
    .B(_0247_));
 sg13g2_a21oi_1 _2080_ (.A1(net269),
    .A2(_0207_),
    .Y(_0252_),
    .B1(net403));
 sg13g2_o21ai_1 _2081_ (.B1(net249),
    .Y(_0253_),
    .A1(_0251_),
    .A2(_0252_));
 sg13g2_a21oi_1 _2082_ (.A1(_0251_),
    .A2(_0252_),
    .Y(_0100_),
    .B1(_0253_));
 sg13g2_nor2_1 _2083_ (.A(net6),
    .B(net5),
    .Y(_0254_));
 sg13g2_and2_2 _2084_ (.A(_0871_),
    .B(_0254_),
    .X(_0255_));
 sg13g2_a21oi_1 _2085_ (.A1(net1),
    .A2(_0255_),
    .Y(_0256_),
    .B1(net227));
 sg13g2_o21ai_1 _2086_ (.B1(_0256_),
    .Y(_0101_),
    .A1(_0489_),
    .A2(_0255_));
 sg13g2_o21ai_1 _2087_ (.B1(net240),
    .Y(_0257_),
    .A1(net375),
    .A2(_0255_));
 sg13g2_a21oi_1 _2088_ (.A1(_0483_),
    .A2(_0255_),
    .Y(_0102_),
    .B1(_0257_));
 sg13g2_o21ai_1 _2089_ (.B1(net240),
    .Y(_0258_),
    .A1(net363),
    .A2(_0255_));
 sg13g2_a21oi_1 _2090_ (.A1(_0481_),
    .A2(_0255_),
    .Y(_0103_),
    .B1(_0258_));
 sg13g2_o21ai_1 _2091_ (.B1(net240),
    .Y(_0259_),
    .A1(net372),
    .A2(_0255_));
 sg13g2_a21oi_1 _2092_ (.A1(_0479_),
    .A2(_0255_),
    .Y(_0104_),
    .B1(_0259_));
 sg13g2_or2_1 _2093_ (.X(_0260_),
    .B(_0670_),
    .A(_0533_));
 sg13g2_nand2_1 _2094_ (.Y(_0261_),
    .A(net243),
    .B(_0260_));
 sg13g2_a21oi_1 _2095_ (.A1(_0533_),
    .A2(_0670_),
    .Y(_0105_),
    .B1(_0261_));
 sg13g2_xnor2_1 _2096_ (.Y(_0262_),
    .A(net493),
    .B(_0663_));
 sg13g2_and2_1 _2097_ (.A(_0260_),
    .B(_0262_),
    .X(_0263_));
 sg13g2_nor2_1 _2098_ (.A(_0260_),
    .B(_0262_),
    .Y(_0264_));
 sg13g2_nor3_1 _2099_ (.A(net228),
    .B(_0263_),
    .C(_0264_),
    .Y(_0106_));
 sg13g2_nand2_1 _2100_ (.Y(_0265_),
    .A(net475),
    .B(_0611_));
 sg13g2_xnor2_1 _2101_ (.Y(_0266_),
    .A(net475),
    .B(_0611_));
 sg13g2_a21oi_1 _2102_ (.A1(\genblk4[3].pwm.accumulator[1] ),
    .A2(_0663_),
    .Y(_0267_),
    .B1(_0264_));
 sg13g2_o21ai_1 _2103_ (.B1(net236),
    .Y(_0268_),
    .A1(_0266_),
    .A2(_0267_));
 sg13g2_a21oi_1 _2104_ (.A1(_0266_),
    .A2(_0267_),
    .Y(_0107_),
    .B1(_0268_));
 sg13g2_xnor2_1 _2105_ (.Y(_0269_),
    .A(net494),
    .B(_0636_));
 sg13g2_o21ai_1 _2106_ (.B1(_0265_),
    .Y(_0270_),
    .A1(_0266_),
    .A2(_0267_));
 sg13g2_and2_1 _2107_ (.A(_0269_),
    .B(_0270_),
    .X(_0271_));
 sg13g2_o21ai_1 _2108_ (.B1(net236),
    .Y(_0272_),
    .A1(_0269_),
    .A2(_0270_));
 sg13g2_nor2_1 _2109_ (.A(_0271_),
    .B(_0272_),
    .Y(_0108_));
 sg13g2_xor2_1 _2110_ (.B(_0681_),
    .A(net501),
    .X(_0273_));
 sg13g2_a21oi_1 _2111_ (.A1(net494),
    .A2(_0637_),
    .Y(_0274_),
    .B1(_0271_));
 sg13g2_and2_1 _2112_ (.A(_0273_),
    .B(_0274_),
    .X(_0275_));
 sg13g2_nor2_1 _2113_ (.A(_0273_),
    .B(_0274_),
    .Y(_0276_));
 sg13g2_nor3_1 _2114_ (.A(net224),
    .B(_0275_),
    .C(_0276_),
    .Y(_0109_));
 sg13g2_a21oi_2 _2115_ (.B1(_0276_),
    .Y(_0277_),
    .A2(_0682_),
    .A1(\genblk4[3].pwm.accumulator[4] ));
 sg13g2_nand2_1 _2116_ (.Y(_0278_),
    .A(\genblk4[3].pwm.accumulator[5] ),
    .B(_0714_));
 sg13g2_nor2_1 _2117_ (.A(\genblk4[3].pwm.accumulator[5] ),
    .B(_0714_),
    .Y(_0279_));
 sg13g2_xnor2_1 _2118_ (.Y(_0280_),
    .A(net486),
    .B(_0714_));
 sg13g2_xnor2_1 _2119_ (.Y(_0281_),
    .A(_0277_),
    .B(_0280_));
 sg13g2_nor2_1 _2120_ (.A(net224),
    .B(net487),
    .Y(_0110_));
 sg13g2_nor2b_1 _2121_ (.A(_0722_),
    .B_N(\genblk4[3].pwm.accumulator[6] ),
    .Y(_0282_));
 sg13g2_xnor2_1 _2122_ (.Y(_0283_),
    .A(net456),
    .B(_0722_));
 sg13g2_o21ai_1 _2123_ (.B1(_0278_),
    .Y(_0284_),
    .A1(_0277_),
    .A2(_0279_));
 sg13g2_o21ai_1 _2124_ (.B1(net234),
    .Y(_0285_),
    .A1(_0283_),
    .A2(_0284_));
 sg13g2_a21oi_1 _2125_ (.A1(_0283_),
    .A2(_0284_),
    .Y(_0111_),
    .B1(_0285_));
 sg13g2_a21oi_1 _2126_ (.A1(_0283_),
    .A2(_0284_),
    .Y(_0286_),
    .B1(_0282_));
 sg13g2_nand2_1 _2127_ (.Y(_0287_),
    .A(net433),
    .B(_0749_));
 sg13g2_xnor2_1 _2128_ (.Y(_0288_),
    .A(net433),
    .B(_0749_));
 sg13g2_or2_1 _2129_ (.X(_0289_),
    .B(_0288_),
    .A(_0286_));
 sg13g2_nand2_1 _2130_ (.Y(_0290_),
    .A(net234),
    .B(_0289_));
 sg13g2_a21oi_1 _2131_ (.A1(_0286_),
    .A2(_0288_),
    .Y(_0112_),
    .B1(_0290_));
 sg13g2_and2_1 _2132_ (.A(_0287_),
    .B(_0289_),
    .X(_0291_));
 sg13g2_xnor2_1 _2133_ (.Y(_0292_),
    .A(net440),
    .B(_0770_));
 sg13g2_nor2_1 _2134_ (.A(_0291_),
    .B(_0292_),
    .Y(_0293_));
 sg13g2_a21oi_1 _2135_ (.A1(_0291_),
    .A2(_0292_),
    .Y(_0294_),
    .B1(net224));
 sg13g2_nor2b_1 _2136_ (.A(_0293_),
    .B_N(_0294_),
    .Y(_0113_));
 sg13g2_nand2_1 _2137_ (.Y(_0295_),
    .A(net359),
    .B(_0791_));
 sg13g2_xnor2_1 _2138_ (.Y(_0296_),
    .A(net359),
    .B(_0791_));
 sg13g2_a21oi_2 _2139_ (.B1(_0293_),
    .Y(_0297_),
    .A2(_0770_),
    .A1(net440));
 sg13g2_o21ai_1 _2140_ (.B1(net234),
    .Y(_0298_),
    .A1(_0296_),
    .A2(_0297_));
 sg13g2_a21oi_1 _2141_ (.A1(_0296_),
    .A2(_0297_),
    .Y(_0114_),
    .B1(_0298_));
 sg13g2_o21ai_1 _2142_ (.B1(net234),
    .Y(_0299_),
    .A1(net359),
    .A2(_0791_));
 sg13g2_a21oi_1 _2143_ (.A1(_0295_),
    .A2(_0297_),
    .Y(_0115_),
    .B1(_0299_));
 sg13g2_o21ai_1 _2144_ (.B1(net237),
    .Y(_0300_),
    .A1(\noise[0].gen.counter[0] ),
    .A2(net199));
 sg13g2_a21oi_1 _2145_ (.A1(_0488_),
    .A2(net199),
    .Y(_0116_),
    .B1(_0300_));
 sg13g2_a21oi_1 _2146_ (.A1(\noise[0].gen.counter[0] ),
    .A2(net199),
    .Y(_0301_),
    .B1(net273));
 sg13g2_nand3_1 _2147_ (.B(\noise[0].gen.counter[0] ),
    .C(net199),
    .A(net273),
    .Y(_0302_));
 sg13g2_nand2_1 _2148_ (.Y(_0303_),
    .A(net237),
    .B(_0302_));
 sg13g2_nor2_1 _2149_ (.A(net274),
    .B(_0303_),
    .Y(_0117_));
 sg13g2_and2_1 _2150_ (.A(_0487_),
    .B(_0302_),
    .X(_0304_));
 sg13g2_nor2_1 _2151_ (.A(_0487_),
    .B(_0302_),
    .Y(_0305_));
 sg13g2_nor3_1 _2152_ (.A(net227),
    .B(net423),
    .C(_0305_),
    .Y(_0118_));
 sg13g2_or2_1 _2153_ (.X(_0306_),
    .B(_0305_),
    .A(net461));
 sg13g2_nand2_1 _2154_ (.Y(_0307_),
    .A(net461),
    .B(_0305_));
 sg13g2_and3_1 _2155_ (.X(_0119_),
    .A(net237),
    .B(_0306_),
    .C(_0307_));
 sg13g2_xor2_1 _2156_ (.B(_0307_),
    .A(net369),
    .X(_0308_));
 sg13g2_nor2_1 _2157_ (.A(net225),
    .B(net370),
    .Y(_0120_));
 sg13g2_nor2_1 _2158_ (.A(_0004_),
    .B(_0307_),
    .Y(_0309_));
 sg13g2_o21ai_1 _2159_ (.B1(net237),
    .Y(_0310_),
    .A1(net299),
    .A2(_0309_));
 sg13g2_a21oi_1 _2160_ (.A1(net299),
    .A2(_0309_),
    .Y(_0121_),
    .B1(_0310_));
 sg13g2_nand4_1 _2161_ (.B(\noise[0].gen.counter[4] ),
    .C(\noise[0].gen.counter[3] ),
    .A(net299),
    .Y(_0311_),
    .D(_0305_));
 sg13g2_o21ai_1 _2162_ (.B1(net237),
    .Y(_0312_),
    .A1(_0486_),
    .A2(_0311_));
 sg13g2_a21oi_1 _2163_ (.A1(_0486_),
    .A2(_0311_),
    .Y(_0122_),
    .B1(_0312_));
 sg13g2_nor2b_1 _2164_ (.A(net349),
    .B_N(_0937_),
    .Y(_0313_));
 sg13g2_nand2b_1 _2165_ (.Y(_0314_),
    .B(_0937_),
    .A_N(net349));
 sg13g2_nor2_1 _2166_ (.A(net354),
    .B(_0314_),
    .Y(_0315_));
 sg13g2_nand2b_1 _2167_ (.Y(_0316_),
    .B(net233),
    .A_N(net341));
 sg13g2_nor2_1 _2168_ (.A(net217),
    .B(net194),
    .Y(_0317_));
 sg13g2_nor3_1 _2169_ (.A(_0315_),
    .B(net215),
    .C(_0317_),
    .Y(_0123_));
 sg13g2_nor2_1 _2170_ (.A(\noise[0].gen.lfsr[2] ),
    .B(net192),
    .Y(_0318_));
 sg13g2_nor2_1 _2171_ (.A(net354),
    .B(net194),
    .Y(_0319_));
 sg13g2_nor3_1 _2172_ (.A(net215),
    .B(_0318_),
    .C(_0319_),
    .Y(_0124_));
 sg13g2_nor2_1 _2173_ (.A(\noise[0].gen.lfsr[2] ),
    .B(net194),
    .Y(_0320_));
 sg13g2_nor2_1 _2174_ (.A(net308),
    .B(net192),
    .Y(_0321_));
 sg13g2_nor3_1 _2175_ (.A(net215),
    .B(_0320_),
    .C(_0321_),
    .Y(_0125_));
 sg13g2_nor2_1 _2176_ (.A(net308),
    .B(net194),
    .Y(_0322_));
 sg13g2_nor2_1 _2177_ (.A(net317),
    .B(net192),
    .Y(_0323_));
 sg13g2_nor3_1 _2178_ (.A(net215),
    .B(_0322_),
    .C(_0323_),
    .Y(_0126_));
 sg13g2_nor2_1 _2179_ (.A(net314),
    .B(net192),
    .Y(_0324_));
 sg13g2_nor2_1 _2180_ (.A(net317),
    .B(net194),
    .Y(_0325_));
 sg13g2_nor3_1 _2181_ (.A(net215),
    .B(_0324_),
    .C(net318),
    .Y(_0127_));
 sg13g2_nor2_1 _2182_ (.A(\noise[0].gen.lfsr[6] ),
    .B(net192),
    .Y(_0326_));
 sg13g2_nor2_1 _2183_ (.A(net314),
    .B(net194),
    .Y(_0327_));
 sg13g2_nor3_1 _2184_ (.A(net215),
    .B(_0326_),
    .C(net315),
    .Y(_0128_));
 sg13g2_nor2_1 _2185_ (.A(net311),
    .B(net192),
    .Y(_0328_));
 sg13g2_nor2_1 _2186_ (.A(net325),
    .B(net193),
    .Y(_0329_));
 sg13g2_nor3_1 _2187_ (.A(net215),
    .B(_0328_),
    .C(net326),
    .Y(_0129_));
 sg13g2_nor2_1 _2188_ (.A(\noise[0].gen.lfsr[8] ),
    .B(net192),
    .Y(_0330_));
 sg13g2_nor2_1 _2189_ (.A(net311),
    .B(net193),
    .Y(_0331_));
 sg13g2_nor3_1 _2190_ (.A(net214),
    .B(_0330_),
    .C(net312),
    .Y(_0130_));
 sg13g2_nor2_1 _2191_ (.A(net328),
    .B(net191),
    .Y(_0332_));
 sg13g2_nor2_1 _2192_ (.A(\noise[0].gen.lfsr[8] ),
    .B(net193),
    .Y(_0333_));
 sg13g2_nor3_1 _2193_ (.A(net214),
    .B(_0332_),
    .C(_0333_),
    .Y(_0131_));
 sg13g2_nor2_1 _2194_ (.A(\noise[0].gen.lfsr[9] ),
    .B(net193),
    .Y(_0334_));
 sg13g2_nor2_1 _2195_ (.A(net301),
    .B(net191),
    .Y(_0335_));
 sg13g2_nor3_1 _2196_ (.A(net214),
    .B(_0334_),
    .C(_0335_),
    .Y(_0132_));
 sg13g2_nor2_1 _2197_ (.A(net303),
    .B(net191),
    .Y(_0336_));
 sg13g2_nor2_1 _2198_ (.A(net301),
    .B(net193),
    .Y(_0337_));
 sg13g2_nor3_1 _2199_ (.A(net214),
    .B(_0336_),
    .C(_0337_),
    .Y(_0133_));
 sg13g2_nor2_1 _2200_ (.A(\noise[0].gen.lfsr[12] ),
    .B(net191),
    .Y(_0338_));
 sg13g2_nor2_1 _2201_ (.A(net303),
    .B(net193),
    .Y(_0339_));
 sg13g2_nor3_1 _2202_ (.A(net214),
    .B(_0338_),
    .C(net304),
    .Y(_0134_));
 sg13g2_nor2_1 _2203_ (.A(\noise[0].gen.lfsr[13] ),
    .B(net191),
    .Y(_0340_));
 sg13g2_nor2_1 _2204_ (.A(net322),
    .B(net193),
    .Y(_0341_));
 sg13g2_nor3_1 _2205_ (.A(net214),
    .B(_0340_),
    .C(net323),
    .Y(_0135_));
 sg13g2_nor2_1 _2206_ (.A(\noise[0].gen.lfsr[14] ),
    .B(net191),
    .Y(_0342_));
 sg13g2_nor2_1 _2207_ (.A(net338),
    .B(net193),
    .Y(_0343_));
 sg13g2_nor3_1 _2208_ (.A(net214),
    .B(_0342_),
    .C(net339),
    .Y(_0136_));
 sg13g2_nand2_1 _2209_ (.Y(_0344_),
    .A(net354),
    .B(\control_noise[0][2] ));
 sg13g2_xor2_1 _2210_ (.B(_0344_),
    .A(net217),
    .X(_0345_));
 sg13g2_a21oi_1 _2211_ (.A1(net366),
    .A2(net191),
    .Y(_0346_),
    .B1(net214));
 sg13g2_o21ai_1 _2212_ (.B1(_0346_),
    .Y(_0137_),
    .A1(net191),
    .A2(_0345_));
 sg13g2_and2_2 _2213_ (.A(_0871_),
    .B(_0932_),
    .X(_0347_));
 sg13g2_a21oi_1 _2214_ (.A1(net1),
    .A2(_0347_),
    .Y(_0348_),
    .B1(net227));
 sg13g2_o21ai_1 _2215_ (.B1(_0348_),
    .Y(_0138_),
    .A1(_0485_),
    .A2(_0347_));
 sg13g2_o21ai_1 _2216_ (.B1(net238),
    .Y(_0349_),
    .A1(net391),
    .A2(_0347_));
 sg13g2_a21oi_1 _2217_ (.A1(_0483_),
    .A2(_0347_),
    .Y(_0139_),
    .B1(_0349_));
 sg13g2_o21ai_1 _2218_ (.B1(net238),
    .Y(_0350_),
    .A1(net383),
    .A2(_0347_));
 sg13g2_a21oi_1 _2219_ (.A1(_0481_),
    .A2(_0347_),
    .Y(_0140_),
    .B1(_0350_));
 sg13g2_o21ai_1 _2220_ (.B1(net238),
    .Y(_0351_),
    .A1(net410),
    .A2(_0347_));
 sg13g2_a21oi_1 _2221_ (.A1(_0479_),
    .A2(_0347_),
    .Y(_0141_),
    .B1(_0351_));
 sg13g2_nand2_2 _2222_ (.Y(_0352_),
    .A(_0899_),
    .B(_0254_));
 sg13g2_a21oi_1 _2223_ (.A1(net396),
    .A2(_0352_),
    .Y(_0353_),
    .B1(net228));
 sg13g2_o21ai_1 _2224_ (.B1(_0353_),
    .Y(_0142_),
    .A1(_0484_),
    .A2(_0352_));
 sg13g2_o21ai_1 _2225_ (.B1(net247),
    .Y(_0354_),
    .A1(net2),
    .A2(_0352_));
 sg13g2_a21oi_1 _2226_ (.A1(_0482_),
    .A2(_0352_),
    .Y(_0143_),
    .B1(_0354_));
 sg13g2_o21ai_1 _2227_ (.B1(net247),
    .Y(_0355_),
    .A1(net3),
    .A2(_0352_));
 sg13g2_a21oi_1 _2228_ (.A1(_0480_),
    .A2(_0352_),
    .Y(_0144_),
    .B1(_0355_));
 sg13g2_o21ai_1 _2229_ (.B1(net246),
    .Y(_0356_),
    .A1(net4),
    .A2(_0352_));
 sg13g2_a21oi_1 _2230_ (.A1(_0478_),
    .A2(_0352_),
    .Y(_0145_),
    .B1(_0356_));
 sg13g2_nand2_1 _2231_ (.Y(_0357_),
    .A(net393),
    .B(_0642_));
 sg13g2_o21ai_1 _2232_ (.B1(net233),
    .Y(_0358_),
    .A1(net393),
    .A2(_0642_));
 sg13g2_nor2b_1 _2233_ (.A(_0358_),
    .B_N(_0357_),
    .Y(_0146_));
 sg13g2_xnor2_1 _2234_ (.Y(_0359_),
    .A(net446),
    .B(_0541_));
 sg13g2_and2_1 _2235_ (.A(_0357_),
    .B(_0359_),
    .X(_0360_));
 sg13g2_nor2_1 _2236_ (.A(_0357_),
    .B(_0359_),
    .Y(_0361_));
 sg13g2_nor3_1 _2237_ (.A(net224),
    .B(_0360_),
    .C(_0361_),
    .Y(_0147_));
 sg13g2_nand2_1 _2238_ (.Y(_0362_),
    .A(net504),
    .B(_0586_));
 sg13g2_xnor2_1 _2239_ (.Y(_0363_),
    .A(\genblk4[0].pwm.accumulator[2] ),
    .B(_0586_));
 sg13g2_a21oi_2 _2240_ (.B1(_0361_),
    .Y(_0364_),
    .A2(_0541_),
    .A1(net446));
 sg13g2_o21ai_1 _2241_ (.B1(net231),
    .Y(_0365_),
    .A1(_0363_),
    .A2(_0364_));
 sg13g2_a21oi_1 _2242_ (.A1(_0363_),
    .A2(_0364_),
    .Y(_0148_),
    .B1(_0365_));
 sg13g2_xnor2_1 _2243_ (.Y(_0366_),
    .A(net436),
    .B(_0626_));
 sg13g2_o21ai_1 _2244_ (.B1(_0362_),
    .Y(_0367_),
    .A1(_0363_),
    .A2(_0364_));
 sg13g2_and2_1 _2245_ (.A(_0366_),
    .B(_0367_),
    .X(_0368_));
 sg13g2_o21ai_1 _2246_ (.B1(net231),
    .Y(_0369_),
    .A1(_0366_),
    .A2(_0367_));
 sg13g2_nor2_1 _2247_ (.A(_0368_),
    .B(_0369_),
    .Y(_0149_));
 sg13g2_nand2_1 _2248_ (.Y(_0370_),
    .A(\genblk4[0].pwm.accumulator[4] ),
    .B(_0685_));
 sg13g2_xor2_1 _2249_ (.B(_0684_),
    .A(\genblk4[0].pwm.accumulator[4] ),
    .X(_0371_));
 sg13g2_a21oi_2 _2250_ (.B1(_0368_),
    .Y(_0372_),
    .A2(_0627_),
    .A1(net436));
 sg13g2_o21ai_1 _2251_ (.B1(net231),
    .Y(_0373_),
    .A1(_0371_),
    .A2(_0372_));
 sg13g2_a21oi_1 _2252_ (.A1(_0371_),
    .A2(_0372_),
    .Y(_0150_),
    .B1(_0373_));
 sg13g2_o21ai_1 _2253_ (.B1(_0370_),
    .Y(_0374_),
    .A1(_0371_),
    .A2(_0372_));
 sg13g2_nor2_1 _2254_ (.A(\genblk4[0].pwm.accumulator[5] ),
    .B(_0701_),
    .Y(_0375_));
 sg13g2_xor2_1 _2255_ (.B(_0701_),
    .A(net477),
    .X(_0376_));
 sg13g2_o21ai_1 _2256_ (.B1(net231),
    .Y(_0377_),
    .A1(_0374_),
    .A2(_0376_));
 sg13g2_a21oi_1 _2257_ (.A1(_0374_),
    .A2(_0376_),
    .Y(_0151_),
    .B1(_0377_));
 sg13g2_nor2b_1 _2258_ (.A(_0729_),
    .B_N(\genblk4[0].pwm.accumulator[6] ),
    .Y(_0378_));
 sg13g2_xnor2_1 _2259_ (.Y(_0379_),
    .A(net462),
    .B(_0729_));
 sg13g2_a21oi_1 _2260_ (.A1(\genblk4[0].pwm.accumulator[5] ),
    .A2(_0701_),
    .Y(_0380_),
    .B1(_0374_));
 sg13g2_nor2_1 _2261_ (.A(_0375_),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_o21ai_1 _2262_ (.B1(net231),
    .Y(_0382_),
    .A1(_0379_),
    .A2(_0381_));
 sg13g2_a21oi_1 _2263_ (.A1(_0379_),
    .A2(_0381_),
    .Y(_0152_),
    .B1(_0382_));
 sg13g2_a21oi_1 _2264_ (.A1(_0379_),
    .A2(_0381_),
    .Y(_0383_),
    .B1(_0378_));
 sg13g2_nand2_1 _2265_ (.Y(_0384_),
    .A(net441),
    .B(_0756_));
 sg13g2_xnor2_1 _2266_ (.Y(_0385_),
    .A(net441),
    .B(_0756_));
 sg13g2_or2_1 _2267_ (.X(_0386_),
    .B(_0385_),
    .A(_0383_));
 sg13g2_nand2_1 _2268_ (.Y(_0387_),
    .A(net235),
    .B(_0386_));
 sg13g2_a21oi_1 _2269_ (.A1(_0383_),
    .A2(_0385_),
    .Y(_0153_),
    .B1(_0387_));
 sg13g2_and2_1 _2270_ (.A(_0384_),
    .B(_0386_),
    .X(_0388_));
 sg13g2_xor2_1 _2271_ (.B(_0774_),
    .A(net445),
    .X(_0389_));
 sg13g2_nor2_1 _2272_ (.A(_0388_),
    .B(_0389_),
    .Y(_0390_));
 sg13g2_a21oi_1 _2273_ (.A1(_0388_),
    .A2(_0389_),
    .Y(_0391_),
    .B1(net224));
 sg13g2_nor2b_1 _2274_ (.A(_0390_),
    .B_N(_0391_),
    .Y(_0154_));
 sg13g2_nand2_1 _2275_ (.Y(_0392_),
    .A(net373),
    .B(_0793_));
 sg13g2_xnor2_1 _2276_ (.Y(_0393_),
    .A(net373),
    .B(_0793_));
 sg13g2_a21oi_2 _2277_ (.B1(_0390_),
    .Y(_0394_),
    .A2(_0775_),
    .A1(net445));
 sg13g2_o21ai_1 _2278_ (.B1(net235),
    .Y(_0395_),
    .A1(_0393_),
    .A2(_0394_));
 sg13g2_a21oi_1 _2279_ (.A1(_0393_),
    .A2(_0394_),
    .Y(_0155_),
    .B1(_0395_));
 sg13g2_o21ai_1 _2280_ (.B1(net234),
    .Y(_0396_),
    .A1(net373),
    .A2(_0793_));
 sg13g2_a21oi_1 _2281_ (.A1(_0392_),
    .A2(_0394_),
    .Y(_0156_),
    .B1(_0396_));
 sg13g2_or2_1 _2282_ (.X(_0397_),
    .B(_0648_),
    .A(_0529_));
 sg13g2_nand2_1 _2283_ (.Y(_0398_),
    .A(net233),
    .B(_0397_));
 sg13g2_a21oi_1 _2284_ (.A1(_0529_),
    .A2(_0648_),
    .Y(_0157_),
    .B1(_0398_));
 sg13g2_nand2_1 _2285_ (.Y(_0399_),
    .A(net464),
    .B(_0552_));
 sg13g2_xor2_1 _2286_ (.B(_0552_),
    .A(net464),
    .X(_0400_));
 sg13g2_inv_1 _2287_ (.Y(_0401_),
    .A(_0400_));
 sg13g2_nand2b_1 _2288_ (.Y(_0402_),
    .B(_0400_),
    .A_N(_0397_));
 sg13g2_nand2_1 _2289_ (.Y(_0403_),
    .A(net232),
    .B(_0402_));
 sg13g2_a21oi_1 _2290_ (.A1(_0397_),
    .A2(_0401_),
    .Y(_0158_),
    .B1(_0403_));
 sg13g2_nand2_1 _2291_ (.Y(_0404_),
    .A(net488),
    .B(_0592_));
 sg13g2_xnor2_1 _2292_ (.Y(_0405_),
    .A(net488),
    .B(_0592_));
 sg13g2_nand3_1 _2293_ (.B(_0402_),
    .C(_0405_),
    .A(_0399_),
    .Y(_0406_));
 sg13g2_a21o_1 _2294_ (.A2(_0402_),
    .A1(_0399_),
    .B1(_0405_),
    .X(_0407_));
 sg13g2_and3_1 _2295_ (.X(_0159_),
    .A(net232),
    .B(_0406_),
    .C(_0407_));
 sg13g2_nand2_1 _2296_ (.Y(_0408_),
    .A(net496),
    .B(_0623_));
 sg13g2_xnor2_1 _2297_ (.Y(_0409_),
    .A(\genblk4[1].pwm.accumulator[3] ),
    .B(_0623_));
 sg13g2_nand3_1 _2298_ (.B(_0407_),
    .C(_0409_),
    .A(_0404_),
    .Y(_0410_));
 sg13g2_a21o_1 _2299_ (.A2(_0407_),
    .A1(_0404_),
    .B1(_0409_),
    .X(_0411_));
 sg13g2_and3_1 _2300_ (.X(_0160_),
    .A(net232),
    .B(net489),
    .C(_0411_));
 sg13g2_nor2b_1 _2301_ (.A(_0686_),
    .B_N(\genblk4[1].pwm.accumulator[4] ),
    .Y(_0412_));
 sg13g2_xnor2_1 _2302_ (.Y(_0413_),
    .A(\genblk4[1].pwm.accumulator[4] ),
    .B(_0686_));
 sg13g2_nand2_1 _2303_ (.Y(_0414_),
    .A(_0408_),
    .B(_0411_));
 sg13g2_nor2_1 _2304_ (.A(_0413_),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_and2_1 _2305_ (.A(_0413_),
    .B(_0414_),
    .X(_0416_));
 sg13g2_nor3_1 _2306_ (.A(net224),
    .B(net497),
    .C(_0416_),
    .Y(_0161_));
 sg13g2_a21oi_1 _2307_ (.A1(_0413_),
    .A2(_0414_),
    .Y(_0417_),
    .B1(_0412_));
 sg13g2_nand2_1 _2308_ (.Y(_0418_),
    .A(net484),
    .B(_0703_));
 sg13g2_nor2_1 _2309_ (.A(\genblk4[1].pwm.accumulator[5] ),
    .B(_0703_),
    .Y(_0419_));
 sg13g2_xnor2_1 _2310_ (.Y(_0420_),
    .A(net484),
    .B(_0703_));
 sg13g2_xnor2_1 _2311_ (.Y(_0421_),
    .A(_0417_),
    .B(_0420_));
 sg13g2_nor2_1 _2312_ (.A(net224),
    .B(net485),
    .Y(_0162_));
 sg13g2_xnor2_1 _2313_ (.Y(_0422_),
    .A(net505),
    .B(_0732_));
 sg13g2_o21ai_1 _2314_ (.B1(_0418_),
    .Y(_0423_),
    .A1(_0417_),
    .A2(_0419_));
 sg13g2_nand2_1 _2315_ (.Y(_0424_),
    .A(_0422_),
    .B(_0423_));
 sg13g2_o21ai_1 _2316_ (.B1(net232),
    .Y(_0425_),
    .A1(_0422_),
    .A2(_0423_));
 sg13g2_nor2b_1 _2317_ (.A(net506),
    .B_N(_0424_),
    .Y(_0163_));
 sg13g2_o21ai_1 _2318_ (.B1(_0424_),
    .Y(_0426_),
    .A1(_0530_),
    .A2(_0732_));
 sg13g2_xor2_1 _2319_ (.B(_0758_),
    .A(net507),
    .X(_0427_));
 sg13g2_and2_1 _2320_ (.A(_0426_),
    .B(_0427_),
    .X(_0428_));
 sg13g2_o21ai_1 _2321_ (.B1(net231),
    .Y(_0429_),
    .A1(_0426_),
    .A2(_0427_));
 sg13g2_nor2_1 _2322_ (.A(_0428_),
    .B(_0429_),
    .Y(_0164_));
 sg13g2_a21oi_2 _2323_ (.B1(_0428_),
    .Y(_0430_),
    .A2(_0758_),
    .A1(net507));
 sg13g2_xor2_1 _2324_ (.B(_0776_),
    .A(net435),
    .X(_0431_));
 sg13g2_nor2_1 _2325_ (.A(_0430_),
    .B(_0431_),
    .Y(_0432_));
 sg13g2_a21oi_1 _2326_ (.A1(_0430_),
    .A2(_0431_),
    .Y(_0433_),
    .B1(net230));
 sg13g2_nor2b_1 _2327_ (.A(_0432_),
    .B_N(_0433_),
    .Y(_0165_));
 sg13g2_nand2_1 _2328_ (.Y(_0434_),
    .A(net364),
    .B(_0794_));
 sg13g2_xnor2_1 _2329_ (.Y(_0435_),
    .A(net364),
    .B(_0794_));
 sg13g2_a21oi_2 _2330_ (.B1(_0432_),
    .Y(_0436_),
    .A2(_0777_),
    .A1(net435));
 sg13g2_o21ai_1 _2331_ (.B1(net235),
    .Y(_0437_),
    .A1(_0435_),
    .A2(_0436_));
 sg13g2_a21oi_1 _2332_ (.A1(_0435_),
    .A2(_0436_),
    .Y(_0166_),
    .B1(_0437_));
 sg13g2_o21ai_1 _2333_ (.B1(net234),
    .Y(_0438_),
    .A1(net364),
    .A2(_0794_));
 sg13g2_a21oi_1 _2334_ (.A1(_0434_),
    .A2(_0436_),
    .Y(_0167_),
    .B1(_0438_));
 sg13g2_nand2_1 _2335_ (.Y(_0439_),
    .A(net368),
    .B(_0655_));
 sg13g2_o21ai_1 _2336_ (.B1(net233),
    .Y(_0440_),
    .A1(net368),
    .A2(_0655_));
 sg13g2_nor2b_1 _2337_ (.A(_0440_),
    .B_N(_0439_),
    .Y(_0168_));
 sg13g2_nand3_1 _2338_ (.B(_0557_),
    .C(_0569_),
    .A(net502),
    .Y(_0441_));
 sg13g2_xor2_1 _2339_ (.B(_0570_),
    .A(net379),
    .X(_0442_));
 sg13g2_o21ai_1 _2340_ (.B1(net231),
    .Y(_0443_),
    .A1(_0439_),
    .A2(_0442_));
 sg13g2_a21oi_1 _2341_ (.A1(_0439_),
    .A2(_0442_),
    .Y(_0169_),
    .B1(_0443_));
 sg13g2_nand2_1 _2342_ (.Y(_0444_),
    .A(net490),
    .B(_0577_));
 sg13g2_xnor2_1 _2343_ (.Y(_0445_),
    .A(net490),
    .B(_0577_));
 sg13g2_o21ai_1 _2344_ (.B1(_0441_),
    .Y(_0446_),
    .A1(_0439_),
    .A2(_0442_));
 sg13g2_nand2b_1 _2345_ (.Y(_0447_),
    .B(_0445_),
    .A_N(_0446_));
 sg13g2_nand2b_1 _2346_ (.Y(_0448_),
    .B(_0446_),
    .A_N(_0445_));
 sg13g2_and3_1 _2347_ (.X(_0170_),
    .A(net232),
    .B(_0447_),
    .C(_0448_));
 sg13g2_nand2_1 _2348_ (.Y(_0449_),
    .A(net491),
    .B(_0620_));
 sg13g2_xor2_1 _2349_ (.B(_0619_),
    .A(\genblk4[2].pwm.accumulator[3] ),
    .X(_0450_));
 sg13g2_nand3_1 _2350_ (.B(_0448_),
    .C(_0450_),
    .A(_0444_),
    .Y(_0451_));
 sg13g2_a21o_1 _2351_ (.A2(_0448_),
    .A1(_0444_),
    .B1(_0450_),
    .X(_0452_));
 sg13g2_and3_1 _2352_ (.X(_0171_),
    .A(net231),
    .B(_0451_),
    .C(_0452_));
 sg13g2_xnor2_1 _2353_ (.Y(_0453_),
    .A(_0531_),
    .B(_0652_));
 sg13g2_nand3_1 _2354_ (.B(_0452_),
    .C(_0453_),
    .A(_0449_),
    .Y(_0454_));
 sg13g2_a21o_1 _2355_ (.A2(_0452_),
    .A1(_0449_),
    .B1(_0453_),
    .X(_0455_));
 sg13g2_and3_1 _2356_ (.X(_0172_),
    .A(net235),
    .B(_0454_),
    .C(_0455_));
 sg13g2_o21ai_1 _2357_ (.B1(_0455_),
    .Y(_0456_),
    .A1(_0531_),
    .A2(_0652_));
 sg13g2_xnor2_1 _2358_ (.Y(_0457_),
    .A(net450),
    .B(_0707_));
 sg13g2_o21ai_1 _2359_ (.B1(net235),
    .Y(_0458_),
    .A1(_0456_),
    .A2(_0457_));
 sg13g2_a21oi_1 _2360_ (.A1(_0456_),
    .A2(_0457_),
    .Y(_0173_),
    .B1(_0458_));
 sg13g2_xor2_1 _2361_ (.B(_0725_),
    .A(net431),
    .X(_0459_));
 sg13g2_a21oi_1 _2362_ (.A1(net450),
    .A2(_0708_),
    .Y(_0460_),
    .B1(_0456_));
 sg13g2_a21oi_1 _2363_ (.A1(_0532_),
    .A2(_0707_),
    .Y(_0461_),
    .B1(_0460_));
 sg13g2_and2_1 _2364_ (.A(_0459_),
    .B(_0461_),
    .X(_0462_));
 sg13g2_o21ai_1 _2365_ (.B1(net235),
    .Y(_0463_),
    .A1(_0459_),
    .A2(_0461_));
 sg13g2_nor2_1 _2366_ (.A(_0462_),
    .B(_0463_),
    .Y(_0174_));
 sg13g2_a21oi_1 _2367_ (.A1(net431),
    .A2(_0725_),
    .Y(_0464_),
    .B1(_0462_));
 sg13g2_nand2_1 _2368_ (.Y(_0465_),
    .A(net495),
    .B(_0754_));
 sg13g2_xor2_1 _2369_ (.B(_0753_),
    .A(\genblk4[2].pwm.accumulator[7] ),
    .X(_0466_));
 sg13g2_or2_1 _2370_ (.X(_0467_),
    .B(_0466_),
    .A(_0464_));
 sg13g2_nand2_1 _2371_ (.Y(_0468_),
    .A(net235),
    .B(_0467_));
 sg13g2_a21oi_1 _2372_ (.A1(_0464_),
    .A2(_0466_),
    .Y(_0175_),
    .B1(_0468_));
 sg13g2_and2_1 _2373_ (.A(_0465_),
    .B(_0467_),
    .X(_0469_));
 sg13g2_xnor2_1 _2374_ (.Y(_0470_),
    .A(net448),
    .B(_0773_));
 sg13g2_nor2_1 _2375_ (.A(_0469_),
    .B(_0470_),
    .Y(_0471_));
 sg13g2_a21oi_1 _2376_ (.A1(_0469_),
    .A2(_0470_),
    .Y(_0472_),
    .B1(net230));
 sg13g2_nor2b_1 _2377_ (.A(_0471_),
    .B_N(_0472_),
    .Y(_0176_));
 sg13g2_nand2_1 _2378_ (.Y(_0473_),
    .A(net356),
    .B(_0653_));
 sg13g2_xnor2_1 _2379_ (.Y(_0474_),
    .A(net356),
    .B(_0653_));
 sg13g2_a21oi_1 _2380_ (.A1(net448),
    .A2(_0773_),
    .Y(_0475_),
    .B1(_0471_));
 sg13g2_o21ai_1 _2381_ (.B1(net234),
    .Y(_0476_),
    .A1(_0474_),
    .A2(_0475_));
 sg13g2_a21oi_1 _2382_ (.A1(_0474_),
    .A2(_0475_),
    .Y(_0177_),
    .B1(_0476_));
 sg13g2_o21ai_1 _2383_ (.B1(net234),
    .Y(_0477_),
    .A1(net356),
    .A2(_0653_));
 sg13g2_a21oi_1 _2384_ (.A1(net357),
    .A2(_0475_),
    .Y(_0178_),
    .B1(_0477_));
 sg13g2_nor2_1 _2385_ (.A(net225),
    .B(_0933_),
    .Y(_0179_));
 sg13g2_dfrbp_1 _2386_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net160),
    .D(_0007_),
    .Q_N(_1188_),
    .Q(\pwm.accumulator[0] ));
 sg13g2_dfrbp_1 _2387_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net150),
    .D(net416),
    .Q_N(_1187_),
    .Q(\pwm.accumulator[1] ));
 sg13g2_dfrbp_1 _2388_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net149),
    .D(net483),
    .Q_N(_1186_),
    .Q(\pwm.accumulator[2] ));
 sg13g2_dfrbp_1 _2389_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net148),
    .D(net470),
    .Q_N(_1185_),
    .Q(\pwm.accumulator[3] ));
 sg13g2_dfrbp_1 _2390_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net147),
    .D(_0011_),
    .Q_N(_1184_),
    .Q(\pwm.accumulator[4] ));
 sg13g2_dfrbp_1 _2391_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net146),
    .D(net466),
    .Q_N(_1183_),
    .Q(\pwm.accumulator[5] ));
 sg13g2_dfrbp_1 _2392_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net145),
    .D(_0013_),
    .Q_N(_1182_),
    .Q(\pwm.accumulator[6] ));
 sg13g2_dfrbp_1 _2393_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net144),
    .D(net459),
    .Q_N(_1181_),
    .Q(\pwm.accumulator[7] ));
 sg13g2_dfrbp_1 _2394_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net143),
    .D(_0015_),
    .Q_N(_1180_),
    .Q(\pwm.accumulator[8] ));
 sg13g2_dfrbp_1 _2395_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net142),
    .D(net453),
    .Q_N(_1179_),
    .Q(\pwm.accumulator[9] ));
 sg13g2_dfrbp_1 _2396_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net141),
    .D(net468),
    .Q_N(_1178_),
    .Q(\pwm.accumulator[10] ));
 sg13g2_dfrbp_1 _2397_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net140),
    .D(_0018_),
    .Q_N(_1177_),
    .Q(\pwm.accumulator[11] ));
 sg13g2_dfrbp_1 _2398_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net139),
    .D(net348),
    .Q_N(_1176_),
    .Q(\pwm.accumulator[12] ));
 sg13g2_dfrbp_1 _2399_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net138),
    .D(_0020_),
    .Q_N(_1175_),
    .Q(\latch_control_reg[0] ));
 sg13g2_dfrbp_1 _2400_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net136),
    .D(_0021_),
    .Q_N(_1174_),
    .Q(\latch_control_reg[1] ));
 sg13g2_dfrbp_1 _2401_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net134),
    .D(_0022_),
    .Q_N(_0003_),
    .Q(\latch_control_reg[2] ));
 sg13g2_dfrbp_1 _2402_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net132),
    .D(_0023_),
    .Q_N(_0006_),
    .Q(\clk_counter[0] ));
 sg13g2_dfrbp_1 _2403_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net131),
    .D(net351),
    .Q_N(_1173_),
    .Q(\clk_counter[1] ));
 sg13g2_dfrbp_1 _2404_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net130),
    .D(net289),
    .Q_N(_1172_),
    .Q(\clk_counter[2] ));
 sg13g2_dfrbp_1 _2405_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net129),
    .D(_0026_),
    .Q_N(_1171_),
    .Q(\clk_counter[3] ));
 sg13g2_dfrbp_1 _2406_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net128),
    .D(_0027_),
    .Q_N(_1170_),
    .Q(\clk_counter[4] ));
 sg13g2_dfrbp_1 _2407_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net127),
    .D(_0028_),
    .Q_N(_1169_),
    .Q(\clk_counter[5] ));
 sg13g2_dfrbp_1 _2408_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net126),
    .D(net353),
    .Q_N(_1168_),
    .Q(\clk_counter[6] ));
 sg13g2_dfrbp_1 _2409_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net125),
    .D(_0030_),
    .Q_N(_1167_),
    .Q(\chan[0].attenuation.control[0] ));
 sg13g2_dfrbp_1 _2410_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net123),
    .D(_0031_),
    .Q_N(_1166_),
    .Q(\chan[0].attenuation.control[1] ));
 sg13g2_dfrbp_1 _2411_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net121),
    .D(_0032_),
    .Q_N(_1165_),
    .Q(\chan[0].attenuation.control[2] ));
 sg13g2_dfrbp_1 _2412_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net119),
    .D(_0033_),
    .Q_N(_1164_),
    .Q(\chan[0].attenuation.control[3] ));
 sg13g2_dfrbp_1 _2413_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net117),
    .D(_0034_),
    .Q_N(_1163_),
    .Q(\chan[1].attenuation.control[0] ));
 sg13g2_dfrbp_1 _2414_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net115),
    .D(_0035_),
    .Q_N(_1162_),
    .Q(\chan[1].attenuation.control[1] ));
 sg13g2_dfrbp_1 _2415_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net113),
    .D(_0036_),
    .Q_N(_1161_),
    .Q(\chan[1].attenuation.control[2] ));
 sg13g2_dfrbp_1 _2416_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net111),
    .D(_0037_),
    .Q_N(_1160_),
    .Q(\chan[1].attenuation.control[3] ));
 sg13g2_dfrbp_1 _2417_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net109),
    .D(_0038_),
    .Q_N(_1159_),
    .Q(\chan[2].attenuation.control[0] ));
 sg13g2_dfrbp_1 _2418_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net107),
    .D(_0039_),
    .Q_N(_1158_),
    .Q(\chan[2].attenuation.control[1] ));
 sg13g2_dfrbp_1 _2419_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net105),
    .D(_0040_),
    .Q_N(_1157_),
    .Q(\chan[2].attenuation.control[2] ));
 sg13g2_dfrbp_1 _2420_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net103),
    .D(_0041_),
    .Q_N(_1156_),
    .Q(\chan[2].attenuation.control[3] ));
 sg13g2_dfrbp_1 _2421_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net101),
    .D(_0042_),
    .Q_N(_1155_),
    .Q(\chan[3].attenuation.control[0] ));
 sg13g2_dfrbp_1 _2422_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net99),
    .D(_0043_),
    .Q_N(_1154_),
    .Q(\chan[3].attenuation.control[1] ));
 sg13g2_dfrbp_1 _2423_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net97),
    .D(_0044_),
    .Q_N(_1153_),
    .Q(\chan[3].attenuation.control[2] ));
 sg13g2_dfrbp_1 _2424_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net95),
    .D(_0045_),
    .Q_N(_1152_),
    .Q(\chan[3].attenuation.control[3] ));
 sg13g2_dfrbp_1 _2425_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net93),
    .D(_0046_),
    .Q_N(_1151_),
    .Q(\control_tone_freq[0][4] ));
 sg13g2_dfrbp_1 _2426_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net91),
    .D(_0047_),
    .Q_N(_1150_),
    .Q(\control_tone_freq[0][5] ));
 sg13g2_dfrbp_1 _2427_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net89),
    .D(_0048_),
    .Q_N(_1149_),
    .Q(\control_tone_freq[0][6] ));
 sg13g2_dfrbp_1 _2428_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net87),
    .D(_0049_),
    .Q_N(_1148_),
    .Q(\control_tone_freq[0][7] ));
 sg13g2_dfrbp_1 _2429_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net85),
    .D(_0050_),
    .Q_N(_1147_),
    .Q(\control_tone_freq[0][8] ));
 sg13g2_dfrbp_1 _2430_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net83),
    .D(_0051_),
    .Q_N(_1146_),
    .Q(\control_tone_freq[0][9] ));
 sg13g2_dfrbp_1 _2431_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net81),
    .D(net280),
    .Q_N(_1145_),
    .Q(\control_tone_freq[1][4] ));
 sg13g2_dfrbp_1 _2432_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net79),
    .D(net282),
    .Q_N(_1144_),
    .Q(\control_tone_freq[1][5] ));
 sg13g2_dfrbp_1 _2433_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net77),
    .D(_0054_),
    .Q_N(_1143_),
    .Q(\control_tone_freq[1][6] ));
 sg13g2_dfrbp_1 _2434_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net75),
    .D(net321),
    .Q_N(_1142_),
    .Q(\control_tone_freq[1][7] ));
 sg13g2_dfrbp_1 _2435_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net73),
    .D(net335),
    .Q_N(_1141_),
    .Q(\control_tone_freq[1][8] ));
 sg13g2_dfrbp_1 _2436_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net71),
    .D(_0057_),
    .Q_N(_1140_),
    .Q(\control_tone_freq[1][9] ));
 sg13g2_dfrbp_1 _2437_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net69),
    .D(net331),
    .Q_N(_1139_),
    .Q(\control_tone_freq[2][4] ));
 sg13g2_dfrbp_1 _2438_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net67),
    .D(net291),
    .Q_N(_1138_),
    .Q(\control_tone_freq[2][5] ));
 sg13g2_dfrbp_1 _2439_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net65),
    .D(net285),
    .Q_N(_1137_),
    .Q(\control_tone_freq[2][6] ));
 sg13g2_dfrbp_1 _2440_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net63),
    .D(net296),
    .Q_N(_1136_),
    .Q(\control_tone_freq[2][7] ));
 sg13g2_dfrbp_1 _2441_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net61),
    .D(net293),
    .Q_N(_1135_),
    .Q(\control_tone_freq[2][8] ));
 sg13g2_dfrbp_1 _2442_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net59),
    .D(net270),
    .Q_N(_1134_),
    .Q(\control_tone_freq[2][9] ));
 sg13g2_dfrbp_1 _2443_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net57),
    .D(_0064_),
    .Q_N(_1133_),
    .Q(\control_noise[0][0] ));
 sg13g2_dfrbp_1 _2444_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net55),
    .D(_0065_),
    .Q_N(_1132_),
    .Q(\control_noise[0][1] ));
 sg13g2_dfrbp_1 _2445_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net53),
    .D(_0066_),
    .Q_N(_1131_),
    .Q(\control_noise[0][2] ));
 sg13g2_dfrbp_1 _2446_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net51),
    .D(_0067_),
    .Q_N(_1130_),
    .Q(\noise[0].gen.signal_edge.previous_signal_state_0 ));
 sg13g2_dfrbp_1 _2447_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net50),
    .D(net265),
    .Q_N(_0000_),
    .Q(\chan[0].attenuation.in ));
 sg13g2_dfrbp_1 _2448_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net48),
    .D(net307),
    .Q_N(_1129_),
    .Q(\tone[0].gen.counter[0] ));
 sg13g2_dfrbp_1 _2449_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net46),
    .D(_0070_),
    .Q_N(_1128_),
    .Q(\tone[0].gen.counter[1] ));
 sg13g2_dfrbp_1 _2450_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net44),
    .D(net382),
    .Q_N(_1127_),
    .Q(\tone[0].gen.counter[2] ));
 sg13g2_dfrbp_1 _2451_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net42),
    .D(_0072_),
    .Q_N(_1126_),
    .Q(\tone[0].gen.counter[3] ));
 sg13g2_dfrbp_1 _2452_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net40),
    .D(_0073_),
    .Q_N(_1125_),
    .Q(\tone[0].gen.counter[4] ));
 sg13g2_dfrbp_1 _2453_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net38),
    .D(_0074_),
    .Q_N(_1124_),
    .Q(\tone[0].gen.counter[5] ));
 sg13g2_dfrbp_1 _2454_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net36),
    .D(net395),
    .Q_N(_1123_),
    .Q(\tone[0].gen.counter[6] ));
 sg13g2_dfrbp_1 _2455_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net34),
    .D(_0076_),
    .Q_N(_1122_),
    .Q(\tone[0].gen.counter[7] ));
 sg13g2_dfrbp_1 _2456_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net32),
    .D(_0077_),
    .Q_N(_1121_),
    .Q(\tone[0].gen.counter[8] ));
 sg13g2_dfrbp_1 _2457_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net30),
    .D(net387),
    .Q_N(_1120_),
    .Q(\tone[0].gen.counter[9] ));
 sg13g2_dfrbp_1 _2458_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net28),
    .D(net263),
    .Q_N(_0001_),
    .Q(\chan[1].attenuation.in ));
 sg13g2_dfrbp_1 _2459_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net26),
    .D(net337),
    .Q_N(_1119_),
    .Q(\tone[1].gen.counter[0] ));
 sg13g2_dfrbp_1 _2460_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net24),
    .D(_0081_),
    .Q_N(_1118_),
    .Q(\tone[1].gen.counter[1] ));
 sg13g2_dfrbp_1 _2461_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net22),
    .D(net398),
    .Q_N(_1117_),
    .Q(\tone[1].gen.counter[2] ));
 sg13g2_dfrbp_1 _2462_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net20),
    .D(net401),
    .Q_N(_1116_),
    .Q(\tone[1].gen.counter[3] ));
 sg13g2_dfrbp_1 _2463_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net18),
    .D(_0084_),
    .Q_N(_1115_),
    .Q(\tone[1].gen.counter[4] ));
 sg13g2_dfrbp_1 _2464_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net189),
    .D(_0085_),
    .Q_N(_1114_),
    .Q(\tone[1].gen.counter[5] ));
 sg13g2_dfrbp_1 _2465_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net187),
    .D(_0086_),
    .Q_N(_1113_),
    .Q(\tone[1].gen.counter[6] ));
 sg13g2_dfrbp_1 _2466_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net185),
    .D(_0087_),
    .Q_N(_1112_),
    .Q(\tone[1].gen.counter[7] ));
 sg13g2_dfrbp_1 _2467_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net183),
    .D(_0088_),
    .Q_N(_1111_),
    .Q(\tone[1].gen.counter[8] ));
 sg13g2_dfrbp_1 _2468_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net181),
    .D(net390),
    .Q_N(_1110_),
    .Q(\tone[1].gen.counter[9] ));
 sg13g2_dfrbp_1 _2469_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net179),
    .D(net261),
    .Q_N(_0002_),
    .Q(\chan[2].attenuation.in ));
 sg13g2_dfrbp_1 _2470_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net177),
    .D(net346),
    .Q_N(_1109_),
    .Q(\tone[2].gen.counter[0] ));
 sg13g2_dfrbp_1 _2471_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net175),
    .D(net378),
    .Q_N(_1108_),
    .Q(\tone[2].gen.counter[1] ));
 sg13g2_dfrbp_1 _2472_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net173),
    .D(_0093_),
    .Q_N(_1107_),
    .Q(\tone[2].gen.counter[2] ));
 sg13g2_dfrbp_1 _2473_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net171),
    .D(_0094_),
    .Q_N(_1106_),
    .Q(\tone[2].gen.counter[3] ));
 sg13g2_dfrbp_1 _2474_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net169),
    .D(net426),
    .Q_N(_1105_),
    .Q(\tone[2].gen.counter[4] ));
 sg13g2_dfrbp_1 _2475_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net167),
    .D(_0096_),
    .Q_N(_1104_),
    .Q(\tone[2].gen.counter[5] ));
 sg13g2_dfrbp_1 _2476_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net165),
    .D(_0097_),
    .Q_N(_1103_),
    .Q(\tone[2].gen.counter[6] ));
 sg13g2_dfrbp_1 _2477_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net163),
    .D(_0098_),
    .Q_N(_1102_),
    .Q(\tone[2].gen.counter[7] ));
 sg13g2_dfrbp_1 _2478_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net161),
    .D(_0099_),
    .Q_N(_1101_),
    .Q(\tone[2].gen.counter[8] ));
 sg13g2_dfrbp_1 _2479_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net159),
    .D(net404),
    .Q_N(_1100_),
    .Q(\tone[2].gen.counter[9] ));
 sg13g2_dfrbp_1 _2480_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net157),
    .D(_0101_),
    .Q_N(_1099_),
    .Q(\control_tone_freq[0][0] ));
 sg13g2_dfrbp_1 _2481_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net155),
    .D(_0102_),
    .Q_N(_1098_),
    .Q(\control_tone_freq[0][1] ));
 sg13g2_dfrbp_1 _2482_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net153),
    .D(_0103_),
    .Q_N(_1097_),
    .Q(\control_tone_freq[0][2] ));
 sg13g2_dfrbp_1 _2483_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net151),
    .D(_0104_),
    .Q_N(_1096_),
    .Q(\control_tone_freq[0][3] ));
 sg13g2_dfrbp_1 _2484_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net135),
    .D(_0105_),
    .Q_N(_1095_),
    .Q(\genblk4[3].pwm.accumulator[0] ));
 sg13g2_dfrbp_1 _2485_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net133),
    .D(_0106_),
    .Q_N(_1094_),
    .Q(\genblk4[3].pwm.accumulator[1] ));
 sg13g2_dfrbp_1 _2486_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net124),
    .D(net476),
    .Q_N(_1093_),
    .Q(\genblk4[3].pwm.accumulator[2] ));
 sg13g2_dfrbp_1 _2487_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net122),
    .D(_0108_),
    .Q_N(_1092_),
    .Q(\genblk4[3].pwm.accumulator[3] ));
 sg13g2_dfrbp_1 _2488_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net120),
    .D(_0109_),
    .Q_N(_1091_),
    .Q(\genblk4[3].pwm.accumulator[4] ));
 sg13g2_dfrbp_1 _2489_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net118),
    .D(_0110_),
    .Q_N(_1090_),
    .Q(\genblk4[3].pwm.accumulator[5] ));
 sg13g2_dfrbp_1 _2490_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net116),
    .D(net457),
    .Q_N(_1089_),
    .Q(\genblk4[3].pwm.accumulator[6] ));
 sg13g2_dfrbp_1 _2491_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net114),
    .D(net434),
    .Q_N(_1088_),
    .Q(\genblk4[3].pwm.accumulator[7] ));
 sg13g2_dfrbp_1 _2492_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net112),
    .D(_0113_),
    .Q_N(_1087_),
    .Q(\genblk4[3].pwm.accumulator[8] ));
 sg13g2_dfrbp_1 _2493_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net110),
    .D(_0114_),
    .Q_N(_1086_),
    .Q(\genblk4[3].pwm.accumulator[9] ));
 sg13g2_dfrbp_1 _2494_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net108),
    .D(net360),
    .Q_N(_1085_),
    .Q(\genblk4[3].pwm.accumulator[10] ));
 sg13g2_dfrbp_1 _2495_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net106),
    .D(net259),
    .Q_N(_0005_),
    .Q(\noise[0].gen.counter[0] ));
 sg13g2_dfrbp_1 _2496_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net102),
    .D(net275),
    .Q_N(_1084_),
    .Q(\noise[0].gen.counter[1] ));
 sg13g2_dfrbp_1 _2497_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net98),
    .D(net424),
    .Q_N(_1083_),
    .Q(\noise[0].gen.counter[2] ));
 sg13g2_dfrbp_1 _2498_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net94),
    .D(_0119_),
    .Q_N(_1082_),
    .Q(\noise[0].gen.counter[3] ));
 sg13g2_dfrbp_1 _2499_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net90),
    .D(_0120_),
    .Q_N(_0004_),
    .Q(\noise[0].gen.counter[4] ));
 sg13g2_dfrbp_1 _2500_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net86),
    .D(net300),
    .Q_N(_1081_),
    .Q(\noise[0].gen.counter[5] ));
 sg13g2_dfrbp_1 _2501_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net82),
    .D(net333),
    .Q_N(_1080_),
    .Q(\noise[0].gen.counter[6] ));
 sg13g2_dfrbp_1 _2502_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net78),
    .D(_0123_),
    .Q_N(_1079_),
    .Q(\chan[3].attenuation.in ));
 sg13g2_dfrbp_1 _2503_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net74),
    .D(net355),
    .Q_N(_1078_),
    .Q(\noise[0].gen.lfsr[1] ));
 sg13g2_dfrbp_1 _2504_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net70),
    .D(net309),
    .Q_N(_1077_),
    .Q(\noise[0].gen.lfsr[2] ));
 sg13g2_dfrbp_1 _2505_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net66),
    .D(net342),
    .Q_N(_1076_),
    .Q(\noise[0].gen.lfsr[3] ));
 sg13g2_dfrbp_1 _2506_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net62),
    .D(net319),
    .Q_N(_1075_),
    .Q(\noise[0].gen.lfsr[4] ));
 sg13g2_dfrbp_1 _2507_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net58),
    .D(net316),
    .Q_N(_1074_),
    .Q(\noise[0].gen.lfsr[5] ));
 sg13g2_dfrbp_1 _2508_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net54),
    .D(net327),
    .Q_N(_1073_),
    .Q(\noise[0].gen.lfsr[6] ));
 sg13g2_dfrbp_1 _2509_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net49),
    .D(net313),
    .Q_N(_1072_),
    .Q(\noise[0].gen.lfsr[7] ));
 sg13g2_dfrbp_1 _2510_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net45),
    .D(net329),
    .Q_N(_1071_),
    .Q(\noise[0].gen.lfsr[8] ));
 sg13g2_dfrbp_1 _2511_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net41),
    .D(net302),
    .Q_N(_1070_),
    .Q(\noise[0].gen.lfsr[9] ));
 sg13g2_dfrbp_1 _2512_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net37),
    .D(_0133_),
    .Q_N(_1069_),
    .Q(\noise[0].gen.lfsr[10] ));
 sg13g2_dfrbp_1 _2513_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net33),
    .D(net305),
    .Q_N(_1068_),
    .Q(\noise[0].gen.lfsr[11] ));
 sg13g2_dfrbp_1 _2514_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net29),
    .D(net324),
    .Q_N(_1067_),
    .Q(\noise[0].gen.lfsr[12] ));
 sg13g2_dfrbp_1 _2515_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net25),
    .D(net340),
    .Q_N(_1066_),
    .Q(\noise[0].gen.lfsr[13] ));
 sg13g2_dfrbp_1 _2516_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net21),
    .D(net367),
    .Q_N(_1065_),
    .Q(\noise[0].gen.lfsr[14] ));
 sg13g2_dfrbp_1 _2517_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net190),
    .D(_0138_),
    .Q_N(_1064_),
    .Q(\control_tone_freq[1][0] ));
 sg13g2_dfrbp_1 _2518_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net186),
    .D(_0139_),
    .Q_N(_1063_),
    .Q(\control_tone_freq[1][1] ));
 sg13g2_dfrbp_1 _2519_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net182),
    .D(_0140_),
    .Q_N(_1062_),
    .Q(\control_tone_freq[1][2] ));
 sg13g2_dfrbp_1 _2520_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net178),
    .D(_0141_),
    .Q_N(_1061_),
    .Q(\control_tone_freq[1][3] ));
 sg13g2_dfrbp_1 _2521_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net174),
    .D(_0142_),
    .Q_N(_1060_),
    .Q(\control_tone_freq[2][0] ));
 sg13g2_dfrbp_1 _2522_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net170),
    .D(_0143_),
    .Q_N(_1059_),
    .Q(\control_tone_freq[2][1] ));
 sg13g2_dfrbp_1 _2523_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net166),
    .D(_0144_),
    .Q_N(_1058_),
    .Q(\control_tone_freq[2][2] ));
 sg13g2_dfrbp_1 _2524_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net162),
    .D(_0145_),
    .Q_N(_1057_),
    .Q(\control_tone_freq[2][3] ));
 sg13g2_dfrbp_1 _2525_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net158),
    .D(_0146_),
    .Q_N(_1056_),
    .Q(\genblk4[0].pwm.accumulator[0] ));
 sg13g2_dfrbp_1 _2526_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net156),
    .D(_0147_),
    .Q_N(_1055_),
    .Q(\genblk4[0].pwm.accumulator[1] ));
 sg13g2_dfrbp_1 _2527_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net154),
    .D(net447),
    .Q_N(_1054_),
    .Q(\genblk4[0].pwm.accumulator[2] ));
 sg13g2_dfrbp_1 _2528_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net152),
    .D(_0149_),
    .Q_N(_1053_),
    .Q(\genblk4[0].pwm.accumulator[3] ));
 sg13g2_dfrbp_1 _2529_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net137),
    .D(net437),
    .Q_N(_1052_),
    .Q(\genblk4[0].pwm.accumulator[4] ));
 sg13g2_dfrbp_1 _2530_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net104),
    .D(net478),
    .Q_N(_1051_),
    .Q(\genblk4[0].pwm.accumulator[5] ));
 sg13g2_dfrbp_1 _2531_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net100),
    .D(net463),
    .Q_N(_1050_),
    .Q(\genblk4[0].pwm.accumulator[6] ));
 sg13g2_dfrbp_1 _2532_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net96),
    .D(net442),
    .Q_N(_1049_),
    .Q(\genblk4[0].pwm.accumulator[7] ));
 sg13g2_dfrbp_1 _2533_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net92),
    .D(_0154_),
    .Q_N(_1048_),
    .Q(\genblk4[0].pwm.accumulator[8] ));
 sg13g2_dfrbp_1 _2534_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net88),
    .D(_0155_),
    .Q_N(_1047_),
    .Q(\genblk4[0].pwm.accumulator[9] ));
 sg13g2_dfrbp_1 _2535_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net84),
    .D(net374),
    .Q_N(_1046_),
    .Q(\genblk4[0].pwm.accumulator[10] ));
 sg13g2_dfrbp_1 _2536_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net80),
    .D(_0157_),
    .Q_N(_1045_),
    .Q(\genblk4[1].pwm.accumulator[0] ));
 sg13g2_dfrbp_1 _2537_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net76),
    .D(_0158_),
    .Q_N(_1044_),
    .Q(\genblk4[1].pwm.accumulator[1] ));
 sg13g2_dfrbp_1 _2538_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net72),
    .D(_0159_),
    .Q_N(_1043_),
    .Q(\genblk4[1].pwm.accumulator[2] ));
 sg13g2_dfrbp_1 _2539_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net68),
    .D(_0160_),
    .Q_N(_1042_),
    .Q(\genblk4[1].pwm.accumulator[3] ));
 sg13g2_dfrbp_1 _2540_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net64),
    .D(net498),
    .Q_N(_1041_),
    .Q(\genblk4[1].pwm.accumulator[4] ));
 sg13g2_dfrbp_1 _2541_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net60),
    .D(_0162_),
    .Q_N(_1040_),
    .Q(\genblk4[1].pwm.accumulator[5] ));
 sg13g2_dfrbp_1 _2542_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net56),
    .D(_0163_),
    .Q_N(_1039_),
    .Q(\genblk4[1].pwm.accumulator[6] ));
 sg13g2_dfrbp_1 _2543_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net52),
    .D(_0164_),
    .Q_N(_1038_),
    .Q(\genblk4[1].pwm.accumulator[7] ));
 sg13g2_dfrbp_1 _2544_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net47),
    .D(_0165_),
    .Q_N(_1037_),
    .Q(\genblk4[1].pwm.accumulator[8] ));
 sg13g2_dfrbp_1 _2545_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net43),
    .D(_0166_),
    .Q_N(_1036_),
    .Q(\genblk4[1].pwm.accumulator[9] ));
 sg13g2_dfrbp_1 _2546_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net39),
    .D(net365),
    .Q_N(_1035_),
    .Q(\genblk4[1].pwm.accumulator[10] ));
 sg13g2_dfrbp_1 _2547_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net35),
    .D(_0168_),
    .Q_N(_1034_),
    .Q(\genblk4[2].pwm.accumulator[0] ));
 sg13g2_dfrbp_1 _2548_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net31),
    .D(_0169_),
    .Q_N(_1033_),
    .Q(\genblk4[2].pwm.accumulator[1] ));
 sg13g2_dfrbp_1 _2549_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net27),
    .D(_0170_),
    .Q_N(_1032_),
    .Q(\genblk4[2].pwm.accumulator[2] ));
 sg13g2_dfrbp_1 _2550_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net23),
    .D(_0171_),
    .Q_N(_1031_),
    .Q(\genblk4[2].pwm.accumulator[3] ));
 sg13g2_dfrbp_1 _2551_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net19),
    .D(_0172_),
    .Q_N(_1030_),
    .Q(\genblk4[2].pwm.accumulator[4] ));
 sg13g2_dfrbp_1 _2552_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net188),
    .D(net451),
    .Q_N(_1029_),
    .Q(\genblk4[2].pwm.accumulator[5] ));
 sg13g2_dfrbp_1 _2553_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net184),
    .D(_0174_),
    .Q_N(_1028_),
    .Q(\genblk4[2].pwm.accumulator[6] ));
 sg13g2_dfrbp_1 _2554_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net180),
    .D(net432),
    .Q_N(_1027_),
    .Q(\genblk4[2].pwm.accumulator[7] ));
 sg13g2_dfrbp_1 _2555_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net176),
    .D(_0176_),
    .Q_N(_1026_),
    .Q(\genblk4[2].pwm.accumulator[8] ));
 sg13g2_dfrbp_1 _2556_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net172),
    .D(_0177_),
    .Q_N(_1025_),
    .Q(\genblk4[2].pwm.accumulator[9] ));
 sg13g2_dfrbp_1 _2557_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net168),
    .D(net358),
    .Q_N(_1024_),
    .Q(\genblk4[2].pwm.accumulator[10] ));
 sg13g2_dfrbp_1 _2558_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net164),
    .D(_0179_),
    .Q_N(_1023_),
    .Q(\noise[0].gen.restart_noise ));
 sg13g2_tiehi _2551__19 (.L_HI(net19));
 sg13g2_tiehi _2462__20 (.L_HI(net20));
 sg13g2_tiehi _2516__21 (.L_HI(net21));
 sg13g2_tiehi _2461__22 (.L_HI(net22));
 sg13g2_tiehi _2550__23 (.L_HI(net23));
 sg13g2_tiehi _2460__24 (.L_HI(net24));
 sg13g2_tiehi _2515__25 (.L_HI(net25));
 sg13g2_tiehi _2459__26 (.L_HI(net26));
 sg13g2_tiehi _2549__27 (.L_HI(net27));
 sg13g2_tiehi _2458__28 (.L_HI(net28));
 sg13g2_tiehi _2514__29 (.L_HI(net29));
 sg13g2_tiehi _2457__30 (.L_HI(net30));
 sg13g2_tiehi _2548__31 (.L_HI(net31));
 sg13g2_tiehi _2456__32 (.L_HI(net32));
 sg13g2_tiehi _2513__33 (.L_HI(net33));
 sg13g2_tiehi _2455__34 (.L_HI(net34));
 sg13g2_tiehi _2547__35 (.L_HI(net35));
 sg13g2_tiehi _2454__36 (.L_HI(net36));
 sg13g2_tiehi _2512__37 (.L_HI(net37));
 sg13g2_tiehi _2453__38 (.L_HI(net38));
 sg13g2_tiehi _2546__39 (.L_HI(net39));
 sg13g2_tiehi _2452__40 (.L_HI(net40));
 sg13g2_tiehi _2511__41 (.L_HI(net41));
 sg13g2_tiehi _2451__42 (.L_HI(net42));
 sg13g2_tiehi _2545__43 (.L_HI(net43));
 sg13g2_tiehi _2450__44 (.L_HI(net44));
 sg13g2_tiehi _2510__45 (.L_HI(net45));
 sg13g2_tiehi _2449__46 (.L_HI(net46));
 sg13g2_tiehi _2544__47 (.L_HI(net47));
 sg13g2_tiehi _2448__48 (.L_HI(net48));
 sg13g2_tiehi _2509__49 (.L_HI(net49));
 sg13g2_tiehi _2447__50 (.L_HI(net50));
 sg13g2_tiehi _2446__51 (.L_HI(net51));
 sg13g2_tiehi _2543__52 (.L_HI(net52));
 sg13g2_tiehi _2445__53 (.L_HI(net53));
 sg13g2_tiehi _2508__54 (.L_HI(net54));
 sg13g2_tiehi _2444__55 (.L_HI(net55));
 sg13g2_tiehi _2542__56 (.L_HI(net56));
 sg13g2_tiehi _2443__57 (.L_HI(net57));
 sg13g2_tiehi _2507__58 (.L_HI(net58));
 sg13g2_tiehi _2442__59 (.L_HI(net59));
 sg13g2_tiehi _2541__60 (.L_HI(net60));
 sg13g2_tiehi _2441__61 (.L_HI(net61));
 sg13g2_tiehi _2506__62 (.L_HI(net62));
 sg13g2_tiehi _2440__63 (.L_HI(net63));
 sg13g2_tiehi _2540__64 (.L_HI(net64));
 sg13g2_tiehi _2439__65 (.L_HI(net65));
 sg13g2_tiehi _2505__66 (.L_HI(net66));
 sg13g2_tiehi _2438__67 (.L_HI(net67));
 sg13g2_tiehi _2539__68 (.L_HI(net68));
 sg13g2_tiehi _2437__69 (.L_HI(net69));
 sg13g2_tiehi _2504__70 (.L_HI(net70));
 sg13g2_tiehi _2436__71 (.L_HI(net71));
 sg13g2_tiehi _2538__72 (.L_HI(net72));
 sg13g2_tiehi _2435__73 (.L_HI(net73));
 sg13g2_tiehi _2503__74 (.L_HI(net74));
 sg13g2_tiehi _2434__75 (.L_HI(net75));
 sg13g2_tiehi _2537__76 (.L_HI(net76));
 sg13g2_tiehi _2433__77 (.L_HI(net77));
 sg13g2_tiehi _2502__78 (.L_HI(net78));
 sg13g2_tiehi _2432__79 (.L_HI(net79));
 sg13g2_tiehi _2536__80 (.L_HI(net80));
 sg13g2_tiehi _2431__81 (.L_HI(net81));
 sg13g2_tiehi _2501__82 (.L_HI(net82));
 sg13g2_tiehi _2430__83 (.L_HI(net83));
 sg13g2_tiehi _2535__84 (.L_HI(net84));
 sg13g2_tiehi _2429__85 (.L_HI(net85));
 sg13g2_tiehi _2500__86 (.L_HI(net86));
 sg13g2_tiehi _2428__87 (.L_HI(net87));
 sg13g2_tiehi _2534__88 (.L_HI(net88));
 sg13g2_tiehi _2427__89 (.L_HI(net89));
 sg13g2_tiehi _2499__90 (.L_HI(net90));
 sg13g2_tiehi _2426__91 (.L_HI(net91));
 sg13g2_tiehi _2533__92 (.L_HI(net92));
 sg13g2_tiehi _2425__93 (.L_HI(net93));
 sg13g2_tiehi _2498__94 (.L_HI(net94));
 sg13g2_tiehi _2424__95 (.L_HI(net95));
 sg13g2_tiehi _2532__96 (.L_HI(net96));
 sg13g2_tiehi _2423__97 (.L_HI(net97));
 sg13g2_tiehi _2497__98 (.L_HI(net98));
 sg13g2_tiehi _2422__99 (.L_HI(net99));
 sg13g2_tiehi _2531__100 (.L_HI(net100));
 sg13g2_tiehi _2421__101 (.L_HI(net101));
 sg13g2_tiehi _2496__102 (.L_HI(net102));
 sg13g2_tiehi _2420__103 (.L_HI(net103));
 sg13g2_tiehi _2530__104 (.L_HI(net104));
 sg13g2_tiehi _2419__105 (.L_HI(net105));
 sg13g2_tiehi _2495__106 (.L_HI(net106));
 sg13g2_tiehi _2418__107 (.L_HI(net107));
 sg13g2_tiehi _2494__108 (.L_HI(net108));
 sg13g2_tiehi _2417__109 (.L_HI(net109));
 sg13g2_tiehi _2493__110 (.L_HI(net110));
 sg13g2_tiehi _2416__111 (.L_HI(net111));
 sg13g2_tiehi _2492__112 (.L_HI(net112));
 sg13g2_tiehi _2415__113 (.L_HI(net113));
 sg13g2_tiehi _2491__114 (.L_HI(net114));
 sg13g2_tiehi _2414__115 (.L_HI(net115));
 sg13g2_tiehi _2490__116 (.L_HI(net116));
 sg13g2_tiehi _2413__117 (.L_HI(net117));
 sg13g2_tiehi _2489__118 (.L_HI(net118));
 sg13g2_tiehi _2412__119 (.L_HI(net119));
 sg13g2_tiehi _2488__120 (.L_HI(net120));
 sg13g2_tiehi _2411__121 (.L_HI(net121));
 sg13g2_tiehi _2487__122 (.L_HI(net122));
 sg13g2_tiehi _2410__123 (.L_HI(net123));
 sg13g2_tiehi _2486__124 (.L_HI(net124));
 sg13g2_tiehi _2409__125 (.L_HI(net125));
 sg13g2_tiehi _2408__126 (.L_HI(net126));
 sg13g2_tiehi _2407__127 (.L_HI(net127));
 sg13g2_tiehi _2406__128 (.L_HI(net128));
 sg13g2_tiehi _2405__129 (.L_HI(net129));
 sg13g2_tiehi _2404__130 (.L_HI(net130));
 sg13g2_tiehi _2403__131 (.L_HI(net131));
 sg13g2_tiehi _2402__132 (.L_HI(net132));
 sg13g2_tiehi _2485__133 (.L_HI(net133));
 sg13g2_tiehi _2401__134 (.L_HI(net134));
 sg13g2_tiehi _2484__135 (.L_HI(net135));
 sg13g2_tiehi _2400__136 (.L_HI(net136));
 sg13g2_tiehi _2529__137 (.L_HI(net137));
 sg13g2_tiehi _2399__138 (.L_HI(net138));
 sg13g2_tiehi _2398__139 (.L_HI(net139));
 sg13g2_tiehi _2397__140 (.L_HI(net140));
 sg13g2_tiehi _2396__141 (.L_HI(net141));
 sg13g2_tiehi _2395__142 (.L_HI(net142));
 sg13g2_tiehi _2394__143 (.L_HI(net143));
 sg13g2_tiehi _2393__144 (.L_HI(net144));
 sg13g2_tiehi _2392__145 (.L_HI(net145));
 sg13g2_tiehi _2391__146 (.L_HI(net146));
 sg13g2_tiehi _2390__147 (.L_HI(net147));
 sg13g2_tiehi _2389__148 (.L_HI(net148));
 sg13g2_tiehi _2388__149 (.L_HI(net149));
 sg13g2_tiehi _2387__150 (.L_HI(net150));
 sg13g2_tiehi _2483__151 (.L_HI(net151));
 sg13g2_tiehi _2528__152 (.L_HI(net152));
 sg13g2_tiehi _2482__153 (.L_HI(net153));
 sg13g2_tiehi _2527__154 (.L_HI(net154));
 sg13g2_tiehi _2481__155 (.L_HI(net155));
 sg13g2_tiehi _2526__156 (.L_HI(net156));
 sg13g2_tiehi _2480__157 (.L_HI(net157));
 sg13g2_tiehi _2525__158 (.L_HI(net158));
 sg13g2_tiehi _2479__159 (.L_HI(net159));
 sg13g2_tiehi _2386__160 (.L_HI(net160));
 sg13g2_tiehi _2478__161 (.L_HI(net161));
 sg13g2_tiehi _2524__162 (.L_HI(net162));
 sg13g2_tiehi _2477__163 (.L_HI(net163));
 sg13g2_tiehi _2558__164 (.L_HI(net164));
 sg13g2_tiehi _2476__165 (.L_HI(net165));
 sg13g2_tiehi _2523__166 (.L_HI(net166));
 sg13g2_tiehi _2475__167 (.L_HI(net167));
 sg13g2_tiehi _2557__168 (.L_HI(net168));
 sg13g2_tiehi _2474__169 (.L_HI(net169));
 sg13g2_tiehi _2522__170 (.L_HI(net170));
 sg13g2_tiehi _2473__171 (.L_HI(net171));
 sg13g2_tiehi _2556__172 (.L_HI(net172));
 sg13g2_tiehi _2472__173 (.L_HI(net173));
 sg13g2_tiehi _2521__174 (.L_HI(net174));
 sg13g2_tiehi _2471__175 (.L_HI(net175));
 sg13g2_tiehi _2555__176 (.L_HI(net176));
 sg13g2_tiehi _2470__177 (.L_HI(net177));
 sg13g2_tiehi _2520__178 (.L_HI(net178));
 sg13g2_tiehi _2469__179 (.L_HI(net179));
 sg13g2_tiehi _2554__180 (.L_HI(net180));
 sg13g2_tiehi _2468__181 (.L_HI(net181));
 sg13g2_tiehi _2519__182 (.L_HI(net182));
 sg13g2_tiehi _2467__183 (.L_HI(net183));
 sg13g2_tiehi _2553__184 (.L_HI(net184));
 sg13g2_tiehi _2466__185 (.L_HI(net185));
 sg13g2_tiehi _2518__186 (.L_HI(net186));
 sg13g2_tiehi _2465__187 (.L_HI(net187));
 sg13g2_tiehi _2552__188 (.L_HI(net188));
 sg13g2_tiehi _2464__189 (.L_HI(net189));
 sg13g2_tiehi _2517__190 (.L_HI(net190));
 sg13g2_tiehi tt_um_rejunity_sn76489_191 (.L_HI(net252));
 sg13g2_tiehi tt_um_rejunity_sn76489_192 (.L_HI(net253));
 sg13g2_tiehi tt_um_rejunity_sn76489_193 (.L_HI(net254));
 sg13g2_tiehi tt_um_rejunity_sn76489_194 (.L_HI(net255));
 sg13g2_tiehi tt_um_rejunity_sn76489_195 (.L_HI(net256));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_rejunity_sn76489_13 (.L_LO(net13));
 sg13g2_tielo tt_um_rejunity_sn76489_14 (.L_LO(net14));
 sg13g2_tielo tt_um_rejunity_sn76489_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rejunity_sn76489_16 (.L_LO(net16));
 sg13g2_tielo tt_um_rejunity_sn76489_17 (.L_LO(net17));
 sg13g2_tiehi _2463__18 (.L_HI(net18));
 sg13g2_buf_1 _2743_ (.A(\genblk4[0].pwm.accumulator[10] ),
    .X(uio_out[3]));
 sg13g2_buf_1 _2744_ (.A(\genblk4[1].pwm.accumulator[10] ),
    .X(uio_out[4]));
 sg13g2_buf_1 _2745_ (.A(\genblk4[2].pwm.accumulator[10] ),
    .X(uio_out[5]));
 sg13g2_buf_1 _2746_ (.A(\genblk4[3].pwm.accumulator[10] ),
    .X(uio_out[6]));
 sg13g2_buf_1 _2747_ (.A(\pwm.accumulator[12] ),
    .X(uio_out[7]));
 sg13g2_buf_2 fanout191 (.A(net192),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_0314_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_0313_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_0313_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_0206_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_0998_),
    .X(net196));
 sg13g2_buf_4 fanout197 (.X(net197),
    .A(_0947_));
 sg13g2_buf_1 fanout198 (.A(_0947_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(net201),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(net202),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(net206),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(net204),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(net206),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(net206),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_0946_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_0941_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_0925_),
    .X(net208));
 sg13g2_buf_1 fanout209 (.A(_0925_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_0918_),
    .X(net210));
 sg13g2_buf_1 fanout211 (.A(_0918_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_0911_),
    .X(net212));
 sg13g2_buf_1 fanout213 (.A(_0911_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_0316_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_0316_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_0545_),
    .X(net216));
 sg13g2_buf_4 fanout217 (.X(net217),
    .A(net371));
 sg13g2_buf_2 fanout218 (.A(net219),
    .X(net218));
 sg13g2_buf_4 fanout219 (.X(net219),
    .A(\chan[2].attenuation.in ));
 sg13g2_buf_2 fanout220 (.A(\chan[1].attenuation.in ),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(\chan[0].attenuation.in ),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(\chan[2].attenuation.control[2] ),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(\chan[0].attenuation.control[0] ),
    .X(net223));
 sg13g2_buf_4 fanout224 (.X(net224),
    .A(net230));
 sg13g2_buf_2 fanout225 (.A(net227),
    .X(net225));
 sg13g2_buf_1 fanout226 (.A(net227),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(net229),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(net229),
    .X(net228));
 sg13g2_buf_1 fanout229 (.A(net230),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_0527_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(net232),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(net233),
    .X(net232));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(net251));
 sg13g2_buf_2 fanout234 (.A(net235),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(net236),
    .X(net235));
 sg13g2_buf_4 fanout236 (.X(net236),
    .A(net251));
 sg13g2_buf_4 fanout237 (.X(net237),
    .A(net243));
 sg13g2_buf_2 fanout238 (.A(net242),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(net242),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net242),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(net242),
    .X(net241));
 sg13g2_buf_1 fanout242 (.A(net243),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(net251),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(net245),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(net250),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(net247),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(net250),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(net249),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(net250),
    .X(net249));
 sg13g2_buf_1 fanout250 (.A(net251),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(rst_n),
    .X(net251));
 sg13g2_buf_4 input1 (.X(net1),
    .A(ui_in[0]));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[1]));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[2]));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[3]));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[4]));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[5]));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_tielo tt_um_rejunity_sn76489_12 (.L_LO(net12));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_29__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0006_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0005_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0116_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0002_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0090_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0001_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0079_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0000_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0068_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold10 (.A(\control_tone_freq[0][8] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold11 (.A(\genblk4[1].pwm.accumulator[0] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold12 (.A(\control_tone_freq[2][1] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold13 (.A(\control_tone_freq[2][9] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0063_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold15 (.A(\control_tone_freq[2][2] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold16 (.A(\control_tone_freq[0][5] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold17 (.A(\noise[0].gen.counter[1] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0301_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0117_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold20 (.A(\control_tone_freq[1][6] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold21 (.A(\control_tone_freq[0][7] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold22 (.A(\genblk4[3].pwm.accumulator[0] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold23 (.A(\control_tone_freq[1][4] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0052_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold25 (.A(\control_tone_freq[1][5] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0053_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold27 (.A(\control_tone_freq[0][4] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold28 (.A(\control_tone_freq[2][6] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0060_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold30 (.A(\control_tone_freq[0][6] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold31 (.A(\clk_counter[2] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0873_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0025_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold34 (.A(\control_tone_freq[2][5] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0059_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold36 (.A(\control_tone_freq[2][8] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0062_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold38 (.A(\control_tone_freq[1][9] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold39 (.A(\control_tone_freq[2][7] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0061_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold41 (.A(\control_tone_freq[2][3] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold42 (.A(\control_tone_freq[0][9] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold43 (.A(\noise[0].gen.counter[5] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0121_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold45 (.A(\noise[0].gen.lfsr[10] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0132_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold47 (.A(\noise[0].gen.lfsr[11] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0339_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0134_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold50 (.A(\tone[0].gen.counter[0] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0069_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold52 (.A(\noise[0].gen.lfsr[3] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0125_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold54 (.A(\control_noise[0][1] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold55 (.A(\noise[0].gen.lfsr[7] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0331_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0130_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold58 (.A(\noise[0].gen.lfsr[5] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0327_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0128_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold61 (.A(\noise[0].gen.lfsr[4] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0325_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0127_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold64 (.A(\control_tone_freq[1][7] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0055_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold66 (.A(\noise[0].gen.lfsr[12] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0341_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0135_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold69 (.A(\noise[0].gen.lfsr[6] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0329_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0129_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold72 (.A(\noise[0].gen.lfsr[9] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0131_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold74 (.A(\control_tone_freq[2][4] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0058_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold76 (.A(\noise[0].gen.counter[6] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0122_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold78 (.A(\control_tone_freq[1][8] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0056_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold80 (.A(\tone[1].gen.counter[0] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0080_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold82 (.A(\noise[0].gen.lfsr[13] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0343_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0136_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold85 (.A(\noise[0].gen.restart_noise ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0126_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold87 (.A(\control_tone_freq[0][0] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold88 (.A(\control_tone_freq[1][0] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold89 (.A(\tone[2].gen.counter[0] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0091_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold91 (.A(\pwm.accumulator[11] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0019_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold93 (.A(\noise[0].gen.signal_edge.previous_signal_state_0 ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold94 (.A(\clk_counter[1] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0024_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold96 (.A(\clk_counter[6] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0029_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold98 (.A(\noise[0].gen.lfsr[1] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0124_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold100 (.A(\genblk4[2].pwm.accumulator[9] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0473_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0178_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold103 (.A(\genblk4[3].pwm.accumulator[9] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0115_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold105 (.A(\latch_control_reg[2] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold106 (.A(\control_noise[0][0] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold107 (.A(\control_tone_freq[0][2] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold108 (.A(\genblk4[1].pwm.accumulator[9] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0167_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold110 (.A(\noise[0].gen.lfsr[14] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0137_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold112 (.A(\genblk4[2].pwm.accumulator[0] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold113 (.A(\noise[0].gen.counter[4] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0308_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold115 (.A(\chan[3].attenuation.in ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold116 (.A(\control_tone_freq[0][3] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold117 (.A(\genblk4[0].pwm.accumulator[9] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0156_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold119 (.A(\control_tone_freq[0][1] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold120 (.A(\control_noise[0][2] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold121 (.A(\tone[2].gen.counter[1] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0092_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold123 (.A(\genblk4[2].pwm.accumulator[1] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold124 (.A(\tone[2].gen.counter[2] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold125 (.A(\tone[0].gen.counter[2] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0071_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold127 (.A(\control_tone_freq[1][2] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold128 (.A(\tone[0].gen.counter[7] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold129 (.A(\tone[1].gen.counter[5] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold130 (.A(\tone[0].gen.counter[9] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0078_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold132 (.A(\tone[1].gen.counter[6] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold133 (.A(\tone[1].gen.counter[9] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0089_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold135 (.A(\control_tone_freq[1][1] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold136 (.A(\tone[0].gen.counter[4] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold137 (.A(\genblk4[0].pwm.accumulator[0] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold138 (.A(\tone[0].gen.counter[6] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0075_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold140 (.A(\control_tone_freq[2][0] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold141 (.A(\tone[1].gen.counter[2] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0082_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold143 (.A(\tone[0].gen.counter[1] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold144 (.A(\tone[1].gen.counter[3] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0083_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold146 (.A(\tone[0].gen.counter[5] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold147 (.A(\tone[2].gen.counter[9] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0100_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold149 (.A(\clk_counter[4] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0879_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold151 (.A(\tone[2].gen.counter[7] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold152 (.A(\tone[1].gen.counter[8] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold153 (.A(\tone[2].gen.counter[8] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold154 (.A(\control_tone_freq[1][3] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold155 (.A(\tone[0].gen.counter[8] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold156 (.A(\tone[2].gen.counter[3] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold157 (.A(\tone[1].gen.counter[1] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold158 (.A(\tone[0].gen.counter[3] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold159 (.A(\pwm.accumulator[0] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0008_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold161 (.A(\tone[1].gen.counter[4] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold162 (.A(\tone[1].gen.counter[7] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold163 (.A(\chan[0].attenuation.control[0] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold164 (.A(\tone[2].gen.counter[6] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold165 (.A(\tone[2].gen.counter[5] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold166 (.A(\noise[0].gen.counter[2] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0304_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0118_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold169 (.A(\tone[2].gen.counter[4] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0095_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold171 (.A(\latch_control_reg[0] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold172 (.A(\chan[2].attenuation.control[2] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold173 (.A(\latch_control_reg[1] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold174 (.A(\chan[1].attenuation.control[1] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold175 (.A(\genblk4[2].pwm.accumulator[6] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0175_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold177 (.A(\genblk4[3].pwm.accumulator[7] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0112_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold179 (.A(\genblk4[1].pwm.accumulator[8] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold180 (.A(\genblk4[0].pwm.accumulator[3] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0150_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold182 (.A(\chan[3].attenuation.control[3] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold183 (.A(\chan[0].attenuation.control[3] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold184 (.A(\genblk4[3].pwm.accumulator[8] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold185 (.A(\genblk4[0].pwm.accumulator[7] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0153_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold187 (.A(\clk_counter[3] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0876_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold189 (.A(\genblk4[0].pwm.accumulator[8] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold190 (.A(\genblk4[0].pwm.accumulator[1] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0148_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold192 (.A(\genblk4[2].pwm.accumulator[8] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold193 (.A(\chan[3].attenuation.control[1] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold194 (.A(\genblk4[2].pwm.accumulator[5] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0173_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold196 (.A(\pwm.accumulator[9] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0016_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold198 (.A(\chan[2].attenuation.control[3] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold199 (.A(\clk_counter[5] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold200 (.A(\genblk4[3].pwm.accumulator[6] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0111_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold202 (.A(\pwm.accumulator[7] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0014_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold204 (.A(\chan[1].attenuation.control[0] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold205 (.A(\noise[0].gen.counter[3] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold206 (.A(\genblk4[0].pwm.accumulator[6] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0152_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold208 (.A(\genblk4[1].pwm.accumulator[1] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold209 (.A(\pwm.accumulator[5] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0012_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold211 (.A(\pwm.accumulator[10] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0017_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold213 (.A(\pwm.accumulator[3] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0010_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold215 (.A(\chan[2].attenuation.control[1] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold216 (.A(\chan[3].attenuation.control[0] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold217 (.A(\chan[3].attenuation.control[2] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold218 (.A(\chan[1].attenuation.control[2] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold219 (.A(\genblk4[3].pwm.accumulator[2] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0107_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold221 (.A(\genblk4[0].pwm.accumulator[5] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0151_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold223 (.A(\chan[0].attenuation.control[1] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold224 (.A(\chan[0].attenuation.control[2] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold225 (.A(\chan[1].attenuation.control[3] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold226 (.A(\pwm.accumulator[1] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0009_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold228 (.A(\genblk4[1].pwm.accumulator[5] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0421_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold230 (.A(\genblk4[3].pwm.accumulator[5] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0281_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold232 (.A(\genblk4[1].pwm.accumulator[2] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0410_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold234 (.A(\genblk4[2].pwm.accumulator[2] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold235 (.A(\genblk4[2].pwm.accumulator[3] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold236 (.A(\chan[2].attenuation.control[0] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold237 (.A(\genblk4[3].pwm.accumulator[1] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold238 (.A(\genblk4[3].pwm.accumulator[3] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold239 (.A(\genblk4[2].pwm.accumulator[7] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold240 (.A(\genblk4[1].pwm.accumulator[3] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0415_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0161_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold243 (.A(\pwm.accumulator[8] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold244 (.A(\noise[0].gen.counter[5] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold245 (.A(\genblk4[3].pwm.accumulator[4] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold246 (.A(\genblk4[2].pwm.accumulator[1] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold247 (.A(\pwm.accumulator[4] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold248 (.A(\genblk4[0].pwm.accumulator[2] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold249 (.A(\genblk4[1].pwm.accumulator[6] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0425_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold251 (.A(\genblk4[1].pwm.accumulator[7] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold252 (.A(\latch_control_reg[1] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold253 (.A(\tone[2].gen.counter[5] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0206_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold255 (.A(\pwm.accumulator[5] ),
    .X(net511));
 sg13g2_antennanp ANTENNA_1 (.A(_0094_));
 sg13g2_antennanp ANTENNA_2 (.A(_0095_));
 sg13g2_antennanp ANTENNA_3 (.A(_0095_));
 sg13g2_antennanp ANTENNA_4 (.A(_0095_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_fill_2 FILLER_0_49 ();
 sg13g2_fill_1 FILLER_0_51 ();
 sg13g2_fill_1 FILLER_0_94 ();
 sg13g2_fill_2 FILLER_0_142 ();
 sg13g2_fill_2 FILLER_0_181 ();
 sg13g2_fill_1 FILLER_0_238 ();
 sg13g2_fill_2 FILLER_0_243 ();
 sg13g2_fill_1 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_fill_2 FILLER_1_87 ();
 sg13g2_fill_1 FILLER_1_186 ();
 sg13g2_fill_1 FILLER_1_192 ();
 sg13g2_fill_1 FILLER_1_202 ();
 sg13g2_decap_4 FILLER_1_229 ();
 sg13g2_fill_2 FILLER_1_264 ();
 sg13g2_fill_1 FILLER_1_266 ();
 sg13g2_fill_1 FILLER_1_294 ();
 sg13g2_fill_2 FILLER_1_304 ();
 sg13g2_decap_8 FILLER_1_332 ();
 sg13g2_decap_8 FILLER_1_339 ();
 sg13g2_decap_8 FILLER_1_346 ();
 sg13g2_decap_8 FILLER_1_353 ();
 sg13g2_decap_8 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_fill_2 FILLER_2_49 ();
 sg13g2_fill_2 FILLER_2_131 ();
 sg13g2_fill_1 FILLER_2_133 ();
 sg13g2_fill_2 FILLER_2_165 ();
 sg13g2_fill_2 FILLER_2_181 ();
 sg13g2_fill_1 FILLER_2_218 ();
 sg13g2_fill_1 FILLER_2_293 ();
 sg13g2_fill_1 FILLER_2_306 ();
 sg13g2_fill_2 FILLER_2_334 ();
 sg13g2_fill_1 FILLER_2_341 ();
 sg13g2_fill_2 FILLER_2_350 ();
 sg13g2_decap_4 FILLER_2_364 ();
 sg13g2_fill_1 FILLER_2_368 ();
 sg13g2_fill_1 FILLER_2_373 ();
 sg13g2_decap_4 FILLER_2_383 ();
 sg13g2_fill_1 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_fill_2 FILLER_3_49 ();
 sg13g2_fill_2 FILLER_3_85 ();
 sg13g2_fill_1 FILLER_3_87 ();
 sg13g2_fill_2 FILLER_3_147 ();
 sg13g2_fill_1 FILLER_3_149 ();
 sg13g2_fill_1 FILLER_3_176 ();
 sg13g2_fill_2 FILLER_3_186 ();
 sg13g2_fill_1 FILLER_3_197 ();
 sg13g2_fill_1 FILLER_3_212 ();
 sg13g2_fill_2 FILLER_3_227 ();
 sg13g2_fill_1 FILLER_3_270 ();
 sg13g2_fill_2 FILLER_3_288 ();
 sg13g2_fill_1 FILLER_3_290 ();
 sg13g2_fill_1 FILLER_3_308 ();
 sg13g2_fill_1 FILLER_3_335 ();
 sg13g2_fill_1 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_402 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_fill_2 FILLER_4_56 ();
 sg13g2_fill_1 FILLER_4_58 ();
 sg13g2_fill_2 FILLER_4_85 ();
 sg13g2_fill_1 FILLER_4_110 ();
 sg13g2_fill_2 FILLER_4_138 ();
 sg13g2_fill_1 FILLER_4_140 ();
 sg13g2_fill_1 FILLER_4_177 ();
 sg13g2_fill_2 FILLER_4_187 ();
 sg13g2_fill_2 FILLER_4_257 ();
 sg13g2_fill_1 FILLER_4_329 ();
 sg13g2_fill_2 FILLER_4_371 ();
 sg13g2_fill_1 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_fill_2 FILLER_5_63 ();
 sg13g2_fill_1 FILLER_5_142 ();
 sg13g2_decap_4 FILLER_5_209 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_fill_2 FILLER_5_289 ();
 sg13g2_fill_1 FILLER_5_291 ();
 sg13g2_fill_1 FILLER_5_303 ();
 sg13g2_fill_1 FILLER_5_355 ();
 sg13g2_fill_2 FILLER_5_376 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_4 FILLER_6_70 ();
 sg13g2_fill_1 FILLER_6_78 ();
 sg13g2_fill_2 FILLER_6_109 ();
 sg13g2_fill_1 FILLER_6_162 ();
 sg13g2_fill_1 FILLER_6_182 ();
 sg13g2_fill_1 FILLER_6_188 ();
 sg13g2_fill_2 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_229 ();
 sg13g2_fill_2 FILLER_6_236 ();
 sg13g2_fill_2 FILLER_6_270 ();
 sg13g2_fill_2 FILLER_6_298 ();
 sg13g2_fill_2 FILLER_6_332 ();
 sg13g2_fill_2 FILLER_6_349 ();
 sg13g2_fill_1 FILLER_6_351 ();
 sg13g2_fill_1 FILLER_6_362 ();
 sg13g2_fill_2 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_fill_1 FILLER_7_58 ();
 sg13g2_fill_1 FILLER_7_72 ();
 sg13g2_fill_2 FILLER_7_100 ();
 sg13g2_fill_1 FILLER_7_145 ();
 sg13g2_fill_1 FILLER_7_185 ();
 sg13g2_fill_2 FILLER_7_212 ();
 sg13g2_decap_4 FILLER_7_280 ();
 sg13g2_fill_2 FILLER_7_324 ();
 sg13g2_fill_1 FILLER_7_398 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_fill_1 FILLER_8_49 ();
 sg13g2_fill_1 FILLER_8_105 ();
 sg13g2_fill_1 FILLER_8_171 ();
 sg13g2_fill_1 FILLER_8_203 ();
 sg13g2_decap_4 FILLER_8_240 ();
 sg13g2_fill_1 FILLER_8_244 ();
 sg13g2_fill_2 FILLER_8_249 ();
 sg13g2_decap_4 FILLER_8_261 ();
 sg13g2_fill_1 FILLER_8_301 ();
 sg13g2_fill_1 FILLER_8_311 ();
 sg13g2_fill_1 FILLER_8_316 ();
 sg13g2_decap_4 FILLER_8_352 ();
 sg13g2_fill_1 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_4 FILLER_9_28 ();
 sg13g2_fill_1 FILLER_9_32 ();
 sg13g2_fill_2 FILLER_9_59 ();
 sg13g2_fill_2 FILLER_9_74 ();
 sg13g2_fill_2 FILLER_9_93 ();
 sg13g2_fill_1 FILLER_9_95 ();
 sg13g2_decap_4 FILLER_9_117 ();
 sg13g2_fill_1 FILLER_9_121 ();
 sg13g2_fill_2 FILLER_9_144 ();
 sg13g2_fill_2 FILLER_9_155 ();
 sg13g2_fill_1 FILLER_9_164 ();
 sg13g2_fill_1 FILLER_9_172 ();
 sg13g2_decap_4 FILLER_9_183 ();
 sg13g2_decap_4 FILLER_9_191 ();
 sg13g2_fill_2 FILLER_9_229 ();
 sg13g2_fill_1 FILLER_9_241 ();
 sg13g2_fill_1 FILLER_9_271 ();
 sg13g2_fill_1 FILLER_9_275 ();
 sg13g2_fill_2 FILLER_9_299 ();
 sg13g2_fill_2 FILLER_9_327 ();
 sg13g2_fill_1 FILLER_9_329 ();
 sg13g2_fill_2 FILLER_9_392 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_25 ();
 sg13g2_fill_1 FILLER_10_32 ();
 sg13g2_fill_2 FILLER_10_45 ();
 sg13g2_fill_2 FILLER_10_84 ();
 sg13g2_fill_2 FILLER_10_91 ();
 sg13g2_fill_1 FILLER_10_93 ();
 sg13g2_fill_2 FILLER_10_128 ();
 sg13g2_fill_2 FILLER_10_156 ();
 sg13g2_decap_4 FILLER_10_176 ();
 sg13g2_fill_1 FILLER_10_180 ();
 sg13g2_fill_2 FILLER_10_207 ();
 sg13g2_fill_2 FILLER_10_223 ();
 sg13g2_fill_1 FILLER_10_251 ();
 sg13g2_decap_4 FILLER_10_275 ();
 sg13g2_fill_2 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_9 ();
 sg13g2_fill_2 FILLER_11_58 ();
 sg13g2_fill_1 FILLER_11_97 ();
 sg13g2_fill_1 FILLER_11_125 ();
 sg13g2_fill_2 FILLER_11_152 ();
 sg13g2_fill_1 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_178 ();
 sg13g2_decap_8 FILLER_11_185 ();
 sg13g2_fill_2 FILLER_11_210 ();
 sg13g2_fill_1 FILLER_11_212 ();
 sg13g2_fill_1 FILLER_11_231 ();
 sg13g2_fill_1 FILLER_11_258 ();
 sg13g2_fill_2 FILLER_11_288 ();
 sg13g2_fill_2 FILLER_11_313 ();
 sg13g2_fill_1 FILLER_11_315 ();
 sg13g2_fill_1 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_18 ();
 sg13g2_fill_1 FILLER_12_81 ();
 sg13g2_decap_4 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_122 ();
 sg13g2_fill_2 FILLER_12_129 ();
 sg13g2_fill_2 FILLER_12_139 ();
 sg13g2_fill_2 FILLER_12_145 ();
 sg13g2_fill_2 FILLER_12_155 ();
 sg13g2_fill_1 FILLER_12_157 ();
 sg13g2_fill_1 FILLER_12_175 ();
 sg13g2_fill_2 FILLER_12_202 ();
 sg13g2_fill_1 FILLER_12_204 ();
 sg13g2_fill_2 FILLER_12_262 ();
 sg13g2_fill_1 FILLER_12_264 ();
 sg13g2_fill_1 FILLER_12_293 ();
 sg13g2_fill_2 FILLER_12_314 ();
 sg13g2_fill_1 FILLER_12_316 ();
 sg13g2_fill_1 FILLER_12_358 ();
 sg13g2_fill_1 FILLER_12_401 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_53 ();
 sg13g2_fill_2 FILLER_13_64 ();
 sg13g2_fill_2 FILLER_13_70 ();
 sg13g2_fill_1 FILLER_13_72 ();
 sg13g2_decap_4 FILLER_13_82 ();
 sg13g2_fill_2 FILLER_13_86 ();
 sg13g2_fill_2 FILLER_13_102 ();
 sg13g2_fill_1 FILLER_13_104 ();
 sg13g2_fill_1 FILLER_13_110 ();
 sg13g2_decap_4 FILLER_13_119 ();
 sg13g2_fill_1 FILLER_13_123 ();
 sg13g2_fill_2 FILLER_13_158 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_fill_2 FILLER_13_200 ();
 sg13g2_fill_1 FILLER_13_225 ();
 sg13g2_decap_8 FILLER_13_235 ();
 sg13g2_fill_1 FILLER_13_242 ();
 sg13g2_decap_8 FILLER_13_247 ();
 sg13g2_fill_1 FILLER_13_254 ();
 sg13g2_fill_2 FILLER_13_281 ();
 sg13g2_fill_1 FILLER_13_321 ();
 sg13g2_fill_1 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_4 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_15 ();
 sg13g2_decap_4 FILLER_14_22 ();
 sg13g2_fill_2 FILLER_14_26 ();
 sg13g2_decap_4 FILLER_14_41 ();
 sg13g2_fill_1 FILLER_14_138 ();
 sg13g2_fill_2 FILLER_14_164 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_fill_2 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_4 FILLER_14_259 ();
 sg13g2_fill_2 FILLER_14_282 ();
 sg13g2_fill_2 FILLER_14_294 ();
 sg13g2_fill_1 FILLER_14_296 ();
 sg13g2_decap_8 FILLER_14_302 ();
 sg13g2_fill_1 FILLER_14_309 ();
 sg13g2_fill_1 FILLER_14_314 ();
 sg13g2_fill_2 FILLER_14_348 ();
 sg13g2_fill_2 FILLER_14_393 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_2 FILLER_15_44 ();
 sg13g2_fill_1 FILLER_15_46 ();
 sg13g2_fill_2 FILLER_15_68 ();
 sg13g2_fill_1 FILLER_15_78 ();
 sg13g2_decap_4 FILLER_15_90 ();
 sg13g2_fill_1 FILLER_15_94 ();
 sg13g2_decap_8 FILLER_15_100 ();
 sg13g2_decap_8 FILLER_15_107 ();
 sg13g2_decap_4 FILLER_15_114 ();
 sg13g2_fill_2 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_204 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_242 ();
 sg13g2_fill_1 FILLER_15_244 ();
 sg13g2_fill_1 FILLER_15_253 ();
 sg13g2_decap_4 FILLER_15_303 ();
 sg13g2_fill_1 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_316 ();
 sg13g2_fill_2 FILLER_15_323 ();
 sg13g2_fill_1 FILLER_15_356 ();
 sg13g2_fill_1 FILLER_15_362 ();
 sg13g2_fill_2 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_fill_1 FILLER_16_76 ();
 sg13g2_fill_2 FILLER_16_82 ();
 sg13g2_decap_8 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_117 ();
 sg13g2_fill_2 FILLER_16_138 ();
 sg13g2_fill_1 FILLER_16_140 ();
 sg13g2_fill_2 FILLER_16_159 ();
 sg13g2_fill_2 FILLER_16_168 ();
 sg13g2_fill_2 FILLER_16_183 ();
 sg13g2_fill_1 FILLER_16_185 ();
 sg13g2_decap_8 FILLER_16_191 ();
 sg13g2_decap_8 FILLER_16_198 ();
 sg13g2_fill_1 FILLER_16_231 ();
 sg13g2_fill_2 FILLER_16_258 ();
 sg13g2_fill_2 FILLER_16_264 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_fill_2 FILLER_16_288 ();
 sg13g2_fill_1 FILLER_16_290 ();
 sg13g2_fill_2 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_361 ();
 sg13g2_fill_2 FILLER_16_394 ();
 sg13g2_fill_2 FILLER_17_53 ();
 sg13g2_fill_1 FILLER_17_55 ();
 sg13g2_fill_2 FILLER_17_97 ();
 sg13g2_fill_1 FILLER_17_99 ();
 sg13g2_decap_4 FILLER_17_128 ();
 sg13g2_fill_1 FILLER_17_132 ();
 sg13g2_decap_8 FILLER_17_159 ();
 sg13g2_fill_2 FILLER_17_166 ();
 sg13g2_fill_1 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_176 ();
 sg13g2_decap_4 FILLER_17_183 ();
 sg13g2_fill_1 FILLER_17_187 ();
 sg13g2_fill_2 FILLER_17_210 ();
 sg13g2_fill_2 FILLER_17_273 ();
 sg13g2_fill_2 FILLER_17_288 ();
 sg13g2_fill_2 FILLER_17_294 ();
 sg13g2_decap_4 FILLER_17_305 ();
 sg13g2_fill_1 FILLER_17_309 ();
 sg13g2_fill_1 FILLER_17_319 ();
 sg13g2_fill_2 FILLER_17_325 ();
 sg13g2_fill_2 FILLER_17_355 ();
 sg13g2_fill_2 FILLER_17_381 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_23 ();
 sg13g2_decap_8 FILLER_18_55 ();
 sg13g2_fill_2 FILLER_18_74 ();
 sg13g2_decap_4 FILLER_18_115 ();
 sg13g2_decap_8 FILLER_18_135 ();
 sg13g2_decap_4 FILLER_18_142 ();
 sg13g2_fill_1 FILLER_18_146 ();
 sg13g2_decap_4 FILLER_18_159 ();
 sg13g2_fill_2 FILLER_18_163 ();
 sg13g2_fill_1 FILLER_18_170 ();
 sg13g2_fill_1 FILLER_18_215 ();
 sg13g2_fill_1 FILLER_18_250 ();
 sg13g2_fill_2 FILLER_18_277 ();
 sg13g2_fill_1 FILLER_18_371 ();
 sg13g2_fill_1 FILLER_19_26 ();
 sg13g2_fill_2 FILLER_19_62 ();
 sg13g2_fill_1 FILLER_19_79 ();
 sg13g2_fill_2 FILLER_19_98 ();
 sg13g2_fill_1 FILLER_19_100 ();
 sg13g2_fill_1 FILLER_19_129 ();
 sg13g2_decap_8 FILLER_19_143 ();
 sg13g2_fill_1 FILLER_19_150 ();
 sg13g2_decap_4 FILLER_19_164 ();
 sg13g2_decap_4 FILLER_19_180 ();
 sg13g2_fill_1 FILLER_19_184 ();
 sg13g2_fill_2 FILLER_19_197 ();
 sg13g2_fill_1 FILLER_19_226 ();
 sg13g2_fill_2 FILLER_19_259 ();
 sg13g2_fill_1 FILLER_19_279 ();
 sg13g2_decap_8 FILLER_19_289 ();
 sg13g2_fill_2 FILLER_19_318 ();
 sg13g2_fill_2 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_9 ();
 sg13g2_fill_2 FILLER_20_45 ();
 sg13g2_fill_1 FILLER_20_47 ();
 sg13g2_decap_8 FILLER_20_71 ();
 sg13g2_decap_4 FILLER_20_78 ();
 sg13g2_fill_2 FILLER_20_82 ();
 sg13g2_fill_2 FILLER_20_92 ();
 sg13g2_decap_8 FILLER_20_103 ();
 sg13g2_decap_4 FILLER_20_110 ();
 sg13g2_fill_2 FILLER_20_114 ();
 sg13g2_fill_1 FILLER_20_137 ();
 sg13g2_fill_2 FILLER_20_151 ();
 sg13g2_fill_1 FILLER_20_153 ();
 sg13g2_fill_2 FILLER_20_167 ();
 sg13g2_fill_1 FILLER_20_169 ();
 sg13g2_fill_2 FILLER_20_175 ();
 sg13g2_fill_1 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_324 ();
 sg13g2_fill_1 FILLER_20_326 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_fill_1 FILLER_21_26 ();
 sg13g2_fill_1 FILLER_21_73 ();
 sg13g2_fill_2 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_131 ();
 sg13g2_fill_2 FILLER_21_138 ();
 sg13g2_decap_4 FILLER_21_153 ();
 sg13g2_fill_2 FILLER_21_170 ();
 sg13g2_fill_1 FILLER_21_172 ();
 sg13g2_fill_2 FILLER_21_190 ();
 sg13g2_fill_1 FILLER_21_192 ();
 sg13g2_decap_8 FILLER_21_197 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_fill_1 FILLER_21_210 ();
 sg13g2_fill_2 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_decap_4 FILLER_21_222 ();
 sg13g2_fill_2 FILLER_21_230 ();
 sg13g2_fill_1 FILLER_21_262 ();
 sg13g2_fill_2 FILLER_21_343 ();
 sg13g2_fill_2 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_15 ();
 sg13g2_fill_2 FILLER_22_48 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_decap_4 FILLER_22_69 ();
 sg13g2_fill_2 FILLER_22_73 ();
 sg13g2_fill_1 FILLER_22_101 ();
 sg13g2_decap_4 FILLER_22_107 ();
 sg13g2_decap_8 FILLER_22_131 ();
 sg13g2_decap_4 FILLER_22_138 ();
 sg13g2_fill_1 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_168 ();
 sg13g2_decap_4 FILLER_22_181 ();
 sg13g2_fill_1 FILLER_22_198 ();
 sg13g2_fill_2 FILLER_22_225 ();
 sg13g2_decap_4 FILLER_22_237 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_fill_1 FILLER_22_266 ();
 sg13g2_fill_1 FILLER_22_293 ();
 sg13g2_fill_2 FILLER_22_331 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_15 ();
 sg13g2_fill_1 FILLER_23_22 ();
 sg13g2_decap_4 FILLER_23_32 ();
 sg13g2_decap_4 FILLER_23_40 ();
 sg13g2_fill_1 FILLER_23_44 ();
 sg13g2_fill_1 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_59 ();
 sg13g2_fill_1 FILLER_23_76 ();
 sg13g2_fill_2 FILLER_23_85 ();
 sg13g2_fill_1 FILLER_23_87 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_fill_1 FILLER_23_138 ();
 sg13g2_decap_4 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_201 ();
 sg13g2_decap_4 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_263 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_fill_1 FILLER_23_315 ();
 sg13g2_fill_2 FILLER_23_320 ();
 sg13g2_fill_2 FILLER_23_363 ();
 sg13g2_fill_1 FILLER_23_373 ();
 sg13g2_fill_1 FILLER_24_60 ();
 sg13g2_fill_1 FILLER_24_75 ();
 sg13g2_fill_2 FILLER_24_83 ();
 sg13g2_fill_1 FILLER_24_85 ();
 sg13g2_fill_1 FILLER_24_90 ();
 sg13g2_decap_4 FILLER_24_101 ();
 sg13g2_decap_4 FILLER_24_117 ();
 sg13g2_decap_8 FILLER_24_131 ();
 sg13g2_decap_8 FILLER_24_138 ();
 sg13g2_fill_2 FILLER_24_145 ();
 sg13g2_fill_1 FILLER_24_147 ();
 sg13g2_fill_2 FILLER_24_160 ();
 sg13g2_decap_8 FILLER_24_219 ();
 sg13g2_fill_2 FILLER_24_226 ();
 sg13g2_fill_1 FILLER_24_264 ();
 sg13g2_fill_2 FILLER_24_286 ();
 sg13g2_fill_2 FILLER_24_310 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_fill_2 FILLER_24_341 ();
 sg13g2_fill_2 FILLER_24_362 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_26 ();
 sg13g2_decap_8 FILLER_25_40 ();
 sg13g2_fill_1 FILLER_25_47 ();
 sg13g2_fill_2 FILLER_25_87 ();
 sg13g2_fill_2 FILLER_25_107 ();
 sg13g2_decap_4 FILLER_25_134 ();
 sg13g2_fill_1 FILLER_25_138 ();
 sg13g2_fill_1 FILLER_25_178 ();
 sg13g2_fill_1 FILLER_25_186 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_224 ();
 sg13g2_fill_1 FILLER_25_226 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_fill_1 FILLER_25_293 ();
 sg13g2_fill_2 FILLER_25_302 ();
 sg13g2_fill_1 FILLER_25_304 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_fill_1 FILLER_25_374 ();
 sg13g2_fill_2 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_1 FILLER_26_75 ();
 sg13g2_decap_8 FILLER_26_81 ();
 sg13g2_decap_4 FILLER_26_88 ();
 sg13g2_fill_1 FILLER_26_92 ();
 sg13g2_fill_2 FILLER_26_97 ();
 sg13g2_fill_1 FILLER_26_99 ();
 sg13g2_decap_8 FILLER_26_113 ();
 sg13g2_fill_1 FILLER_26_120 ();
 sg13g2_fill_1 FILLER_26_161 ();
 sg13g2_fill_2 FILLER_26_171 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_fill_1 FILLER_26_195 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_decap_4 FILLER_26_223 ();
 sg13g2_fill_2 FILLER_26_227 ();
 sg13g2_fill_2 FILLER_26_248 ();
 sg13g2_fill_1 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_359 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_20 ();
 sg13g2_fill_2 FILLER_27_44 ();
 sg13g2_fill_1 FILLER_27_46 ();
 sg13g2_fill_2 FILLER_27_76 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_114 ();
 sg13g2_decap_8 FILLER_27_121 ();
 sg13g2_decap_4 FILLER_27_128 ();
 sg13g2_decap_8 FILLER_27_171 ();
 sg13g2_fill_2 FILLER_27_190 ();
 sg13g2_fill_2 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_264 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_decap_4 FILLER_28_52 ();
 sg13g2_fill_1 FILLER_28_56 ();
 sg13g2_fill_2 FILLER_28_65 ();
 sg13g2_fill_1 FILLER_28_67 ();
 sg13g2_fill_1 FILLER_28_108 ();
 sg13g2_decap_8 FILLER_28_135 ();
 sg13g2_decap_4 FILLER_28_142 ();
 sg13g2_decap_8 FILLER_28_162 ();
 sg13g2_decap_8 FILLER_28_169 ();
 sg13g2_fill_2 FILLER_28_176 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_fill_1 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_236 ();
 sg13g2_fill_2 FILLER_28_251 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_278 ();
 sg13g2_fill_2 FILLER_28_293 ();
 sg13g2_fill_1 FILLER_28_295 ();
 sg13g2_fill_2 FILLER_28_300 ();
 sg13g2_fill_1 FILLER_28_312 ();
 sg13g2_fill_1 FILLER_28_361 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_24 ();
 sg13g2_fill_1 FILLER_29_36 ();
 sg13g2_decap_8 FILLER_29_66 ();
 sg13g2_fill_1 FILLER_29_73 ();
 sg13g2_decap_4 FILLER_29_88 ();
 sg13g2_fill_1 FILLER_29_100 ();
 sg13g2_fill_1 FILLER_29_106 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_139 ();
 sg13g2_decap_4 FILLER_29_153 ();
 sg13g2_fill_1 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_171 ();
 sg13g2_fill_2 FILLER_29_192 ();
 sg13g2_fill_1 FILLER_29_215 ();
 sg13g2_fill_1 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_fill_2 FILLER_29_377 ();
 sg13g2_fill_2 FILLER_29_388 ();
 sg13g2_fill_2 FILLER_30_34 ();
 sg13g2_fill_1 FILLER_30_122 ();
 sg13g2_fill_2 FILLER_30_136 ();
 sg13g2_fill_1 FILLER_30_158 ();
 sg13g2_fill_2 FILLER_30_179 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_decap_4 FILLER_30_192 ();
 sg13g2_fill_1 FILLER_30_196 ();
 sg13g2_fill_2 FILLER_30_205 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_220 ();
 sg13g2_fill_2 FILLER_30_260 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_fill_1 FILLER_30_273 ();
 sg13g2_fill_2 FILLER_30_284 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_1 FILLER_30_311 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_fill_2 FILLER_31_22 ();
 sg13g2_fill_1 FILLER_31_24 ();
 sg13g2_fill_1 FILLER_31_39 ();
 sg13g2_fill_2 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_51 ();
 sg13g2_fill_1 FILLER_31_73 ();
 sg13g2_decap_4 FILLER_31_82 ();
 sg13g2_fill_1 FILLER_31_105 ();
 sg13g2_fill_1 FILLER_31_118 ();
 sg13g2_fill_2 FILLER_31_132 ();
 sg13g2_fill_2 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_145 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_fill_2 FILLER_31_187 ();
 sg13g2_fill_1 FILLER_31_189 ();
 sg13g2_fill_2 FILLER_31_253 ();
 sg13g2_fill_1 FILLER_31_255 ();
 sg13g2_fill_2 FILLER_31_300 ();
 sg13g2_fill_1 FILLER_31_333 ();
 sg13g2_fill_2 FILLER_31_381 ();
 sg13g2_fill_2 FILLER_32_110 ();
 sg13g2_fill_2 FILLER_32_129 ();
 sg13g2_fill_1 FILLER_32_159 ();
 sg13g2_fill_2 FILLER_32_165 ();
 sg13g2_fill_1 FILLER_32_215 ();
 sg13g2_fill_2 FILLER_32_225 ();
 sg13g2_fill_2 FILLER_32_275 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_15 ();
 sg13g2_fill_1 FILLER_33_38 ();
 sg13g2_decap_8 FILLER_33_67 ();
 sg13g2_fill_2 FILLER_33_92 ();
 sg13g2_fill_2 FILLER_33_103 ();
 sg13g2_decap_4 FILLER_33_124 ();
 sg13g2_fill_2 FILLER_33_128 ();
 sg13g2_fill_2 FILLER_33_140 ();
 sg13g2_fill_2 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_179 ();
 sg13g2_fill_2 FILLER_33_188 ();
 sg13g2_fill_1 FILLER_33_190 ();
 sg13g2_fill_2 FILLER_33_206 ();
 sg13g2_fill_1 FILLER_33_208 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_fill_2 FILLER_33_300 ();
 sg13g2_fill_1 FILLER_33_345 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_fill_2 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_57 ();
 sg13g2_fill_2 FILLER_34_64 ();
 sg13g2_fill_2 FILLER_34_97 ();
 sg13g2_fill_2 FILLER_34_133 ();
 sg13g2_fill_1 FILLER_34_169 ();
 sg13g2_fill_1 FILLER_34_191 ();
 sg13g2_fill_2 FILLER_34_366 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_fill_1 FILLER_35_40 ();
 sg13g2_fill_1 FILLER_35_55 ();
 sg13g2_fill_1 FILLER_35_82 ();
 sg13g2_fill_2 FILLER_35_100 ();
 sg13g2_fill_2 FILLER_35_106 ();
 sg13g2_fill_1 FILLER_35_108 ();
 sg13g2_fill_1 FILLER_35_114 ();
 sg13g2_fill_2 FILLER_35_123 ();
 sg13g2_decap_8 FILLER_35_130 ();
 sg13g2_fill_1 FILLER_35_137 ();
 sg13g2_fill_1 FILLER_35_162 ();
 sg13g2_fill_1 FILLER_35_196 ();
 sg13g2_fill_2 FILLER_35_207 ();
 sg13g2_fill_2 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_251 ();
 sg13g2_fill_1 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_292 ();
 sg13g2_fill_1 FILLER_35_342 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_fill_2 FILLER_36_23 ();
 sg13g2_fill_1 FILLER_36_25 ();
 sg13g2_fill_2 FILLER_36_34 ();
 sg13g2_fill_1 FILLER_36_36 ();
 sg13g2_fill_1 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_81 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_fill_2 FILLER_36_110 ();
 sg13g2_fill_2 FILLER_36_116 ();
 sg13g2_fill_1 FILLER_36_158 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_fill_2 FILLER_36_335 ();
 sg13g2_fill_1 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_30 ();
 sg13g2_fill_1 FILLER_37_36 ();
 sg13g2_fill_1 FILLER_37_62 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_fill_1 FILLER_37_69 ();
 sg13g2_fill_2 FILLER_37_115 ();
 sg13g2_fill_2 FILLER_37_148 ();
 sg13g2_fill_2 FILLER_37_185 ();
 sg13g2_fill_1 FILLER_37_191 ();
 sg13g2_fill_1 FILLER_37_197 ();
 sg13g2_fill_2 FILLER_37_206 ();
 sg13g2_fill_1 FILLER_37_208 ();
 sg13g2_fill_2 FILLER_37_230 ();
 sg13g2_fill_2 FILLER_37_255 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_fill_2 FILLER_37_285 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_fill_1 FILLER_37_298 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_45 ();
 sg13g2_fill_1 FILLER_38_47 ();
 sg13g2_fill_1 FILLER_38_202 ();
 sg13g2_fill_2 FILLER_38_234 ();
 sg13g2_fill_1 FILLER_38_236 ();
 sg13g2_fill_2 FILLER_38_268 ();
 sg13g2_fill_2 FILLER_38_296 ();
 sg13g2_fill_1 FILLER_38_298 ();
 sg13g2_fill_2 FILLER_38_330 ();
 sg13g2_fill_1 FILLER_38_332 ();
 sg13g2_fill_2 FILLER_38_359 ();
 assign uio_oe[0] = net12;
 assign uio_oe[1] = net13;
 assign uio_oe[2] = net14;
 assign uio_oe[3] = net252;
 assign uio_oe[4] = net253;
 assign uio_oe[5] = net254;
 assign uio_oe[6] = net255;
 assign uio_oe[7] = net256;
 assign uio_out[0] = net15;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
endmodule

module tt_um_Qwendu_spi_fpu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire clknet_leaf_0_clk;
 wire \main.SPI_input_data[0] ;
 wire \main.SPI_input_data[1] ;
 wire \main.SPI_input_data[2] ;
 wire \main.SPI_input_data[3] ;
 wire \main.SPI_input_data[4] ;
 wire \main.SPI_input_data[5] ;
 wire \main.SPI_input_data[6] ;
 wire \main.SPI_input_data[7] ;
 wire \main.SPI_input_data_valid ;
 wire \main.SPI_out ;
 wire \main.SPI_output_data_ready ;
 wire \main.adder.in_valid ;
 wire \main.adder.out[0] ;
 wire \main.adder.out[10] ;
 wire \main.adder.out[11] ;
 wire \main.adder.out[12] ;
 wire \main.adder.out[13] ;
 wire \main.adder.out[14] ;
 wire \main.adder.out[15] ;
 wire \main.adder.out[16] ;
 wire \main.adder.out[17] ;
 wire \main.adder.out[18] ;
 wire \main.adder.out[19] ;
 wire \main.adder.out[1] ;
 wire \main.adder.out[20] ;
 wire \main.adder.out[21] ;
 wire \main.adder.out[22] ;
 wire \main.adder.out[23] ;
 wire \main.adder.out[24] ;
 wire \main.adder.out[25] ;
 wire \main.adder.out[26] ;
 wire \main.adder.out[27] ;
 wire \main.adder.out[28] ;
 wire \main.adder.out[29] ;
 wire \main.adder.out[2] ;
 wire \main.adder.out[30] ;
 wire \main.adder.out[31] ;
 wire \main.adder.out[3] ;
 wire \main.adder.out[4] ;
 wire \main.adder.out[5] ;
 wire \main.adder.out[6] ;
 wire \main.adder.out[7] ;
 wire \main.adder.out[8] ;
 wire \main.adder.out[9] ;
 wire \main.adder.out_valid ;
 wire \main.adder.s1_exp_diff[0] ;
 wire \main.adder.s1_exp_diff[1] ;
 wire \main.adder.s1_exp_diff[2] ;
 wire \main.adder.s1_exp_diff[3] ;
 wire \main.adder.s1_exp_diff[4] ;
 wire \main.adder.s1_exp_diff[5] ;
 wire \main.adder.s1_exp_diff[6] ;
 wire \main.adder.s1_exp_diff[7] ;
 wire \main.adder.s1_exp_diff[8] ;
 wire \main.adder.s1_exp_diff[9] ;
 wire \main.adder.s1_inf ;
 wire \main.adder.s1_larger[0] ;
 wire \main.adder.s1_larger[10] ;
 wire \main.adder.s1_larger[11] ;
 wire \main.adder.s1_larger[12] ;
 wire \main.adder.s1_larger[13] ;
 wire \main.adder.s1_larger[14] ;
 wire \main.adder.s1_larger[15] ;
 wire \main.adder.s1_larger[16] ;
 wire \main.adder.s1_larger[17] ;
 wire \main.adder.s1_larger[18] ;
 wire \main.adder.s1_larger[19] ;
 wire \main.adder.s1_larger[1] ;
 wire \main.adder.s1_larger[20] ;
 wire \main.adder.s1_larger[21] ;
 wire \main.adder.s1_larger[22] ;
 wire \main.adder.s1_larger[23] ;
 wire \main.adder.s1_larger[24] ;
 wire \main.adder.s1_larger[25] ;
 wire \main.adder.s1_larger[26] ;
 wire \main.adder.s1_larger[27] ;
 wire \main.adder.s1_larger[28] ;
 wire \main.adder.s1_larger[29] ;
 wire \main.adder.s1_larger[2] ;
 wire \main.adder.s1_larger[30] ;
 wire \main.adder.s1_larger[31] ;
 wire \main.adder.s1_larger[3] ;
 wire \main.adder.s1_larger[4] ;
 wire \main.adder.s1_larger[5] ;
 wire \main.adder.s1_larger[6] ;
 wire \main.adder.s1_larger[7] ;
 wire \main.adder.s1_larger[8] ;
 wire \main.adder.s1_larger[9] ;
 wire \main.adder.s1_nan ;
 wire \main.adder.s1_rs.levels[0][23] ;
 wire \main.adder.s1_rs.levels[0][24] ;
 wire \main.adder.s1_rs.levels[0][25] ;
 wire \main.adder.s1_rs.levels[0][26] ;
 wire \main.adder.s1_rs.levels[0][27] ;
 wire \main.adder.s1_rs.levels[0][28] ;
 wire \main.adder.s1_rs.levels[0][29] ;
 wire \main.adder.s1_rs.levels[0][30] ;
 wire \main.adder.s1_rs.levels[0][31] ;
 wire \main.adder.s1_rs.levels[0][32] ;
 wire \main.adder.s1_rs.levels[0][33] ;
 wire \main.adder.s1_rs.levels[0][34] ;
 wire \main.adder.s1_rs.levels[0][35] ;
 wire \main.adder.s1_rs.levels[0][36] ;
 wire \main.adder.s1_rs.levels[0][37] ;
 wire \main.adder.s1_rs.levels[0][38] ;
 wire \main.adder.s1_rs.levels[0][39] ;
 wire \main.adder.s1_rs.levels[0][40] ;
 wire \main.adder.s1_rs.levels[0][41] ;
 wire \main.adder.s1_rs.levels[0][42] ;
 wire \main.adder.s1_rs.levels[0][43] ;
 wire \main.adder.s1_rs.levels[0][44] ;
 wire \main.adder.s1_rs.levels[0][45] ;
 wire \main.adder.s1_smaler[23] ;
 wire \main.adder.s1_smaler[24] ;
 wire \main.adder.s1_smaler[25] ;
 wire \main.adder.s1_smaler[26] ;
 wire \main.adder.s1_smaler[27] ;
 wire \main.adder.s1_smaler[28] ;
 wire \main.adder.s1_smaler[29] ;
 wire \main.adder.s1_smaler[30] ;
 wire \main.adder.s1_smaler[31] ;
 wire \main.adder.s1_valid ;
 wire \main.adder.s2_exponent[0] ;
 wire \main.adder.s2_exponent[1] ;
 wire \main.adder.s2_exponent[2] ;
 wire \main.adder.s2_exponent[3] ;
 wire \main.adder.s2_exponent[4] ;
 wire \main.adder.s2_exponent[5] ;
 wire \main.adder.s2_exponent[6] ;
 wire \main.adder.s2_exponent[7] ;
 wire \main.adder.s2_flip_sign ;
 wire \main.adder.s2_inf ;
 wire \main.adder.s2_larger[23] ;
 wire \main.adder.s2_larger[24] ;
 wire \main.adder.s2_larger[25] ;
 wire \main.adder.s2_larger[26] ;
 wire \main.adder.s2_larger[27] ;
 wire \main.adder.s2_larger[28] ;
 wire \main.adder.s2_larger[29] ;
 wire \main.adder.s2_larger[30] ;
 wire \main.adder.s2_larger[31] ;
 wire \main.adder.s2_larger[32] ;
 wire \main.adder.s2_larger[33] ;
 wire \main.adder.s2_larger[34] ;
 wire \main.adder.s2_larger[35] ;
 wire \main.adder.s2_larger[36] ;
 wire \main.adder.s2_larger[37] ;
 wire \main.adder.s2_larger[38] ;
 wire \main.adder.s2_larger[39] ;
 wire \main.adder.s2_larger[40] ;
 wire \main.adder.s2_larger[41] ;
 wire \main.adder.s2_larger[42] ;
 wire \main.adder.s2_larger[43] ;
 wire \main.adder.s2_larger[44] ;
 wire \main.adder.s2_larger[45] ;
 wire \main.adder.s2_larger[46] ;
 wire \main.adder.s2_nan ;
 wire \main.adder.s2_shared_sign ;
 wire \main.adder.s2_smaler[0] ;
 wire \main.adder.s2_smaler[10] ;
 wire \main.adder.s2_smaler[11] ;
 wire \main.adder.s2_smaler[12] ;
 wire \main.adder.s2_smaler[13] ;
 wire \main.adder.s2_smaler[14] ;
 wire \main.adder.s2_smaler[15] ;
 wire \main.adder.s2_smaler[16] ;
 wire \main.adder.s2_smaler[17] ;
 wire \main.adder.s2_smaler[18] ;
 wire \main.adder.s2_smaler[19] ;
 wire \main.adder.s2_smaler[1] ;
 wire \main.adder.s2_smaler[20] ;
 wire \main.adder.s2_smaler[21] ;
 wire \main.adder.s2_smaler[22] ;
 wire \main.adder.s2_smaler[23] ;
 wire \main.adder.s2_smaler[24] ;
 wire \main.adder.s2_smaler[25] ;
 wire \main.adder.s2_smaler[26] ;
 wire \main.adder.s2_smaler[27] ;
 wire \main.adder.s2_smaler[28] ;
 wire \main.adder.s2_smaler[29] ;
 wire \main.adder.s2_smaler[2] ;
 wire \main.adder.s2_smaler[30] ;
 wire \main.adder.s2_smaler[31] ;
 wire \main.adder.s2_smaler[32] ;
 wire \main.adder.s2_smaler[33] ;
 wire \main.adder.s2_smaler[34] ;
 wire \main.adder.s2_smaler[35] ;
 wire \main.adder.s2_smaler[36] ;
 wire \main.adder.s2_smaler[37] ;
 wire \main.adder.s2_smaler[38] ;
 wire \main.adder.s2_smaler[39] ;
 wire \main.adder.s2_smaler[3] ;
 wire \main.adder.s2_smaler[40] ;
 wire \main.adder.s2_smaler[41] ;
 wire \main.adder.s2_smaler[42] ;
 wire \main.adder.s2_smaler[43] ;
 wire \main.adder.s2_smaler[44] ;
 wire \main.adder.s2_smaler[45] ;
 wire \main.adder.s2_smaler[46] ;
 wire \main.adder.s2_smaler[4] ;
 wire \main.adder.s2_smaler[5] ;
 wire \main.adder.s2_smaler[6] ;
 wire \main.adder.s2_smaler[7] ;
 wire \main.adder.s2_smaler[8] ;
 wire \main.adder.s2_smaler[9] ;
 wire \main.adder.s2_valid ;
 wire \main.adder.s3_exponent[0] ;
 wire \main.adder.s3_exponent[1] ;
 wire \main.adder.s3_exponent[2] ;
 wire \main.adder.s3_exponent[3] ;
 wire \main.adder.s3_exponent[4] ;
 wire \main.adder.s3_exponent[5] ;
 wire \main.adder.s3_exponent[6] ;
 wire \main.adder.s3_exponent[7] ;
 wire \main.adder.s3_flipped ;
 wire \main.adder.s3_inf ;
 wire \main.adder.s3_nan ;
 wire \main.adder.s3_shared_sign ;
 wire \main.adder.s3_sum[0] ;
 wire \main.adder.s3_sum[10] ;
 wire \main.adder.s3_sum[11] ;
 wire \main.adder.s3_sum[12] ;
 wire \main.adder.s3_sum[13] ;
 wire \main.adder.s3_sum[14] ;
 wire \main.adder.s3_sum[15] ;
 wire \main.adder.s3_sum[16] ;
 wire \main.adder.s3_sum[17] ;
 wire \main.adder.s3_sum[18] ;
 wire \main.adder.s3_sum[19] ;
 wire \main.adder.s3_sum[1] ;
 wire \main.adder.s3_sum[20] ;
 wire \main.adder.s3_sum[21] ;
 wire \main.adder.s3_sum[22] ;
 wire \main.adder.s3_sum[23] ;
 wire \main.adder.s3_sum[24] ;
 wire \main.adder.s3_sum[25] ;
 wire \main.adder.s3_sum[26] ;
 wire \main.adder.s3_sum[27] ;
 wire \main.adder.s3_sum[28] ;
 wire \main.adder.s3_sum[29] ;
 wire \main.adder.s3_sum[2] ;
 wire \main.adder.s3_sum[30] ;
 wire \main.adder.s3_sum[31] ;
 wire \main.adder.s3_sum[32] ;
 wire \main.adder.s3_sum[33] ;
 wire \main.adder.s3_sum[34] ;
 wire \main.adder.s3_sum[35] ;
 wire \main.adder.s3_sum[36] ;
 wire \main.adder.s3_sum[37] ;
 wire \main.adder.s3_sum[38] ;
 wire \main.adder.s3_sum[39] ;
 wire \main.adder.s3_sum[3] ;
 wire \main.adder.s3_sum[40] ;
 wire \main.adder.s3_sum[41] ;
 wire \main.adder.s3_sum[42] ;
 wire \main.adder.s3_sum[43] ;
 wire \main.adder.s3_sum[44] ;
 wire \main.adder.s3_sum[45] ;
 wire \main.adder.s3_sum[46] ;
 wire \main.adder.s3_sum[47] ;
 wire \main.adder.s3_sum[48] ;
 wire \main.adder.s3_sum[4] ;
 wire \main.adder.s3_sum[5] ;
 wire \main.adder.s3_sum[6] ;
 wire \main.adder.s3_sum[7] ;
 wire \main.adder.s3_sum[8] ;
 wire \main.adder.s3_sum[9] ;
 wire \main.adder.s3_valid ;
 wire \main.adder.s4_exponent[0] ;
 wire \main.adder.s4_exponent[1] ;
 wire \main.adder.s4_exponent[2] ;
 wire \main.adder.s4_exponent[3] ;
 wire \main.adder.s4_exponent[4] ;
 wire \main.adder.s4_exponent[5] ;
 wire \main.adder.s4_exponent[6] ;
 wire \main.adder.s4_exponent[7] ;
 wire \main.adder.s4_exponent_adjust[0] ;
 wire \main.adder.s4_exponent_adjust[1] ;
 wire \main.adder.s4_exponent_adjust[2] ;
 wire \main.adder.s4_exponent_adjust[3] ;
 wire \main.adder.s4_exponent_adjust[4] ;
 wire \main.adder.s4_exponent_adjust[5] ;
 wire \main.adder.s4_exponent_adjust[6] ;
 wire \main.adder.s4_exponent_adjust[7] ;
 wire \main.adder.s4_exponent_adjust[8] ;
 wire \main.adder.s4_exponent_adjust[9] ;
 wire \main.adder.s4_flipped ;
 wire \main.adder.s4_inf ;
 wire \main.adder.s4_mant[0] ;
 wire \main.adder.s4_mant[10] ;
 wire \main.adder.s4_mant[11] ;
 wire \main.adder.s4_mant[12] ;
 wire \main.adder.s4_mant[13] ;
 wire \main.adder.s4_mant[14] ;
 wire \main.adder.s4_mant[15] ;
 wire \main.adder.s4_mant[16] ;
 wire \main.adder.s4_mant[17] ;
 wire \main.adder.s4_mant[18] ;
 wire \main.adder.s4_mant[19] ;
 wire \main.adder.s4_mant[1] ;
 wire \main.adder.s4_mant[20] ;
 wire \main.adder.s4_mant[21] ;
 wire \main.adder.s4_mant[22] ;
 wire \main.adder.s4_mant[23] ;
 wire \main.adder.s4_mant[24] ;
 wire \main.adder.s4_mant[25] ;
 wire \main.adder.s4_mant[26] ;
 wire \main.adder.s4_mant[27] ;
 wire \main.adder.s4_mant[28] ;
 wire \main.adder.s4_mant[29] ;
 wire \main.adder.s4_mant[2] ;
 wire \main.adder.s4_mant[30] ;
 wire \main.adder.s4_mant[31] ;
 wire \main.adder.s4_mant[32] ;
 wire \main.adder.s4_mant[33] ;
 wire \main.adder.s4_mant[34] ;
 wire \main.adder.s4_mant[35] ;
 wire \main.adder.s4_mant[36] ;
 wire \main.adder.s4_mant[37] ;
 wire \main.adder.s4_mant[38] ;
 wire \main.adder.s4_mant[39] ;
 wire \main.adder.s4_mant[3] ;
 wire \main.adder.s4_mant[40] ;
 wire \main.adder.s4_mant[41] ;
 wire \main.adder.s4_mant[42] ;
 wire \main.adder.s4_mant[43] ;
 wire \main.adder.s4_mant[44] ;
 wire \main.adder.s4_mant[45] ;
 wire \main.adder.s4_mant[46] ;
 wire \main.adder.s4_mant[47] ;
 wire \main.adder.s4_mant[4] ;
 wire \main.adder.s4_mant[5] ;
 wire \main.adder.s4_mant[6] ;
 wire \main.adder.s4_mant[7] ;
 wire \main.adder.s4_mant[8] ;
 wire \main.adder.s4_mant[9] ;
 wire \main.adder.s4_nan ;
 wire \main.adder.s4_shared_sign ;
 wire \main.adder.s4_sum[48] ;
 wire \main.adder.s4_valid ;
 wire \main.adder.s5_R ;
 wire \main.adder.s5_S ;
 wire \main.adder.s5_exponent[0] ;
 wire \main.adder.s5_exponent[1] ;
 wire \main.adder.s5_exponent[2] ;
 wire \main.adder.s5_exponent[3] ;
 wire \main.adder.s5_exponent[4] ;
 wire \main.adder.s5_exponent[5] ;
 wire \main.adder.s5_exponent[6] ;
 wire \main.adder.s5_exponent[7] ;
 wire \main.adder.s5_exponent[8] ;
 wire \main.adder.s5_exponent[9] ;
 wire \main.adder.s5_inf ;
 wire \main.adder.s5_mant[0] ;
 wire \main.adder.s5_mant[10] ;
 wire \main.adder.s5_mant[11] ;
 wire \main.adder.s5_mant[12] ;
 wire \main.adder.s5_mant[13] ;
 wire \main.adder.s5_mant[14] ;
 wire \main.adder.s5_mant[15] ;
 wire \main.adder.s5_mant[16] ;
 wire \main.adder.s5_mant[17] ;
 wire \main.adder.s5_mant[18] ;
 wire \main.adder.s5_mant[19] ;
 wire \main.adder.s5_mant[1] ;
 wire \main.adder.s5_mant[20] ;
 wire \main.adder.s5_mant[21] ;
 wire \main.adder.s5_mant[22] ;
 wire \main.adder.s5_mant[23] ;
 wire \main.adder.s5_mant[2] ;
 wire \main.adder.s5_mant[3] ;
 wire \main.adder.s5_mant[4] ;
 wire \main.adder.s5_mant[5] ;
 wire \main.adder.s5_mant[6] ;
 wire \main.adder.s5_mant[7] ;
 wire \main.adder.s5_mant[8] ;
 wire \main.adder.s5_mant[9] ;
 wire \main.adder.s5_nan ;
 wire \main.adder.s5_sign ;
 wire \main.adder.s5_valid ;
 wire \main.byte_counter[0] ;
 wire \main.byte_counter[1] ;
 wire \main.float_registers[0][0] ;
 wire \main.float_registers[0][10] ;
 wire \main.float_registers[0][11] ;
 wire \main.float_registers[0][12] ;
 wire \main.float_registers[0][13] ;
 wire \main.float_registers[0][14] ;
 wire \main.float_registers[0][15] ;
 wire \main.float_registers[0][16] ;
 wire \main.float_registers[0][17] ;
 wire \main.float_registers[0][18] ;
 wire \main.float_registers[0][19] ;
 wire \main.float_registers[0][1] ;
 wire \main.float_registers[0][20] ;
 wire \main.float_registers[0][21] ;
 wire \main.float_registers[0][22] ;
 wire \main.float_registers[0][23] ;
 wire \main.float_registers[0][24] ;
 wire \main.float_registers[0][25] ;
 wire \main.float_registers[0][26] ;
 wire \main.float_registers[0][27] ;
 wire \main.float_registers[0][28] ;
 wire \main.float_registers[0][29] ;
 wire \main.float_registers[0][2] ;
 wire \main.float_registers[0][30] ;
 wire \main.float_registers[0][31] ;
 wire \main.float_registers[0][3] ;
 wire \main.float_registers[0][4] ;
 wire \main.float_registers[0][5] ;
 wire \main.float_registers[0][6] ;
 wire \main.float_registers[0][7] ;
 wire \main.float_registers[0][8] ;
 wire \main.float_registers[0][9] ;
 wire \main.float_registers[1][0] ;
 wire \main.float_registers[1][10] ;
 wire \main.float_registers[1][11] ;
 wire \main.float_registers[1][12] ;
 wire \main.float_registers[1][13] ;
 wire \main.float_registers[1][14] ;
 wire \main.float_registers[1][15] ;
 wire \main.float_registers[1][16] ;
 wire \main.float_registers[1][17] ;
 wire \main.float_registers[1][18] ;
 wire \main.float_registers[1][19] ;
 wire \main.float_registers[1][1] ;
 wire \main.float_registers[1][20] ;
 wire \main.float_registers[1][21] ;
 wire \main.float_registers[1][22] ;
 wire \main.float_registers[1][23] ;
 wire \main.float_registers[1][24] ;
 wire \main.float_registers[1][25] ;
 wire \main.float_registers[1][26] ;
 wire \main.float_registers[1][27] ;
 wire \main.float_registers[1][28] ;
 wire \main.float_registers[1][29] ;
 wire \main.float_registers[1][2] ;
 wire \main.float_registers[1][30] ;
 wire \main.float_registers[1][31] ;
 wire \main.float_registers[1][3] ;
 wire \main.float_registers[1][4] ;
 wire \main.float_registers[1][5] ;
 wire \main.float_registers[1][6] ;
 wire \main.float_registers[1][7] ;
 wire \main.float_registers[1][8] ;
 wire \main.float_registers[1][9] ;
 wire \main.float_registers[2][0] ;
 wire \main.float_registers[2][10] ;
 wire \main.float_registers[2][11] ;
 wire \main.float_registers[2][12] ;
 wire \main.float_registers[2][13] ;
 wire \main.float_registers[2][14] ;
 wire \main.float_registers[2][15] ;
 wire \main.float_registers[2][16] ;
 wire \main.float_registers[2][17] ;
 wire \main.float_registers[2][18] ;
 wire \main.float_registers[2][19] ;
 wire \main.float_registers[2][1] ;
 wire \main.float_registers[2][20] ;
 wire \main.float_registers[2][21] ;
 wire \main.float_registers[2][22] ;
 wire \main.float_registers[2][23] ;
 wire \main.float_registers[2][24] ;
 wire \main.float_registers[2][25] ;
 wire \main.float_registers[2][26] ;
 wire \main.float_registers[2][27] ;
 wire \main.float_registers[2][28] ;
 wire \main.float_registers[2][29] ;
 wire \main.float_registers[2][2] ;
 wire \main.float_registers[2][30] ;
 wire \main.float_registers[2][31] ;
 wire \main.float_registers[2][3] ;
 wire \main.float_registers[2][4] ;
 wire \main.float_registers[2][5] ;
 wire \main.float_registers[2][6] ;
 wire \main.float_registers[2][7] ;
 wire \main.float_registers[2][8] ;
 wire \main.float_registers[2][9] ;
 wire \main.float_registers[3][0] ;
 wire \main.float_registers[3][10] ;
 wire \main.float_registers[3][11] ;
 wire \main.float_registers[3][12] ;
 wire \main.float_registers[3][13] ;
 wire \main.float_registers[3][14] ;
 wire \main.float_registers[3][15] ;
 wire \main.float_registers[3][16] ;
 wire \main.float_registers[3][17] ;
 wire \main.float_registers[3][18] ;
 wire \main.float_registers[3][19] ;
 wire \main.float_registers[3][1] ;
 wire \main.float_registers[3][20] ;
 wire \main.float_registers[3][21] ;
 wire \main.float_registers[3][22] ;
 wire \main.float_registers[3][23] ;
 wire \main.float_registers[3][24] ;
 wire \main.float_registers[3][25] ;
 wire \main.float_registers[3][26] ;
 wire \main.float_registers[3][27] ;
 wire \main.float_registers[3][28] ;
 wire \main.float_registers[3][29] ;
 wire \main.float_registers[3][2] ;
 wire \main.float_registers[3][30] ;
 wire \main.float_registers[3][31] ;
 wire \main.float_registers[3][3] ;
 wire \main.float_registers[3][4] ;
 wire \main.float_registers[3][5] ;
 wire \main.float_registers[3][6] ;
 wire \main.float_registers[3][7] ;
 wire \main.float_registers[3][8] ;
 wire \main.float_registers[3][9] ;
 wire \main.read_command[0] ;
 wire \main.read_command[1] ;
 wire \main.register_id_input_a[0] ;
 wire \main.register_id_input_a[1] ;
 wire \main.register_id_input_b[0] ;
 wire \main.register_id_input_b[1] ;
 wire \main.register_id_result[0] ;
 wire \main.register_id_result[1] ;
 wire \main.spi.SPI_clock_sampled ;
 wire \main.spi.SPI_clock_sampler.sample_register[0] ;
 wire \main.spi.SPI_in_sampled ;
 wire \main.spi.SPI_in_sampler.sample_register[0] ;
 wire \main.spi.SPI_not_chip_select_sampled ;
 wire \main.spi.SPI_not_chip_select_sampler.sample_register[0] ;
 wire \main.spi.in_bit_counter[0] ;
 wire \main.spi.in_bit_counter[1] ;
 wire \main.spi.in_bit_counter[2] ;
 wire \main.spi.out_bit_counter[0] ;
 wire \main.spi.out_bit_counter[1] ;
 wire \main.spi.out_bit_counter[2] ;
 wire \main.spi.out_data_r[0] ;
 wire \main.spi.out_data_r[1] ;
 wire \main.spi.out_data_r[2] ;
 wire \main.spi.out_data_r[3] ;
 wire \main.spi.out_data_r[4] ;
 wire \main.spi.out_data_r[5] ;
 wire \main.spi.out_data_r[6] ;
 wire \main.spi.out_data_r[7] ;
 wire \main.spi.state[0] ;
 wire \main.state[0] ;
 wire \main.state[1] ;
 wire \main.state[2] ;
 wire \main.state[4] ;
 wire \main.state[6] ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;

 sg13g2_inv_2 _3833_ (.Y(_0664_),
    .A(net702));
 sg13g2_inv_1 _3834_ (.Y(_0665_),
    .A(\main.register_id_result[0] ));
 sg13g2_inv_2 _3835_ (.Y(_0666_),
    .A(net665));
 sg13g2_inv_1 _3836_ (.Y(_0667_),
    .A(net712));
 sg13g2_inv_1 _3837_ (.Y(_0668_),
    .A(net713));
 sg13g2_inv_1 _3838_ (.Y(_0669_),
    .A(net692));
 sg13g2_inv_1 _3839_ (.Y(_0670_),
    .A(net627));
 sg13g2_inv_1 _3840_ (.Y(_0671_),
    .A(net1555));
 sg13g2_inv_1 _3841_ (.Y(_0672_),
    .A(net1531));
 sg13g2_inv_1 _3842_ (.Y(_0673_),
    .A(net1573));
 sg13g2_inv_1 _3843_ (.Y(_0674_),
    .A(net1537));
 sg13g2_inv_1 _3844_ (.Y(_0675_),
    .A(net1544));
 sg13g2_inv_1 _3845_ (.Y(_0676_),
    .A(net615));
 sg13g2_inv_1 _3846_ (.Y(_0677_),
    .A(net582));
 sg13g2_inv_1 _3847_ (.Y(_0678_),
    .A(net1429));
 sg13g2_inv_1 _3848_ (.Y(_0679_),
    .A(net1592));
 sg13g2_inv_1 _3849_ (.Y(_0680_),
    .A(\main.spi.out_bit_counter[0] ));
 sg13g2_inv_1 _3850_ (.Y(_0681_),
    .A(\main.adder.s3_sum[15] ));
 sg13g2_inv_1 _3851_ (.Y(_0682_),
    .A(\main.adder.s3_sum[12] ));
 sg13g2_inv_1 _3852_ (.Y(_0683_),
    .A(\main.adder.s3_sum[7] ));
 sg13g2_inv_1 _3853_ (.Y(_0684_),
    .A(net953));
 sg13g2_inv_1 _3854_ (.Y(_0685_),
    .A(\main.adder.s3_sum[30] ));
 sg13g2_inv_1 _3855_ (.Y(_0686_),
    .A(\main.adder.s3_sum[32] ));
 sg13g2_inv_2 _3856_ (.Y(_0687_),
    .A(net1618));
 sg13g2_inv_1 _3857_ (.Y(_0688_),
    .A(\main.adder.s3_sum[47] ));
 sg13g2_inv_1 _3858_ (.Y(_0689_),
    .A(net1568));
 sg13g2_inv_1 _3859_ (.Y(_0690_),
    .A(net1600));
 sg13g2_inv_1 _3860_ (.Y(_0691_),
    .A(net1548));
 sg13g2_inv_1 _3861_ (.Y(_0692_),
    .A(net1571));
 sg13g2_inv_1 _3862_ (.Y(_0693_),
    .A(net1543));
 sg13g2_inv_1 _3863_ (.Y(_0694_),
    .A(net1580));
 sg13g2_inv_1 _3864_ (.Y(_0695_),
    .A(_0022_));
 sg13g2_inv_1 _3865_ (.Y(_0696_),
    .A(_0030_));
 sg13g2_inv_1 _3866_ (.Y(_0697_),
    .A(net1273));
 sg13g2_inv_1 _3867_ (.Y(_0698_),
    .A(net1590));
 sg13g2_inv_1 _3868_ (.Y(_0699_),
    .A(net1527));
 sg13g2_inv_1 _3869_ (.Y(_0700_),
    .A(net1345));
 sg13g2_inv_1 _3870_ (.Y(_0701_),
    .A(net588));
 sg13g2_inv_1 _3871_ (.Y(_0702_),
    .A(\main.state[4] ));
 sg13g2_inv_1 _3872_ (.Y(_0703_),
    .A(\main.adder.s5_R ));
 sg13g2_inv_2 _3873_ (.Y(_0704_),
    .A(net1508));
 sg13g2_inv_1 _3874_ (.Y(_0705_),
    .A(net805));
 sg13g2_inv_1 _3875_ (.Y(_0706_),
    .A(net1561));
 sg13g2_inv_2 _3876_ (.Y(_0707_),
    .A(net1513));
 sg13g2_inv_1 _3877_ (.Y(_0708_),
    .A(net1461));
 sg13g2_inv_1 _3878_ (.Y(_0709_),
    .A(net1474));
 sg13g2_inv_2 _3879_ (.Y(_0710_),
    .A(\main.adder.s5_mant[13] ));
 sg13g2_inv_1 _3880_ (.Y(_0711_),
    .A(net1597));
 sg13g2_inv_1 _3881_ (.Y(_0712_),
    .A(net1401));
 sg13g2_inv_1 _3882_ (.Y(_0713_),
    .A(net962));
 sg13g2_inv_1 _3883_ (.Y(_0714_),
    .A(\main.adder.s4_exponent_adjust[6] ));
 sg13g2_inv_2 _3884_ (.Y(_0715_),
    .A(net1282));
 sg13g2_inv_2 _3885_ (.Y(_0716_),
    .A(net1281));
 sg13g2_inv_1 _3886_ (.Y(_0717_),
    .A(_0061_));
 sg13g2_inv_1 _3887_ (.Y(_0718_),
    .A(_0062_));
 sg13g2_inv_1 _3888_ (.Y(_0719_),
    .A(_0063_));
 sg13g2_inv_1 _3889_ (.Y(_0720_),
    .A(_0065_));
 sg13g2_inv_1 _3890_ (.Y(_0721_),
    .A(_0066_));
 sg13g2_inv_1 _3891_ (.Y(_0722_),
    .A(_0067_));
 sg13g2_inv_1 _3892_ (.Y(_0723_),
    .A(_0069_));
 sg13g2_inv_1 _3893_ (.Y(_0724_),
    .A(_0070_));
 sg13g2_inv_1 _3894_ (.Y(_0725_),
    .A(_0071_));
 sg13g2_inv_2 _3895_ (.Y(_0726_),
    .A(\main.adder.s3_exponent[3] ));
 sg13g2_inv_2 _3896_ (.Y(_0727_),
    .A(\main.adder.s3_exponent[6] ));
 sg13g2_inv_1 _3897_ (.Y(_0728_),
    .A(net1574));
 sg13g2_inv_1 _3898_ (.Y(_0729_),
    .A(\main.adder.out[16] ));
 sg13g2_inv_1 _3899_ (.Y(_0730_),
    .A(\main.adder.out[17] ));
 sg13g2_inv_1 _3900_ (.Y(_0731_),
    .A(\main.adder.out[18] ));
 sg13g2_inv_1 _3901_ (.Y(_0732_),
    .A(\main.adder.out[19] ));
 sg13g2_inv_1 _3902_ (.Y(_0733_),
    .A(\main.adder.out[20] ));
 sg13g2_inv_1 _3903_ (.Y(_0734_),
    .A(\main.adder.out[21] ));
 sg13g2_inv_1 _3904_ (.Y(_0735_),
    .A(\main.adder.out[22] ));
 sg13g2_inv_1 _3905_ (.Y(_0736_),
    .A(net946));
 sg13g2_inv_1 _3906_ (.Y(_0737_),
    .A(net886));
 sg13g2_inv_1 _3907_ (.Y(_0738_),
    .A(net758));
 sg13g2_inv_1 _3908_ (.Y(_0739_),
    .A(net1022));
 sg13g2_inv_1 _3909_ (.Y(_0740_),
    .A(net1004));
 sg13g2_inv_1 _3910_ (.Y(_0741_),
    .A(net916));
 sg13g2_inv_1 _3911_ (.Y(_0742_),
    .A(net1398));
 sg13g2_inv_1 _3912_ (.Y(_0743_),
    .A(net968));
 sg13g2_inv_1 _3913_ (.Y(_0744_),
    .A(\main.adder.out[31] ));
 sg13g2_inv_1 _3914_ (.Y(_0745_),
    .A(_0075_));
 sg13g2_inv_2 _3915_ (.Y(_0746_),
    .A(net1441));
 sg13g2_inv_1 _3916_ (.Y(_0747_),
    .A(\main.adder.s2_larger[26] ));
 sg13g2_inv_1 _3917_ (.Y(_0748_),
    .A(net801));
 sg13g2_inv_1 _3918_ (.Y(_0749_),
    .A(net1041));
 sg13g2_inv_1 _3919_ (.Y(_0750_),
    .A(net1557));
 sg13g2_inv_1 _3920_ (.Y(_0751_),
    .A(net899));
 sg13g2_inv_1 _3921_ (.Y(_0752_),
    .A(net748));
 sg13g2_inv_1 _3922_ (.Y(_0753_),
    .A(net885));
 sg13g2_inv_1 _3923_ (.Y(_0754_),
    .A(net1001));
 sg13g2_inv_1 _3924_ (.Y(_0755_),
    .A(net1581));
 sg13g2_inv_1 _3925_ (.Y(_0756_),
    .A(net959));
 sg13g2_inv_1 _3926_ (.Y(_0757_),
    .A(net688));
 sg13g2_inv_1 _3927_ (.Y(_0758_),
    .A(net1028));
 sg13g2_inv_1 _3928_ (.Y(_0759_),
    .A(net686));
 sg13g2_inv_1 _3929_ (.Y(_0760_),
    .A(net1554));
 sg13g2_inv_1 _3930_ (.Y(_0761_),
    .A(net807));
 sg13g2_inv_1 _3931_ (.Y(_0762_),
    .A(net715));
 sg13g2_inv_1 _3932_ (.Y(_0763_),
    .A(net732));
 sg13g2_nor2_1 _3933_ (.A(_0697_),
    .B(\main.spi.SPI_not_chip_select_sampled ),
    .Y(_0764_));
 sg13g2_nor2_1 _3934_ (.A(\main.spi.SPI_not_chip_select_sampled ),
    .B(net1300),
    .Y(_0765_));
 sg13g2_inv_1 _3935_ (.Y(_0006_),
    .A(net1225));
 sg13g2_nand3_1 _3936_ (.B(net1273),
    .C(net1225),
    .A(net749),
    .Y(_0766_));
 sg13g2_nor2_1 _3937_ (.A(\main.read_command[0] ),
    .B(_0699_),
    .Y(_0767_));
 sg13g2_nand2_1 _3938_ (.Y(_0768_),
    .A(_0698_),
    .B(\main.read_command[1] ));
 sg13g2_nor2_1 _3939_ (.A(\main.SPI_output_data_ready ),
    .B(_0768_),
    .Y(_0769_));
 sg13g2_and2_2 _3940_ (.A(net1292),
    .B(net1283),
    .X(_0770_));
 sg13g2_inv_1 _3941_ (.Y(_0771_),
    .A(_0770_));
 sg13g2_o21ai_1 _3942_ (.B1(_0770_),
    .Y(_0772_),
    .A1(net1273),
    .A2(\main.read_command[1] ));
 sg13g2_a21oi_1 _3943_ (.A1(_0698_),
    .A2(_0772_),
    .Y(_0773_),
    .B1(_0769_));
 sg13g2_nand2_1 _3944_ (.Y(_0774_),
    .A(net851),
    .B(net1225));
 sg13g2_o21ai_1 _3945_ (.B1(_0766_),
    .Y(_0011_),
    .A1(_0773_),
    .A2(_0774_));
 sg13g2_and2_1 _3946_ (.A(net1338),
    .B(net879),
    .X(_0523_));
 sg13g2_nand2_1 _3947_ (.Y(_0775_),
    .A(\main.adder.in_valid ),
    .B(_0765_));
 sg13g2_nand2_1 _3948_ (.Y(_0776_),
    .A(net1274),
    .B(net1225));
 sg13g2_nor2b_2 _3949_ (.A(net1283),
    .B_N(net1292),
    .Y(_0777_));
 sg13g2_nand2b_1 _3950_ (.Y(_0778_),
    .B(net1292),
    .A_N(net1283));
 sg13g2_nand4_1 _3951_ (.B(net1274),
    .C(net1225),
    .A(net1273),
    .Y(_0779_),
    .D(_0777_));
 sg13g2_o21ai_1 _3952_ (.B1(_0779_),
    .Y(_0010_),
    .A1(net709),
    .A2(_0775_));
 sg13g2_nand2_1 _3953_ (.Y(_0780_),
    .A(_0697_),
    .B(\main.state[4] ));
 sg13g2_a21oi_1 _3954_ (.A1(_0701_),
    .A2(_0780_),
    .Y(_0009_),
    .B1(_0006_));
 sg13g2_nand3_1 _3955_ (.B(\main.state[4] ),
    .C(net1225),
    .A(net1273),
    .Y(_0781_));
 sg13g2_nor2_1 _3956_ (.A(net1246),
    .B(_0781_),
    .Y(_0782_));
 sg13g2_nand3_1 _3957_ (.B(_0697_),
    .C(net1225),
    .A(net749),
    .Y(_0783_));
 sg13g2_o21ai_1 _3958_ (.B1(_0783_),
    .Y(_0008_),
    .A1(net1246),
    .A2(_0781_));
 sg13g2_nor2_1 _3959_ (.A(net702),
    .B(_0781_),
    .Y(_0784_));
 sg13g2_a21oi_1 _3960_ (.A1(net1273),
    .A2(net1292),
    .Y(_0785_),
    .B1(_0776_));
 sg13g2_a21o_1 _3961_ (.A2(_0784_),
    .A1(net1246),
    .B1(_0785_),
    .X(_0007_));
 sg13g2_mux2_1 _3962_ (.A0(net1),
    .A1(net1498),
    .S(net1345),
    .X(_0012_));
 sg13g2_mux2_1 _3963_ (.A0(net2),
    .A1(net577),
    .S(net1344),
    .X(_0014_));
 sg13g2_mux2_1 _3964_ (.A0(net3),
    .A1(net764),
    .S(net1345),
    .X(_0013_));
 sg13g2_nor2_1 _3965_ (.A(net1274),
    .B(net851),
    .Y(_0786_));
 sg13g2_o21ai_1 _3966_ (.B1(\main.state[6] ),
    .Y(_0787_),
    .A1(\main.read_command[0] ),
    .A2(_0769_));
 sg13g2_nand3b_1 _3967_ (.B(_0031_),
    .C(_0702_),
    .Y(_0788_),
    .A_N(net1274));
 sg13g2_nand4_1 _3968_ (.B(_0780_),
    .C(_0787_),
    .A(net1225),
    .Y(_0789_),
    .D(_0788_));
 sg13g2_a21oi_1 _3969_ (.A1(net1622),
    .A2(_0767_),
    .Y(_0790_),
    .B1(net1273));
 sg13g2_nor2_1 _3970_ (.A(_0789_),
    .B(_0790_),
    .Y(_0791_));
 sg13g2_nor2_2 _3971_ (.A(net1292),
    .B(net1283),
    .Y(_0792_));
 sg13g2_nor2b_1 _3972_ (.A(net1292),
    .B_N(net1283),
    .Y(_0793_));
 sg13g2_nand2b_1 _3973_ (.Y(_0794_),
    .B(net1283),
    .A_N(net1292));
 sg13g2_nor2_1 _3974_ (.A(_0770_),
    .B(_0792_),
    .Y(_0795_));
 sg13g2_o21ai_1 _3975_ (.B1(_0697_),
    .Y(_0796_),
    .A1(net1274),
    .A2(_0768_));
 sg13g2_nor3_1 _3976_ (.A(net1291),
    .B(_0789_),
    .C(_0796_),
    .Y(_0797_));
 sg13g2_a21oi_1 _3977_ (.A1(_0791_),
    .A2(_0795_),
    .Y(_0798_),
    .B1(_0797_));
 sg13g2_nand2_1 _3978_ (.Y(_0799_),
    .A(net1292),
    .B(_0789_));
 sg13g2_o21ai_1 _3979_ (.B1(_0799_),
    .Y(_0126_),
    .A1(_0786_),
    .A2(net1607));
 sg13g2_a21oi_1 _3980_ (.A1(net1283),
    .A2(_0796_),
    .Y(_0800_),
    .B1(_0786_));
 sg13g2_nor2_1 _3981_ (.A(_0789_),
    .B(_0800_),
    .Y(_0801_));
 sg13g2_nor2_1 _3982_ (.A(net1283),
    .B(_0791_),
    .Y(_0802_));
 sg13g2_nor2_1 _3983_ (.A(_0801_),
    .B(_0802_),
    .Y(_0127_));
 sg13g2_nor4_2 _3984_ (.A(\main.read_command[0] ),
    .B(\main.read_command[1] ),
    .C(_0031_),
    .Y(_0803_),
    .D(_0006_));
 sg13g2_nand2_2 _3985_ (.Y(_0804_),
    .A(\main.SPI_input_data_valid ),
    .B(_0803_));
 sg13g2_nor3_1 _3986_ (.A(net1296),
    .B(net1284),
    .C(_0032_),
    .Y(_0805_));
 sg13g2_and3_1 _3987_ (.X(_0806_),
    .A(\main.adder.in_valid ),
    .B(\main.adder.out_valid ),
    .C(_0765_));
 sg13g2_nand3_1 _3988_ (.B(\main.adder.out_valid ),
    .C(_0765_),
    .A(\main.adder.in_valid ),
    .Y(_0807_));
 sg13g2_a21oi_1 _3989_ (.A1(_0803_),
    .A2(_0805_),
    .Y(_0808_),
    .B1(net1217));
 sg13g2_o21ai_1 _3990_ (.B1(_0808_),
    .Y(_0809_),
    .A1(_0792_),
    .A2(_0804_));
 sg13g2_nand2_1 _3991_ (.Y(_0810_),
    .A(_0665_),
    .B(net1124));
 sg13g2_nand3_1 _3992_ (.B(_0665_),
    .C(net1124),
    .A(\main.register_id_result[1] ),
    .Y(_0811_));
 sg13g2_nand2_1 _3993_ (.Y(_0812_),
    .A(net1341),
    .B(_0811_));
 sg13g2_nor2_1 _3994_ (.A(net1300),
    .B(net1217),
    .Y(_0813_));
 sg13g2_o21ai_1 _3995_ (.B1(_0813_),
    .Y(_0814_),
    .A1(_0771_),
    .A2(_0804_));
 sg13g2_and2_1 _3996_ (.A(_0812_),
    .B(_0814_),
    .X(_0815_));
 sg13g2_nor2_1 _3997_ (.A(net1486),
    .B(net1105),
    .Y(_0816_));
 sg13g2_nand4_1 _3998_ (.B(net1294),
    .C(net1286),
    .A(\main.SPI_input_data[6] ),
    .Y(_0817_),
    .D(net1215));
 sg13g2_o21ai_1 _3999_ (.B1(_0817_),
    .Y(_0818_),
    .A1(_0743_),
    .A2(net1215));
 sg13g2_nand2_2 _4000_ (.Y(_0819_),
    .A(net1125),
    .B(_0818_));
 sg13g2_a21oi_1 _4001_ (.A1(net1105),
    .A2(_0819_),
    .Y(_0128_),
    .B1(_0816_));
 sg13g2_and2_1 _4002_ (.A(net1339),
    .B(_0808_),
    .X(_0820_));
 sg13g2_nand2b_1 _4003_ (.Y(_0821_),
    .B(net1124),
    .A_N(\main.register_id_result[1] ));
 sg13g2_nand2_2 _4004_ (.Y(_0822_),
    .A(_0810_),
    .B(_0821_));
 sg13g2_nor2_1 _4005_ (.A(_0820_),
    .B(_0822_),
    .Y(_0823_));
 sg13g2_nor2_1 _4006_ (.A(_0674_),
    .B(net1286),
    .Y(_0824_));
 sg13g2_a21o_1 _4007_ (.A2(_0824_),
    .A1(net1290),
    .B1(_0806_),
    .X(_0825_));
 sg13g2_o21ai_1 _4008_ (.B1(_0825_),
    .Y(_0826_),
    .A1(\main.adder.out[3] ),
    .A2(net1213));
 sg13g2_nand2b_2 _4009_ (.Y(_0827_),
    .B(net1125),
    .A_N(_0826_));
 sg13g2_nor2_1 _4010_ (.A(net1489),
    .B(net1104),
    .Y(_0828_));
 sg13g2_a21oi_1 _4011_ (.A1(net1104),
    .A2(_0827_),
    .Y(_0129_),
    .B1(_0828_));
 sg13g2_nor2_1 _4012_ (.A(_0673_),
    .B(net1288),
    .Y(_0829_));
 sg13g2_a21o_1 _4013_ (.A2(_0829_),
    .A1(net1290),
    .B1(_0806_),
    .X(_0830_));
 sg13g2_o21ai_1 _4014_ (.B1(_0830_),
    .Y(_0831_),
    .A1(\main.adder.out[4] ),
    .A2(net1209));
 sg13g2_nand2b_2 _4015_ (.Y(_0832_),
    .B(net1126),
    .A_N(_0831_));
 sg13g2_nor2_1 _4016_ (.A(net1514),
    .B(net1103),
    .Y(_0833_));
 sg13g2_a21oi_1 _4017_ (.A1(net1103),
    .A2(_0832_),
    .Y(_0130_),
    .B1(_0833_));
 sg13g2_o21ai_1 _4018_ (.B1(_0813_),
    .Y(_0834_),
    .A1(_0794_),
    .A2(_0804_));
 sg13g2_nor2b_1 _4019_ (.A(_0822_),
    .B_N(_0834_),
    .Y(_0835_));
 sg13g2_nor2_1 _4020_ (.A(net1026),
    .B(net1101),
    .Y(_0836_));
 sg13g2_nand3_1 _4021_ (.B(net1288),
    .C(net1290),
    .A(net1246),
    .Y(_0837_));
 sg13g2_nor2_1 _4022_ (.A(\main.adder.out[8] ),
    .B(net1214),
    .Y(_0838_));
 sg13g2_a21oi_2 _4023_ (.B1(_0838_),
    .Y(_0839_),
    .A2(_0837_),
    .A1(net1209));
 sg13g2_nand2_2 _4024_ (.Y(_0840_),
    .A(net1123),
    .B(_0839_));
 sg13g2_a21oi_1 _4025_ (.A1(net1101),
    .A2(_0840_),
    .Y(_0131_),
    .B1(_0836_));
 sg13g2_o21ai_1 _4026_ (.B1(net1341),
    .Y(_0841_),
    .A1(\main.register_id_result[0] ),
    .A2(_0821_));
 sg13g2_nand2b_1 _4027_ (.Y(_0842_),
    .B(_0841_),
    .A_N(_0820_));
 sg13g2_nor2b_1 _4028_ (.A(net1285),
    .B_N(\main.SPI_input_data[7] ),
    .Y(_0843_));
 sg13g2_a21o_1 _4029_ (.A2(_0843_),
    .A1(net1290),
    .B1(net1217),
    .X(_0844_));
 sg13g2_o21ai_1 _4030_ (.B1(_0844_),
    .Y(_0845_),
    .A1(\main.adder.out[7] ),
    .A2(net1211));
 sg13g2_nand2b_2 _4031_ (.Y(_0846_),
    .B(net1126),
    .A_N(_0845_));
 sg13g2_nand2_1 _4032_ (.Y(_0847_),
    .A(net839),
    .B(net1100));
 sg13g2_o21ai_1 _4033_ (.B1(_0847_),
    .Y(_0132_),
    .A1(net1100),
    .A2(_0846_));
 sg13g2_nor2_1 _4034_ (.A(_0671_),
    .B(net1285),
    .Y(_0848_));
 sg13g2_a21o_1 _4035_ (.A2(_0848_),
    .A1(net1290),
    .B1(net1217),
    .X(_0849_));
 sg13g2_o21ai_1 _4036_ (.B1(_0849_),
    .Y(_0850_),
    .A1(\main.adder.out[6] ),
    .A2(net1212));
 sg13g2_nand2b_2 _4037_ (.Y(_0851_),
    .B(net1126),
    .A_N(_0850_));
 sg13g2_nand2_1 _4038_ (.Y(_0852_),
    .A(net853),
    .B(net1100));
 sg13g2_o21ai_1 _4039_ (.B1(_0852_),
    .Y(_0133_),
    .A1(net1100),
    .A2(_0851_));
 sg13g2_o21ai_1 _4040_ (.B1(_0813_),
    .Y(_0853_),
    .A1(_0778_),
    .A2(_0804_));
 sg13g2_nand2_1 _4041_ (.Y(_0854_),
    .A(_0841_),
    .B(_0853_));
 sg13g2_nor2_1 _4042_ (.A(_0666_),
    .B(net1284),
    .Y(_0855_));
 sg13g2_nand3_1 _4043_ (.B(net1210),
    .C(_0855_),
    .A(net1296),
    .Y(_0856_));
 sg13g2_o21ai_1 _4044_ (.B1(_0856_),
    .Y(_0857_),
    .A1(_0729_),
    .A2(net1210));
 sg13g2_nand2_2 _4045_ (.Y(_0858_),
    .A(net1122),
    .B(_0857_));
 sg13g2_nand2_1 _4046_ (.Y(_0859_),
    .A(net815),
    .B(net1097));
 sg13g2_o21ai_1 _4047_ (.B1(_0859_),
    .Y(_0134_),
    .A1(net1096),
    .A2(_0858_));
 sg13g2_nor2_1 _4048_ (.A(_0672_),
    .B(net1287),
    .Y(_0860_));
 sg13g2_a21o_1 _4049_ (.A2(_0860_),
    .A1(net1289),
    .B1(net1217),
    .X(_0861_));
 sg13g2_o21ai_1 _4050_ (.B1(_0861_),
    .Y(_0862_),
    .A1(\main.adder.out[5] ),
    .A2(net1209));
 sg13g2_nand2b_2 _4051_ (.Y(_0863_),
    .B(net1126),
    .A_N(_0862_));
 sg13g2_nand2_1 _4052_ (.Y(_0864_),
    .A(net821),
    .B(net1099));
 sg13g2_o21ai_1 _4053_ (.B1(_0864_),
    .Y(_0135_),
    .A1(net1099),
    .A2(_0863_));
 sg13g2_nand2_1 _4054_ (.Y(_0865_),
    .A(net970),
    .B(net1099));
 sg13g2_o21ai_1 _4055_ (.B1(_0865_),
    .Y(_0136_),
    .A1(_0832_),
    .A2(net1099));
 sg13g2_nand2_1 _4056_ (.Y(_0866_),
    .A(_0834_),
    .B(_0841_));
 sg13g2_nand3_1 _4057_ (.B(net1285),
    .C(net1289),
    .A(\main.SPI_input_data[7] ),
    .Y(_0867_));
 sg13g2_nor2_1 _4058_ (.A(\main.adder.out[15] ),
    .B(net1214),
    .Y(_0868_));
 sg13g2_a21oi_2 _4059_ (.B1(_0868_),
    .Y(_0869_),
    .A2(_0867_),
    .A1(net1214));
 sg13g2_nand2_2 _4060_ (.Y(_0870_),
    .A(net1122),
    .B(_0869_));
 sg13g2_nand2_1 _4061_ (.Y(_0871_),
    .A(net878),
    .B(net1094));
 sg13g2_o21ai_1 _4062_ (.B1(_0871_),
    .Y(_0137_),
    .A1(net1094),
    .A2(_0870_));
 sg13g2_nand2_1 _4063_ (.Y(_0872_),
    .A(net932),
    .B(net1100));
 sg13g2_o21ai_1 _4064_ (.B1(_0872_),
    .Y(_0138_),
    .A1(_0827_),
    .A2(net1100));
 sg13g2_nand3_1 _4065_ (.B(net1284),
    .C(net1291),
    .A(\main.SPI_input_data[1] ),
    .Y(_0873_));
 sg13g2_nor2_1 _4066_ (.A(\main.adder.out[9] ),
    .B(net1216),
    .Y(_0874_));
 sg13g2_a21oi_2 _4067_ (.B1(_0874_),
    .Y(_0875_),
    .A2(_0873_),
    .A1(net1210));
 sg13g2_nand2_2 _4068_ (.Y(_0876_),
    .A(net1122),
    .B(_0875_));
 sg13g2_nand2_1 _4069_ (.Y(_0877_),
    .A(net862),
    .B(net1095));
 sg13g2_o21ai_1 _4070_ (.B1(_0877_),
    .Y(_0139_),
    .A1(net1095),
    .A2(_0876_));
 sg13g2_nand2_1 _4071_ (.Y(_0878_),
    .A(net915),
    .B(net1094));
 sg13g2_o21ai_1 _4072_ (.B1(_0878_),
    .Y(_0140_),
    .A1(_0840_),
    .A2(net1094));
 sg13g2_nand3_1 _4073_ (.B(net1214),
    .C(_0843_),
    .A(net1293),
    .Y(_0879_));
 sg13g2_o21ai_1 _4074_ (.B1(_0879_),
    .Y(_0880_),
    .A1(_0736_),
    .A2(net1214));
 sg13g2_nand2_2 _4075_ (.Y(_0881_),
    .A(net1124),
    .B(_0880_));
 sg13g2_nand2_1 _4076_ (.Y(_0882_),
    .A(net855),
    .B(net1098));
 sg13g2_o21ai_1 _4077_ (.B1(_0882_),
    .Y(_0141_),
    .A1(net1098),
    .A2(_0881_));
 sg13g2_nand3_1 _4078_ (.B(net1213),
    .C(_0848_),
    .A(net1293),
    .Y(_0883_));
 sg13g2_o21ai_1 _4079_ (.B1(_0883_),
    .Y(_0884_),
    .A1(_0735_),
    .A2(net1211));
 sg13g2_nand2_2 _4080_ (.Y(_0885_),
    .A(net1122),
    .B(_0884_));
 sg13g2_nand2_1 _4081_ (.Y(_0886_),
    .A(net840),
    .B(net1098));
 sg13g2_o21ai_1 _4082_ (.B1(_0886_),
    .Y(_0142_),
    .A1(net1098),
    .A2(_0885_));
 sg13g2_nand3_1 _4083_ (.B(net1287),
    .C(net1289),
    .A(\main.SPI_input_data[4] ),
    .Y(_0887_));
 sg13g2_nor2_1 _4084_ (.A(net841),
    .B(net1211),
    .Y(_0888_));
 sg13g2_a21oi_2 _4085_ (.B1(_0888_),
    .Y(_0889_),
    .A2(_0887_),
    .A1(net1212));
 sg13g2_nand2_2 _4086_ (.Y(_0890_),
    .A(net1122),
    .B(_0889_));
 sg13g2_nand2_1 _4087_ (.Y(_0891_),
    .A(net812),
    .B(net1095));
 sg13g2_o21ai_1 _4088_ (.B1(_0891_),
    .Y(_0143_),
    .A1(net1095),
    .A2(_0890_));
 sg13g2_nand3_1 _4089_ (.B(net1285),
    .C(net1289),
    .A(net1623),
    .Y(_0892_));
 sg13g2_nor2_1 _4090_ (.A(\main.adder.out[11] ),
    .B(net1214),
    .Y(_0893_));
 sg13g2_a21oi_2 _4091_ (.B1(_0893_),
    .Y(_0894_),
    .A2(_0892_),
    .A1(net1211));
 sg13g2_nand2_2 _4092_ (.Y(_0895_),
    .A(net1123),
    .B(_0894_));
 sg13g2_nand2_1 _4093_ (.Y(_0896_),
    .A(net832),
    .B(net1094));
 sg13g2_o21ai_1 _4094_ (.B1(_0896_),
    .Y(_0144_),
    .A1(net1094),
    .A2(_0895_));
 sg13g2_nand3_1 _4095_ (.B(net1288),
    .C(net1289),
    .A(\main.SPI_input_data[2] ),
    .Y(_0897_));
 sg13g2_nor2_1 _4096_ (.A(net796),
    .B(net1212),
    .Y(_0898_));
 sg13g2_a21oi_2 _4097_ (.B1(_0898_),
    .Y(_0899_),
    .A2(_0897_),
    .A1(net1209));
 sg13g2_nand2_2 _4098_ (.Y(_0900_),
    .A(net1123),
    .B(_0899_));
 sg13g2_nand2_1 _4099_ (.Y(_0901_),
    .A(net912),
    .B(net1095));
 sg13g2_o21ai_1 _4100_ (.B1(_0901_),
    .Y(_0145_),
    .A1(net1095),
    .A2(_0900_));
 sg13g2_nand3_1 _4101_ (.B(net1212),
    .C(_0860_),
    .A(net1294),
    .Y(_0902_));
 sg13g2_o21ai_1 _4102_ (.B1(_0902_),
    .Y(_0903_),
    .A1(_0734_),
    .A2(net1212));
 sg13g2_nand2_2 _4103_ (.Y(_0904_),
    .A(net1123),
    .B(_0903_));
 sg13g2_nand2_1 _4104_ (.Y(_0905_),
    .A(net848),
    .B(net1097));
 sg13g2_o21ai_1 _4105_ (.B1(_0905_),
    .Y(_0146_),
    .A1(net1096),
    .A2(_0904_));
 sg13g2_nand3_1 _4106_ (.B(net1210),
    .C(_0829_),
    .A(net1295),
    .Y(_0906_));
 sg13g2_o21ai_1 _4107_ (.B1(_0906_),
    .Y(_0907_),
    .A1(_0733_),
    .A2(net1209));
 sg13g2_nand2_2 _4108_ (.Y(_0908_),
    .A(net1123),
    .B(_0907_));
 sg13g2_nand2_1 _4109_ (.Y(_0909_),
    .A(net811),
    .B(net1096));
 sg13g2_o21ai_1 _4110_ (.B1(_0909_),
    .Y(_0147_),
    .A1(net1096),
    .A2(_0908_));
 sg13g2_nand3_1 _4111_ (.B(net1213),
    .C(_0824_),
    .A(net1293),
    .Y(_0910_));
 sg13g2_o21ai_1 _4112_ (.B1(_0910_),
    .Y(_0911_),
    .A1(_0732_),
    .A2(net1211));
 sg13g2_nand2_2 _4113_ (.Y(_0912_),
    .A(net1124),
    .B(_0911_));
 sg13g2_nand2_1 _4114_ (.Y(_0913_),
    .A(net845),
    .B(net1097));
 sg13g2_o21ai_1 _4115_ (.B1(_0913_),
    .Y(_0148_),
    .A1(net1097),
    .A2(_0912_));
 sg13g2_nor2_1 _4116_ (.A(_0675_),
    .B(net1287),
    .Y(_0914_));
 sg13g2_nand3_1 _4117_ (.B(net1212),
    .C(_0914_),
    .A(net1294),
    .Y(_0915_));
 sg13g2_o21ai_1 _4118_ (.B1(_0915_),
    .Y(_0916_),
    .A1(_0731_),
    .A2(net1211));
 sg13g2_nand2_2 _4119_ (.Y(_0917_),
    .A(net1122),
    .B(_0916_));
 sg13g2_nand2_1 _4120_ (.Y(_0918_),
    .A(net925),
    .B(net1096));
 sg13g2_o21ai_1 _4121_ (.B1(_0918_),
    .Y(_0149_),
    .A1(net1096),
    .A2(_0917_));
 sg13g2_nor2_1 _4122_ (.A(_0664_),
    .B(net1288),
    .Y(_0919_));
 sg13g2_nand3_1 _4123_ (.B(net1209),
    .C(_0919_),
    .A(net1295),
    .Y(_0920_));
 sg13g2_o21ai_1 _4124_ (.B1(_0920_),
    .Y(_0921_),
    .A1(_0730_),
    .A2(net1209));
 sg13g2_nand2_2 _4125_ (.Y(_0922_),
    .A(net1122),
    .B(_0921_));
 sg13g2_nand2_1 _4126_ (.Y(_0923_),
    .A(net849),
    .B(net1096));
 sg13g2_o21ai_1 _4127_ (.B1(_0923_),
    .Y(_0150_),
    .A1(net1096),
    .A2(_0922_));
 sg13g2_a21o_1 _4128_ (.A2(_0914_),
    .A1(net1289),
    .B1(net1217),
    .X(_0924_));
 sg13g2_o21ai_1 _4129_ (.B1(_0924_),
    .Y(_0925_),
    .A1(\main.adder.out[2] ),
    .A2(net1213));
 sg13g2_nand2b_2 _4130_ (.Y(_0926_),
    .B(net1125),
    .A_N(_0925_));
 sg13g2_nand2_1 _4131_ (.Y(_0927_),
    .A(net846),
    .B(net1100));
 sg13g2_o21ai_1 _4132_ (.B1(_0927_),
    .Y(_0151_),
    .A1(net1100),
    .A2(_0926_));
 sg13g2_a21o_1 _4133_ (.A2(_0855_),
    .A1(net1291),
    .B1(net1217),
    .X(_0928_));
 sg13g2_o21ai_1 _4134_ (.B1(_0928_),
    .Y(_0929_),
    .A1(\main.adder.out[0] ),
    .A2(net1210));
 sg13g2_nand2b_2 _4135_ (.Y(_0930_),
    .B(net1124),
    .A_N(_0929_));
 sg13g2_nand2_1 _4136_ (.Y(_0931_),
    .A(net882),
    .B(net1099));
 sg13g2_o21ai_1 _4137_ (.B1(_0931_),
    .Y(_0152_),
    .A1(net1099),
    .A2(_0930_));
 sg13g2_nand3_1 _4138_ (.B(net1287),
    .C(net1289),
    .A(net1624),
    .Y(_0932_));
 sg13g2_nor2_1 _4139_ (.A(\main.adder.out[13] ),
    .B(net1211),
    .Y(_0933_));
 sg13g2_a21oi_2 _4140_ (.B1(_0933_),
    .Y(_0934_),
    .A2(_0932_),
    .A1(net1212));
 sg13g2_nand2_2 _4141_ (.Y(_0935_),
    .A(net1122),
    .B(_0934_));
 sg13g2_nand2_1 _4142_ (.Y(_0936_),
    .A(net827),
    .B(net1095));
 sg13g2_o21ai_1 _4143_ (.B1(_0936_),
    .Y(_0153_),
    .A1(net1095),
    .A2(_0935_));
 sg13g2_nand3_1 _4144_ (.B(net1285),
    .C(net1289),
    .A(\main.SPI_input_data[6] ),
    .Y(_0937_));
 sg13g2_nor2_1 _4145_ (.A(\main.adder.out[14] ),
    .B(net1214),
    .Y(_0938_));
 sg13g2_a21oi_2 _4146_ (.B1(_0938_),
    .Y(_0939_),
    .A2(_0937_),
    .A1(net1211));
 sg13g2_nand2_2 _4147_ (.Y(_0940_),
    .A(net1123),
    .B(_0939_));
 sg13g2_nand2_1 _4148_ (.Y(_0941_),
    .A(net817),
    .B(net1094));
 sg13g2_o21ai_1 _4149_ (.B1(_0941_),
    .Y(_0154_),
    .A1(net1094),
    .A2(_0940_));
 sg13g2_nand2_1 _4150_ (.Y(_0942_),
    .A(_0814_),
    .B(_0841_));
 sg13g2_nand4_1 _4151_ (.B(net1295),
    .C(net1288),
    .A(\main.SPI_input_data[1] ),
    .Y(_0943_),
    .D(net1210));
 sg13g2_o21ai_1 _4152_ (.B1(_0943_),
    .Y(_0944_),
    .A1(_0738_),
    .A2(net1210));
 sg13g2_nand2_2 _4153_ (.Y(_0945_),
    .A(net1126),
    .B(_0944_));
 sg13g2_nand2_1 _4154_ (.Y(_0946_),
    .A(net880),
    .B(net1093));
 sg13g2_o21ai_1 _4155_ (.B1(_0946_),
    .Y(_0155_),
    .A1(net1093),
    .A2(_0945_));
 sg13g2_nand4_1 _4156_ (.B(net1293),
    .C(net1285),
    .A(net1627),
    .Y(_0947_),
    .D(net1215));
 sg13g2_o21ai_1 _4157_ (.B1(_0947_),
    .Y(_0948_),
    .A1(_0739_),
    .A2(net1216));
 sg13g2_nand2_2 _4158_ (.Y(_0949_),
    .A(net1126),
    .B(_0948_));
 sg13g2_nand2_1 _4159_ (.Y(_0950_),
    .A(net854),
    .B(net1092));
 sg13g2_o21ai_1 _4160_ (.B1(_0950_),
    .Y(_0156_),
    .A1(net1092),
    .A2(_0949_));
 sg13g2_nand4_1 _4161_ (.B(net1293),
    .C(net1286),
    .A(net1623),
    .Y(_0951_),
    .D(net1215));
 sg13g2_o21ai_1 _4162_ (.B1(_0951_),
    .Y(_0952_),
    .A1(_0740_),
    .A2(net1215));
 sg13g2_nand2_2 _4163_ (.Y(_0953_),
    .A(net1125),
    .B(_0952_));
 sg13g2_nand2_1 _4164_ (.Y(_0954_),
    .A(net895),
    .B(net1093));
 sg13g2_o21ai_1 _4165_ (.B1(_0954_),
    .Y(_0157_),
    .A1(_0942_),
    .A2(_0953_));
 sg13g2_nand4_1 _4166_ (.B(net1293),
    .C(net1286),
    .A(net1625),
    .Y(_0955_),
    .D(net1215));
 sg13g2_o21ai_1 _4167_ (.B1(_0955_),
    .Y(_0956_),
    .A1(_0741_),
    .A2(net1216));
 sg13g2_nand2_2 _4168_ (.Y(_0957_),
    .A(net1125),
    .B(_0956_));
 sg13g2_nand2_1 _4169_ (.Y(_0958_),
    .A(net803),
    .B(net1093));
 sg13g2_o21ai_1 _4170_ (.B1(_0958_),
    .Y(_0158_),
    .A1(net1093),
    .A2(_0957_));
 sg13g2_nand4_1 _4171_ (.B(net1293),
    .C(net1285),
    .A(\main.SPI_input_data[5] ),
    .Y(_0959_),
    .D(net1215));
 sg13g2_o21ai_1 _4172_ (.B1(_0959_),
    .Y(_0960_),
    .A1(_0742_),
    .A2(net1215));
 sg13g2_nand2_2 _4173_ (.Y(_0961_),
    .A(net1125),
    .B(_0960_));
 sg13g2_nand2_1 _4174_ (.Y(_0962_),
    .A(net948),
    .B(net1092));
 sg13g2_o21ai_1 _4175_ (.B1(_0962_),
    .Y(_0159_),
    .A1(net1092),
    .A2(_0961_));
 sg13g2_nand2_1 _4176_ (.Y(_0963_),
    .A(net890),
    .B(net1092));
 sg13g2_o21ai_1 _4177_ (.B1(_0963_),
    .Y(_0160_),
    .A1(_0819_),
    .A2(net1092));
 sg13g2_nand4_1 _4178_ (.B(net1293),
    .C(net1285),
    .A(\main.SPI_input_data[7] ),
    .Y(_0964_),
    .D(net1214));
 sg13g2_o21ai_1 _4179_ (.B1(_0964_),
    .Y(_0965_),
    .A1(_0744_),
    .A2(net1216));
 sg13g2_nand2_2 _4180_ (.Y(_0966_),
    .A(net1125),
    .B(_0965_));
 sg13g2_nand2_1 _4181_ (.Y(_0967_),
    .A(net871),
    .B(net1092));
 sg13g2_o21ai_1 _4182_ (.B1(_0967_),
    .Y(_0161_),
    .A1(net1092),
    .A2(_0966_));
 sg13g2_a21o_1 _4183_ (.A2(_0919_),
    .A1(net1290),
    .B1(net1217),
    .X(_0968_));
 sg13g2_o21ai_1 _4184_ (.B1(_0968_),
    .Y(_0969_),
    .A1(\main.adder.out[1] ),
    .A2(net1209));
 sg13g2_nand2b_2 _4185_ (.Y(_0970_),
    .B(net1126),
    .A_N(_0969_));
 sg13g2_nand2_1 _4186_ (.Y(_0971_),
    .A(net996),
    .B(net1099));
 sg13g2_o21ai_1 _4187_ (.B1(_0971_),
    .Y(_0162_),
    .A1(net1099),
    .A2(_0970_));
 sg13g2_o21ai_1 _4188_ (.B1(net1341),
    .Y(_0972_),
    .A1(_0665_),
    .A2(_0821_));
 sg13g2_nor2b_1 _4189_ (.A(_0820_),
    .B_N(_0972_),
    .Y(_0973_));
 sg13g2_nor2_1 _4190_ (.A(net892),
    .B(net1090),
    .Y(_0974_));
 sg13g2_a21oi_1 _4191_ (.A1(_0970_),
    .A2(net1090),
    .Y(_0163_),
    .B1(_0974_));
 sg13g2_nor2_1 _4192_ (.A(net992),
    .B(net1091),
    .Y(_0975_));
 sg13g2_a21oi_1 _4193_ (.A1(_0926_),
    .A2(net1091),
    .Y(_0164_),
    .B1(_0975_));
 sg13g2_nor2_1 _4194_ (.A(net734),
    .B(net1091),
    .Y(_0976_));
 sg13g2_a21oi_1 _4195_ (.A1(_0827_),
    .A2(net1091),
    .Y(_0165_),
    .B1(_0976_));
 sg13g2_nor2_1 _4196_ (.A(net1433),
    .B(net1090),
    .Y(_0977_));
 sg13g2_a21oi_1 _4197_ (.A1(_0832_),
    .A2(net1090),
    .Y(_0166_),
    .B1(_0977_));
 sg13g2_nor2_1 _4198_ (.A(net978),
    .B(net1090),
    .Y(_0978_));
 sg13g2_a21oi_1 _4199_ (.A1(_0863_),
    .A2(net1090),
    .Y(_0167_),
    .B1(_0978_));
 sg13g2_nor2_1 _4200_ (.A(net991),
    .B(net1091),
    .Y(_0979_));
 sg13g2_a21oi_1 _4201_ (.A1(_0851_),
    .A2(net1091),
    .Y(_0168_),
    .B1(_0979_));
 sg13g2_nor2_1 _4202_ (.A(net1012),
    .B(net1091),
    .Y(_0980_));
 sg13g2_a21oi_1 _4203_ (.A1(_0846_),
    .A2(net1091),
    .Y(_0169_),
    .B1(_0980_));
 sg13g2_and2_1 _4204_ (.A(_0834_),
    .B(_0972_),
    .X(_0981_));
 sg13g2_nor2_1 _4205_ (.A(net1018),
    .B(net1088),
    .Y(_0982_));
 sg13g2_a21oi_1 _4206_ (.A1(_0840_),
    .A2(net1088),
    .Y(_0170_),
    .B1(_0982_));
 sg13g2_nor2_1 _4207_ (.A(net1494),
    .B(net1089),
    .Y(_0983_));
 sg13g2_a21oi_1 _4208_ (.A1(_0876_),
    .A2(net1089),
    .Y(_0171_),
    .B1(_0983_));
 sg13g2_nor2_1 _4209_ (.A(net1413),
    .B(net1089),
    .Y(_0984_));
 sg13g2_a21oi_1 _4210_ (.A1(_0900_),
    .A2(net1089),
    .Y(_0172_),
    .B1(_0984_));
 sg13g2_nor2_1 _4211_ (.A(net957),
    .B(net1088),
    .Y(_0985_));
 sg13g2_a21oi_1 _4212_ (.A1(_0895_),
    .A2(net1088),
    .Y(_0173_),
    .B1(_0985_));
 sg13g2_nor2_1 _4213_ (.A(net1447),
    .B(net1089),
    .Y(_0986_));
 sg13g2_a21oi_1 _4214_ (.A1(_0890_),
    .A2(net1089),
    .Y(_0174_),
    .B1(_0986_));
 sg13g2_nor2_1 _4215_ (.A(net1008),
    .B(net1089),
    .Y(_0987_));
 sg13g2_a21oi_1 _4216_ (.A1(_0935_),
    .A2(net1089),
    .Y(_0175_),
    .B1(_0987_));
 sg13g2_nor2_1 _4217_ (.A(net1511),
    .B(net1088),
    .Y(_0988_));
 sg13g2_a21oi_1 _4218_ (.A1(_0940_),
    .A2(net1088),
    .Y(_0176_),
    .B1(_0988_));
 sg13g2_nor2_1 _4219_ (.A(net1032),
    .B(net1088),
    .Y(_0989_));
 sg13g2_a21oi_1 _4220_ (.A1(_0870_),
    .A2(net1088),
    .Y(_0177_),
    .B1(_0989_));
 sg13g2_and2_1 _4221_ (.A(_0853_),
    .B(_0972_),
    .X(_0990_));
 sg13g2_nor2_1 _4222_ (.A(net1421),
    .B(net1085),
    .Y(_0991_));
 sg13g2_a21oi_1 _4223_ (.A1(_0858_),
    .A2(net1085),
    .Y(_0178_),
    .B1(_0991_));
 sg13g2_nor2_1 _4224_ (.A(net1408),
    .B(net1085),
    .Y(_0992_));
 sg13g2_a21oi_1 _4225_ (.A1(_0922_),
    .A2(net1085),
    .Y(_0179_),
    .B1(_0992_));
 sg13g2_nor2_1 _4226_ (.A(net972),
    .B(net1086),
    .Y(_0993_));
 sg13g2_a21oi_1 _4227_ (.A1(_0917_),
    .A2(net1085),
    .Y(_0180_),
    .B1(_0993_));
 sg13g2_nor2_1 _4228_ (.A(net1434),
    .B(net1087),
    .Y(_0994_));
 sg13g2_a21oi_1 _4229_ (.A1(_0912_),
    .A2(net1087),
    .Y(_0181_),
    .B1(_0994_));
 sg13g2_nor2_1 _4230_ (.A(net986),
    .B(net1085),
    .Y(_0995_));
 sg13g2_a21oi_1 _4231_ (.A1(_0908_),
    .A2(net1085),
    .Y(_0182_),
    .B1(_0995_));
 sg13g2_nor2_1 _4232_ (.A(net773),
    .B(net1087),
    .Y(_0996_));
 sg13g2_a21oi_1 _4233_ (.A1(_0904_),
    .A2(net1085),
    .Y(_0183_),
    .B1(_0996_));
 sg13g2_nor2_1 _4234_ (.A(net1035),
    .B(net1086),
    .Y(_0997_));
 sg13g2_a21oi_1 _4235_ (.A1(_0885_),
    .A2(net1086),
    .Y(_0184_),
    .B1(_0997_));
 sg13g2_nor2_1 _4236_ (.A(net1448),
    .B(net1087),
    .Y(_0998_));
 sg13g2_a21oi_1 _4237_ (.A1(_0881_),
    .A2(net1087),
    .Y(_0185_),
    .B1(_0998_));
 sg13g2_and2_1 _4238_ (.A(_0814_),
    .B(_0972_),
    .X(_0999_));
 sg13g2_nor2_1 _4239_ (.A(net1439),
    .B(net1084),
    .Y(_1000_));
 sg13g2_nand4_1 _4240_ (.B(net1294),
    .C(net1287),
    .A(net1246),
    .Y(_1001_),
    .D(net1213));
 sg13g2_o21ai_1 _4241_ (.B1(_1001_),
    .Y(_1002_),
    .A1(_0737_),
    .A2(net1213));
 sg13g2_nand2_2 _4242_ (.Y(_1003_),
    .A(net1125),
    .B(_1002_));
 sg13g2_a21oi_1 _4243_ (.A1(net1084),
    .A2(_1003_),
    .Y(_0186_),
    .B1(_1000_));
 sg13g2_nor2_1 _4244_ (.A(net1427),
    .B(net1084),
    .Y(_1004_));
 sg13g2_a21oi_1 _4245_ (.A1(_0945_),
    .A2(net1084),
    .Y(_0187_),
    .B1(_1004_));
 sg13g2_nor2_1 _4246_ (.A(net1462),
    .B(net1083),
    .Y(_1005_));
 sg13g2_a21oi_1 _4247_ (.A1(_0949_),
    .A2(net1083),
    .Y(_0188_),
    .B1(_1005_));
 sg13g2_nor2_1 _4248_ (.A(net1446),
    .B(net1084),
    .Y(_1006_));
 sg13g2_a21oi_1 _4249_ (.A1(_0953_),
    .A2(_0999_),
    .Y(_0189_),
    .B1(_1006_));
 sg13g2_nor2_1 _4250_ (.A(net1036),
    .B(net1084),
    .Y(_1007_));
 sg13g2_a21oi_1 _4251_ (.A1(_0957_),
    .A2(net1084),
    .Y(_0190_),
    .B1(_1007_));
 sg13g2_nor2_1 _4252_ (.A(net973),
    .B(net1083),
    .Y(_1008_));
 sg13g2_a21oi_1 _4253_ (.A1(_0961_),
    .A2(net1083),
    .Y(_0191_),
    .B1(_1008_));
 sg13g2_nor2_1 _4254_ (.A(net1019),
    .B(net1083),
    .Y(_1009_));
 sg13g2_a21oi_1 _4255_ (.A1(_0819_),
    .A2(net1083),
    .Y(_0192_),
    .B1(_1009_));
 sg13g2_nor2_1 _4256_ (.A(net1013),
    .B(net1083),
    .Y(_1010_));
 sg13g2_a21oi_1 _4257_ (.A1(_0966_),
    .A2(net1083),
    .Y(_0193_),
    .B1(_1010_));
 sg13g2_a21oi_1 _4258_ (.A1(net1341),
    .A2(_0811_),
    .Y(_1011_),
    .B1(_0820_));
 sg13g2_nor2_1 _4259_ (.A(net1515),
    .B(net1110),
    .Y(_1012_));
 sg13g2_a21oi_1 _4260_ (.A1(_0970_),
    .A2(net1110),
    .Y(_0194_),
    .B1(_1012_));
 sg13g2_nor2_1 _4261_ (.A(net971),
    .B(net1111),
    .Y(_1013_));
 sg13g2_a21oi_1 _4262_ (.A1(_0926_),
    .A2(net1111),
    .Y(_0195_),
    .B1(_1013_));
 sg13g2_nor2_1 _4263_ (.A(net977),
    .B(net1111),
    .Y(_1014_));
 sg13g2_a21oi_1 _4264_ (.A1(_0827_),
    .A2(net1111),
    .Y(_0196_),
    .B1(_1014_));
 sg13g2_nor2_1 _4265_ (.A(net1466),
    .B(net1110),
    .Y(_1015_));
 sg13g2_a21oi_1 _4266_ (.A1(_0832_),
    .A2(net1110),
    .Y(_0197_),
    .B1(_1015_));
 sg13g2_nor2_1 _4267_ (.A(net990),
    .B(net1110),
    .Y(_1016_));
 sg13g2_a21oi_1 _4268_ (.A1(_0863_),
    .A2(net1110),
    .Y(_0198_),
    .B1(_1016_));
 sg13g2_nor2_1 _4269_ (.A(net1049),
    .B(net1111),
    .Y(_1017_));
 sg13g2_a21oi_1 _4270_ (.A1(_0851_),
    .A2(net1111),
    .Y(_0199_),
    .B1(_1017_));
 sg13g2_nor2_1 _4271_ (.A(net1024),
    .B(net1111),
    .Y(_1018_));
 sg13g2_a21oi_1 _4272_ (.A1(_0846_),
    .A2(net1111),
    .Y(_0200_),
    .B1(_1018_));
 sg13g2_and2_1 _4273_ (.A(_0812_),
    .B(_0834_),
    .X(_1019_));
 sg13g2_nor2_1 _4274_ (.A(net1431),
    .B(net1081),
    .Y(_1020_));
 sg13g2_a21oi_1 _4275_ (.A1(_0840_),
    .A2(net1081),
    .Y(_0201_),
    .B1(_1020_));
 sg13g2_nor2_1 _4276_ (.A(net1524),
    .B(net1082),
    .Y(_1021_));
 sg13g2_a21oi_1 _4277_ (.A1(_0876_),
    .A2(net1082),
    .Y(_0202_),
    .B1(_1021_));
 sg13g2_nor2_1 _4278_ (.A(net1417),
    .B(net1082),
    .Y(_1022_));
 sg13g2_a21oi_1 _4279_ (.A1(_0900_),
    .A2(net1082),
    .Y(_0203_),
    .B1(_1022_));
 sg13g2_nor2_1 _4280_ (.A(net1027),
    .B(net1081),
    .Y(_1023_));
 sg13g2_a21oi_1 _4281_ (.A1(_0895_),
    .A2(net1081),
    .Y(_0204_),
    .B1(_1023_));
 sg13g2_nor2_1 _4282_ (.A(net1039),
    .B(net1082),
    .Y(_1024_));
 sg13g2_a21oi_1 _4283_ (.A1(_0890_),
    .A2(net1082),
    .Y(_0205_),
    .B1(_1024_));
 sg13g2_nor2_1 _4284_ (.A(net1457),
    .B(net1082),
    .Y(_1025_));
 sg13g2_a21oi_1 _4285_ (.A1(_0935_),
    .A2(net1082),
    .Y(_0206_),
    .B1(_1025_));
 sg13g2_nor2_1 _4286_ (.A(net1491),
    .B(net1081),
    .Y(_1026_));
 sg13g2_a21oi_1 _4287_ (.A1(_0940_),
    .A2(net1081),
    .Y(_0207_),
    .B1(_1026_));
 sg13g2_nor2_1 _4288_ (.A(net1440),
    .B(net1081),
    .Y(_1027_));
 sg13g2_a21oi_1 _4289_ (.A1(_0870_),
    .A2(net1081),
    .Y(_0208_),
    .B1(_1027_));
 sg13g2_and2_1 _4290_ (.A(_0812_),
    .B(_0853_),
    .X(_1028_));
 sg13g2_nor2_1 _4291_ (.A(net1044),
    .B(net1078),
    .Y(_1029_));
 sg13g2_a21oi_1 _4292_ (.A1(_0858_),
    .A2(net1078),
    .Y(_0209_),
    .B1(_1029_));
 sg13g2_nor2_1 _4293_ (.A(net1437),
    .B(net1078),
    .Y(_1030_));
 sg13g2_a21oi_1 _4294_ (.A1(_0922_),
    .A2(net1078),
    .Y(_0210_),
    .B1(_1030_));
 sg13g2_nor2_1 _4295_ (.A(net1438),
    .B(net1078),
    .Y(_1031_));
 sg13g2_a21oi_1 _4296_ (.A1(_0917_),
    .A2(net1078),
    .Y(_0211_),
    .B1(_1031_));
 sg13g2_nor2_1 _4297_ (.A(net1501),
    .B(net1079),
    .Y(_1032_));
 sg13g2_a21oi_1 _4298_ (.A1(_0912_),
    .A2(net1079),
    .Y(_0212_),
    .B1(_1032_));
 sg13g2_nor2_1 _4299_ (.A(net1432),
    .B(net1078),
    .Y(_1033_));
 sg13g2_a21oi_1 _4300_ (.A1(_0908_),
    .A2(net1078),
    .Y(_0213_),
    .B1(_1033_));
 sg13g2_nor2_1 _4301_ (.A(net1043),
    .B(net1079),
    .Y(_1034_));
 sg13g2_a21oi_1 _4302_ (.A1(_0904_),
    .A2(net1079),
    .Y(_0214_),
    .B1(_1034_));
 sg13g2_nor2_1 _4303_ (.A(net1040),
    .B(net1079),
    .Y(_1035_));
 sg13g2_a21oi_1 _4304_ (.A1(_0885_),
    .A2(net1080),
    .Y(_0215_),
    .B1(_1035_));
 sg13g2_nor2_1 _4305_ (.A(net1042),
    .B(net1080),
    .Y(_1036_));
 sg13g2_a21oi_1 _4306_ (.A1(_0881_),
    .A2(net1080),
    .Y(_0216_),
    .B1(_1036_));
 sg13g2_nor2_1 _4307_ (.A(net1449),
    .B(net1106),
    .Y(_1037_));
 sg13g2_a21oi_1 _4308_ (.A1(net1106),
    .A2(_1003_),
    .Y(_0217_),
    .B1(_1037_));
 sg13g2_nor2_1 _4309_ (.A(net1002),
    .B(net1106),
    .Y(_1038_));
 sg13g2_a21oi_1 _4310_ (.A1(net1106),
    .A2(_0945_),
    .Y(_0218_),
    .B1(_1038_));
 sg13g2_nor2_1 _4311_ (.A(net1025),
    .B(net1105),
    .Y(_1039_));
 sg13g2_a21oi_1 _4312_ (.A1(net1105),
    .A2(_0949_),
    .Y(_0219_),
    .B1(_1039_));
 sg13g2_nor2_1 _4313_ (.A(net1017),
    .B(net1106),
    .Y(_1040_));
 sg13g2_a21oi_1 _4314_ (.A1(_0815_),
    .A2(_0953_),
    .Y(_0220_),
    .B1(_1040_));
 sg13g2_nor2_1 _4315_ (.A(net1010),
    .B(net1106),
    .Y(_1041_));
 sg13g2_a21oi_1 _4316_ (.A1(net1106),
    .A2(_0957_),
    .Y(_0221_),
    .B1(_1041_));
 sg13g2_nor2_1 _4317_ (.A(net1458),
    .B(net1105),
    .Y(_1042_));
 sg13g2_a21oi_1 _4318_ (.A1(net1105),
    .A2(_0961_),
    .Y(_0222_),
    .B1(_1042_));
 sg13g2_nor2b_2 _4319_ (.A(_0822_),
    .B_N(_0814_),
    .Y(_1043_));
 sg13g2_nor2_1 _4320_ (.A(net1442),
    .B(net1076),
    .Y(_1044_));
 sg13g2_a21oi_1 _4321_ (.A1(_0966_),
    .A2(net1076),
    .Y(_0223_),
    .B1(_1044_));
 sg13g2_nor2_1 _4322_ (.A(net1015),
    .B(net1076),
    .Y(_1045_));
 sg13g2_a21oi_1 _4323_ (.A1(_0819_),
    .A2(net1076),
    .Y(_0224_),
    .B1(_1045_));
 sg13g2_nand2_1 _4324_ (.Y(_1046_),
    .A(net1321),
    .B(\main.adder.s4_exponent_adjust[0] ));
 sg13g2_or3_1 _4325_ (.A(\main.adder.s3_sum[2] ),
    .B(\main.adder.s3_sum[0] ),
    .C(\main.adder.s3_sum[1] ),
    .X(_1047_));
 sg13g2_or4_1 _4326_ (.A(\main.adder.s3_sum[3] ),
    .B(\main.adder.s3_sum[2] ),
    .C(\main.adder.s3_sum[0] ),
    .D(\main.adder.s3_sum[1] ),
    .X(_1048_));
 sg13g2_or2_1 _4327_ (.X(_1049_),
    .B(_1048_),
    .A(\main.adder.s3_sum[4] ));
 sg13g2_nor4_2 _4328_ (.A(\main.adder.s3_sum[6] ),
    .B(\main.adder.s3_sum[5] ),
    .C(\main.adder.s3_sum[4] ),
    .Y(_1050_),
    .D(_1048_));
 sg13g2_nand2_1 _4329_ (.Y(_1051_),
    .A(_0683_),
    .B(_1050_));
 sg13g2_or2_1 _4330_ (.X(_1052_),
    .B(_1051_),
    .A(\main.adder.s3_sum[8] ));
 sg13g2_or3_1 _4331_ (.A(\main.adder.s3_sum[10] ),
    .B(\main.adder.s3_sum[9] ),
    .C(_1052_),
    .X(_1053_));
 sg13g2_nor4_1 _4332_ (.A(\main.adder.s3_sum[11] ),
    .B(\main.adder.s3_sum[10] ),
    .C(\main.adder.s3_sum[9] ),
    .D(\main.adder.s3_sum[8] ),
    .Y(_1054_));
 sg13g2_and4_2 _4333_ (.A(_0682_),
    .B(_0683_),
    .C(_1050_),
    .D(_1054_),
    .X(_1055_));
 sg13g2_nand4_1 _4334_ (.B(_0683_),
    .C(_1050_),
    .A(_0682_),
    .Y(_1056_),
    .D(_1054_));
 sg13g2_nor3_1 _4335_ (.A(\main.adder.s3_sum[14] ),
    .B(\main.adder.s3_sum[13] ),
    .C(_1056_),
    .Y(_1057_));
 sg13g2_nor3_2 _4336_ (.A(\main.adder.s3_sum[15] ),
    .B(\main.adder.s3_sum[14] ),
    .C(\main.adder.s3_sum[13] ),
    .Y(_1058_));
 sg13g2_and2_1 _4337_ (.A(_1055_),
    .B(_1058_),
    .X(_1059_));
 sg13g2_nand2_1 _4338_ (.Y(_1060_),
    .A(_1055_),
    .B(_1058_));
 sg13g2_nor4_1 _4339_ (.A(\main.adder.s3_sum[23] ),
    .B(\main.adder.s3_sum[22] ),
    .C(\main.adder.s3_sum[21] ),
    .D(\main.adder.s3_sum[20] ),
    .Y(_1061_));
 sg13g2_nor4_2 _4340_ (.A(\main.adder.s3_sum[19] ),
    .B(\main.adder.s3_sum[18] ),
    .C(\main.adder.s3_sum[17] ),
    .Y(_1062_),
    .D(\main.adder.s3_sum[16] ));
 sg13g2_and2_1 _4341_ (.A(_1061_),
    .B(_1062_),
    .X(_1063_));
 sg13g2_nor2_1 _4342_ (.A(\main.adder.s3_sum[25] ),
    .B(\main.adder.s3_sum[24] ),
    .Y(_1064_));
 sg13g2_and4_2 _4343_ (.A(_1055_),
    .B(_1058_),
    .C(_1063_),
    .D(_1064_),
    .X(_1065_));
 sg13g2_nand4_1 _4344_ (.B(_1058_),
    .C(_1063_),
    .A(_1055_),
    .Y(_1066_),
    .D(_1064_));
 sg13g2_nor4_2 _4345_ (.A(\main.adder.s3_sum[29] ),
    .B(\main.adder.s3_sum[28] ),
    .C(\main.adder.s3_sum[27] ),
    .Y(_1067_),
    .D(\main.adder.s3_sum[26] ));
 sg13g2_nand3_1 _4346_ (.B(_0685_),
    .C(_1067_),
    .A(_0684_),
    .Y(_1068_));
 sg13g2_inv_1 _4347_ (.Y(_1069_),
    .A(_1068_));
 sg13g2_nor2_2 _4348_ (.A(net1127),
    .B(_1068_),
    .Y(_1070_));
 sg13g2_nor2_1 _4349_ (.A(\main.adder.s3_sum[37] ),
    .B(\main.adder.s3_sum[36] ),
    .Y(_1071_));
 sg13g2_nor3_1 _4350_ (.A(\main.adder.s3_sum[38] ),
    .B(\main.adder.s3_sum[37] ),
    .C(\main.adder.s3_sum[36] ),
    .Y(_1072_));
 sg13g2_nor3_1 _4351_ (.A(\main.adder.s3_sum[32] ),
    .B(\main.adder.s3_sum[34] ),
    .C(\main.adder.s3_sum[33] ),
    .Y(_1073_));
 sg13g2_nand3_1 _4352_ (.B(_0693_),
    .C(_0694_),
    .A(_0686_),
    .Y(_1074_));
 sg13g2_nor2_1 _4353_ (.A(\main.adder.s3_sum[39] ),
    .B(\main.adder.s3_sum[35] ),
    .Y(_1075_));
 sg13g2_nand3_1 _4354_ (.B(_1073_),
    .C(_1075_),
    .A(_1072_),
    .Y(_1076_));
 sg13g2_inv_1 _4355_ (.Y(_1077_),
    .A(_1076_));
 sg13g2_nor2_1 _4356_ (.A(\main.adder.s3_sum[41] ),
    .B(\main.adder.s3_sum[40] ),
    .Y(_1078_));
 sg13g2_nor4_2 _4357_ (.A(\main.adder.s3_sum[43] ),
    .B(\main.adder.s3_sum[42] ),
    .C(\main.adder.s3_sum[41] ),
    .Y(_1079_),
    .D(\main.adder.s3_sum[40] ));
 sg13g2_nor2_1 _4358_ (.A(\main.adder.s3_sum[45] ),
    .B(\main.adder.s3_sum[44] ),
    .Y(_1080_));
 sg13g2_nand2b_1 _4359_ (.Y(_1081_),
    .B(_1080_),
    .A_N(\main.adder.s3_sum[46] ));
 sg13g2_nand2_1 _4360_ (.Y(_1082_),
    .A(_0688_),
    .B(_1079_));
 sg13g2_nor3_1 _4361_ (.A(_1076_),
    .B(_1081_),
    .C(_1082_),
    .Y(_1083_));
 sg13g2_nand3_1 _4362_ (.B(_1069_),
    .C(_1083_),
    .A(_1065_),
    .Y(_1084_));
 sg13g2_xnor2_1 _4363_ (.Y(_1085_),
    .A(net1262),
    .B(net1121));
 sg13g2_and2_1 _4364_ (.A(\main.adder.s3_sum[48] ),
    .B(_1085_),
    .X(_1086_));
 sg13g2_nand2_1 _4365_ (.Y(_1087_),
    .A(\main.adder.s3_sum[48] ),
    .B(_1085_));
 sg13g2_and4_1 _4366_ (.A(_0687_),
    .B(_1065_),
    .C(_1069_),
    .D(_1083_),
    .X(_1088_));
 sg13g2_a21oi_2 _4367_ (.B1(net1119),
    .Y(_1089_),
    .A2(net1121),
    .A1(net1261));
 sg13g2_a21o_1 _4368_ (.A2(net1120),
    .A1(net1261),
    .B1(net1118),
    .X(_1090_));
 sg13g2_nor3_2 _4369_ (.A(net1127),
    .B(_1068_),
    .C(_1076_),
    .Y(_1091_));
 sg13g2_and2_1 _4370_ (.A(_1079_),
    .B(_1091_),
    .X(_1092_));
 sg13g2_a221oi_1 _4371_ (.B2(_1079_),
    .C1(net1119),
    .B1(_1091_),
    .A1(net1262),
    .Y(_1093_),
    .A2(net1121));
 sg13g2_a21o_1 _4372_ (.A2(net1115),
    .A1(_1081_),
    .B1(_1093_),
    .X(_1094_));
 sg13g2_xnor2_1 _4373_ (.Y(_1095_),
    .A(\main.adder.s3_sum[47] ),
    .B(_1094_));
 sg13g2_xnor2_1 _4374_ (.Y(_1096_),
    .A(_0688_),
    .B(_1094_));
 sg13g2_and4_1 _4375_ (.A(_1065_),
    .B(_1069_),
    .C(_1077_),
    .D(_1078_),
    .X(_1097_));
 sg13g2_a221oi_1 _4376_ (.B2(_1078_),
    .C1(net1119),
    .B1(_1091_),
    .A1(net1261),
    .Y(_1098_),
    .A2(net1120));
 sg13g2_a221oi_1 _4377_ (.B2(_0689_),
    .C1(net1118),
    .B1(_1097_),
    .A1(net1260),
    .Y(_1099_),
    .A2(net1120));
 sg13g2_xnor2_1 _4378_ (.Y(_1100_),
    .A(\main.adder.s3_sum[43] ),
    .B(_1099_));
 sg13g2_nor3_1 _4379_ (.A(net1127),
    .B(_1068_),
    .C(_1074_),
    .Y(_1101_));
 sg13g2_nor4_2 _4380_ (.A(\main.adder.s3_sum[35] ),
    .B(net1127),
    .C(_1068_),
    .Y(_1102_),
    .D(_1074_));
 sg13g2_a221oi_1 _4381_ (.B2(_0692_),
    .C1(net1118),
    .B1(_1101_),
    .A1(net1260),
    .Y(_1103_),
    .A2(net1120));
 sg13g2_xnor2_1 _4382_ (.Y(_1104_),
    .A(\main.adder.s3_sum[36] ),
    .B(_1103_));
 sg13g2_xnor2_1 _4383_ (.Y(_1105_),
    .A(\main.adder.s3_sum[44] ),
    .B(_1093_));
 sg13g2_xnor2_1 _4384_ (.Y(_1106_),
    .A(\main.adder.s3_sum[42] ),
    .B(_1098_));
 sg13g2_inv_1 _4385_ (.Y(_1107_),
    .A(_1106_));
 sg13g2_a21oi_1 _4386_ (.A1(_1071_),
    .A2(_1102_),
    .Y(_1108_),
    .B1(net1112));
 sg13g2_a21oi_1 _4387_ (.A1(_1072_),
    .A2(_1102_),
    .Y(_1109_),
    .B1(net1112));
 sg13g2_xor2_1 _4388_ (.B(_1109_),
    .A(\main.adder.s3_sum[39] ),
    .X(_1110_));
 sg13g2_a21o_1 _4389_ (.A2(_1089_),
    .A1(\main.adder.s3_sum[44] ),
    .B1(_1093_),
    .X(_1111_));
 sg13g2_xnor2_1 _4390_ (.Y(_1112_),
    .A(\main.adder.s3_sum[45] ),
    .B(_1111_));
 sg13g2_a21oi_1 _4391_ (.A1(_1080_),
    .A2(_1092_),
    .Y(_1113_),
    .B1(net1113));
 sg13g2_xnor2_1 _4392_ (.Y(_1114_),
    .A(\main.adder.s3_sum[46] ),
    .B(_1113_));
 sg13g2_nor3_1 _4393_ (.A(\main.adder.s3_sum[32] ),
    .B(net1127),
    .C(_1068_),
    .Y(_1115_));
 sg13g2_a221oi_1 _4394_ (.B2(net1260),
    .C1(net1118),
    .B1(net1120),
    .A1(_0686_),
    .Y(_1116_),
    .A2(_1070_));
 sg13g2_xnor2_1 _4395_ (.Y(_1117_),
    .A(\main.adder.s3_sum[33] ),
    .B(_1116_));
 sg13g2_a221oi_1 _4396_ (.B2(_0691_),
    .C1(net1118),
    .B1(_1102_),
    .A1(net1260),
    .Y(_1118_),
    .A2(net1120));
 sg13g2_xnor2_1 _4397_ (.Y(_1119_),
    .A(\main.adder.s3_sum[37] ),
    .B(_1118_));
 sg13g2_nor2_1 _4398_ (.A(net1260),
    .B(_1070_),
    .Y(_1120_));
 sg13g2_xnor2_1 _4399_ (.Y(_1121_),
    .A(\main.adder.s3_sum[32] ),
    .B(_1120_));
 sg13g2_a21oi_1 _4400_ (.A1(_1070_),
    .A2(_1077_),
    .Y(_1122_),
    .B1(net1260));
 sg13g2_xnor2_1 _4401_ (.Y(_1123_),
    .A(\main.adder.s3_sum[40] ),
    .B(_1122_));
 sg13g2_a221oi_1 _4402_ (.B2(net1260),
    .C1(net1118),
    .B1(net1120),
    .A1(_1070_),
    .Y(_1124_),
    .A2(_1073_));
 sg13g2_xnor2_1 _4403_ (.Y(_1125_),
    .A(\main.adder.s3_sum[35] ),
    .B(_1124_));
 sg13g2_a221oi_1 _4404_ (.B2(_0690_),
    .C1(net1118),
    .B1(_1091_),
    .A1(net1261),
    .Y(_1126_),
    .A2(net1121));
 sg13g2_xnor2_1 _4405_ (.Y(_1127_),
    .A(\main.adder.s3_sum[41] ),
    .B(_1126_));
 sg13g2_xnor2_1 _4406_ (.Y(_1128_),
    .A(\main.adder.s3_sum[38] ),
    .B(_1108_));
 sg13g2_a221oi_1 _4407_ (.B2(_0694_),
    .C1(net1118),
    .B1(_1115_),
    .A1(net1260),
    .Y(_1129_),
    .A2(net1120));
 sg13g2_xnor2_1 _4408_ (.Y(_1130_),
    .A(net1626),
    .B(_1129_));
 sg13g2_nand4_1 _4409_ (.B(_1117_),
    .C(_1121_),
    .A(_1104_),
    .Y(_1131_),
    .D(_1130_));
 sg13g2_and4_2 _4410_ (.A(_1095_),
    .B(_1112_),
    .C(_1114_),
    .D(_1128_),
    .X(_1132_));
 sg13g2_nand4_1 _4411_ (.B(_1105_),
    .C(_1106_),
    .A(_1087_),
    .Y(_1133_),
    .D(_1119_));
 sg13g2_nand4_1 _4412_ (.B(_1123_),
    .C(_1125_),
    .A(_1100_),
    .Y(_1134_),
    .D(_1127_));
 sg13g2_nor4_2 _4413_ (.A(_1110_),
    .B(_1131_),
    .C(_1133_),
    .Y(_1135_),
    .D(_1134_));
 sg13g2_and2_2 _4414_ (.A(_1132_),
    .B(_1135_),
    .X(_1136_));
 sg13g2_nand2_1 _4415_ (.Y(_1137_),
    .A(_1132_),
    .B(_1135_));
 sg13g2_nor2_1 _4416_ (.A(_0021_),
    .B(net1116),
    .Y(_1138_));
 sg13g2_nor3_2 _4417_ (.A(\main.adder.s3_sum[17] ),
    .B(\main.adder.s3_sum[16] ),
    .C(_1060_),
    .Y(_1139_));
 sg13g2_nor2b_1 _4418_ (.A(\main.adder.s3_sum[18] ),
    .B_N(_1139_),
    .Y(_1140_));
 sg13g2_nand3_1 _4419_ (.B(_1058_),
    .C(_1062_),
    .A(_1055_),
    .Y(_1141_));
 sg13g2_nor3_2 _4420_ (.A(\main.adder.s3_sum[21] ),
    .B(\main.adder.s3_sum[20] ),
    .C(_1141_),
    .Y(_1142_));
 sg13g2_nand2b_1 _4421_ (.Y(_1143_),
    .B(_1142_),
    .A_N(\main.adder.s3_sum[22] ));
 sg13g2_xnor2_1 _4422_ (.Y(_1144_),
    .A(\main.adder.s3_sum[22] ),
    .B(_1142_));
 sg13g2_a21oi_2 _4423_ (.B1(_1138_),
    .Y(_1145_),
    .A2(_1144_),
    .A1(net1117));
 sg13g2_nor2_1 _4424_ (.A(_0029_),
    .B(net1114),
    .Y(_1146_));
 sg13g2_nor3_1 _4425_ (.A(\main.adder.s3_sum[27] ),
    .B(\main.adder.s3_sum[26] ),
    .C(net1127),
    .Y(_1147_));
 sg13g2_nor4_1 _4426_ (.A(\main.adder.s3_sum[28] ),
    .B(\main.adder.s3_sum[27] ),
    .C(\main.adder.s3_sum[26] ),
    .D(net1127),
    .Y(_1148_));
 sg13g2_nand2_1 _4427_ (.Y(_1149_),
    .A(_1065_),
    .B(_1067_));
 sg13g2_xnor2_1 _4428_ (.Y(_1150_),
    .A(_0685_),
    .B(_1149_));
 sg13g2_a21oi_2 _4429_ (.B1(_1146_),
    .Y(_1151_),
    .A2(_1150_),
    .A1(net1117));
 sg13g2_a221oi_1 _4430_ (.B2(net1262),
    .C1(net1119),
    .B1(net1121),
    .A1(_1059_),
    .Y(_1152_),
    .A2(_1063_));
 sg13g2_xor2_1 _4431_ (.B(_1152_),
    .A(_0023_),
    .X(_1153_));
 sg13g2_inv_1 _4432_ (.Y(_1154_),
    .A(_1153_));
 sg13g2_o21ai_1 _4433_ (.B1(\main.adder.s3_sum[31] ),
    .Y(_1155_),
    .A1(\main.adder.s3_sum[30] ),
    .A2(_1149_));
 sg13g2_a22oi_1 _4434_ (.Y(_1156_),
    .B1(_1120_),
    .B2(_1155_),
    .A2(net1112),
    .A1(_0696_));
 sg13g2_a221oi_1 _4435_ (.B2(net1262),
    .C1(net1119),
    .B1(net1121),
    .A1(_0681_),
    .Y(_1157_),
    .A2(_1057_));
 sg13g2_xnor2_1 _4436_ (.Y(_1158_),
    .A(\main.adder.s3_sum[16] ),
    .B(_1157_));
 sg13g2_nand2_1 _4437_ (.Y(_1159_),
    .A(_1156_),
    .B(_1158_));
 sg13g2_nand2_1 _4438_ (.Y(_1160_),
    .A(\main.adder.s3_sum[23] ),
    .B(_1143_));
 sg13g2_a22oi_1 _4439_ (.Y(_1161_),
    .B1(_1152_),
    .B2(_1160_),
    .A2(net1112),
    .A1(_0695_));
 sg13g2_nor2_1 _4440_ (.A(_0018_),
    .B(net1114),
    .Y(_1162_));
 sg13g2_xnor2_1 _4441_ (.Y(_1163_),
    .A(\main.adder.s3_sum[19] ),
    .B(_1140_));
 sg13g2_a21oi_2 _4442_ (.B1(_1162_),
    .Y(_1164_),
    .A2(_1163_),
    .A1(net1114));
 sg13g2_nand3_1 _4443_ (.B(_1059_),
    .C(_1063_),
    .A(_0023_),
    .Y(_1165_));
 sg13g2_xnor2_1 _4444_ (.Y(_1166_),
    .A(net963),
    .B(_1165_));
 sg13g2_mux2_2 _4445_ (.A0(_0024_),
    .A1(_1166_),
    .S(net1114),
    .X(_1167_));
 sg13g2_xor2_1 _4446_ (.B(_1147_),
    .A(\main.adder.s3_sum[28] ),
    .X(_1168_));
 sg13g2_mux2_2 _4447_ (.A0(_0027_),
    .A1(_1168_),
    .S(net1116),
    .X(_1169_));
 sg13g2_xnor2_1 _4448_ (.Y(_1170_),
    .A(\main.adder.s3_sum[26] ),
    .B(_1066_));
 sg13g2_mux2_2 _4449_ (.A0(_0025_),
    .A1(_1170_),
    .S(net1116),
    .X(_1171_));
 sg13g2_nor2_1 _4450_ (.A(_0019_),
    .B(net1116),
    .Y(_1172_));
 sg13g2_xor2_1 _4451_ (.B(_1141_),
    .A(\main.adder.s3_sum[20] ),
    .X(_1173_));
 sg13g2_a21oi_2 _4452_ (.B1(_1172_),
    .Y(_1174_),
    .A2(_1173_),
    .A1(net1116));
 sg13g2_inv_1 _4453_ (.Y(_1175_),
    .A(_1174_));
 sg13g2_xor2_1 _4454_ (.B(_1148_),
    .A(\main.adder.s3_sum[29] ),
    .X(_1176_));
 sg13g2_mux2_2 _4455_ (.A0(_0028_),
    .A1(_1176_),
    .S(net1116),
    .X(_1177_));
 sg13g2_nor2_1 _4456_ (.A(_0026_),
    .B(net1116),
    .Y(_1178_));
 sg13g2_o21ai_1 _4457_ (.B1(\main.adder.s3_sum[27] ),
    .Y(_1179_),
    .A1(\main.adder.s3_sum[26] ),
    .A2(net1127));
 sg13g2_nor2b_1 _4458_ (.A(_1147_),
    .B_N(_1179_),
    .Y(_1180_));
 sg13g2_a21oi_2 _4459_ (.B1(_1178_),
    .Y(_1181_),
    .A2(_1180_),
    .A1(net1116));
 sg13g2_xor2_1 _4460_ (.B(_1139_),
    .A(\main.adder.s3_sum[18] ),
    .X(_1182_));
 sg13g2_mux2_2 _4461_ (.A0(_0017_),
    .A1(_1182_),
    .S(net1114),
    .X(_1183_));
 sg13g2_o21ai_1 _4462_ (.B1(\main.adder.s3_sum[21] ),
    .Y(_1184_),
    .A1(\main.adder.s3_sum[20] ),
    .A2(_1141_));
 sg13g2_nand2b_1 _4463_ (.Y(_1185_),
    .B(_1184_),
    .A_N(_1142_));
 sg13g2_mux2_2 _4464_ (.A0(_0020_),
    .A1(_1185_),
    .S(net1117),
    .X(_1186_));
 sg13g2_o21ai_1 _4465_ (.B1(\main.adder.s3_sum[17] ),
    .Y(_1187_),
    .A1(\main.adder.s3_sum[16] ),
    .A2(_1060_));
 sg13g2_nand2b_1 _4466_ (.Y(_1188_),
    .B(_1187_),
    .A_N(_1139_));
 sg13g2_mux2_2 _4467_ (.A0(_0016_),
    .A1(_1188_),
    .S(net1114),
    .X(_1189_));
 sg13g2_nand4_1 _4468_ (.B(_1171_),
    .C(_1183_),
    .A(_1167_),
    .Y(_1190_),
    .D(_1189_));
 sg13g2_and4_1 _4469_ (.A(_1151_),
    .B(_1164_),
    .C(_1174_),
    .D(_1181_),
    .X(_1191_));
 sg13g2_nand4_1 _4470_ (.B(_1169_),
    .C(_1177_),
    .A(_1153_),
    .Y(_1192_),
    .D(_1186_));
 sg13g2_nor3_1 _4471_ (.A(_1159_),
    .B(_1190_),
    .C(_1192_),
    .Y(_1193_));
 sg13g2_and4_1 _4472_ (.A(_1145_),
    .B(_1161_),
    .C(_1191_),
    .D(_1193_),
    .X(_1194_));
 sg13g2_nand4_1 _4473_ (.B(_1161_),
    .C(_1191_),
    .A(_1145_),
    .Y(_1195_),
    .D(_1193_));
 sg13g2_a21oi_2 _4474_ (.B1(net1107),
    .Y(_1196_),
    .A2(_1195_),
    .A1(net1072));
 sg13g2_o21ai_1 _4475_ (.B1(_1087_),
    .Y(_1197_),
    .A1(net1071),
    .A2(_1194_));
 sg13g2_o21ai_1 _4476_ (.B1(_1157_),
    .Y(_1198_),
    .A1(_0681_),
    .A2(_1057_));
 sg13g2_o21ai_1 _4477_ (.B1(_1198_),
    .Y(_1199_),
    .A1(_0072_),
    .A2(net1114));
 sg13g2_nor2_1 _4478_ (.A(net1071),
    .B(_1156_),
    .Y(_1200_));
 sg13g2_nor3_2 _4479_ (.A(net1107),
    .B(net1071),
    .C(_1195_),
    .Y(_1201_));
 sg13g2_a221oi_1 _4480_ (.B2(_1201_),
    .C1(_1200_),
    .B1(_1199_),
    .A1(_1096_),
    .Y(_1202_),
    .A2(_1196_));
 sg13g2_o21ai_1 _4481_ (.B1(net1114),
    .Y(_1203_),
    .A1(\main.adder.s3_sum[13] ),
    .A2(_1056_));
 sg13g2_xnor2_1 _4482_ (.Y(_1204_),
    .A(\main.adder.s3_sum[14] ),
    .B(_1203_));
 sg13g2_nand2_1 _4483_ (.Y(_1205_),
    .A(_1201_),
    .B(_1204_));
 sg13g2_nor3_1 _4484_ (.A(net1070),
    .B(_1151_),
    .C(_1194_),
    .Y(_1206_));
 sg13g2_a221oi_1 _4485_ (.B2(_1195_),
    .C1(_1114_),
    .B1(net1072),
    .A1(\main.adder.s3_sum[48] ),
    .Y(_1207_),
    .A2(_1085_));
 sg13g2_nor2_1 _4486_ (.A(_1206_),
    .B(_1207_),
    .Y(_1208_));
 sg13g2_nand3_1 _4487_ (.B(_1205_),
    .C(_1208_),
    .A(_1202_),
    .Y(_1209_));
 sg13g2_o21ai_1 _4488_ (.B1(net1115),
    .Y(_1210_),
    .A1(\main.adder.s3_sum[9] ),
    .A2(_1052_));
 sg13g2_xor2_1 _4489_ (.B(_1210_),
    .A(\main.adder.s3_sum[10] ),
    .X(_1211_));
 sg13g2_inv_1 _4490_ (.Y(_1212_),
    .A(_1211_));
 sg13g2_nor2_1 _4491_ (.A(net1070),
    .B(_1171_),
    .Y(_1213_));
 sg13g2_a221oi_1 _4492_ (.B2(_1212_),
    .C1(_1213_),
    .B1(_1201_),
    .A1(_1107_),
    .Y(_1214_),
    .A2(_1196_));
 sg13g2_inv_1 _4493_ (.Y(_1215_),
    .A(_1214_));
 sg13g2_nor2_1 _4494_ (.A(net1070),
    .B(_1167_),
    .Y(_1216_));
 sg13g2_a21oi_1 _4495_ (.A1(\main.adder.s3_sum[9] ),
    .A2(_1052_),
    .Y(_1217_),
    .B1(_1210_));
 sg13g2_a21oi_2 _4496_ (.B1(_1217_),
    .Y(_1218_),
    .A2(net1113),
    .A1(_0723_));
 sg13g2_nand3b_1 _4497_ (.B(_1135_),
    .C(_1132_),
    .Y(_1219_),
    .A_N(_1218_));
 sg13g2_a221oi_1 _4498_ (.B2(_1127_),
    .C1(net1107),
    .B1(_1219_),
    .A1(net1072),
    .Y(_1220_),
    .A2(_1195_));
 sg13g2_nor2_1 _4499_ (.A(net1070),
    .B(_1181_),
    .Y(_1221_));
 sg13g2_o21ai_1 _4500_ (.B1(net1115),
    .Y(_1222_),
    .A1(\main.adder.s3_sum[11] ),
    .A2(_1053_));
 sg13g2_a21oi_1 _4501_ (.A1(\main.adder.s3_sum[11] ),
    .A2(_1053_),
    .Y(_1223_),
    .B1(_1222_));
 sg13g2_a21oi_2 _4502_ (.B1(_1223_),
    .Y(_1224_),
    .A2(net1113),
    .A1(_0724_));
 sg13g2_nand3b_1 _4503_ (.B(_1135_),
    .C(_1132_),
    .Y(_1225_),
    .A_N(_1224_));
 sg13g2_a221oi_1 _4504_ (.B2(_1100_),
    .C1(net1107),
    .B1(_1225_),
    .A1(net1072),
    .Y(_1226_),
    .A2(_1195_));
 sg13g2_or2_1 _4505_ (.X(_1227_),
    .B(_1226_),
    .A(_1221_));
 sg13g2_nor4_1 _4506_ (.A(_1216_),
    .B(_1220_),
    .C(_1221_),
    .D(_1226_),
    .Y(_1228_));
 sg13g2_nor2_1 _4507_ (.A(net1070),
    .B(_1177_),
    .Y(_1229_));
 sg13g2_a21oi_1 _4508_ (.A1(\main.adder.s3_sum[13] ),
    .A2(_1056_),
    .Y(_1230_),
    .B1(_1203_));
 sg13g2_a21oi_2 _4509_ (.B1(_1230_),
    .Y(_1231_),
    .A2(net1113),
    .A1(_0725_));
 sg13g2_nand3b_1 _4510_ (.B(_1135_),
    .C(_1132_),
    .Y(_1232_),
    .A_N(_1231_));
 sg13g2_a221oi_1 _4511_ (.B2(_1112_),
    .C1(net1107),
    .B1(_1232_),
    .A1(net1072),
    .Y(_1233_),
    .A2(_1195_));
 sg13g2_nor2_1 _4512_ (.A(net1070),
    .B(_1169_),
    .Y(_1234_));
 sg13g2_xnor2_1 _4513_ (.Y(_1235_),
    .A(_0682_),
    .B(_1222_));
 sg13g2_nand3b_1 _4514_ (.B(_1135_),
    .C(_1132_),
    .Y(_1236_),
    .A_N(_1235_));
 sg13g2_a221oi_1 _4515_ (.B2(_1105_),
    .C1(net1107),
    .B1(_1236_),
    .A1(net1072),
    .Y(_1237_),
    .A2(_1195_));
 sg13g2_nor4_2 _4516_ (.A(_1229_),
    .B(_1233_),
    .C(_1234_),
    .Y(_1238_),
    .D(_1237_));
 sg13g2_nand2_1 _4517_ (.Y(_1239_),
    .A(_1051_),
    .B(net1115));
 sg13g2_xor2_1 _4518_ (.B(_1239_),
    .A(\main.adder.s3_sum[8] ),
    .X(_1240_));
 sg13g2_and3_1 _4519_ (.X(_1241_),
    .A(_1132_),
    .B(_1135_),
    .C(_1240_));
 sg13g2_a221oi_1 _4520_ (.B2(_1195_),
    .C1(_1241_),
    .B1(net1072),
    .A1(\main.adder.s3_sum[48] ),
    .Y(_1242_),
    .A2(_1085_));
 sg13g2_a21oi_1 _4521_ (.A1(_1123_),
    .A2(net1070),
    .Y(_1243_),
    .B1(net1107));
 sg13g2_o21ai_1 _4522_ (.B1(_1243_),
    .Y(_1244_),
    .A1(_1154_),
    .A2(_1242_));
 sg13g2_and4_1 _4523_ (.A(_1214_),
    .B(_1228_),
    .C(_1238_),
    .D(_1244_),
    .X(_1245_));
 sg13g2_nand4_1 _4524_ (.B(_1228_),
    .C(_1238_),
    .A(_1214_),
    .Y(_1246_),
    .D(_1244_));
 sg13g2_nor2_1 _4525_ (.A(_0683_),
    .B(_1050_),
    .Y(_1247_));
 sg13g2_nand2b_1 _4526_ (.Y(_1248_),
    .B(net1112),
    .A_N(_0068_));
 sg13g2_o21ai_1 _4527_ (.B1(_1248_),
    .Y(_1249_),
    .A1(_1239_),
    .A2(_1247_));
 sg13g2_nor2_1 _4528_ (.A(net1071),
    .B(_1161_),
    .Y(_1250_));
 sg13g2_a221oi_1 _4529_ (.B2(_1249_),
    .C1(_1250_),
    .B1(_1201_),
    .A1(_1110_),
    .Y(_1251_),
    .A2(_1196_));
 sg13g2_o21ai_1 _4530_ (.B1(net1115),
    .Y(_1252_),
    .A1(\main.adder.s3_sum[5] ),
    .A2(_1049_));
 sg13g2_xor2_1 _4531_ (.B(_1252_),
    .A(\main.adder.s3_sum[6] ),
    .X(_1253_));
 sg13g2_nor2_1 _4532_ (.A(net1071),
    .B(_1145_),
    .Y(_1254_));
 sg13g2_o21ai_1 _4533_ (.B1(_1128_),
    .Y(_1255_),
    .A1(net1071),
    .A2(_1253_));
 sg13g2_a21oi_1 _4534_ (.A1(_1196_),
    .A2(_1255_),
    .Y(_1256_),
    .B1(_1254_));
 sg13g2_nand2_1 _4535_ (.Y(_1257_),
    .A(_1251_),
    .B(_1256_));
 sg13g2_nor2_2 _4536_ (.A(_1209_),
    .B(_1246_),
    .Y(_1258_));
 sg13g2_a21oi_1 _4537_ (.A1(_1245_),
    .A2(_1257_),
    .Y(_1259_),
    .B1(_1209_));
 sg13g2_nand2_1 _4538_ (.Y(_1260_),
    .A(_1048_),
    .B(net1115));
 sg13g2_xnor2_1 _4539_ (.Y(_1261_),
    .A(\main.adder.s3_sum[4] ),
    .B(_1260_));
 sg13g2_mux2_1 _4540_ (.A0(_1175_),
    .A1(_1261_),
    .S(_1196_),
    .X(_1262_));
 sg13g2_o21ai_1 _4541_ (.B1(_1137_),
    .Y(_1263_),
    .A1(net1108),
    .A2(_1119_));
 sg13g2_a21oi_1 _4542_ (.A1(\main.adder.s3_sum[5] ),
    .A2(_1049_),
    .Y(_1264_),
    .B1(_1252_));
 sg13g2_a21oi_1 _4543_ (.A1(_0722_),
    .A2(net1112),
    .Y(_1265_),
    .B1(_1264_));
 sg13g2_and2_1 _4544_ (.A(_1136_),
    .B(_1265_),
    .X(_1266_));
 sg13g2_o21ai_1 _4545_ (.B1(_1186_),
    .Y(_1267_),
    .A1(_1197_),
    .A2(_1266_));
 sg13g2_nand2_1 _4546_ (.Y(_1268_),
    .A(_1263_),
    .B(_1267_));
 sg13g2_nor2_1 _4547_ (.A(net1108),
    .B(_1104_),
    .Y(_1269_));
 sg13g2_a221oi_1 _4548_ (.B2(_1267_),
    .C1(_1269_),
    .B1(_1263_),
    .A1(net1072),
    .Y(_1270_),
    .A2(_1262_));
 sg13g2_nor3_1 _4549_ (.A(_1209_),
    .B(_1246_),
    .C(_1270_),
    .Y(_1271_));
 sg13g2_nor3_1 _4550_ (.A(_1209_),
    .B(_1246_),
    .C(_1268_),
    .Y(_1272_));
 sg13g2_nand2b_1 _4551_ (.Y(_1273_),
    .B(_1238_),
    .A_N(_1271_));
 sg13g2_nor2_1 _4552_ (.A(_1125_),
    .B(_1197_),
    .Y(_1274_));
 sg13g2_a21oi_1 _4553_ (.A1(\main.adder.s3_sum[3] ),
    .A2(_1047_),
    .Y(_1275_),
    .B1(_1260_));
 sg13g2_a21oi_2 _4554_ (.B1(_1275_),
    .Y(_1276_),
    .A2(net1112),
    .A1(_0721_));
 sg13g2_nor2b_1 _4555_ (.A(_1276_),
    .B_N(_1201_),
    .Y(_1277_));
 sg13g2_nor2_1 _4556_ (.A(_1137_),
    .B(_1164_),
    .Y(_1278_));
 sg13g2_nor3_1 _4557_ (.A(_1274_),
    .B(_1277_),
    .C(_1278_),
    .Y(_1279_));
 sg13g2_nor3_1 _4558_ (.A(_1209_),
    .B(_1246_),
    .C(_1279_),
    .Y(_1280_));
 sg13g2_nor2_1 _4559_ (.A(_1227_),
    .B(_1280_),
    .Y(_1281_));
 sg13g2_nor2_1 _4560_ (.A(net1107),
    .B(_1130_),
    .Y(_1282_));
 sg13g2_nand2_1 _4561_ (.Y(_1283_),
    .A(_1183_),
    .B(_1197_));
 sg13g2_o21ai_1 _4562_ (.B1(net1115),
    .Y(_1284_),
    .A1(\main.adder.s3_sum[0] ),
    .A2(\main.adder.s3_sum[1] ));
 sg13g2_xor2_1 _4563_ (.B(_1284_),
    .A(\main.adder.s3_sum[2] ),
    .X(_1285_));
 sg13g2_a21oi_1 _4564_ (.A1(_1196_),
    .A2(_1285_),
    .Y(_1286_),
    .B1(net1071));
 sg13g2_a21oi_1 _4565_ (.A1(_1283_),
    .A2(_1286_),
    .Y(_1287_),
    .B1(_1282_));
 sg13g2_nor3_1 _4566_ (.A(_1209_),
    .B(_1246_),
    .C(_1287_),
    .Y(_1288_));
 sg13g2_nor4_1 _4567_ (.A(_1215_),
    .B(_1227_),
    .C(_1280_),
    .D(_1288_),
    .Y(_1289_));
 sg13g2_o21ai_1 _4568_ (.B1(_1259_),
    .Y(_1290_),
    .A1(_1273_),
    .A2(_1289_));
 sg13g2_nand3b_1 _4569_ (.B(_1259_),
    .C(_1238_),
    .Y(_1291_),
    .A_N(_1271_));
 sg13g2_a21oi_1 _4570_ (.A1(\main.adder.s3_sum[0] ),
    .A2(\main.adder.s3_sum[1] ),
    .Y(_1292_),
    .B1(_1284_));
 sg13g2_a21oi_2 _4571_ (.B1(_1292_),
    .Y(_1293_),
    .A2(net1112),
    .A1(_0720_));
 sg13g2_nor2b_1 _4572_ (.A(_1293_),
    .B_N(_1201_),
    .Y(_1294_));
 sg13g2_nor2_1 _4573_ (.A(net1070),
    .B(_1189_),
    .Y(_1295_));
 sg13g2_nor2_1 _4574_ (.A(_1117_),
    .B(_1197_),
    .Y(_1296_));
 sg13g2_nor3_1 _4575_ (.A(_1294_),
    .B(_1295_),
    .C(_1296_),
    .Y(_1297_));
 sg13g2_nor3_1 _4576_ (.A(_1209_),
    .B(_1246_),
    .C(_1297_),
    .Y(_1298_));
 sg13g2_nor3_1 _4577_ (.A(_1216_),
    .B(_1220_),
    .C(_1298_),
    .Y(_1299_));
 sg13g2_nor3_1 _4578_ (.A(_1229_),
    .B(_1233_),
    .C(_1272_),
    .Y(_1300_));
 sg13g2_o21ai_1 _4579_ (.B1(_1300_),
    .Y(_1301_),
    .A1(_1291_),
    .A2(_1299_));
 sg13g2_nand2b_1 _4580_ (.Y(_1302_),
    .B(_1301_),
    .A_N(_1290_));
 sg13g2_nor3_1 _4581_ (.A(_1209_),
    .B(_1246_),
    .C(_1251_),
    .Y(_1303_));
 sg13g2_o21ai_1 _4582_ (.B1(_1202_),
    .Y(_1304_),
    .A1(_1281_),
    .A2(_1291_));
 sg13g2_nor2_2 _4583_ (.A(_1303_),
    .B(_1304_),
    .Y(_1305_));
 sg13g2_nand2_1 _4584_ (.Y(_1306_),
    .A(_0745_),
    .B(_1290_));
 sg13g2_nand4_1 _4585_ (.B(_1302_),
    .C(_1305_),
    .A(_0076_),
    .Y(_1307_),
    .D(_1306_));
 sg13g2_nand2_1 _4586_ (.Y(_1308_),
    .A(_0726_),
    .B(_1258_));
 sg13g2_xnor2_1 _4587_ (.Y(_1309_),
    .A(_0726_),
    .B(_1258_));
 sg13g2_xor2_1 _4588_ (.B(_1291_),
    .A(\main.adder.s3_exponent[2] ),
    .X(_1310_));
 sg13g2_o21ai_1 _4589_ (.B1(_1310_),
    .Y(_1311_),
    .A1(_0745_),
    .A2(_1290_));
 sg13g2_nor2_1 _4590_ (.A(_1309_),
    .B(_1311_),
    .Y(_1312_));
 sg13g2_nand3_1 _4591_ (.B(_1291_),
    .C(_1308_),
    .A(\main.adder.s3_exponent[2] ),
    .Y(_1313_));
 sg13g2_o21ai_1 _4592_ (.B1(_1313_),
    .Y(_1314_),
    .A1(_0726_),
    .A2(_1258_));
 sg13g2_a21o_1 _4593_ (.A2(_1312_),
    .A1(_1307_),
    .B1(_1314_),
    .X(_1315_));
 sg13g2_nor2_2 _4594_ (.A(net1108),
    .B(_1201_),
    .Y(_1316_));
 sg13g2_nor2b_1 _4595_ (.A(\main.adder.s3_exponent[6] ),
    .B_N(_0074_),
    .Y(_1317_));
 sg13g2_nor2_1 _4596_ (.A(_0727_),
    .B(_0074_),
    .Y(_1318_));
 sg13g2_mux2_1 _4597_ (.A0(_1317_),
    .A1(_1318_),
    .S(net1109),
    .X(_1319_));
 sg13g2_o21ai_1 _4598_ (.B1(_1319_),
    .Y(_1320_),
    .A1(\main.adder.s3_exponent[5] ),
    .A2(_1316_));
 sg13g2_a22oi_1 _4599_ (.Y(_1321_),
    .B1(_1316_),
    .B2(\main.adder.s3_exponent[5] ),
    .A2(_1196_),
    .A1(\main.adder.s3_exponent[4] ));
 sg13g2_o21ai_1 _4600_ (.B1(_1321_),
    .Y(_1322_),
    .A1(\main.adder.s3_exponent[4] ),
    .A2(_1196_));
 sg13g2_nor2_1 _4601_ (.A(_1320_),
    .B(_1322_),
    .Y(_1323_));
 sg13g2_o21ai_1 _4602_ (.B1(_1317_),
    .Y(_1324_),
    .A1(_1320_),
    .A2(_1321_));
 sg13g2_a21oi_2 _4603_ (.B1(_1324_),
    .Y(_1325_),
    .A2(_1323_),
    .A1(_1315_));
 sg13g2_nor2_2 _4604_ (.A(net1109),
    .B(_1325_),
    .Y(_1326_));
 sg13g2_a221oi_1 _4605_ (.B2(_1305_),
    .C1(_1325_),
    .B1(_1302_),
    .A1(\main.adder.s3_sum[48] ),
    .Y(_1327_),
    .A2(_1085_));
 sg13g2_o21ai_1 _4606_ (.B1(net1390),
    .Y(_1328_),
    .A1(net1550),
    .A2(net1055));
 sg13g2_o21ai_1 _4607_ (.B1(_1046_),
    .Y(_0225_),
    .A1(_1327_),
    .A2(_1328_));
 sg13g2_xor2_1 _4608_ (.B(\main.adder.s3_exponent[0] ),
    .A(\main.adder.s3_exponent[1] ),
    .X(_1329_));
 sg13g2_o21ai_1 _4609_ (.B1(net1383),
    .Y(_1330_),
    .A1(net1055),
    .A2(_1329_));
 sg13g2_a21oi_1 _4610_ (.A1(_1290_),
    .A2(net1055),
    .Y(_1331_),
    .B1(_1330_));
 sg13g2_a21o_1 _4611_ (.A2(net1613),
    .A1(net1314),
    .B1(_1331_),
    .X(_0226_));
 sg13g2_nand3_1 _4612_ (.B(\main.adder.s3_exponent[0] ),
    .C(\main.adder.s3_exponent[2] ),
    .A(\main.adder.s3_exponent[1] ),
    .Y(_1332_));
 sg13g2_a21o_1 _4613_ (.A2(\main.adder.s3_exponent[0] ),
    .A1(\main.adder.s3_exponent[1] ),
    .B1(\main.adder.s3_exponent[2] ),
    .X(_1333_));
 sg13g2_and2_1 _4614_ (.A(_1332_),
    .B(_1333_),
    .X(_1334_));
 sg13g2_o21ai_1 _4615_ (.B1(net1391),
    .Y(_1335_),
    .A1(net1055),
    .A2(_1334_));
 sg13g2_a21o_1 _4616_ (.A2(net1055),
    .A1(_1291_),
    .B1(_1335_),
    .X(_1336_));
 sg13g2_o21ai_1 _4617_ (.B1(_1336_),
    .Y(_0227_),
    .A1(net1391),
    .A2(_0715_));
 sg13g2_nand2_1 _4618_ (.Y(_1337_),
    .A(net1321),
    .B(net1281));
 sg13g2_nor2_1 _4619_ (.A(_0726_),
    .B(_1332_),
    .Y(_1338_));
 sg13g2_xnor2_1 _4620_ (.Y(_1339_),
    .A(\main.adder.s3_exponent[3] ),
    .B(_1332_));
 sg13g2_nor3_1 _4621_ (.A(net1109),
    .B(_1258_),
    .C(_1325_),
    .Y(_1340_));
 sg13g2_o21ai_1 _4622_ (.B1(net1391),
    .Y(_1341_),
    .A1(net1055),
    .A2(_1339_));
 sg13g2_o21ai_1 _4623_ (.B1(_1337_),
    .Y(_0228_),
    .A1(_1340_),
    .A2(_1341_));
 sg13g2_nand2_1 _4624_ (.Y(_1342_),
    .A(net1321),
    .B(net1277));
 sg13g2_xor2_1 _4625_ (.B(_1338_),
    .A(\main.adder.s3_exponent[4] ),
    .X(_1343_));
 sg13g2_nor2_1 _4626_ (.A(net1055),
    .B(_1343_),
    .Y(_1344_));
 sg13g2_nor2_1 _4627_ (.A(_1197_),
    .B(_1325_),
    .Y(_1345_));
 sg13g2_o21ai_1 _4628_ (.B1(net1391),
    .Y(_1346_),
    .A1(_1197_),
    .A2(_1325_));
 sg13g2_o21ai_1 _4629_ (.B1(_1342_),
    .Y(_0229_),
    .A1(_1344_),
    .A2(_1346_));
 sg13g2_nor2_1 _4630_ (.A(net1391),
    .B(net1608),
    .Y(_1347_));
 sg13g2_nand3_1 _4631_ (.B(\main.adder.s3_exponent[4] ),
    .C(_1338_),
    .A(\main.adder.s3_exponent[5] ),
    .Y(_1348_));
 sg13g2_a21o_1 _4632_ (.A2(_1338_),
    .A1(\main.adder.s3_exponent[4] ),
    .B1(\main.adder.s3_exponent[5] ),
    .X(_1349_));
 sg13g2_nand2_1 _4633_ (.Y(_1350_),
    .A(_1348_),
    .B(_1349_));
 sg13g2_nor2_1 _4634_ (.A(net1055),
    .B(_1350_),
    .Y(_1351_));
 sg13g2_a21oi_1 _4635_ (.A1(_1136_),
    .A2(_1345_),
    .Y(_1352_),
    .B1(_1351_));
 sg13g2_a21oi_1 _4636_ (.A1(net1391),
    .A2(_1352_),
    .Y(_0230_),
    .B1(_1347_));
 sg13g2_nand2_1 _4637_ (.Y(_1353_),
    .A(net1316),
    .B(net1521));
 sg13g2_or2_1 _4638_ (.X(_1354_),
    .B(_1348_),
    .A(_0727_));
 sg13g2_a21oi_1 _4639_ (.A1(_0727_),
    .A2(_1348_),
    .Y(_1355_),
    .B1(net1316));
 sg13g2_nand2_1 _4640_ (.Y(_1356_),
    .A(_1354_),
    .B(_1355_));
 sg13g2_o21ai_1 _4641_ (.B1(_1353_),
    .Y(_0231_),
    .A1(_1326_),
    .A2(_1356_));
 sg13g2_xor2_1 _4642_ (.B(_1354_),
    .A(net1405),
    .X(_1357_));
 sg13g2_nor3_1 _4643_ (.A(net1315),
    .B(_1326_),
    .C(_1357_),
    .Y(_1358_));
 sg13g2_a21o_1 _4644_ (.A2(net1584),
    .A1(net1315),
    .B1(_1358_),
    .X(_0232_));
 sg13g2_nand2_1 _4645_ (.Y(_1359_),
    .A(net1392),
    .B(net1405));
 sg13g2_nor3_1 _4646_ (.A(_1326_),
    .B(_1354_),
    .C(_1359_),
    .Y(_1360_));
 sg13g2_a21o_1 _4647_ (.A2(net1575),
    .A1(net1316),
    .B1(_1360_),
    .X(_0233_));
 sg13g2_nor2b_1 _4648_ (.A(_0822_),
    .B_N(_0853_),
    .Y(_1361_));
 sg13g2_nor2_1 _4649_ (.A(net987),
    .B(net1073),
    .Y(_1362_));
 sg13g2_a21oi_1 _4650_ (.A1(_0922_),
    .A2(net1073),
    .Y(_0234_),
    .B1(_1362_));
 sg13g2_nor2_1 _4651_ (.A(net1411),
    .B(net1074),
    .Y(_1363_));
 sg13g2_a21oi_1 _4652_ (.A1(_0858_),
    .A2(net1074),
    .Y(_0235_),
    .B1(_1363_));
 sg13g2_nor2_1 _4653_ (.A(net1410),
    .B(net1075),
    .Y(_1364_));
 sg13g2_a21oi_1 _4654_ (.A1(_0885_),
    .A2(net1075),
    .Y(_0236_),
    .B1(_1364_));
 sg13g2_nor2_1 _4655_ (.A(net1047),
    .B(net1075),
    .Y(_1365_));
 sg13g2_a21oi_1 _4656_ (.A1(_0881_),
    .A2(net1075),
    .Y(_0237_),
    .B1(_1365_));
 sg13g2_nor2_1 _4657_ (.A(net984),
    .B(net1102),
    .Y(_1366_));
 sg13g2_a21oi_1 _4658_ (.A1(net1102),
    .A2(_0876_),
    .Y(_0238_),
    .B1(_1366_));
 sg13g2_nor2_1 _4659_ (.A(net1419),
    .B(net1077),
    .Y(_1367_));
 sg13g2_a21oi_1 _4660_ (.A1(_0961_),
    .A2(_1043_),
    .Y(_0239_),
    .B1(_1367_));
 sg13g2_nor2_1 _4661_ (.A(net988),
    .B(net1103),
    .Y(_1368_));
 sg13g2_a21oi_1 _4662_ (.A1(net1103),
    .A2(_0930_),
    .Y(_0240_),
    .B1(_1368_));
 sg13g2_a21o_1 _4663_ (.A2(net1339),
    .A1(\main.spi.state[0] ),
    .B1(_0697_),
    .X(_1369_));
 sg13g2_nor2b_1 _4664_ (.A(net1488),
    .B_N(\main.spi.SPI_clock_sampler.sample_register[0] ),
    .Y(_1370_));
 sg13g2_nand2_1 _4665_ (.Y(_1371_),
    .A(\main.spi.state[0] ),
    .B(net1220));
 sg13g2_nand4_1 _4666_ (.B(net1477),
    .C(\main.spi.in_bit_counter[0] ),
    .A(net700),
    .Y(_1372_),
    .D(net1339));
 sg13g2_o21ai_1 _4667_ (.B1(_1369_),
    .Y(_0241_),
    .A1(_1371_),
    .A2(net1478));
 sg13g2_nor2_1 _4668_ (.A(net1406),
    .B(net1103),
    .Y(_1373_));
 sg13g2_a21oi_1 _4669_ (.A1(net1103),
    .A2(_0863_),
    .Y(_0242_),
    .B1(_1373_));
 sg13g2_nor2_1 _4670_ (.A(net1000),
    .B(net1104),
    .Y(_1374_));
 sg13g2_a21oi_1 _4671_ (.A1(net1104),
    .A2(_0926_),
    .Y(_0243_),
    .B1(_1374_));
 sg13g2_nor2_1 _4672_ (.A(net993),
    .B(net1073),
    .Y(_1375_));
 sg13g2_a21oi_1 _4673_ (.A1(_0904_),
    .A2(net1073),
    .Y(_0244_),
    .B1(_1375_));
 sg13g2_mux2_1 _4674_ (.A0(net826),
    .A1(net771),
    .S(net1383),
    .X(_0245_));
 sg13g2_mux2_1 _4675_ (.A0(\main.adder.s3_exponent[1] ),
    .A1(net737),
    .S(net1383),
    .X(_0246_));
 sg13g2_mux2_1 _4676_ (.A0(net808),
    .A1(net765),
    .S(net1384),
    .X(_0247_));
 sg13g2_nand2_1 _4677_ (.Y(_1376_),
    .A(net1383),
    .B(net601));
 sg13g2_o21ai_1 _4678_ (.B1(_1376_),
    .Y(_0248_),
    .A1(net1385),
    .A2(_0726_));
 sg13g2_mux2_1 _4679_ (.A0(net867),
    .A1(net822),
    .S(net1384),
    .X(_0249_));
 sg13g2_mux2_1 _4680_ (.A0(net958),
    .A1(net922),
    .S(net1384),
    .X(_0250_));
 sg13g2_nand2_1 _4681_ (.Y(_1377_),
    .A(net1384),
    .B(net788));
 sg13g2_o21ai_1 _4682_ (.B1(_1377_),
    .Y(_0251_),
    .A1(net1384),
    .A2(_0727_));
 sg13g2_mux2_1 _4683_ (.A0(net1405),
    .A1(net819),
    .S(net1384),
    .X(_0252_));
 sg13g2_mux2_1 _4684_ (.A0(net950),
    .A1(net826),
    .S(net1385),
    .X(_0253_));
 sg13g2_mux2_1 _4685_ (.A0(net994),
    .A1(\main.adder.s3_exponent[1] ),
    .S(net1384),
    .X(_0254_));
 sg13g2_mux2_1 _4686_ (.A0(net1029),
    .A1(net808),
    .S(net1384),
    .X(_0255_));
 sg13g2_nor2_1 _4687_ (.A(net1391),
    .B(net809),
    .Y(_1378_));
 sg13g2_a21oi_1 _4688_ (.A1(net1391),
    .A2(_0726_),
    .Y(_0256_),
    .B1(_1378_));
 sg13g2_mux2_1 _4689_ (.A0(net967),
    .A1(net867),
    .S(net1387),
    .X(_0257_));
 sg13g2_mux2_1 _4690_ (.A0(net961),
    .A1(net958),
    .S(net1392),
    .X(_0258_));
 sg13g2_nor2_1 _4691_ (.A(net1392),
    .B(net951),
    .Y(_1379_));
 sg13g2_a21oi_1 _4692_ (.A1(net1392),
    .A2(_0727_),
    .Y(_0259_),
    .B1(_1379_));
 sg13g2_mux2_1 _4693_ (.A0(net1006),
    .A1(\main.adder.s3_exponent[7] ),
    .S(net1392),
    .X(_0260_));
 sg13g2_nand2_1 _4694_ (.Y(_1380_),
    .A(net1302),
    .B(net965));
 sg13g2_nand2b_1 _4695_ (.Y(_1381_),
    .B(\main.adder.s5_S ),
    .A_N(_0033_));
 sg13g2_o21ai_1 _4696_ (.B1(_1381_),
    .Y(_1382_),
    .A1(_0703_),
    .A2(\main.adder.s5_S ));
 sg13g2_and2_1 _4697_ (.A(\main.adder.s5_mant[0] ),
    .B(_1382_),
    .X(_1383_));
 sg13g2_and2_1 _4698_ (.A(\main.adder.s5_mant[1] ),
    .B(_1383_),
    .X(_1384_));
 sg13g2_nand3_1 _4699_ (.B(\main.adder.s5_mant[2] ),
    .C(_1384_),
    .A(\main.adder.s5_mant[3] ),
    .Y(_1385_));
 sg13g2_and4_1 _4700_ (.A(\main.adder.s5_mant[3] ),
    .B(\main.adder.s5_mant[2] ),
    .C(\main.adder.s5_mant[4] ),
    .D(_1384_),
    .X(_1386_));
 sg13g2_nand3_1 _4701_ (.B(\main.adder.s5_mant[5] ),
    .C(_1386_),
    .A(\main.adder.s5_mant[6] ),
    .Y(_1387_));
 sg13g2_and4_1 _4702_ (.A(\main.adder.s5_mant[7] ),
    .B(\main.adder.s5_mant[6] ),
    .C(\main.adder.s5_mant[5] ),
    .D(_1386_),
    .X(_1388_));
 sg13g2_nand3_1 _4703_ (.B(\main.adder.s5_mant[8] ),
    .C(_1388_),
    .A(\main.adder.s5_mant[9] ),
    .Y(_1389_));
 sg13g2_nor2_1 _4704_ (.A(_0709_),
    .B(_1389_),
    .Y(_1390_));
 sg13g2_nand3_1 _4705_ (.B(\main.adder.s5_mant[12] ),
    .C(_1390_),
    .A(\main.adder.s5_mant[11] ),
    .Y(_1391_));
 sg13g2_nor2_1 _4706_ (.A(_0710_),
    .B(_1391_),
    .Y(_1392_));
 sg13g2_nand3_1 _4707_ (.B(\main.adder.s5_mant[14] ),
    .C(_1392_),
    .A(\main.adder.s5_mant[15] ),
    .Y(_1393_));
 sg13g2_nor2_1 _4708_ (.A(_0707_),
    .B(_1393_),
    .Y(_1394_));
 sg13g2_nand3_1 _4709_ (.B(\main.adder.s5_mant[17] ),
    .C(_1394_),
    .A(\main.adder.s5_mant[18] ),
    .Y(_1395_));
 sg13g2_nor2_1 _4710_ (.A(_0704_),
    .B(_1395_),
    .Y(_1396_));
 sg13g2_and2_1 _4711_ (.A(\main.adder.s5_mant[20] ),
    .B(_1396_),
    .X(_1397_));
 sg13g2_nand2_1 _4712_ (.Y(_1398_),
    .A(\main.adder.s5_mant[21] ),
    .B(_1397_));
 sg13g2_nand4_1 _4713_ (.B(\main.adder.s5_mant[22] ),
    .C(\main.adder.s5_mant[21] ),
    .A(\main.adder.s5_mant[23] ),
    .Y(_1399_),
    .D(_1397_));
 sg13g2_nand2_2 _4714_ (.Y(_1400_),
    .A(\main.adder.s5_exponent[1] ),
    .B(\main.adder.s5_exponent[0] ));
 sg13g2_nand2_1 _4715_ (.Y(_1401_),
    .A(\main.adder.s5_exponent[3] ),
    .B(\main.adder.s5_exponent[2] ));
 sg13g2_nor2_1 _4716_ (.A(_1400_),
    .B(_1401_),
    .Y(_1402_));
 sg13g2_nor2b_1 _4717_ (.A(net1057),
    .B_N(_1402_),
    .Y(_1403_));
 sg13g2_xor2_1 _4718_ (.B(_1403_),
    .A(_0038_),
    .X(_1404_));
 sg13g2_nand4_1 _4719_ (.B(\main.adder.s5_exponent[6] ),
    .C(\main.adder.s5_exponent[5] ),
    .A(\main.adder.s5_exponent[7] ),
    .Y(_1405_),
    .D(\main.adder.s5_exponent[4] ));
 sg13g2_nand2b_1 _4720_ (.Y(_1406_),
    .B(\main.adder.s5_exponent[1] ),
    .A_N(\main.adder.s5_exponent[0] ));
 sg13g2_nor4_1 _4721_ (.A(\main.adder.s5_exponent[9] ),
    .B(\main.adder.s5_exponent[8] ),
    .C(_1401_),
    .D(_1406_),
    .Y(_1407_));
 sg13g2_nand2b_1 _4722_ (.Y(_1408_),
    .B(_1407_),
    .A_N(_1405_));
 sg13g2_o21ai_1 _4723_ (.B1(_1404_),
    .Y(_1409_),
    .A1(net1056),
    .A2(_1408_));
 sg13g2_mux2_1 _4724_ (.A0(\main.adder.s5_exponent[0] ),
    .A1(_0034_),
    .S(net1056),
    .X(_1410_));
 sg13g2_inv_1 _4725_ (.Y(_1411_),
    .A(_1410_));
 sg13g2_nand2_1 _4726_ (.Y(_1412_),
    .A(_0041_),
    .B(net1057));
 sg13g2_nand2_1 _4727_ (.Y(_1413_),
    .A(\main.adder.s5_exponent[4] ),
    .B(_1402_));
 sg13g2_nand3_1 _4728_ (.B(\main.adder.s5_exponent[4] ),
    .C(_1402_),
    .A(\main.adder.s5_exponent[5] ),
    .Y(_1414_));
 sg13g2_nor2_1 _4729_ (.A(_0040_),
    .B(_1414_),
    .Y(_1415_));
 sg13g2_xor2_1 _4730_ (.B(_1415_),
    .A(\main.adder.s5_exponent[7] ),
    .X(_1416_));
 sg13g2_o21ai_1 _4731_ (.B1(_1412_),
    .Y(_1417_),
    .A1(net1057),
    .A2(_1416_));
 sg13g2_inv_1 _4732_ (.Y(_1418_),
    .A(_1417_));
 sg13g2_xnor2_1 _4733_ (.Y(_1419_),
    .A(\main.adder.s5_exponent[2] ),
    .B(_1400_));
 sg13g2_nand2_1 _4734_ (.Y(_1420_),
    .A(_0036_),
    .B(net1056));
 sg13g2_o21ai_1 _4735_ (.B1(_1420_),
    .Y(_1421_),
    .A1(net1056),
    .A2(_1419_));
 sg13g2_inv_1 _4736_ (.Y(_1422_),
    .A(_1421_));
 sg13g2_nand2_1 _4737_ (.Y(_1423_),
    .A(_0039_),
    .B(net1057));
 sg13g2_xnor2_1 _4738_ (.Y(_1424_),
    .A(\main.adder.s5_exponent[5] ),
    .B(_1413_));
 sg13g2_o21ai_1 _4739_ (.B1(_1423_),
    .Y(_1425_),
    .A1(net1057),
    .A2(_1424_));
 sg13g2_inv_1 _4740_ (.Y(_1426_),
    .A(_1425_));
 sg13g2_xnor2_1 _4741_ (.Y(_1427_),
    .A(\main.adder.s5_exponent[6] ),
    .B(_1414_));
 sg13g2_nor2_1 _4742_ (.A(net1057),
    .B(_1427_),
    .Y(_1428_));
 sg13g2_a21oi_2 _4743_ (.B1(_1428_),
    .Y(_1429_),
    .A2(net1057),
    .A1(_0040_));
 sg13g2_xnor2_1 _4744_ (.Y(_1430_),
    .A(\main.adder.s5_exponent[1] ),
    .B(\main.adder.s5_exponent[0] ));
 sg13g2_mux2_1 _4745_ (.A0(_1430_),
    .A1(_0035_),
    .S(net1056),
    .X(_1431_));
 sg13g2_inv_1 _4746_ (.Y(_1432_),
    .A(_1431_));
 sg13g2_nor2_1 _4747_ (.A(_0036_),
    .B(_1400_),
    .Y(_1433_));
 sg13g2_xor2_1 _4748_ (.B(_1433_),
    .A(\main.adder.s5_exponent[3] ),
    .X(_1434_));
 sg13g2_nor2_1 _4749_ (.A(net1056),
    .B(_1434_),
    .Y(_1435_));
 sg13g2_a21oi_1 _4750_ (.A1(_0037_),
    .A2(net1056),
    .Y(_1436_),
    .B1(_1435_));
 sg13g2_nor4_1 _4751_ (.A(_1417_),
    .B(_1421_),
    .C(_1425_),
    .D(_1431_),
    .Y(_1437_));
 sg13g2_nand3_1 _4752_ (.B(_1429_),
    .C(_1436_),
    .A(_1411_),
    .Y(_1438_));
 sg13g2_nand3b_1 _4753_ (.B(_1409_),
    .C(_1437_),
    .Y(_1439_),
    .A_N(_1438_));
 sg13g2_nor4_1 _4754_ (.A(net1056),
    .B(_1400_),
    .C(_1401_),
    .D(_1405_),
    .Y(_1440_));
 sg13g2_xnor2_1 _4755_ (.Y(_1441_),
    .A(\main.adder.s5_exponent[8] ),
    .B(_1440_));
 sg13g2_a21oi_1 _4756_ (.A1(_1439_),
    .A2(_1441_),
    .Y(_1442_),
    .B1(net1520));
 sg13g2_nor2_1 _4757_ (.A(net828),
    .B(net1312),
    .Y(_1443_));
 sg13g2_or4_1 _4758_ (.A(\main.adder.s5_nan ),
    .B(net1312),
    .C(\main.adder.s5_inf ),
    .D(_1442_),
    .X(_1444_));
 sg13g2_xnor2_1 _4759_ (.Y(_1445_),
    .A(\main.adder.s5_mant[1] ),
    .B(_1383_));
 sg13g2_o21ai_1 _4760_ (.B1(_1380_),
    .Y(_0261_),
    .A1(net1054),
    .A2(_1445_));
 sg13g2_nand2_1 _4761_ (.Y(_1446_),
    .A(net1312),
    .B(net908));
 sg13g2_xnor2_1 _4762_ (.Y(_1447_),
    .A(\main.adder.s5_mant[2] ),
    .B(_1384_));
 sg13g2_o21ai_1 _4763_ (.B1(_1446_),
    .Y(_0262_),
    .A1(net1052),
    .A2(_1447_));
 sg13g2_nand2_1 _4764_ (.Y(_1448_),
    .A(net1302),
    .B(net998));
 sg13g2_a21o_1 _4765_ (.A2(_1384_),
    .A1(\main.adder.s5_mant[2] ),
    .B1(\main.adder.s5_mant[3] ),
    .X(_1449_));
 sg13g2_nand2_1 _4766_ (.Y(_1450_),
    .A(_1385_),
    .B(_1449_));
 sg13g2_o21ai_1 _4767_ (.B1(_1448_),
    .Y(_0263_),
    .A1(net1054),
    .A2(_1450_));
 sg13g2_nand2_1 _4768_ (.Y(_1451_),
    .A(net1312),
    .B(net1503));
 sg13g2_xor2_1 _4769_ (.B(_1385_),
    .A(\main.adder.s5_mant[4] ),
    .X(_1452_));
 sg13g2_o21ai_1 _4770_ (.B1(_1451_),
    .Y(_0264_),
    .A1(net1051),
    .A2(_1452_));
 sg13g2_nand2_1 _4771_ (.Y(_1453_),
    .A(net1302),
    .B(net920));
 sg13g2_xnor2_1 _4772_ (.Y(_1454_),
    .A(\main.adder.s5_mant[5] ),
    .B(_1386_));
 sg13g2_o21ai_1 _4773_ (.B1(_1453_),
    .Y(_0265_),
    .A1(net1054),
    .A2(_1454_));
 sg13g2_nand2_1 _4774_ (.Y(_1455_),
    .A(net1301),
    .B(net735));
 sg13g2_a21o_1 _4775_ (.A2(_1386_),
    .A1(\main.adder.s5_mant[5] ),
    .B1(\main.adder.s5_mant[6] ),
    .X(_1456_));
 sg13g2_nand2_1 _4776_ (.Y(_1457_),
    .A(_1387_),
    .B(_1456_));
 sg13g2_o21ai_1 _4777_ (.B1(_1455_),
    .Y(_0266_),
    .A1(net1050),
    .A2(_1457_));
 sg13g2_nand2_1 _4778_ (.Y(_1458_),
    .A(net1301),
    .B(net703));
 sg13g2_xor2_1 _4779_ (.B(_1387_),
    .A(\main.adder.s5_mant[7] ),
    .X(_1459_));
 sg13g2_o21ai_1 _4780_ (.B1(_1458_),
    .Y(_0267_),
    .A1(net1050),
    .A2(_1459_));
 sg13g2_nand2_1 _4781_ (.Y(_1460_),
    .A(net1301),
    .B(net672));
 sg13g2_xnor2_1 _4782_ (.Y(_1461_),
    .A(\main.adder.s5_mant[8] ),
    .B(_1388_));
 sg13g2_o21ai_1 _4783_ (.B1(_1460_),
    .Y(_0268_),
    .A1(net1050),
    .A2(_1461_));
 sg13g2_nand2_1 _4784_ (.Y(_1462_),
    .A(net1301),
    .B(net774));
 sg13g2_a21o_1 _4785_ (.A2(_1388_),
    .A1(\main.adder.s5_mant[8] ),
    .B1(\main.adder.s5_mant[9] ),
    .X(_1463_));
 sg13g2_nand2_1 _4786_ (.Y(_1464_),
    .A(_1389_),
    .B(_1463_));
 sg13g2_o21ai_1 _4787_ (.B1(_1462_),
    .Y(_0269_),
    .A1(net1050),
    .A2(_1464_));
 sg13g2_nand2_1 _4788_ (.Y(_1465_),
    .A(net1301),
    .B(net796));
 sg13g2_xnor2_1 _4789_ (.Y(_1466_),
    .A(_0709_),
    .B(_1389_));
 sg13g2_o21ai_1 _4790_ (.B1(_1465_),
    .Y(_0270_),
    .A1(net1050),
    .A2(_1466_));
 sg13g2_nand2_1 _4791_ (.Y(_1467_),
    .A(net1311),
    .B(net893));
 sg13g2_xnor2_1 _4792_ (.Y(_1468_),
    .A(\main.adder.s5_mant[11] ),
    .B(_1390_));
 sg13g2_o21ai_1 _4793_ (.B1(_1467_),
    .Y(_0271_),
    .A1(net1053),
    .A2(_1468_));
 sg13g2_nand2_1 _4794_ (.Y(_1469_),
    .A(net1301),
    .B(net841));
 sg13g2_a21o_1 _4795_ (.A2(_1390_),
    .A1(\main.adder.s5_mant[11] ),
    .B1(\main.adder.s5_mant[12] ),
    .X(_1470_));
 sg13g2_nand2_1 _4796_ (.Y(_1471_),
    .A(_1391_),
    .B(_1470_));
 sg13g2_o21ai_1 _4797_ (.B1(_1469_),
    .Y(_0272_),
    .A1(net1050),
    .A2(_1471_));
 sg13g2_nand2_1 _4798_ (.Y(_1472_),
    .A(net1311),
    .B(net837));
 sg13g2_xnor2_1 _4799_ (.Y(_1473_),
    .A(_0710_),
    .B(_1391_));
 sg13g2_o21ai_1 _4800_ (.B1(_1472_),
    .Y(_0273_),
    .A1(net1053),
    .A2(_1473_));
 sg13g2_nand2_1 _4801_ (.Y(_1474_),
    .A(net1311),
    .B(net941));
 sg13g2_xnor2_1 _4802_ (.Y(_1475_),
    .A(\main.adder.s5_mant[14] ),
    .B(_1392_));
 sg13g2_o21ai_1 _4803_ (.B1(_1474_),
    .Y(_0274_),
    .A1(net1053),
    .A2(_1475_));
 sg13g2_nand2_1 _4804_ (.Y(_1476_),
    .A(net1301),
    .B(net754));
 sg13g2_a21o_1 _4805_ (.A2(_1392_),
    .A1(\main.adder.s5_mant[14] ),
    .B1(\main.adder.s5_mant[15] ),
    .X(_1477_));
 sg13g2_nand2_1 _4806_ (.Y(_1478_),
    .A(_1393_),
    .B(_1477_));
 sg13g2_o21ai_1 _4807_ (.B1(_1476_),
    .Y(_0275_),
    .A1(net1050),
    .A2(_1478_));
 sg13g2_nand2_1 _4808_ (.Y(_1479_),
    .A(net1311),
    .B(net690));
 sg13g2_xnor2_1 _4809_ (.Y(_1480_),
    .A(_0707_),
    .B(_1393_));
 sg13g2_o21ai_1 _4810_ (.B1(_1479_),
    .Y(_0276_),
    .A1(net1053),
    .A2(_1480_));
 sg13g2_nand2_1 _4811_ (.Y(_1481_),
    .A(net1311),
    .B(net683));
 sg13g2_xnor2_1 _4812_ (.Y(_1482_),
    .A(\main.adder.s5_mant[17] ),
    .B(_1394_));
 sg13g2_o21ai_1 _4813_ (.B1(_1481_),
    .Y(_0277_),
    .A1(net1053),
    .A2(_1482_));
 sg13g2_nand2_1 _4814_ (.Y(_1483_),
    .A(net1301),
    .B(net656));
 sg13g2_a21o_1 _4815_ (.A2(_1394_),
    .A1(\main.adder.s5_mant[17] ),
    .B1(\main.adder.s5_mant[18] ),
    .X(_1484_));
 sg13g2_nand2_1 _4816_ (.Y(_1485_),
    .A(_1395_),
    .B(_1484_));
 sg13g2_o21ai_1 _4817_ (.B1(_1483_),
    .Y(_0278_),
    .A1(net1053),
    .A2(_1485_));
 sg13g2_nand2_1 _4818_ (.Y(_1486_),
    .A(net1311),
    .B(net653));
 sg13g2_xnor2_1 _4819_ (.Y(_1487_),
    .A(_0704_),
    .B(_1395_));
 sg13g2_o21ai_1 _4820_ (.B1(_1486_),
    .Y(_0279_),
    .A1(net1053),
    .A2(_1487_));
 sg13g2_nand2_1 _4821_ (.Y(_1488_),
    .A(net1312),
    .B(net676));
 sg13g2_xnor2_1 _4822_ (.Y(_1489_),
    .A(\main.adder.s5_mant[20] ),
    .B(_1396_));
 sg13g2_o21ai_1 _4823_ (.B1(_1488_),
    .Y(_0280_),
    .A1(net1051),
    .A2(_1489_));
 sg13g2_nand2_1 _4824_ (.Y(_1490_),
    .A(net1311),
    .B(net674));
 sg13g2_xnor2_1 _4825_ (.Y(_1491_),
    .A(\main.adder.s5_mant[21] ),
    .B(_1397_));
 sg13g2_o21ai_1 _4826_ (.B1(_1490_),
    .Y(_0281_),
    .A1(net1053),
    .A2(_1491_));
 sg13g2_nand2_1 _4827_ (.Y(_1492_),
    .A(net1302),
    .B(net695));
 sg13g2_xnor2_1 _4828_ (.Y(_1493_),
    .A(_0708_),
    .B(_1398_));
 sg13g2_o21ai_1 _4829_ (.B1(_1492_),
    .Y(_0282_),
    .A1(net1050),
    .A2(_1493_));
 sg13g2_nand2_1 _4830_ (.Y(_1494_),
    .A(net1319),
    .B(net1545));
 sg13g2_nor4_2 _4831_ (.A(\main.adder.s4_exponent_adjust[9] ),
    .B(\main.adder.s4_exponent_adjust[8] ),
    .C(\main.adder.s4_exponent_adjust[7] ),
    .Y(_1495_),
    .D(\main.adder.s4_exponent_adjust[6] ));
 sg13g2_or4_2 _4832_ (.A(\main.adder.s4_exponent_adjust[9] ),
    .B(\main.adder.s4_exponent_adjust[8] ),
    .C(\main.adder.s4_exponent_adjust[7] ),
    .D(\main.adder.s4_exponent_adjust[6] ),
    .X(_1496_));
 sg13g2_nor2_2 _4833_ (.A(\main.adder.s4_exponent_adjust[5] ),
    .B(_1496_),
    .Y(_1497_));
 sg13g2_nand2b_2 _4834_ (.Y(_1498_),
    .B(_1495_),
    .A_N(\main.adder.s4_exponent_adjust[5] ));
 sg13g2_nor2_2 _4835_ (.A(net1317),
    .B(_1498_),
    .Y(_1499_));
 sg13g2_nand2_1 _4836_ (.Y(_1500_),
    .A(net1394),
    .B(_1497_));
 sg13g2_nor2_1 _4837_ (.A(net1275),
    .B(_1496_),
    .Y(_1501_));
 sg13g2_nand2b_1 _4838_ (.Y(_1502_),
    .B(_1495_),
    .A_N(net1275));
 sg13g2_nor2_1 _4839_ (.A(net1319),
    .B(net1204),
    .Y(_1503_));
 sg13g2_nor2_1 _4840_ (.A(net1282),
    .B(_1496_),
    .Y(_1504_));
 sg13g2_nand2_1 _4841_ (.Y(_1505_),
    .A(_0715_),
    .B(_1495_));
 sg13g2_nor2_2 _4842_ (.A(\main.adder.s4_exponent_adjust[0] ),
    .B(_1496_),
    .Y(_1506_));
 sg13g2_nand2b_1 _4843_ (.Y(_1507_),
    .B(_1495_),
    .A_N(\main.adder.s4_exponent_adjust[0] ));
 sg13g2_nor3_2 _4844_ (.A(_0042_),
    .B(\main.adder.s4_exponent_adjust[1] ),
    .C(net1184),
    .Y(_1508_));
 sg13g2_and3_1 _4845_ (.X(_1509_),
    .A(_0716_),
    .B(net1196),
    .C(_1508_));
 sg13g2_a21oi_1 _4846_ (.A1(_1503_),
    .A2(_1509_),
    .Y(_1510_),
    .B1(_1499_));
 sg13g2_nor2_1 _4847_ (.A(\main.adder.s4_exponent_adjust[1] ),
    .B(_1496_),
    .Y(_1511_));
 sg13g2_nand2b_1 _4848_ (.Y(_1512_),
    .B(_1495_),
    .A_N(\main.adder.s4_exponent_adjust[1] ));
 sg13g2_mux4_1 _4849_ (.S0(net1190),
    .A0(\main.adder.s4_mant[21] ),
    .A1(\main.adder.s4_mant[22] ),
    .A2(\main.adder.s4_mant[23] ),
    .A3(\main.adder.s4_mant[24] ),
    .S1(net1177),
    .X(_1513_));
 sg13g2_nor2_1 _4850_ (.A(net1194),
    .B(_1513_),
    .Y(_1514_));
 sg13g2_mux4_1 _4851_ (.S0(net1191),
    .A0(_0059_),
    .A1(_0060_),
    .A2(_0061_),
    .A3(_0062_),
    .S1(net1177),
    .X(_1515_));
 sg13g2_a21oi_1 _4852_ (.A1(net1195),
    .A2(_1515_),
    .Y(_1516_),
    .B1(_1514_));
 sg13g2_nor2_1 _4853_ (.A(net1281),
    .B(_1496_),
    .Y(_1517_));
 sg13g2_nand2_1 _4854_ (.Y(_1518_),
    .A(_0716_),
    .B(_1495_));
 sg13g2_mux2_1 _4855_ (.A0(\main.adder.s4_mant[26] ),
    .A1(\main.adder.s4_mant[25] ),
    .S(net1182),
    .X(_1519_));
 sg13g2_nor2_1 _4856_ (.A(net1178),
    .B(_1519_),
    .Y(_1520_));
 sg13g2_and2_1 _4857_ (.A(\main.adder.s4_mant[28] ),
    .B(net1190),
    .X(_1521_));
 sg13g2_a21oi_1 _4858_ (.A1(\main.adder.s4_mant[27] ),
    .A2(net1183),
    .Y(_1522_),
    .B1(_1521_));
 sg13g2_a21oi_1 _4859_ (.A1(net1178),
    .A2(_1522_),
    .Y(_1523_),
    .B1(_1520_));
 sg13g2_mux2_1 _4860_ (.A0(\main.adder.s4_mant[30] ),
    .A1(\main.adder.s4_mant[29] ),
    .S(net1182),
    .X(_1524_));
 sg13g2_mux2_1 _4861_ (.A0(\main.adder.s4_mant[32] ),
    .A1(\main.adder.s4_mant[31] ),
    .S(net1182),
    .X(_1525_));
 sg13g2_mux2_1 _4862_ (.A0(_1524_),
    .A1(_1525_),
    .S(net1178),
    .X(_1526_));
 sg13g2_mux2_1 _4863_ (.A0(_1523_),
    .A1(_1526_),
    .S(net1198),
    .X(_1527_));
 sg13g2_and2_1 _4864_ (.A(_0048_),
    .B(net1185),
    .X(_1528_));
 sg13g2_a21oi_1 _4865_ (.A1(_0047_),
    .A2(net1184),
    .Y(_1529_),
    .B1(_1528_));
 sg13g2_mux2_1 _4866_ (.A0(_0049_),
    .A1(_0050_),
    .S(net1185),
    .X(_1530_));
 sg13g2_nor2_1 _4867_ (.A(net1171),
    .B(_1530_),
    .Y(_1531_));
 sg13g2_a21oi_2 _4868_ (.B1(_1531_),
    .Y(_1532_),
    .A2(_1529_),
    .A1(net1171));
 sg13g2_mux2_1 _4869_ (.A0(_0043_),
    .A1(_0044_),
    .S(net1186),
    .X(_1533_));
 sg13g2_mux2_1 _4870_ (.A0(_0045_),
    .A1(_0046_),
    .S(net1185),
    .X(_1534_));
 sg13g2_mux2_1 _4871_ (.A0(_1533_),
    .A1(_1534_),
    .S(net1181),
    .X(_1535_));
 sg13g2_mux2_1 _4872_ (.A0(_1532_),
    .A1(_1535_),
    .S(net1192),
    .X(_1536_));
 sg13g2_mux4_1 _4873_ (.S0(_1506_),
    .A0(_0055_),
    .A1(_0056_),
    .A2(_0057_),
    .A3(_0058_),
    .S1(net1175),
    .X(_1537_));
 sg13g2_mux4_1 _4874_ (.S0(net1187),
    .A0(_0051_),
    .A1(_0052_),
    .A2(_0053_),
    .A3(_0054_),
    .S1(net1175),
    .X(_1538_));
 sg13g2_mux2_1 _4875_ (.A0(_1537_),
    .A1(_1538_),
    .S(net1192),
    .X(_1539_));
 sg13g2_or2_1 _4876_ (.X(_1540_),
    .B(_1539_),
    .A(net1161));
 sg13g2_o21ai_1 _4877_ (.B1(_1540_),
    .Y(_1541_),
    .A1(net1166),
    .A2(_1536_));
 sg13g2_a22oi_1 _4878_ (.Y(_1542_),
    .B1(net1167),
    .B2(_1527_),
    .A2(_1516_),
    .A1(net1279));
 sg13g2_o21ai_1 _4879_ (.B1(_1497_),
    .Y(_1543_),
    .A1(net1275),
    .A2(_1542_));
 sg13g2_a21oi_1 _4880_ (.A1(net1275),
    .A2(_1541_),
    .Y(_1544_),
    .B1(_1543_));
 sg13g2_o21ai_1 _4881_ (.B1(_1494_),
    .Y(_0283_),
    .A1(_1510_),
    .A2(_1544_));
 sg13g2_nand2_1 _4882_ (.Y(_1545_),
    .A(net1319),
    .B(net940));
 sg13g2_mux2_1 _4883_ (.A0(_0042_),
    .A1(_0043_),
    .S(net1186),
    .X(_1546_));
 sg13g2_nor2_1 _4884_ (.A(net1171),
    .B(_1546_),
    .Y(_1547_));
 sg13g2_nor4_2 _4885_ (.A(net1281),
    .B(net1192),
    .C(net1171),
    .Y(_1548_),
    .D(_1546_));
 sg13g2_a21oi_1 _4886_ (.A1(_1503_),
    .A2(_1548_),
    .Y(_1549_),
    .B1(_1499_));
 sg13g2_mux4_1 _4887_ (.S0(net1177),
    .A0(\main.adder.s4_mant[22] ),
    .A1(\main.adder.s4_mant[24] ),
    .A2(\main.adder.s4_mant[23] ),
    .A3(\main.adder.s4_mant[25] ),
    .S1(net1189),
    .X(_1550_));
 sg13g2_nor2_1 _4888_ (.A(net1194),
    .B(_1550_),
    .Y(_1551_));
 sg13g2_mux4_1 _4889_ (.S0(net1191),
    .A0(_0060_),
    .A1(_0061_),
    .A2(_0062_),
    .A3(_0063_),
    .S1(net1177),
    .X(_1552_));
 sg13g2_a21oi_2 _4890_ (.B1(_1551_),
    .Y(_1553_),
    .A2(_1552_),
    .A1(net1194));
 sg13g2_mux2_1 _4891_ (.A0(\main.adder.s4_mant[26] ),
    .A1(\main.adder.s4_mant[27] ),
    .S(net1189),
    .X(_1554_));
 sg13g2_nor2_1 _4892_ (.A(net1178),
    .B(_1554_),
    .Y(_1555_));
 sg13g2_and2_1 _4893_ (.A(\main.adder.s4_mant[29] ),
    .B(net1189),
    .X(_1556_));
 sg13g2_a21oi_1 _4894_ (.A1(\main.adder.s4_mant[28] ),
    .A2(net1183),
    .Y(_1557_),
    .B1(_1556_));
 sg13g2_a21oi_1 _4895_ (.A1(net1178),
    .A2(_1557_),
    .Y(_1558_),
    .B1(_1555_));
 sg13g2_mux2_1 _4896_ (.A0(\main.adder.s4_mant[30] ),
    .A1(\main.adder.s4_mant[31] ),
    .S(net1189),
    .X(_1559_));
 sg13g2_mux2_1 _4897_ (.A0(\main.adder.s4_mant[32] ),
    .A1(\main.adder.s4_mant[33] ),
    .S(net1189),
    .X(_1560_));
 sg13g2_mux2_1 _4898_ (.A0(_1559_),
    .A1(_1560_),
    .S(net1178),
    .X(_1561_));
 sg13g2_mux2_1 _4899_ (.A0(_1558_),
    .A1(_1561_),
    .S(net1198),
    .X(_1562_));
 sg13g2_a22oi_1 _4900_ (.Y(_1563_),
    .B1(_1562_),
    .B2(net1167),
    .A2(_1553_),
    .A1(net1279));
 sg13g2_nor2_1 _4901_ (.A(net1276),
    .B(_1563_),
    .Y(_1564_));
 sg13g2_and2_1 _4902_ (.A(_0049_),
    .B(net1185),
    .X(_1565_));
 sg13g2_a21oi_1 _4903_ (.A1(_0048_),
    .A2(net1184),
    .Y(_1566_),
    .B1(_1565_));
 sg13g2_mux2_1 _4904_ (.A0(_0050_),
    .A1(_0051_),
    .S(net1185),
    .X(_1567_));
 sg13g2_nor2_1 _4905_ (.A(net1171),
    .B(_1567_),
    .Y(_1568_));
 sg13g2_a21oi_1 _4906_ (.A1(net1171),
    .A2(_1566_),
    .Y(_1569_),
    .B1(_1568_));
 sg13g2_mux2_1 _4907_ (.A0(_0044_),
    .A1(_0045_),
    .S(net1186),
    .X(_1570_));
 sg13g2_mux2_1 _4908_ (.A0(_0046_),
    .A1(_0047_),
    .S(net1185),
    .X(_1571_));
 sg13g2_mux2_1 _4909_ (.A0(_1570_),
    .A1(_1571_),
    .S(net1181),
    .X(_1572_));
 sg13g2_mux2_1 _4910_ (.A0(_1569_),
    .A1(_1572_),
    .S(net1192),
    .X(_1573_));
 sg13g2_mux4_1 _4911_ (.S0(net1188),
    .A0(_0056_),
    .A1(_0057_),
    .A2(_0058_),
    .A3(_0059_),
    .S1(net1175),
    .X(_1574_));
 sg13g2_mux4_1 _4912_ (.S0(net1187),
    .A0(_0052_),
    .A1(_0053_),
    .A2(_0054_),
    .A3(_0055_),
    .S1(net1175),
    .X(_1575_));
 sg13g2_mux2_1 _4913_ (.A0(_1574_),
    .A1(_1575_),
    .S(net1193),
    .X(_1576_));
 sg13g2_mux2_1 _4914_ (.A0(_1573_),
    .A1(_1576_),
    .S(net1166),
    .X(_1577_));
 sg13g2_o21ai_1 _4915_ (.B1(_1497_),
    .Y(_1578_),
    .A1(net1207),
    .A2(_1577_));
 sg13g2_nor2_1 _4916_ (.A(_1564_),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_o21ai_1 _4917_ (.B1(_1545_),
    .Y(_0284_),
    .A1(_1549_),
    .A2(_1579_));
 sg13g2_nand3b_1 _4918_ (.B(\main.adder.s4_exponent_adjust[1] ),
    .C(net1186),
    .Y(_1580_),
    .A_N(_0042_));
 sg13g2_o21ai_1 _4919_ (.B1(_1580_),
    .Y(_1581_),
    .A1(net1171),
    .A2(_1533_));
 sg13g2_and2_1 _4920_ (.A(net1197),
    .B(_1581_),
    .X(_1582_));
 sg13g2_and2_1 _4921_ (.A(_0716_),
    .B(_1582_),
    .X(_1583_));
 sg13g2_a21o_1 _4922_ (.A2(_1583_),
    .A1(_1503_),
    .B1(_1499_),
    .X(_1584_));
 sg13g2_mux4_1 _4923_ (.S0(net1173),
    .A0(\main.adder.s4_mant[26] ),
    .A1(\main.adder.s4_mant[24] ),
    .A2(\main.adder.s4_mant[25] ),
    .A3(\main.adder.s4_mant[23] ),
    .S1(net1182),
    .X(_1585_));
 sg13g2_mux4_1 _4924_ (.S0(net1191),
    .A0(_0717_),
    .A1(_0718_),
    .A2(\main.adder.s4_mant[21] ),
    .A3(\main.adder.s4_mant[22] ),
    .S1(net1177),
    .X(_1586_));
 sg13g2_mux2_1 _4925_ (.A0(_1585_),
    .A1(_1586_),
    .S(net1195),
    .X(_1587_));
 sg13g2_nor2_1 _4926_ (.A(net1173),
    .B(_1524_),
    .Y(_1588_));
 sg13g2_a21oi_1 _4927_ (.A1(net1172),
    .A2(_1522_),
    .Y(_1589_),
    .B1(_1588_));
 sg13g2_mux2_1 _4928_ (.A0(\main.adder.s4_mant[34] ),
    .A1(\main.adder.s4_mant[33] ),
    .S(net1182),
    .X(_1590_));
 sg13g2_mux2_1 _4929_ (.A0(_1525_),
    .A1(_1590_),
    .S(net1179),
    .X(_1591_));
 sg13g2_mux2_1 _4930_ (.A0(_1589_),
    .A1(_1591_),
    .S(net1200),
    .X(_1592_));
 sg13g2_a22oi_1 _4931_ (.Y(_1593_),
    .B1(_1592_),
    .B2(net1168),
    .A2(_1587_),
    .A1(net1279));
 sg13g2_nor2_1 _4932_ (.A(net1276),
    .B(_1593_),
    .Y(_1594_));
 sg13g2_mux4_1 _4933_ (.S0(net1185),
    .A0(_0049_),
    .A1(_0050_),
    .A2(_0051_),
    .A3(_0052_),
    .S1(net1175),
    .X(_1595_));
 sg13g2_and2_1 _4934_ (.A(net1197),
    .B(_1595_),
    .X(_1596_));
 sg13g2_nor2_1 _4935_ (.A(net1181),
    .B(_1534_),
    .Y(_1597_));
 sg13g2_a21oi_1 _4936_ (.A1(net1176),
    .A2(_1529_),
    .Y(_1598_),
    .B1(_1597_));
 sg13g2_a21oi_1 _4937_ (.A1(net1192),
    .A2(_1598_),
    .Y(_1599_),
    .B1(_1596_));
 sg13g2_mux4_1 _4938_ (.S0(net1188),
    .A0(_0057_),
    .A1(_0058_),
    .A2(_0059_),
    .A3(_0060_),
    .S1(net1175),
    .X(_1600_));
 sg13g2_mux4_1 _4939_ (.S0(net1187),
    .A0(_0053_),
    .A1(_0054_),
    .A2(_0055_),
    .A3(_0056_),
    .S1(net1175),
    .X(_1601_));
 sg13g2_mux2_1 _4940_ (.A0(_1600_),
    .A1(_1601_),
    .S(net1193),
    .X(_1602_));
 sg13g2_nor2_1 _4941_ (.A(net1161),
    .B(_1602_),
    .Y(_1603_));
 sg13g2_a21oi_1 _4942_ (.A1(net1161),
    .A2(_1599_),
    .Y(_1604_),
    .B1(_1603_));
 sg13g2_o21ai_1 _4943_ (.B1(_1497_),
    .Y(_1605_),
    .A1(net1207),
    .A2(_1604_));
 sg13g2_o21ai_1 _4944_ (.B1(_1584_),
    .Y(_1606_),
    .A1(_1594_),
    .A2(_1605_));
 sg13g2_o21ai_1 _4945_ (.B1(_1606_),
    .Y(_0285_),
    .A1(net1392),
    .A2(_0709_));
 sg13g2_mux4_1 _4946_ (.S0(net1190),
    .A0(_0718_),
    .A1(_0719_),
    .A2(\main.adder.s4_mant[22] ),
    .A3(\main.adder.s4_mant[23] ),
    .S1(net1177),
    .X(_1607_));
 sg13g2_mux4_1 _4947_ (.S0(net1189),
    .A0(\main.adder.s4_mant[26] ),
    .A1(\main.adder.s4_mant[27] ),
    .A2(\main.adder.s4_mant[24] ),
    .A3(\main.adder.s4_mant[25] ),
    .S1(net1173),
    .X(_1608_));
 sg13g2_mux2_1 _4948_ (.A0(_1607_),
    .A1(_1608_),
    .S(net1200),
    .X(_1609_));
 sg13g2_nor2_1 _4949_ (.A(net1172),
    .B(_1559_),
    .Y(_1610_));
 sg13g2_a21oi_1 _4950_ (.A1(net1173),
    .A2(_1557_),
    .Y(_1611_),
    .B1(_1610_));
 sg13g2_mux2_1 _4951_ (.A0(\main.adder.s4_mant[34] ),
    .A1(\main.adder.s4_mant[35] ),
    .S(net1190),
    .X(_1612_));
 sg13g2_mux2_1 _4952_ (.A0(_1560_),
    .A1(_1612_),
    .S(net1178),
    .X(_1613_));
 sg13g2_mux2_1 _4953_ (.A0(_1611_),
    .A1(_1613_),
    .S(net1200),
    .X(_1614_));
 sg13g2_nand2_1 _4954_ (.Y(_1615_),
    .A(net1168),
    .B(_1614_));
 sg13g2_a21oi_1 _4955_ (.A1(net1279),
    .A2(_1609_),
    .Y(_1616_),
    .B1(net1202));
 sg13g2_mux4_1 _4956_ (.S0(net1185),
    .A0(_0050_),
    .A1(_0051_),
    .A2(_0052_),
    .A3(_0053_),
    .S1(net1175),
    .X(_1617_));
 sg13g2_and2_1 _4957_ (.A(net1197),
    .B(_1617_),
    .X(_1618_));
 sg13g2_nor2_1 _4958_ (.A(net1176),
    .B(_1571_),
    .Y(_1619_));
 sg13g2_a21oi_2 _4959_ (.B1(_1619_),
    .Y(_1620_),
    .A2(_1566_),
    .A1(net1176));
 sg13g2_a21oi_2 _4960_ (.B1(_1618_),
    .Y(_1621_),
    .A2(_1620_),
    .A1(net1192));
 sg13g2_mux4_1 _4961_ (.S0(net1188),
    .A0(_0058_),
    .A1(_0059_),
    .A2(_0060_),
    .A3(_0061_),
    .S1(net1177),
    .X(_1622_));
 sg13g2_mux4_1 _4962_ (.S0(net1188),
    .A0(_0054_),
    .A1(_0055_),
    .A2(_0056_),
    .A3(_0057_),
    .S1(net1176),
    .X(_1623_));
 sg13g2_mux2_1 _4963_ (.A0(_1622_),
    .A1(_1623_),
    .S(net1194),
    .X(_1624_));
 sg13g2_nor2_1 _4964_ (.A(net1162),
    .B(_1624_),
    .Y(_1625_));
 sg13g2_a21oi_1 _4965_ (.A1(net1162),
    .A2(_1621_),
    .Y(_1626_),
    .B1(_1625_));
 sg13g2_a221oi_1 _4966_ (.B2(net1202),
    .C1(net1132),
    .B1(_1626_),
    .A1(_1615_),
    .Y(_1627_),
    .A2(_1616_));
 sg13g2_nand2_1 _4967_ (.Y(_1628_),
    .A(net1317),
    .B(net1621));
 sg13g2_mux2_1 _4968_ (.A0(_1546_),
    .A1(_1570_),
    .S(net1176),
    .X(_1629_));
 sg13g2_nor2_1 _4969_ (.A(net1192),
    .B(_1629_),
    .Y(_1630_));
 sg13g2_nand2_1 _4970_ (.Y(_1631_),
    .A(_0716_),
    .B(_1630_));
 sg13g2_nand2_2 _4971_ (.Y(_1632_),
    .A(\main.adder.s4_exponent_adjust[5] ),
    .B(net1207));
 sg13g2_nor2_1 _4972_ (.A(net1317),
    .B(_1632_),
    .Y(_1633_));
 sg13g2_nand3_1 _4973_ (.B(\main.adder.s4_exponent_adjust[5] ),
    .C(net1207),
    .A(net1393),
    .Y(_1634_));
 sg13g2_o21ai_1 _4974_ (.B1(_1628_),
    .Y(_1635_),
    .A1(_1631_),
    .A2(_1634_));
 sg13g2_or2_1 _4975_ (.X(_0286_),
    .B(_1635_),
    .A(_1627_));
 sg13g2_mux2_1 _4976_ (.A0(_1513_),
    .A1(_1523_),
    .S(net1198),
    .X(_1636_));
 sg13g2_a21oi_1 _4977_ (.A1(net1278),
    .A2(_1636_),
    .Y(_1637_),
    .B1(net1203));
 sg13g2_or2_1 _4978_ (.X(_1638_),
    .B(_1526_),
    .A(net1198));
 sg13g2_mux2_1 _4979_ (.A0(\main.adder.s4_mant[36] ),
    .A1(\main.adder.s4_mant[35] ),
    .S(net1182),
    .X(_1639_));
 sg13g2_mux2_1 _4980_ (.A0(_1590_),
    .A1(_1639_),
    .S(net1179),
    .X(_1640_));
 sg13g2_o21ai_1 _4981_ (.B1(_1638_),
    .Y(_1641_),
    .A1(net1195),
    .A2(_1640_));
 sg13g2_o21ai_1 _4982_ (.B1(_1637_),
    .Y(_1642_),
    .A1(net1278),
    .A2(_1641_));
 sg13g2_mux2_1 _4983_ (.A0(_1532_),
    .A1(_1538_),
    .S(net1197),
    .X(_1643_));
 sg13g2_mux2_1 _4984_ (.A0(_1515_),
    .A1(_1537_),
    .S(net1193),
    .X(_1644_));
 sg13g2_mux2_1 _4985_ (.A0(_1643_),
    .A1(_1644_),
    .S(net1164),
    .X(_1645_));
 sg13g2_a21oi_1 _4986_ (.A1(net1202),
    .A2(_1645_),
    .Y(_1646_),
    .B1(net1132));
 sg13g2_nor2_1 _4987_ (.A(net1196),
    .B(_1508_),
    .Y(_1647_));
 sg13g2_a21oi_1 _4988_ (.A1(net1196),
    .A2(_1535_),
    .Y(_1648_),
    .B1(_1647_));
 sg13g2_nand2_1 _4989_ (.Y(_1649_),
    .A(net1165),
    .B(_1648_));
 sg13g2_a22oi_1 _4990_ (.Y(_1650_),
    .B1(_1642_),
    .B2(_1646_),
    .A2(net1598),
    .A1(net1321));
 sg13g2_o21ai_1 _4991_ (.B1(_1650_),
    .Y(_0287_),
    .A1(_1634_),
    .A2(_1649_));
 sg13g2_mux2_1 _4992_ (.A0(_1550_),
    .A1(_1558_),
    .S(net1198),
    .X(_1651_));
 sg13g2_a21oi_1 _4993_ (.A1(net1278),
    .A2(_1651_),
    .Y(_1652_),
    .B1(net1203));
 sg13g2_or2_1 _4994_ (.X(_1653_),
    .B(_1561_),
    .A(net1198));
 sg13g2_mux2_1 _4995_ (.A0(\main.adder.s4_mant[36] ),
    .A1(\main.adder.s4_mant[37] ),
    .S(net1189),
    .X(_1654_));
 sg13g2_mux2_1 _4996_ (.A0(_1612_),
    .A1(_1654_),
    .S(net1179),
    .X(_1655_));
 sg13g2_o21ai_1 _4997_ (.B1(_1653_),
    .Y(_1656_),
    .A1(net1195),
    .A2(_1655_));
 sg13g2_o21ai_1 _4998_ (.B1(_1652_),
    .Y(_1657_),
    .A1(net1278),
    .A2(_1656_));
 sg13g2_mux2_1 _4999_ (.A0(_1569_),
    .A1(_1575_),
    .S(net1197),
    .X(_1658_));
 sg13g2_mux2_1 _5000_ (.A0(_1552_),
    .A1(_1574_),
    .S(net1194),
    .X(_1659_));
 sg13g2_mux2_1 _5001_ (.A0(_1658_),
    .A1(_1659_),
    .S(net1165),
    .X(_1660_));
 sg13g2_a21oi_1 _5002_ (.A1(net1202),
    .A2(_1660_),
    .Y(_1661_),
    .B1(net1132));
 sg13g2_nand2_1 _5003_ (.Y(_1662_),
    .A(net1196),
    .B(_1572_));
 sg13g2_o21ai_1 _5004_ (.B1(_1662_),
    .Y(_1663_),
    .A1(net1196),
    .A2(_1547_));
 sg13g2_or2_1 _5005_ (.X(_1664_),
    .B(_1663_),
    .A(net1162));
 sg13g2_a22oi_1 _5006_ (.Y(_1665_),
    .B1(_1657_),
    .B2(_1661_),
    .A2(net1572),
    .A1(net1321));
 sg13g2_o21ai_1 _5007_ (.B1(_1665_),
    .Y(_0288_),
    .A1(_1634_),
    .A2(_1664_));
 sg13g2_mux2_1 _5008_ (.A0(_1585_),
    .A1(_1589_),
    .S(net1200),
    .X(_1666_));
 sg13g2_mux2_1 _5009_ (.A0(\main.adder.s4_mant[38] ),
    .A1(\main.adder.s4_mant[37] ),
    .S(net1182),
    .X(_1667_));
 sg13g2_mux2_1 _5010_ (.A0(_1639_),
    .A1(_1667_),
    .S(net1179),
    .X(_1668_));
 sg13g2_mux2_1 _5011_ (.A0(_1591_),
    .A1(_1668_),
    .S(net1201),
    .X(_1669_));
 sg13g2_nand2_1 _5012_ (.Y(_1670_),
    .A(net1168),
    .B(_1669_));
 sg13g2_a21oi_1 _5013_ (.A1(net1278),
    .A2(_1666_),
    .Y(_1671_),
    .B1(net1202));
 sg13g2_mux2_1 _5014_ (.A0(_1595_),
    .A1(_1601_),
    .S(net1197),
    .X(_1672_));
 sg13g2_nand2_1 _5015_ (.Y(_1673_),
    .A(net1194),
    .B(_1600_));
 sg13g2_o21ai_1 _5016_ (.B1(_1673_),
    .Y(_1674_),
    .A1(net1195),
    .A2(_1586_));
 sg13g2_mux2_1 _5017_ (.A0(_1672_),
    .A1(_1674_),
    .S(net1164),
    .X(_1675_));
 sg13g2_a221oi_1 _5018_ (.B2(net1202),
    .C1(net1132),
    .B1(_1675_),
    .A1(_1670_),
    .Y(_1676_),
    .A2(_1671_));
 sg13g2_nand2_1 _5019_ (.Y(_1677_),
    .A(net1317),
    .B(net1620));
 sg13g2_nor2_1 _5020_ (.A(net1196),
    .B(_1581_),
    .Y(_1678_));
 sg13g2_a21oi_1 _5021_ (.A1(net1196),
    .A2(_1598_),
    .Y(_1679_),
    .B1(_1678_));
 sg13g2_nand2_1 _5022_ (.Y(_1680_),
    .A(net1165),
    .B(_1679_));
 sg13g2_o21ai_1 _5023_ (.B1(_1677_),
    .Y(_1681_),
    .A1(_1634_),
    .A2(_1680_));
 sg13g2_or2_1 _5024_ (.X(_0289_),
    .B(_1681_),
    .A(_1676_));
 sg13g2_mux2_1 _5025_ (.A0(_1608_),
    .A1(_1611_),
    .S(net1200),
    .X(_1682_));
 sg13g2_mux2_1 _5026_ (.A0(\main.adder.s4_mant[38] ),
    .A1(\main.adder.s4_mant[39] ),
    .S(net1189),
    .X(_1683_));
 sg13g2_mux2_1 _5027_ (.A0(_1654_),
    .A1(_1683_),
    .S(net1178),
    .X(_1684_));
 sg13g2_mux2_1 _5028_ (.A0(_1613_),
    .A1(_1684_),
    .S(net1200),
    .X(_1685_));
 sg13g2_mux2_1 _5029_ (.A0(_1682_),
    .A1(_1685_),
    .S(net1168),
    .X(_1686_));
 sg13g2_mux2_1 _5030_ (.A0(_1617_),
    .A1(_1623_),
    .S(net1197),
    .X(_1687_));
 sg13g2_nand2b_1 _5031_ (.Y(_1688_),
    .B(net1162),
    .A_N(_1687_));
 sg13g2_nand2_1 _5032_ (.Y(_1689_),
    .A(net1194),
    .B(_1622_));
 sg13g2_o21ai_1 _5033_ (.B1(_1689_),
    .Y(_1690_),
    .A1(net1195),
    .A2(_1607_));
 sg13g2_o21ai_1 _5034_ (.B1(_1688_),
    .Y(_1691_),
    .A1(net1162),
    .A2(_1690_));
 sg13g2_nor2_1 _5035_ (.A(net1208),
    .B(_1691_),
    .Y(_1692_));
 sg13g2_o21ai_1 _5036_ (.B1(_1499_),
    .Y(_1693_),
    .A1(net1205),
    .A2(_1686_));
 sg13g2_mux2_1 _5037_ (.A0(_1620_),
    .A1(_1629_),
    .S(net1192),
    .X(_1694_));
 sg13g2_nor2_2 _5038_ (.A(net1161),
    .B(_1694_),
    .Y(_1695_));
 sg13g2_a22oi_1 _5039_ (.Y(_1696_),
    .B1(_1633_),
    .B2(_1695_),
    .A2(net1599),
    .A1(net1317));
 sg13g2_o21ai_1 _5040_ (.B1(_1696_),
    .Y(_0290_),
    .A1(_1692_),
    .A2(_1693_));
 sg13g2_nor2_1 _5041_ (.A(net1177),
    .B(_1667_),
    .Y(_1697_));
 sg13g2_and2_1 _5042_ (.A(\main.adder.s4_mant[40] ),
    .B(net1190),
    .X(_1698_));
 sg13g2_a21oi_1 _5043_ (.A1(\main.adder.s4_mant[39] ),
    .A2(net1182),
    .Y(_1699_),
    .B1(_1698_));
 sg13g2_a21oi_1 _5044_ (.A1(net1179),
    .A2(_1699_),
    .Y(_1700_),
    .B1(_1697_));
 sg13g2_nor2_1 _5045_ (.A(net1198),
    .B(_1640_),
    .Y(_1701_));
 sg13g2_o21ai_1 _5046_ (.B1(net1169),
    .Y(_1702_),
    .A1(\main.adder.s4_exponent_adjust[2] ),
    .A2(_1700_));
 sg13g2_a21oi_1 _5047_ (.A1(net1163),
    .A2(_1527_),
    .Y(_1703_),
    .B1(net1203));
 sg13g2_o21ai_1 _5048_ (.B1(_1703_),
    .Y(_1704_),
    .A1(_1701_),
    .A2(_1702_));
 sg13g2_nor2_1 _5049_ (.A(net1164),
    .B(_1539_),
    .Y(_1705_));
 sg13g2_a21oi_2 _5050_ (.B1(_1705_),
    .Y(_1706_),
    .A2(net1164),
    .A1(_1516_));
 sg13g2_a21oi_1 _5051_ (.A1(net1275),
    .A2(_1706_),
    .Y(_1707_),
    .B1(_1498_));
 sg13g2_nand2_1 _5052_ (.Y(_1708_),
    .A(_1704_),
    .B(_1707_));
 sg13g2_nand3_1 _5053_ (.B(net1196),
    .C(_1508_),
    .A(net1280),
    .Y(_1709_));
 sg13g2_o21ai_1 _5054_ (.B1(_1709_),
    .Y(_1710_),
    .A1(net1161),
    .A2(_1536_));
 sg13g2_nor2b_1 _5055_ (.A(_1632_),
    .B_N(_1710_),
    .Y(_1711_));
 sg13g2_nor2_1 _5056_ (.A(net1317),
    .B(_1711_),
    .Y(_1712_));
 sg13g2_a22oi_1 _5057_ (.Y(_0291_),
    .B1(_1708_),
    .B2(_1712_),
    .A2(_0707_),
    .A1(net1318));
 sg13g2_nor2_1 _5058_ (.A(net1180),
    .B(_1683_),
    .Y(_1713_));
 sg13g2_and2_1 _5059_ (.A(\main.adder.s4_mant[41] ),
    .B(net1191),
    .X(_1714_));
 sg13g2_a21oi_1 _5060_ (.A1(\main.adder.s4_mant[40] ),
    .A2(net1183),
    .Y(_1715_),
    .B1(_1714_));
 sg13g2_a21oi_1 _5061_ (.A1(net1179),
    .A2(_1715_),
    .Y(_1716_),
    .B1(_1713_));
 sg13g2_nor2_1 _5062_ (.A(net1198),
    .B(_1655_),
    .Y(_1717_));
 sg13g2_o21ai_1 _5063_ (.B1(net1169),
    .Y(_1718_),
    .A1(net1282),
    .A2(_1716_));
 sg13g2_a21oi_1 _5064_ (.A1(net1162),
    .A2(_1562_),
    .Y(_1719_),
    .B1(net1203));
 sg13g2_o21ai_1 _5065_ (.B1(_1719_),
    .Y(_1720_),
    .A1(_1717_),
    .A2(_1718_));
 sg13g2_nor2_1 _5066_ (.A(net1166),
    .B(_1576_),
    .Y(_1721_));
 sg13g2_a21oi_2 _5067_ (.B1(_1721_),
    .Y(_1722_),
    .A2(_1553_),
    .A1(net1164));
 sg13g2_a21oi_1 _5068_ (.A1(net1276),
    .A2(_1722_),
    .Y(_1723_),
    .B1(_1498_));
 sg13g2_nand2_1 _5069_ (.Y(_1724_),
    .A(_1720_),
    .B(_1723_));
 sg13g2_nand3_1 _5070_ (.B(net1201),
    .C(_1547_),
    .A(net1280),
    .Y(_1725_));
 sg13g2_o21ai_1 _5071_ (.B1(_1725_),
    .Y(_1726_),
    .A1(net1161),
    .A2(_1573_));
 sg13g2_nor2b_1 _5072_ (.A(_1632_),
    .B_N(_1726_),
    .Y(_1727_));
 sg13g2_nor2_1 _5073_ (.A(net1319),
    .B(_1727_),
    .Y(_1728_));
 sg13g2_a22oi_1 _5074_ (.Y(_0292_),
    .B1(_1724_),
    .B2(_1728_),
    .A2(_0706_),
    .A1(net1319));
 sg13g2_nand2_1 _5075_ (.Y(_1729_),
    .A(net1172),
    .B(_1699_));
 sg13g2_mux2_1 _5076_ (.A0(\main.adder.s4_mant[42] ),
    .A1(\main.adder.s4_mant[41] ),
    .S(net1183),
    .X(_1730_));
 sg13g2_o21ai_1 _5077_ (.B1(_1729_),
    .Y(_1731_),
    .A1(net1172),
    .A2(_1730_));
 sg13g2_a21oi_1 _5078_ (.A1(_0715_),
    .A2(_1731_),
    .Y(_1732_),
    .B1(net1162));
 sg13g2_o21ai_1 _5079_ (.B1(_1732_),
    .Y(_1733_),
    .A1(net1200),
    .A2(_1668_));
 sg13g2_a21oi_1 _5080_ (.A1(net1163),
    .A2(_1592_),
    .Y(_1734_),
    .B1(net1202));
 sg13g2_nor2_1 _5081_ (.A(net1164),
    .B(_1602_),
    .Y(_1735_));
 sg13g2_a21oi_2 _5082_ (.B1(_1735_),
    .Y(_1736_),
    .A2(_1587_),
    .A1(net1164));
 sg13g2_a221oi_1 _5083_ (.B2(net1275),
    .C1(_1498_),
    .B1(_1736_),
    .A1(_1733_),
    .Y(_1737_),
    .A2(_1734_));
 sg13g2_a22oi_1 _5084_ (.Y(_1738_),
    .B1(_1599_),
    .B2(net1166),
    .A2(_1582_),
    .A1(net1280));
 sg13g2_o21ai_1 _5085_ (.B1(net1393),
    .Y(_1739_),
    .A1(_1632_),
    .A2(_1738_));
 sg13g2_nor2_1 _5086_ (.A(_1737_),
    .B(_1739_),
    .Y(_1740_));
 sg13g2_a21oi_1 _5087_ (.A1(net1313),
    .A2(_0705_),
    .Y(_0293_),
    .B1(_1740_));
 sg13g2_mux2_1 _5088_ (.A0(\main.adder.s4_mant[42] ),
    .A1(\main.adder.s4_mant[43] ),
    .S(net1191),
    .X(_1741_));
 sg13g2_nor2_1 _5089_ (.A(net1172),
    .B(_1741_),
    .Y(_1742_));
 sg13g2_a21oi_1 _5090_ (.A1(net1172),
    .A2(_1715_),
    .Y(_1743_),
    .B1(_1742_));
 sg13g2_nor2_1 _5091_ (.A(net1199),
    .B(_1684_),
    .Y(_1744_));
 sg13g2_o21ai_1 _5092_ (.B1(net1169),
    .Y(_1745_),
    .A1(net1282),
    .A2(_1743_));
 sg13g2_a21oi_1 _5093_ (.A1(net1163),
    .A2(_1614_),
    .Y(_1746_),
    .B1(net1203));
 sg13g2_o21ai_1 _5094_ (.B1(_1746_),
    .Y(_1747_),
    .A1(_1744_),
    .A2(_1745_));
 sg13g2_nor2_1 _5095_ (.A(net1167),
    .B(_1624_),
    .Y(_1748_));
 sg13g2_a21oi_1 _5096_ (.A1(net1168),
    .A2(_1609_),
    .Y(_1749_),
    .B1(_1748_));
 sg13g2_a21oi_1 _5097_ (.A1(net1275),
    .A2(_1749_),
    .Y(_1750_),
    .B1(_1498_));
 sg13g2_nand2_1 _5098_ (.Y(_1751_),
    .A(_1747_),
    .B(_1750_));
 sg13g2_a22oi_1 _5099_ (.Y(_1752_),
    .B1(_1630_),
    .B2(net1280),
    .A2(_1621_),
    .A1(net1166));
 sg13g2_nor2_1 _5100_ (.A(_1632_),
    .B(_1752_),
    .Y(_1753_));
 sg13g2_nor2_1 _5101_ (.A(net1317),
    .B(_1753_),
    .Y(_1754_));
 sg13g2_a22oi_1 _5102_ (.Y(_0294_),
    .B1(_1751_),
    .B2(_1754_),
    .A2(_0704_),
    .A1(net1318));
 sg13g2_nor2_1 _5103_ (.A(net1167),
    .B(_1644_),
    .Y(_1755_));
 sg13g2_a21oi_2 _5104_ (.B1(_1755_),
    .Y(_1756_),
    .A2(_1636_),
    .A1(net1167));
 sg13g2_nor2_1 _5105_ (.A(net1180),
    .B(_1730_),
    .Y(_1757_));
 sg13g2_mux2_1 _5106_ (.A0(\main.adder.s4_mant[44] ),
    .A1(\main.adder.s4_mant[43] ),
    .S(net1184),
    .X(_1758_));
 sg13g2_o21ai_1 _5107_ (.B1(net1199),
    .Y(_1759_),
    .A1(net1172),
    .A2(_1758_));
 sg13g2_o21ai_1 _5108_ (.B1(net1169),
    .Y(_1760_),
    .A1(_1757_),
    .A2(_1759_));
 sg13g2_a21oi_1 _5109_ (.A1(net1282),
    .A2(_1700_),
    .Y(_1761_),
    .B1(_1760_));
 sg13g2_a21oi_1 _5110_ (.A1(net1278),
    .A2(_1641_),
    .Y(_1762_),
    .B1(_1761_));
 sg13g2_nor2_1 _5111_ (.A(net1202),
    .B(_1762_),
    .Y(_1763_));
 sg13g2_a21oi_1 _5112_ (.A1(net1205),
    .A2(_1756_),
    .Y(_1764_),
    .B1(_1763_));
 sg13g2_nand2_1 _5113_ (.Y(_1765_),
    .A(net1164),
    .B(_1643_));
 sg13g2_o21ai_1 _5114_ (.B1(_1765_),
    .Y(_1766_),
    .A1(net1166),
    .A2(_1648_));
 sg13g2_a22oi_1 _5115_ (.Y(_1767_),
    .B1(_1499_),
    .B2(_1764_),
    .A2(net1602),
    .A1(net1317));
 sg13g2_o21ai_1 _5116_ (.B1(_1767_),
    .Y(_0295_),
    .A1(_1634_),
    .A2(_1766_));
 sg13g2_nor2_1 _5117_ (.A(net1167),
    .B(_1659_),
    .Y(_1768_));
 sg13g2_a21oi_1 _5118_ (.A1(net1168),
    .A2(_1651_),
    .Y(_1769_),
    .B1(_1768_));
 sg13g2_nor2_1 _5119_ (.A(net1180),
    .B(_1741_),
    .Y(_1770_));
 sg13g2_mux2_1 _5120_ (.A0(\main.adder.s4_mant[44] ),
    .A1(\main.adder.s4_mant[45] ),
    .S(net1188),
    .X(_1771_));
 sg13g2_o21ai_1 _5121_ (.B1(net1199),
    .Y(_1772_),
    .A1(net1172),
    .A2(_1771_));
 sg13g2_o21ai_1 _5122_ (.B1(net1169),
    .Y(_1773_),
    .A1(_1770_),
    .A2(_1772_));
 sg13g2_a21oi_1 _5123_ (.A1(net1282),
    .A2(_1716_),
    .Y(_1774_),
    .B1(_1773_));
 sg13g2_a21oi_1 _5124_ (.A1(net1278),
    .A2(_1656_),
    .Y(_1775_),
    .B1(_1774_));
 sg13g2_a21oi_1 _5125_ (.A1(net1205),
    .A2(_1769_),
    .Y(_1776_),
    .B1(net1132));
 sg13g2_o21ai_1 _5126_ (.B1(_1776_),
    .Y(_1777_),
    .A1(net1205),
    .A2(_1775_));
 sg13g2_mux2_1 _5127_ (.A0(_1658_),
    .A1(_1663_),
    .S(net1161),
    .X(_1778_));
 sg13g2_o21ai_1 _5128_ (.B1(_1777_),
    .Y(_1779_),
    .A1(_1634_),
    .A2(_1778_));
 sg13g2_a21o_1 _5129_ (.A2(net1569),
    .A1(net1313),
    .B1(_1779_),
    .X(_0296_));
 sg13g2_nor2_1 _5130_ (.A(net1167),
    .B(_1674_),
    .Y(_1780_));
 sg13g2_a21oi_2 _5131_ (.B1(_1780_),
    .Y(_1781_),
    .A2(_1666_),
    .A1(net1167));
 sg13g2_nand2_1 _5132_ (.Y(_1782_),
    .A(net1194),
    .B(_1731_));
 sg13g2_nor2_1 _5133_ (.A(\main.adder.s4_mant[46] ),
    .B(net1184),
    .Y(_1783_));
 sg13g2_o21ai_1 _5134_ (.B1(net1176),
    .Y(_1784_),
    .A1(\main.adder.s4_mant[45] ),
    .A2(net1188));
 sg13g2_a21oi_1 _5135_ (.A1(net1174),
    .A2(_1758_),
    .Y(_1785_),
    .B1(net1193));
 sg13g2_o21ai_1 _5136_ (.B1(_1785_),
    .Y(_1786_),
    .A1(_1783_),
    .A2(_1784_));
 sg13g2_nand3_1 _5137_ (.B(_1782_),
    .C(_1786_),
    .A(net1170),
    .Y(_1787_));
 sg13g2_a21oi_1 _5138_ (.A1(net1163),
    .A2(_1669_),
    .Y(_1788_),
    .B1(net1203));
 sg13g2_a22oi_1 _5139_ (.Y(_1789_),
    .B1(_1787_),
    .B2(_1788_),
    .A2(_1781_),
    .A1(net1206));
 sg13g2_nand2_1 _5140_ (.Y(_1790_),
    .A(net1166),
    .B(_1672_));
 sg13g2_o21ai_1 _5141_ (.B1(_1790_),
    .Y(_1791_),
    .A1(net1166),
    .A2(_1679_));
 sg13g2_o21ai_1 _5142_ (.B1(net1393),
    .Y(_1792_),
    .A1(_1632_),
    .A2(_1791_));
 sg13g2_a21oi_1 _5143_ (.A1(_1497_),
    .A2(_1789_),
    .Y(_1793_),
    .B1(_1792_));
 sg13g2_a21oi_1 _5144_ (.A1(net1313),
    .A2(_0708_),
    .Y(_0297_),
    .B1(_1793_));
 sg13g2_mux2_1 _5145_ (.A0(_1687_),
    .A1(_1694_),
    .S(net1161),
    .X(_1794_));
 sg13g2_nor2_1 _5146_ (.A(_1632_),
    .B(_1794_),
    .Y(_1795_));
 sg13g2_nor2_1 _5147_ (.A(net1168),
    .B(_1690_),
    .Y(_1796_));
 sg13g2_a21oi_2 _5148_ (.B1(_1796_),
    .Y(_1797_),
    .A2(_1682_),
    .A1(net1169));
 sg13g2_nand2_1 _5149_ (.Y(_1798_),
    .A(\main.adder.s4_mant[47] ),
    .B(net1188));
 sg13g2_a21oi_1 _5150_ (.A1(\main.adder.s4_exponent_adjust[0] ),
    .A2(\main.adder.s4_mant[46] ),
    .Y(_1799_),
    .B1(net1171));
 sg13g2_o21ai_1 _5151_ (.B1(net1197),
    .Y(_1800_),
    .A1(net1176),
    .A2(_1771_));
 sg13g2_a21oi_1 _5152_ (.A1(_1798_),
    .A2(_1799_),
    .Y(_1801_),
    .B1(_1800_));
 sg13g2_a21oi_1 _5153_ (.A1(net1282),
    .A2(_1743_),
    .Y(_1802_),
    .B1(_1801_));
 sg13g2_a21oi_1 _5154_ (.A1(net1278),
    .A2(_1685_),
    .Y(_1803_),
    .B1(net1203));
 sg13g2_o21ai_1 _5155_ (.B1(_1803_),
    .Y(_1804_),
    .A1(net1279),
    .A2(_1802_));
 sg13g2_a21oi_1 _5156_ (.A1(net1276),
    .A2(_1797_),
    .Y(_1805_),
    .B1(_1498_));
 sg13g2_a21oi_2 _5157_ (.B1(_1795_),
    .Y(_1806_),
    .A2(_1805_),
    .A1(_1804_));
 sg13g2_nor2_1 _5158_ (.A(net1387),
    .B(net1031),
    .Y(_1807_));
 sg13g2_a21oi_1 _5159_ (.A1(net1387),
    .A2(_1806_),
    .Y(_0298_),
    .B1(_1807_));
 sg13g2_mux2_1 _5160_ (.A0(\main.adder.s2_larger[23] ),
    .A1(net728),
    .S(net1331),
    .X(_0299_));
 sg13g2_mux2_1 _5161_ (.A0(\main.adder.s2_larger[24] ),
    .A1(net868),
    .S(net1331),
    .X(_0300_));
 sg13g2_mux2_1 _5162_ (.A0(net830),
    .A1(net752),
    .S(net1331),
    .X(_0301_));
 sg13g2_nand2_1 _5163_ (.Y(_1808_),
    .A(net1331),
    .B(net639));
 sg13g2_o21ai_1 _5164_ (.B1(_1808_),
    .Y(_0302_),
    .A1(net1331),
    .A2(_0747_));
 sg13g2_nand2_1 _5165_ (.Y(_1809_),
    .A(net1326),
    .B(net753));
 sg13g2_o21ai_1 _5166_ (.B1(_1809_),
    .Y(_0303_),
    .A1(net1331),
    .A2(_0748_));
 sg13g2_mux2_1 _5167_ (.A0(net873),
    .A1(\main.adder.s1_larger[5] ),
    .S(net1329),
    .X(_0304_));
 sg13g2_mux2_1 _5168_ (.A0(net816),
    .A1(net770),
    .S(net1329),
    .X(_0305_));
 sg13g2_mux2_1 _5169_ (.A0(\main.adder.s2_larger[30] ),
    .A1(net784),
    .S(net1329),
    .X(_0306_));
 sg13g2_mux2_1 _5170_ (.A0(net956),
    .A1(net914),
    .S(net1324),
    .X(_0307_));
 sg13g2_mux2_1 _5171_ (.A0(net870),
    .A1(net857),
    .S(net1325),
    .X(_0308_));
 sg13g2_mux2_1 _5172_ (.A0(net802),
    .A1(net794),
    .S(net1325),
    .X(_0309_));
 sg13g2_mux2_1 _5173_ (.A0(net931),
    .A1(net843),
    .S(net1324),
    .X(_0310_));
 sg13g2_mux2_1 _5174_ (.A0(net858),
    .A1(net798),
    .S(net1327),
    .X(_0311_));
 sg13g2_mux2_1 _5175_ (.A0(net918),
    .A1(net891),
    .S(net1324),
    .X(_0312_));
 sg13g2_mux2_1 _5176_ (.A0(\main.adder.s2_larger[37] ),
    .A1(net698),
    .S(net1329),
    .X(_0313_));
 sg13g2_mux2_1 _5177_ (.A0(\main.adder.s2_larger[38] ),
    .A1(net859),
    .S(net1330),
    .X(_0314_));
 sg13g2_mux2_1 _5178_ (.A0(\main.adder.s2_larger[39] ),
    .A1(net746),
    .S(net1330),
    .X(_0315_));
 sg13g2_mux2_1 _5179_ (.A0(net1422),
    .A1(\main.adder.s1_larger[17] ),
    .S(net1330),
    .X(_0316_));
 sg13g2_mux2_1 _5180_ (.A0(\main.adder.s2_larger[41] ),
    .A1(net901),
    .S(net1329),
    .X(_0317_));
 sg13g2_mux2_1 _5181_ (.A0(net806),
    .A1(net739),
    .S(net1329),
    .X(_0318_));
 sg13g2_mux2_1 _5182_ (.A0(net975),
    .A1(\main.adder.s1_larger[20] ),
    .S(net1332),
    .X(_0319_));
 sg13g2_mux2_1 _5183_ (.A0(\main.adder.s2_larger[44] ),
    .A1(net723),
    .S(net1333),
    .X(_0320_));
 sg13g2_mux2_1 _5184_ (.A0(net933),
    .A1(net847),
    .S(net1333),
    .X(_0321_));
 sg13g2_or2_1 _5185_ (.X(_1810_),
    .B(net844),
    .A(net876));
 sg13g2_nor4_2 _5186_ (.A(net1314),
    .B(net742),
    .C(net711),
    .Y(_1811_),
    .D(net1436));
 sg13g2_nor4_2 _5187_ (.A(net1493),
    .B(net1038),
    .C(net943),
    .Y(_1812_),
    .D(_1810_));
 sg13g2_a22oi_1 _5188_ (.Y(_0322_),
    .B1(_1811_),
    .B2(_1812_),
    .A2(_0755_),
    .A1(net1309));
 sg13g2_nor4_2 _5189_ (.A(\main.adder.s1_exp_diff[9] ),
    .B(\main.adder.s1_exp_diff[8] ),
    .C(\main.adder.s1_exp_diff[7] ),
    .Y(_1813_),
    .D(\main.adder.s1_exp_diff[6] ));
 sg13g2_or4_2 _5190_ (.A(\main.adder.s1_exp_diff[9] ),
    .B(\main.adder.s1_exp_diff[8] ),
    .C(\main.adder.s1_exp_diff[7] ),
    .D(\main.adder.s1_exp_diff[6] ),
    .X(_1814_));
 sg13g2_nor2_2 _5191_ (.A(net1247),
    .B(_1814_),
    .Y(_1815_));
 sg13g2_nand2b_2 _5192_ (.Y(_1816_),
    .B(_1813_),
    .A_N(net1247));
 sg13g2_nor2_1 _5193_ (.A(net1305),
    .B(_1816_),
    .Y(_1817_));
 sg13g2_nand2_2 _5194_ (.Y(_1818_),
    .A(net1348),
    .B(_1815_));
 sg13g2_and2_2 _5195_ (.A(net1249),
    .B(_1815_),
    .X(_1819_));
 sg13g2_nand2_2 _5196_ (.Y(_1820_),
    .A(net1249),
    .B(_1815_));
 sg13g2_nor2_2 _5197_ (.A(net1305),
    .B(_1820_),
    .Y(_1821_));
 sg13g2_nand2_2 _5198_ (.Y(_1822_),
    .A(net1249),
    .B(net1131));
 sg13g2_nor2_1 _5199_ (.A(net1250),
    .B(_1814_),
    .Y(_1823_));
 sg13g2_nand2b_1 _5200_ (.Y(_1824_),
    .B(_1813_),
    .A_N(net1250));
 sg13g2_nor2_1 _5201_ (.A(\main.adder.s1_exp_diff[2] ),
    .B(_1814_),
    .Y(_1825_));
 sg13g2_nand2b_1 _5202_ (.Y(_1826_),
    .B(_1813_),
    .A_N(\main.adder.s1_exp_diff[2] ));
 sg13g2_nor2_1 _5203_ (.A(\main.adder.s1_exp_diff[1] ),
    .B(_1814_),
    .Y(_1827_));
 sg13g2_nand2_1 _5204_ (.Y(_1828_),
    .A(_0746_),
    .B(_1813_));
 sg13g2_nor2_2 _5205_ (.A(\main.adder.s1_exp_diff[0] ),
    .B(_1814_),
    .Y(_1829_));
 sg13g2_nand2_1 _5206_ (.Y(_1830_),
    .A(_0097_),
    .B(net1142));
 sg13g2_nor4_2 _5207_ (.A(\main.adder.s1_smaler[28] ),
    .B(\main.adder.s1_smaler[27] ),
    .C(\main.adder.s1_smaler[30] ),
    .Y(_1831_),
    .D(\main.adder.s1_smaler[29] ));
 sg13g2_nor4_1 _5208_ (.A(\main.adder.s1_smaler[24] ),
    .B(\main.adder.s1_smaler[23] ),
    .C(\main.adder.s1_smaler[26] ),
    .D(\main.adder.s1_smaler[25] ),
    .Y(_1832_));
 sg13g2_nand2_2 _5209_ (.Y(_1833_),
    .A(_1831_),
    .B(_1832_));
 sg13g2_o21ai_1 _5210_ (.B1(_1830_),
    .Y(_1834_),
    .A1(net1142),
    .A2(_1833_));
 sg13g2_nor2_1 _5211_ (.A(net1148),
    .B(_1834_),
    .Y(_1835_));
 sg13g2_nor2b_1 _5212_ (.A(net1142),
    .B_N(_0098_),
    .Y(_1836_));
 sg13g2_a21oi_2 _5213_ (.B1(_1836_),
    .Y(_1837_),
    .A2(_1829_),
    .A1(_0095_));
 sg13g2_a21oi_2 _5214_ (.B1(_1835_),
    .Y(_1838_),
    .A2(_1837_),
    .A1(net1148));
 sg13g2_mux2_1 _5215_ (.A0(_0096_),
    .A1(_0093_),
    .S(net1138),
    .X(_1839_));
 sg13g2_mux2_1 _5216_ (.A0(_0094_),
    .A1(_0091_),
    .S(net1138),
    .X(_1840_));
 sg13g2_mux2_1 _5217_ (.A0(_1839_),
    .A1(_1840_),
    .S(net1146),
    .X(_1841_));
 sg13g2_mux2_1 _5218_ (.A0(_1838_),
    .A1(_1841_),
    .S(net1154),
    .X(_1842_));
 sg13g2_nor2b_1 _5219_ (.A(net1139),
    .B_N(_0092_),
    .Y(_1843_));
 sg13g2_a21oi_1 _5220_ (.A1(_0089_),
    .A2(net1138),
    .Y(_1844_),
    .B1(_1843_));
 sg13g2_mux2_1 _5221_ (.A0(_0090_),
    .A1(_0087_),
    .S(net1139),
    .X(_1845_));
 sg13g2_nor2_1 _5222_ (.A(net1143),
    .B(_1845_),
    .Y(_1846_));
 sg13g2_a21oi_1 _5223_ (.A1(net1143),
    .A2(_1844_),
    .Y(_1847_),
    .B1(_1846_));
 sg13g2_nor2b_1 _5224_ (.A(net1140),
    .B_N(_0088_),
    .Y(_1848_));
 sg13g2_a221oi_1 _5225_ (.B2(_0085_),
    .C1(_1848_),
    .B1(net1140),
    .A1(_0746_),
    .Y(_1849_),
    .A2(_1813_));
 sg13g2_nor2b_1 _5226_ (.A(net1139),
    .B_N(_0086_),
    .Y(_1850_));
 sg13g2_a21oi_1 _5227_ (.A1(_0083_),
    .A2(net1140),
    .Y(_1851_),
    .B1(_1850_));
 sg13g2_a21oi_1 _5228_ (.A1(net1146),
    .A2(_1851_),
    .Y(_1852_),
    .B1(_1849_));
 sg13g2_mux2_1 _5229_ (.A0(_1847_),
    .A1(_1852_),
    .S(net1153),
    .X(_1853_));
 sg13g2_mux2_1 _5230_ (.A0(_1842_),
    .A1(_1853_),
    .S(net1160),
    .X(_1854_));
 sg13g2_mux2_1 _5231_ (.A0(_0080_),
    .A1(_0077_),
    .S(net1141),
    .X(_1855_));
 sg13g2_mux2_1 _5232_ (.A0(\main.adder.s1_rs.levels[0][24] ),
    .A1(\main.adder.s1_rs.levels[0][23] ),
    .S(net1142),
    .X(_1856_));
 sg13g2_nand2_1 _5233_ (.Y(_1857_),
    .A(net1148),
    .B(_1856_));
 sg13g2_o21ai_1 _5234_ (.B1(_1857_),
    .Y(_1858_),
    .A1(net1148),
    .A2(_1855_));
 sg13g2_nor2_1 _5235_ (.A(net1150),
    .B(_1858_),
    .Y(_1859_));
 sg13g2_mux2_1 _5236_ (.A0(_0084_),
    .A1(_0081_),
    .S(net1141),
    .X(_1860_));
 sg13g2_mux2_1 _5237_ (.A0(_0082_),
    .A1(_0079_),
    .S(net1142),
    .X(_1861_));
 sg13g2_mux2_1 _5238_ (.A0(_1860_),
    .A1(_1861_),
    .S(net1147),
    .X(_1862_));
 sg13g2_a21oi_2 _5239_ (.B1(_1859_),
    .Y(_1863_),
    .A2(_1862_),
    .A1(net1150));
 sg13g2_nor2_1 _5240_ (.A(net1249),
    .B(_1814_),
    .Y(_1864_));
 sg13g2_nand2b_2 _5241_ (.Y(_1865_),
    .B(_1813_),
    .A_N(net1249));
 sg13g2_nand2_2 _5242_ (.Y(_1866_),
    .A(net1250),
    .B(net1134));
 sg13g2_nor2_1 _5243_ (.A(_1818_),
    .B(_1866_),
    .Y(_1867_));
 sg13g2_a22oi_1 _5244_ (.Y(_1868_),
    .B1(_1863_),
    .B2(_1867_),
    .A2(net927),
    .A1(net1305));
 sg13g2_o21ai_1 _5245_ (.B1(_1868_),
    .Y(_0323_),
    .A1(_1822_),
    .A2(_1854_));
 sg13g2_mux2_1 _5246_ (.A0(_0095_),
    .A1(_0096_),
    .S(net1139),
    .X(_1869_));
 sg13g2_mux2_1 _5247_ (.A0(_0093_),
    .A1(_0094_),
    .S(net1138),
    .X(_1870_));
 sg13g2_mux2_1 _5248_ (.A0(_1869_),
    .A1(_1870_),
    .S(net1146),
    .X(_1871_));
 sg13g2_nand2_2 _5249_ (.Y(_1872_),
    .A(net1142),
    .B(_1833_));
 sg13g2_mux2_1 _5250_ (.A0(_0097_),
    .A1(_0098_),
    .S(_1829_),
    .X(_1873_));
 sg13g2_mux2_1 _5251_ (.A0(_1872_),
    .A1(_1873_),
    .S(net1148),
    .X(_1874_));
 sg13g2_mux2_1 _5252_ (.A0(_1871_),
    .A1(_1874_),
    .S(net1151),
    .X(_1875_));
 sg13g2_mux4_1 _5253_ (.S0(net1138),
    .A0(_0085_),
    .A1(_0086_),
    .A2(_0087_),
    .A3(_0088_),
    .S1(net1144),
    .X(_1876_));
 sg13g2_nor2b_1 _5254_ (.A(net1138),
    .B_N(_0091_),
    .Y(_1877_));
 sg13g2_a21oi_2 _5255_ (.B1(_1877_),
    .Y(_1878_),
    .A2(net1139),
    .A1(_0092_));
 sg13g2_mux2_1 _5256_ (.A0(_0089_),
    .A1(_0090_),
    .S(net1138),
    .X(_1879_));
 sg13g2_nor2_1 _5257_ (.A(net1143),
    .B(_1879_),
    .Y(_1880_));
 sg13g2_a21oi_1 _5258_ (.A1(net1143),
    .A2(_1878_),
    .Y(_1881_),
    .B1(_1880_));
 sg13g2_mux2_1 _5259_ (.A0(_1876_),
    .A1(_1881_),
    .S(net1150),
    .X(_1882_));
 sg13g2_mux2_1 _5260_ (.A0(_1875_),
    .A1(_1882_),
    .S(net1160),
    .X(_1883_));
 sg13g2_nor2_1 _5261_ (.A(net1297),
    .B(net1249),
    .Y(_1884_));
 sg13g2_nand2b_1 _5262_ (.Y(_1885_),
    .B(net1348),
    .A_N(net1249));
 sg13g2_nor2_2 _5263_ (.A(_1816_),
    .B(_1885_),
    .Y(_1886_));
 sg13g2_nand2_1 _5264_ (.Y(_1887_),
    .A(_1815_),
    .B(_1884_));
 sg13g2_nor2b_1 _5265_ (.A(net1141),
    .B_N(_0083_),
    .Y(_1888_));
 sg13g2_a221oi_1 _5266_ (.B2(_0084_),
    .C1(_1888_),
    .B1(net1141),
    .A1(_0746_),
    .Y(_1889_),
    .A2(_1813_));
 sg13g2_nor2b_1 _5267_ (.A(net1141),
    .B_N(_0081_),
    .Y(_1890_));
 sg13g2_a21oi_1 _5268_ (.A1(_0082_),
    .A2(net1141),
    .Y(_1891_),
    .B1(_1890_));
 sg13g2_a21oi_1 _5269_ (.A1(net1147),
    .A2(_1891_),
    .Y(_1892_),
    .B1(_1889_));
 sg13g2_mux2_1 _5270_ (.A0(_0079_),
    .A1(_0080_),
    .S(net1141),
    .X(_1893_));
 sg13g2_mux2_1 _5271_ (.A0(_0077_),
    .A1(_0078_),
    .S(net1142),
    .X(_1894_));
 sg13g2_mux2_1 _5272_ (.A0(_1893_),
    .A1(_1894_),
    .S(net1149),
    .X(_1895_));
 sg13g2_mux2_1 _5273_ (.A0(_1892_),
    .A1(_1895_),
    .S(net1154),
    .X(_1896_));
 sg13g2_o21ai_1 _5274_ (.B1(\main.adder.s1_rs.levels[0][23] ),
    .Y(_1897_),
    .A1(\main.adder.s1_exp_diff[0] ),
    .A2(_1814_));
 sg13g2_nor3_2 _5275_ (.A(_1825_),
    .B(net1148),
    .C(_1897_),
    .Y(_1898_));
 sg13g2_nor2_1 _5276_ (.A(net1157),
    .B(_1898_),
    .Y(_1899_));
 sg13g2_a21oi_2 _5277_ (.B1(_1899_),
    .Y(_1900_),
    .A2(_1896_),
    .A1(net1156));
 sg13g2_a22oi_1 _5278_ (.Y(_1901_),
    .B1(_1886_),
    .B2(_1900_),
    .A2(net906),
    .A1(net1306));
 sg13g2_o21ai_1 _5279_ (.B1(_1901_),
    .Y(_0324_),
    .A1(_1822_),
    .A2(_1883_));
 sg13g2_nor2_1 _5280_ (.A(net1145),
    .B(_1834_),
    .Y(_1902_));
 sg13g2_nor2_1 _5281_ (.A(net1155),
    .B(_1902_),
    .Y(_1903_));
 sg13g2_nor2_1 _5282_ (.A(net1143),
    .B(_1839_),
    .Y(_1904_));
 sg13g2_a21oi_2 _5283_ (.B1(_1904_),
    .Y(_1905_),
    .A2(_1837_),
    .A1(net1144));
 sg13g2_a21oi_2 _5284_ (.B1(_1903_),
    .Y(_1906_),
    .A2(_1905_),
    .A1(net1155));
 sg13g2_mux4_1 _5285_ (.S0(net1146),
    .A0(_0090_),
    .A1(_0088_),
    .A2(_0087_),
    .A3(_0085_),
    .S1(net1140),
    .X(_1907_));
 sg13g2_nor2_1 _5286_ (.A(net1146),
    .B(_1840_),
    .Y(_1908_));
 sg13g2_a21oi_1 _5287_ (.A1(net1146),
    .A2(_1844_),
    .Y(_1909_),
    .B1(_1908_));
 sg13g2_mux2_1 _5288_ (.A0(_1907_),
    .A1(_1909_),
    .S(net1150),
    .X(_1910_));
 sg13g2_nor2_1 _5289_ (.A(net1156),
    .B(_1910_),
    .Y(_1911_));
 sg13g2_a21oi_2 _5290_ (.B1(_1911_),
    .Y(_1912_),
    .A2(_1906_),
    .A1(net1156));
 sg13g2_nor2_1 _5291_ (.A(net1143),
    .B(_1860_),
    .Y(_1913_));
 sg13g2_a21oi_1 _5292_ (.A1(net1144),
    .A2(_1851_),
    .Y(_1914_),
    .B1(_1913_));
 sg13g2_mux2_1 _5293_ (.A0(_1855_),
    .A1(_1861_),
    .S(net1144),
    .X(_1915_));
 sg13g2_mux2_1 _5294_ (.A0(_1914_),
    .A1(_1915_),
    .S(net1153),
    .X(_1916_));
 sg13g2_nand3_1 _5295_ (.B(net1145),
    .C(_1856_),
    .A(net1150),
    .Y(_1917_));
 sg13g2_and2_1 _5296_ (.A(net1158),
    .B(_1917_),
    .X(_1918_));
 sg13g2_a21oi_2 _5297_ (.B1(_1918_),
    .Y(_1919_),
    .A2(_1916_),
    .A1(net1156));
 sg13g2_a22oi_1 _5298_ (.Y(_1920_),
    .B1(_1886_),
    .B2(_1919_),
    .A2(net1020),
    .A1(net1306));
 sg13g2_o21ai_1 _5299_ (.B1(_1920_),
    .Y(_0325_),
    .A1(_1822_),
    .A2(_1912_));
 sg13g2_nor2_1 _5300_ (.A(net1146),
    .B(_1870_),
    .Y(_1921_));
 sg13g2_a21oi_2 _5301_ (.B1(_1921_),
    .Y(_1922_),
    .A2(_1878_),
    .A1(net1146));
 sg13g2_mux4_1 _5302_ (.S0(net1138),
    .A0(_0087_),
    .A1(_0088_),
    .A2(_0089_),
    .A3(_0090_),
    .S1(net1143),
    .X(_1923_));
 sg13g2_mux2_1 _5303_ (.A0(_1922_),
    .A1(_1923_),
    .S(net1153),
    .X(_1924_));
 sg13g2_nand2_1 _5304_ (.Y(_1925_),
    .A(net1159),
    .B(_1924_));
 sg13g2_mux2_1 _5305_ (.A0(_1869_),
    .A1(_1873_),
    .S(net1145),
    .X(_1926_));
 sg13g2_nor2_1 _5306_ (.A(\main.adder.s1_exp_diff[1] ),
    .B(_1872_),
    .Y(_1927_));
 sg13g2_nand2_1 _5307_ (.Y(_1928_),
    .A(net1152),
    .B(_1927_));
 sg13g2_o21ai_1 _5308_ (.B1(_1928_),
    .Y(_1929_),
    .A1(net1152),
    .A2(_1926_));
 sg13g2_o21ai_1 _5309_ (.B1(_1925_),
    .Y(_1930_),
    .A1(net1159),
    .A2(_1929_));
 sg13g2_mux4_1 _5310_ (.S0(net1139),
    .A0(_0083_),
    .A1(_0084_),
    .A2(_0085_),
    .A3(_0086_),
    .S1(net1143),
    .X(_1931_));
 sg13g2_nand2_1 _5311_ (.Y(_1932_),
    .A(net1147),
    .B(_1893_));
 sg13g2_o21ai_1 _5312_ (.B1(_1932_),
    .Y(_1933_),
    .A1(net1147),
    .A2(_1891_));
 sg13g2_mux2_1 _5313_ (.A0(_1931_),
    .A1(_1933_),
    .S(net1154),
    .X(_1934_));
 sg13g2_mux2_1 _5314_ (.A0(_1894_),
    .A1(_1897_),
    .S(net1148),
    .X(_1935_));
 sg13g2_nand3b_1 _5315_ (.B(net1158),
    .C(net1151),
    .Y(_1936_),
    .A_N(_1935_));
 sg13g2_o21ai_1 _5316_ (.B1(_1936_),
    .Y(_1937_),
    .A1(net1158),
    .A2(_1934_));
 sg13g2_a22oi_1 _5317_ (.Y(_1938_),
    .B1(_1886_),
    .B2(_1937_),
    .A2(net982),
    .A1(net1306));
 sg13g2_o21ai_1 _5318_ (.B1(_1938_),
    .Y(_0326_),
    .A1(_1822_),
    .A2(_1930_));
 sg13g2_nand3b_1 _5319_ (.B(net1155),
    .C(net1250),
    .Y(_1939_),
    .A_N(_1838_));
 sg13g2_mux2_1 _5320_ (.A0(_1841_),
    .A1(_1847_),
    .S(net1153),
    .X(_1940_));
 sg13g2_o21ai_1 _5321_ (.B1(_1939_),
    .Y(_1941_),
    .A1(net1156),
    .A2(_1940_));
 sg13g2_mux2_1 _5322_ (.A0(_1852_),
    .A1(_1862_),
    .S(net1153),
    .X(_1942_));
 sg13g2_and2_1 _5323_ (.A(net1156),
    .B(_1942_),
    .X(_1943_));
 sg13g2_nand2_1 _5324_ (.Y(_1944_),
    .A(net1151),
    .B(_1858_));
 sg13g2_a21oi_2 _5325_ (.B1(_1943_),
    .Y(_1945_),
    .A2(_1944_),
    .A1(net1159));
 sg13g2_a22oi_1 _5326_ (.Y(_1946_),
    .B1(_1945_),
    .B2(_1886_),
    .A2(_1941_),
    .A1(_1821_));
 sg13g2_o21ai_1 _5327_ (.B1(_1946_),
    .Y(_0327_),
    .A1(net1350),
    .A2(_0757_));
 sg13g2_nor2_1 _5328_ (.A(net1151),
    .B(_1874_),
    .Y(_1947_));
 sg13g2_and2_1 _5329_ (.A(net1153),
    .B(_1881_),
    .X(_1948_));
 sg13g2_a21oi_2 _5330_ (.B1(_1948_),
    .Y(_1949_),
    .A2(_1871_),
    .A1(net1150));
 sg13g2_a22oi_1 _5331_ (.Y(_1950_),
    .B1(_1949_),
    .B2(net1158),
    .A2(_1947_),
    .A1(net1251));
 sg13g2_nor2_1 _5332_ (.A(net1154),
    .B(_1895_),
    .Y(_1951_));
 sg13g2_nor3_1 _5333_ (.A(net1152),
    .B(net1148),
    .C(_1897_),
    .Y(_1952_));
 sg13g2_nor2_1 _5334_ (.A(_1951_),
    .B(_1952_),
    .Y(_1953_));
 sg13g2_mux2_1 _5335_ (.A0(_1876_),
    .A1(_1892_),
    .S(net1154),
    .X(_1954_));
 sg13g2_mux2_1 _5336_ (.A0(_1953_),
    .A1(_1954_),
    .S(net1157),
    .X(_1955_));
 sg13g2_nor2_1 _5337_ (.A(net1130),
    .B(_1955_),
    .Y(_1956_));
 sg13g2_a21oi_1 _5338_ (.A1(net1305),
    .A2(net1566),
    .Y(_1957_),
    .B1(_1956_));
 sg13g2_o21ai_1 _5339_ (.B1(_1957_),
    .Y(_0328_),
    .A1(_1822_),
    .A2(_1950_));
 sg13g2_nand3_1 _5340_ (.B(net1155),
    .C(_1902_),
    .A(net1250),
    .Y(_1958_));
 sg13g2_mux2_1 _5341_ (.A0(_1905_),
    .A1(_1909_),
    .S(net1153),
    .X(_1959_));
 sg13g2_o21ai_1 _5342_ (.B1(_1958_),
    .Y(_1960_),
    .A1(net1156),
    .A2(_1959_));
 sg13g2_a21oi_1 _5343_ (.A1(net1145),
    .A2(_1856_),
    .Y(_1961_),
    .B1(net1150));
 sg13g2_a21oi_1 _5344_ (.A1(net1150),
    .A2(_1915_),
    .Y(_1962_),
    .B1(_1961_));
 sg13g2_mux2_1 _5345_ (.A0(_1907_),
    .A1(_1914_),
    .S(net1153),
    .X(_1963_));
 sg13g2_nand2_1 _5346_ (.Y(_1964_),
    .A(net1156),
    .B(_1963_));
 sg13g2_o21ai_1 _5347_ (.B1(_1964_),
    .Y(_1965_),
    .A1(net1157),
    .A2(_1962_));
 sg13g2_nor2_1 _5348_ (.A(net1130),
    .B(_1965_),
    .Y(_1966_));
 sg13g2_a21oi_1 _5349_ (.A1(_1821_),
    .A2(_1960_),
    .Y(_1967_),
    .B1(_1966_));
 sg13g2_o21ai_1 _5350_ (.B1(_1967_),
    .Y(_0329_),
    .A1(net1350),
    .A2(_0758_));
 sg13g2_nand3_1 _5351_ (.B(net1155),
    .C(_1927_),
    .A(net1250),
    .Y(_1968_));
 sg13g2_mux2_1 _5352_ (.A0(_1922_),
    .A1(_1926_),
    .S(net1152),
    .X(_1969_));
 sg13g2_o21ai_1 _5353_ (.B1(_1968_),
    .Y(_1970_),
    .A1(net1157),
    .A2(_1969_));
 sg13g2_mux2_1 _5354_ (.A0(_1933_),
    .A1(_1935_),
    .S(net1155),
    .X(_1971_));
 sg13g2_mux2_1 _5355_ (.A0(_1923_),
    .A1(_1931_),
    .S(net1154),
    .X(_1972_));
 sg13g2_mux2_1 _5356_ (.A0(_1971_),
    .A1(_1972_),
    .S(net1157),
    .X(_1973_));
 sg13g2_nor2_1 _5357_ (.A(net1130),
    .B(_1973_),
    .Y(_1974_));
 sg13g2_a21oi_2 _5358_ (.B1(_1974_),
    .Y(_1975_),
    .A2(_1970_),
    .A1(_1821_));
 sg13g2_o21ai_1 _5359_ (.B1(_1975_),
    .Y(_0330_),
    .A1(net1364),
    .A2(_0759_));
 sg13g2_nand2b_2 _5360_ (.Y(_1976_),
    .B(net1160),
    .A_N(_1842_));
 sg13g2_nand2_1 _5361_ (.Y(_1977_),
    .A(net1160),
    .B(_1863_));
 sg13g2_o21ai_1 _5362_ (.B1(_1977_),
    .Y(_1978_),
    .A1(net1160),
    .A2(_1853_));
 sg13g2_a22oi_1 _5363_ (.Y(_1979_),
    .B1(_1886_),
    .B2(_1978_),
    .A2(net1559),
    .A1(net1305));
 sg13g2_o21ai_1 _5364_ (.B1(_1979_),
    .Y(_0331_),
    .A1(_1822_),
    .A2(_1976_));
 sg13g2_or2_2 _5365_ (.X(_1980_),
    .B(_1875_),
    .A(net1157));
 sg13g2_nor2_1 _5366_ (.A(_1822_),
    .B(_1980_),
    .Y(_1981_));
 sg13g2_a21oi_1 _5367_ (.A1(net1297),
    .A2(net1552),
    .Y(_1982_),
    .B1(_1981_));
 sg13g2_mux2_1 _5368_ (.A0(_1882_),
    .A1(_1896_),
    .S(net1158),
    .X(_1983_));
 sg13g2_o21ai_1 _5369_ (.B1(_1982_),
    .Y(_0332_),
    .A1(net1129),
    .A2(_1983_));
 sg13g2_nand2_2 _5370_ (.Y(_1984_),
    .A(net1159),
    .B(_1906_));
 sg13g2_mux2_1 _5371_ (.A0(_1910_),
    .A1(_1916_),
    .S(net1159),
    .X(_1985_));
 sg13g2_nor2_1 _5372_ (.A(net1129),
    .B(_1985_),
    .Y(_1986_));
 sg13g2_a21oi_1 _5373_ (.A1(net1297),
    .A2(net1576),
    .Y(_1987_),
    .B1(_1986_));
 sg13g2_o21ai_1 _5374_ (.B1(_1987_),
    .Y(_0333_),
    .A1(_1822_),
    .A2(_1984_));
 sg13g2_and2_2 _5375_ (.A(net1159),
    .B(_1929_),
    .X(_1988_));
 sg13g2_a22oi_1 _5376_ (.Y(_1989_),
    .B1(_1821_),
    .B2(_1988_),
    .A2(net1539),
    .A1(net1297));
 sg13g2_mux2_1 _5377_ (.A0(_1924_),
    .A1(_1934_),
    .S(net1158),
    .X(_1990_));
 sg13g2_o21ai_1 _5378_ (.B1(_1989_),
    .Y(_0334_),
    .A1(net1129),
    .A2(_1990_));
 sg13g2_mux2_1 _5379_ (.A0(_1940_),
    .A1(_1942_),
    .S(net1159),
    .X(_1991_));
 sg13g2_nor3_2 _5380_ (.A(net1250),
    .B(net1151),
    .C(_1838_),
    .Y(_1992_));
 sg13g2_a22oi_1 _5381_ (.Y(_1993_),
    .B1(_1821_),
    .B2(_1992_),
    .A2(net1586),
    .A1(net1297));
 sg13g2_o21ai_1 _5382_ (.B1(_1993_),
    .Y(_0335_),
    .A1(net1129),
    .A2(_1991_));
 sg13g2_nand2_1 _5383_ (.Y(_1994_),
    .A(net1158),
    .B(_1954_));
 sg13g2_o21ai_1 _5384_ (.B1(_1994_),
    .Y(_1995_),
    .A1(net1158),
    .A2(_1949_));
 sg13g2_nor3_2 _5385_ (.A(net1251),
    .B(net1151),
    .C(_1874_),
    .Y(_1996_));
 sg13g2_a22oi_1 _5386_ (.Y(_1997_),
    .B1(_1821_),
    .B2(_1996_),
    .A2(net1570),
    .A1(net1298));
 sg13g2_o21ai_1 _5387_ (.B1(_1997_),
    .Y(_0336_),
    .A1(net1129),
    .A2(_1995_));
 sg13g2_mux2_1 _5388_ (.A0(_1959_),
    .A1(_1963_),
    .S(net1159),
    .X(_1998_));
 sg13g2_nor4_2 _5389_ (.A(net1250),
    .B(net1151),
    .C(net1145),
    .Y(_1999_),
    .D(_1834_));
 sg13g2_a22oi_1 _5390_ (.Y(_2000_),
    .B1(_1821_),
    .B2(_1999_),
    .A2(net1585),
    .A1(net1297));
 sg13g2_o21ai_1 _5391_ (.B1(_2000_),
    .Y(_0337_),
    .A1(net1129),
    .A2(_1998_));
 sg13g2_mux2_1 _5392_ (.A0(_1969_),
    .A1(_1972_),
    .S(net1160),
    .X(_2001_));
 sg13g2_nor4_2 _5393_ (.A(net1441),
    .B(net1251),
    .C(net1151),
    .Y(_2002_),
    .D(_1872_));
 sg13g2_a22oi_1 _5394_ (.Y(_2003_),
    .B1(_1821_),
    .B2(_2002_),
    .A2(net1553),
    .A1(net1305));
 sg13g2_o21ai_1 _5395_ (.B1(_2003_),
    .Y(_0338_),
    .A1(net1130),
    .A2(_2001_));
 sg13g2_nor2_1 _5396_ (.A(_1865_),
    .B(_1883_),
    .Y(_2004_));
 sg13g2_nor3_1 _5397_ (.A(_1818_),
    .B(_1865_),
    .C(_1883_),
    .Y(_2005_));
 sg13g2_a21o_1 _5398_ (.A2(net1526),
    .A1(net1307),
    .B1(_2005_),
    .X(_0339_));
 sg13g2_nor2_1 _5399_ (.A(_1865_),
    .B(_1912_),
    .Y(_2006_));
 sg13g2_nor3_1 _5400_ (.A(_1818_),
    .B(_1865_),
    .C(_1912_),
    .Y(_2007_));
 sg13g2_a21o_1 _5401_ (.A2(net1456),
    .A1(net1307),
    .B1(_2007_),
    .X(_0340_));
 sg13g2_nor2_1 _5402_ (.A(_1865_),
    .B(_1930_),
    .Y(_2008_));
 sg13g2_nor3_1 _5403_ (.A(_1818_),
    .B(_1865_),
    .C(_1930_),
    .Y(_2009_));
 sg13g2_a21o_1 _5404_ (.A2(net1516),
    .A1(net1308),
    .B1(_2009_),
    .X(_0341_));
 sg13g2_nand3_1 _5405_ (.B(net1136),
    .C(_1941_),
    .A(_1817_),
    .Y(_2010_));
 sg13g2_o21ai_1 _5406_ (.B1(_2010_),
    .Y(_0342_),
    .A1(net1349),
    .A2(_0749_));
 sg13g2_nor3_1 _5407_ (.A(_1818_),
    .B(_1865_),
    .C(_1950_),
    .Y(_2011_));
 sg13g2_a21o_1 _5408_ (.A2(net1484),
    .A1(net1307),
    .B1(_2011_),
    .X(_0343_));
 sg13g2_nand3_1 _5409_ (.B(net1136),
    .C(_1960_),
    .A(_1817_),
    .Y(_2012_));
 sg13g2_o21ai_1 _5410_ (.B1(_2012_),
    .Y(_0344_),
    .A1(net1347),
    .A2(_0750_));
 sg13g2_nand3_1 _5411_ (.B(net1136),
    .C(_1970_),
    .A(net1131),
    .Y(_2013_));
 sg13g2_o21ai_1 _5412_ (.B1(_2013_),
    .Y(_0345_),
    .A1(net1347),
    .A2(_0751_));
 sg13g2_nand2_1 _5413_ (.Y(_2014_),
    .A(net1307),
    .B(net1426));
 sg13g2_nor2_1 _5414_ (.A(net1249),
    .B(_1976_),
    .Y(_2015_));
 sg13g2_o21ai_1 _5415_ (.B1(_2014_),
    .Y(_0346_),
    .A1(net1130),
    .A2(_1976_));
 sg13g2_nand2_1 _5416_ (.Y(_2016_),
    .A(net1297),
    .B(net875));
 sg13g2_o21ai_1 _5417_ (.B1(_2016_),
    .Y(_0347_),
    .A1(net1129),
    .A2(_1980_));
 sg13g2_nand2_1 _5418_ (.Y(_2017_),
    .A(net1297),
    .B(net725));
 sg13g2_o21ai_1 _5419_ (.B1(_2017_),
    .Y(_0348_),
    .A1(net1129),
    .A2(_1984_));
 sg13g2_nor2b_1 _5420_ (.A(net1347),
    .B_N(net1601),
    .Y(_2018_));
 sg13g2_a21o_1 _5421_ (.A2(_1988_),
    .A1(_1886_),
    .B1(_2018_),
    .X(_0349_));
 sg13g2_nand3_1 _5422_ (.B(net1134),
    .C(_1992_),
    .A(net1131),
    .Y(_2019_));
 sg13g2_o21ai_1 _5423_ (.B1(_2019_),
    .Y(_0350_),
    .A1(net1332),
    .A2(_0752_));
 sg13g2_nand3_1 _5424_ (.B(net1134),
    .C(_1996_),
    .A(net1131),
    .Y(_2020_));
 sg13g2_o21ai_1 _5425_ (.B1(_2020_),
    .Y(_0351_),
    .A1(net1352),
    .A2(_0753_));
 sg13g2_nand3_1 _5426_ (.B(net1135),
    .C(_1999_),
    .A(net1131),
    .Y(_2021_));
 sg13g2_o21ai_1 _5427_ (.B1(_2021_),
    .Y(_0352_),
    .A1(net1352),
    .A2(_0754_));
 sg13g2_nand3_1 _5428_ (.B(net1137),
    .C(_2002_),
    .A(net1131),
    .Y(_2022_));
 sg13g2_o21ai_1 _5429_ (.B1(_2022_),
    .Y(_0353_),
    .A1(net1352),
    .A2(_0756_));
 sg13g2_nor2_1 _5430_ (.A(net1452),
    .B(net1074),
    .Y(_2023_));
 sg13g2_a21oi_1 _5431_ (.A1(_0912_),
    .A2(net1074),
    .Y(_0354_),
    .B1(_2023_));
 sg13g2_nor2_1 _5432_ (.A(net1480),
    .B(net1077),
    .Y(_2024_));
 sg13g2_a21oi_1 _5433_ (.A1(_0957_),
    .A2(net1077),
    .Y(_0355_),
    .B1(_2024_));
 sg13g2_nor2_1 _5434_ (.A(net1400),
    .B(net1103),
    .Y(_2025_));
 sg13g2_a21oi_1 _5435_ (.A1(net1103),
    .A2(_0970_),
    .Y(_0356_),
    .B1(_2025_));
 sg13g2_nor2_1 _5436_ (.A(net1460),
    .B(net1073),
    .Y(_2026_));
 sg13g2_a21oi_1 _5437_ (.A1(_0908_),
    .A2(net1073),
    .Y(_0357_),
    .B1(_2026_));
 sg13g2_nor2_1 _5438_ (.A(net1045),
    .B(net1102),
    .Y(_2027_));
 sg13g2_a21oi_1 _5439_ (.A1(net1102),
    .A2(_0890_),
    .Y(_0358_),
    .B1(_2027_));
 sg13g2_nor2_1 _5440_ (.A(net1412),
    .B(net1073),
    .Y(_2028_));
 sg13g2_a21oi_1 _5441_ (.A1(_0917_),
    .A2(net1073),
    .Y(_0359_),
    .B1(_2028_));
 sg13g2_nor2_1 _5442_ (.A(net1502),
    .B(net1102),
    .Y(_2029_));
 sg13g2_a21oi_1 _5443_ (.A1(net1102),
    .A2(_0935_),
    .Y(_0360_),
    .B1(_2029_));
 sg13g2_nand3_1 _5444_ (.B(\main.state[1] ),
    .C(_0778_),
    .A(net1273),
    .Y(_2030_));
 sg13g2_o21ai_1 _5445_ (.B1(_0764_),
    .Y(_2031_),
    .A1(\main.state[2] ),
    .A2(net1274));
 sg13g2_nor2b_2 _5446_ (.A(_2031_),
    .B_N(_2030_),
    .Y(_2032_));
 sg13g2_o21ai_1 _5447_ (.B1(net1339),
    .Y(_2033_),
    .A1(net1546),
    .A2(_2032_));
 sg13g2_a21oi_1 _5448_ (.A1(_0666_),
    .A2(_2032_),
    .Y(_0361_),
    .B1(_2033_));
 sg13g2_o21ai_1 _5449_ (.B1(net1339),
    .Y(_2034_),
    .A1(net1594),
    .A2(_2032_));
 sg13g2_a21oi_1 _5450_ (.A1(_0664_),
    .A2(_2032_),
    .Y(_0362_),
    .B1(_2034_));
 sg13g2_nor2_1 _5451_ (.A(net1469),
    .B(net1102),
    .Y(_2035_));
 sg13g2_a21oi_1 _5452_ (.A1(net1102),
    .A2(_0900_),
    .Y(_0363_),
    .B1(_2035_));
 sg13g2_nor2_1 _5453_ (.A(net1030),
    .B(net1104),
    .Y(_2036_));
 sg13g2_a21oi_1 _5454_ (.A1(net1104),
    .A2(_0851_),
    .Y(_0364_),
    .B1(_2036_));
 sg13g2_and2_1 _5455_ (.A(net1340),
    .B(net581),
    .X(_0365_));
 sg13g2_nor2b_2 _5456_ (.A(net1483),
    .B_N(_1381_),
    .Y(_2037_));
 sg13g2_or4_1 _5457_ (.A(net833),
    .B(_1383_),
    .C(_1442_),
    .D(_2037_),
    .X(_2038_));
 sg13g2_a22oi_1 _5458_ (.Y(_0366_),
    .B1(_1443_),
    .B2(_2038_),
    .A2(_0728_),
    .A1(net1311));
 sg13g2_nand3b_1 _5459_ (.B(\main.adder.s5_mant[22] ),
    .C(_1382_),
    .Y(_2039_),
    .A_N(_2037_));
 sg13g2_xor2_1 _5460_ (.B(_2039_),
    .A(\main.adder.s5_mant[23] ),
    .X(_2040_));
 sg13g2_o21ai_1 _5461_ (.B1(_1445_),
    .Y(_2041_),
    .A1(_1383_),
    .A2(_2037_));
 sg13g2_nor2b_1 _5462_ (.A(_2041_),
    .B_N(_1447_),
    .Y(_2042_));
 sg13g2_and4_1 _5463_ (.A(_1450_),
    .B(_1452_),
    .C(_1454_),
    .D(_2042_),
    .X(_2043_));
 sg13g2_and4_1 _5464_ (.A(_1457_),
    .B(_1461_),
    .C(_2040_),
    .D(_2043_),
    .X(_2044_));
 sg13g2_and4_1 _5465_ (.A(_1459_),
    .B(_1464_),
    .C(_1466_),
    .D(_2044_),
    .X(_2045_));
 sg13g2_and4_1 _5466_ (.A(_1468_),
    .B(_1471_),
    .C(_1473_),
    .D(_2045_),
    .X(_2046_));
 sg13g2_and4_1 _5467_ (.A(_1475_),
    .B(_1478_),
    .C(_1480_),
    .D(_2046_),
    .X(_2047_));
 sg13g2_and4_1 _5468_ (.A(_1482_),
    .B(_1485_),
    .C(_1487_),
    .D(_2047_),
    .X(_2048_));
 sg13g2_nand4_1 _5469_ (.B(_1491_),
    .C(_1493_),
    .A(_1489_),
    .Y(_2049_),
    .D(_2048_));
 sg13g2_a21oi_1 _5470_ (.A1(_1411_),
    .A2(_2049_),
    .Y(_2050_),
    .B1(net1051));
 sg13g2_a21oi_1 _5471_ (.A1(net1303),
    .A2(_0736_),
    .Y(_0367_),
    .B1(_2050_));
 sg13g2_a21oi_1 _5472_ (.A1(_1432_),
    .A2(_2049_),
    .Y(_2051_),
    .B1(net1052));
 sg13g2_a21oi_1 _5473_ (.A1(net1303),
    .A2(_0737_),
    .Y(_0368_),
    .B1(_2051_));
 sg13g2_a21oi_2 _5474_ (.B1(net1052),
    .Y(_2052_),
    .A2(_2049_),
    .A1(_1422_));
 sg13g2_a21oi_1 _5475_ (.A1(net1304),
    .A2(_0738_),
    .Y(_0369_),
    .B1(_2052_));
 sg13g2_a21oi_1 _5476_ (.A1(_1436_),
    .A2(_2049_),
    .Y(_2053_),
    .B1(net1051));
 sg13g2_a21oi_1 _5477_ (.A1(net1303),
    .A2(_0739_),
    .Y(_0370_),
    .B1(_2053_));
 sg13g2_a21oi_1 _5478_ (.A1(_1409_),
    .A2(_2049_),
    .Y(_2054_),
    .B1(net1051));
 sg13g2_a21oi_1 _5479_ (.A1(net1302),
    .A2(_0740_),
    .Y(_0371_),
    .B1(_2054_));
 sg13g2_a21oi_1 _5480_ (.A1(_1426_),
    .A2(_2049_),
    .Y(_2055_),
    .B1(net1051));
 sg13g2_a21oi_1 _5481_ (.A1(net1303),
    .A2(_0741_),
    .Y(_0372_),
    .B1(_2055_));
 sg13g2_a21oi_1 _5482_ (.A1(_1429_),
    .A2(_2049_),
    .Y(_2056_),
    .B1(net1051));
 sg13g2_a21oi_1 _5483_ (.A1(net1302),
    .A2(_0742_),
    .Y(_0373_),
    .B1(_2056_));
 sg13g2_a21oi_1 _5484_ (.A1(_1418_),
    .A2(_2049_),
    .Y(_2057_),
    .B1(net1051));
 sg13g2_a21oi_1 _5485_ (.A1(net1302),
    .A2(_0743_),
    .Y(_0374_),
    .B1(_2057_));
 sg13g2_nand2_1 _5486_ (.Y(_2058_),
    .A(net1388),
    .B(net631));
 sg13g2_o21ai_1 _5487_ (.B1(_2058_),
    .Y(_0375_),
    .A1(net1388),
    .A2(_0744_));
 sg13g2_and2_1 _5488_ (.A(net1340),
    .B(net579),
    .X(_0376_));
 sg13g2_o21ai_1 _5489_ (.B1(_1499_),
    .Y(_2059_),
    .A1(net1208),
    .A2(_1710_));
 sg13g2_a21oi_1 _5490_ (.A1(_1501_),
    .A2(_1706_),
    .Y(_2060_),
    .B1(_2059_));
 sg13g2_a21o_1 _5491_ (.A2(net1483),
    .A1(net1320),
    .B1(_2060_),
    .X(_0377_));
 sg13g2_o21ai_1 _5492_ (.B1(_1499_),
    .Y(_2061_),
    .A1(net1208),
    .A2(_1726_));
 sg13g2_a21oi_2 _5493_ (.B1(_2061_),
    .Y(_2062_),
    .A2(_1722_),
    .A1(net1207));
 sg13g2_a21o_1 _5494_ (.A2(net1536),
    .A1(net1315),
    .B1(_2062_),
    .X(_0378_));
 sg13g2_nor2b_1 _5495_ (.A(net1393),
    .B_N(net1616),
    .Y(_2063_));
 sg13g2_nand2_1 _5496_ (.Y(_2064_),
    .A(net1204),
    .B(_1738_));
 sg13g2_a21oi_1 _5497_ (.A1(net1207),
    .A2(_1736_),
    .Y(_2065_),
    .B1(net1133));
 sg13g2_a21o_1 _5498_ (.A2(_2065_),
    .A1(_2064_),
    .B1(_2063_),
    .X(_0379_));
 sg13g2_nor2b_1 _5499_ (.A(net1393),
    .B_N(net1615),
    .Y(_2066_));
 sg13g2_nand2_1 _5500_ (.Y(_2067_),
    .A(net1204),
    .B(_1752_));
 sg13g2_a21oi_1 _5501_ (.A1(net1208),
    .A2(_1749_),
    .Y(_2068_),
    .B1(net1133));
 sg13g2_a21o_1 _5502_ (.A2(_2068_),
    .A1(_2067_),
    .B1(_2066_),
    .X(_0380_));
 sg13g2_nor2b_1 _5503_ (.A(net1393),
    .B_N(net1614),
    .Y(_2069_));
 sg13g2_nand2_1 _5504_ (.Y(_2070_),
    .A(net1204),
    .B(_1766_));
 sg13g2_a21oi_1 _5505_ (.A1(net1208),
    .A2(_1756_),
    .Y(_2071_),
    .B1(net1132));
 sg13g2_a21o_1 _5506_ (.A2(_2071_),
    .A1(_2070_),
    .B1(_2069_),
    .X(_0381_));
 sg13g2_nor2b_1 _5507_ (.A(net1393),
    .B_N(net1617),
    .Y(_2072_));
 sg13g2_nand2_1 _5508_ (.Y(_2073_),
    .A(net1204),
    .B(_1778_));
 sg13g2_a21oi_1 _5509_ (.A1(net1208),
    .A2(_1769_),
    .Y(_2074_),
    .B1(net1132));
 sg13g2_a21o_1 _5510_ (.A2(_2074_),
    .A1(_2073_),
    .B1(_2072_),
    .X(_0382_));
 sg13g2_nor2b_1 _5511_ (.A(net1393),
    .B_N(net1611),
    .Y(_2075_));
 sg13g2_nand2_1 _5512_ (.Y(_2076_),
    .A(net1204),
    .B(_1791_));
 sg13g2_a21oi_1 _5513_ (.A1(net1207),
    .A2(_1781_),
    .Y(_2077_),
    .B1(net1133));
 sg13g2_a21o_1 _5514_ (.A2(_2077_),
    .A1(_2076_),
    .B1(_2075_),
    .X(_0383_));
 sg13g2_a21o_1 _5515_ (.A2(_1794_),
    .A1(net1204),
    .B1(net1132),
    .X(_2078_));
 sg13g2_a21oi_1 _5516_ (.A1(net1208),
    .A2(_1797_),
    .Y(_2079_),
    .B1(_2078_));
 sg13g2_a21o_1 _5517_ (.A2(net1583),
    .A1(net1318),
    .B1(_2079_),
    .X(_0384_));
 sg13g2_nand2_1 _5518_ (.Y(_2080_),
    .A(net1319),
    .B(net679));
 sg13g2_a22oi_1 _5519_ (.Y(_2081_),
    .B1(_1695_),
    .B2(net1275),
    .A2(_1691_),
    .A1(net1207));
 sg13g2_o21ai_1 _5520_ (.B1(_2080_),
    .Y(_0385_),
    .A1(net1133),
    .A2(_2081_));
 sg13g2_nor2_1 _5521_ (.A(net1380),
    .B(net631),
    .Y(_2082_));
 sg13g2_nor2b_1 _5522_ (.A(\main.adder.s4_sum[48] ),
    .B_N(\main.adder.s4_flipped ),
    .Y(_2083_));
 sg13g2_xnor2_1 _5523_ (.Y(_2084_),
    .A(net658),
    .B(_2083_));
 sg13g2_a21oi_1 _5524_ (.A1(net1381),
    .A2(net659),
    .Y(_0386_),
    .B1(_2082_));
 sg13g2_nand4_1 _5525_ (.B(_1645_),
    .C(_1660_),
    .A(_1626_),
    .Y(_2085_),
    .D(_1675_));
 sg13g2_nand2_1 _5526_ (.Y(_2086_),
    .A(_1577_),
    .B(_1604_));
 sg13g2_nor4_1 _5527_ (.A(_1541_),
    .B(_1695_),
    .C(_2085_),
    .D(_2086_),
    .Y(_2087_));
 sg13g2_nand2_1 _5528_ (.Y(_2088_),
    .A(_1738_),
    .B(_1752_));
 sg13g2_nand4_1 _5529_ (.B(_1778_),
    .C(_1791_),
    .A(_1766_),
    .Y(_2089_),
    .D(_1794_));
 sg13g2_nor4_1 _5530_ (.A(_1710_),
    .B(_1726_),
    .C(_2088_),
    .D(_2089_),
    .Y(_2090_));
 sg13g2_a21o_1 _5531_ (.A2(_2090_),
    .A1(_2087_),
    .B1(net1204),
    .X(_2091_));
 sg13g2_nand4_1 _5532_ (.B(_1649_),
    .C(_1664_),
    .A(_1631_),
    .Y(_2092_),
    .D(_1680_));
 sg13g2_nor4_1 _5533_ (.A(_1509_),
    .B(_1548_),
    .C(_1583_),
    .D(_2092_),
    .Y(_2093_));
 sg13g2_a21oi_1 _5534_ (.A1(_2091_),
    .A2(_2093_),
    .Y(_2094_),
    .B1(net1133));
 sg13g2_a21o_1 _5535_ (.A2(net1435),
    .A1(net1320),
    .B1(_2094_),
    .X(_0387_));
 sg13g2_mux2_1 _5536_ (.A0(net828),
    .A1(net780),
    .S(net1388),
    .X(_0388_));
 sg13g2_mux2_1 _5537_ (.A0(net833),
    .A1(net793),
    .S(net1388),
    .X(_0389_));
 sg13g2_nor2_1 _5538_ (.A(net1386),
    .B(net1475),
    .Y(_2095_));
 sg13g2_nand2b_1 _5539_ (.Y(_2096_),
    .B(\main.adder.s4_exponent_adjust[0] ),
    .A_N(\main.adder.s4_exponent[0] ));
 sg13g2_xnor2_1 _5540_ (.Y(_2097_),
    .A(\main.adder.s4_exponent_adjust[0] ),
    .B(\main.adder.s4_exponent[0] ));
 sg13g2_nor4_1 _5541_ (.A(\main.adder.s3_exponent[1] ),
    .B(\main.adder.s3_exponent[0] ),
    .C(\main.adder.s3_exponent[3] ),
    .D(\main.adder.s3_exponent[2] ),
    .Y(_2098_));
 sg13g2_nor4_1 _5542_ (.A(\main.adder.s3_exponent[5] ),
    .B(\main.adder.s3_exponent[4] ),
    .C(\main.adder.s3_exponent[7] ),
    .D(\main.adder.s3_exponent[6] ),
    .Y(_2099_));
 sg13g2_nand3b_1 _5543_ (.B(_2098_),
    .C(_2099_),
    .Y(_2100_),
    .A_N(_1806_));
 sg13g2_nand2_1 _5544_ (.Y(_2101_),
    .A(_2097_),
    .B(_2100_));
 sg13g2_xor2_1 _5545_ (.B(_2100_),
    .A(_2097_),
    .X(_2102_));
 sg13g2_a21oi_1 _5546_ (.A1(net1386),
    .A2(_2102_),
    .Y(_0390_),
    .B1(_2095_));
 sg13g2_nor2b_1 _5547_ (.A(\main.adder.s4_exponent_adjust[1] ),
    .B_N(\main.adder.s4_exponent[1] ),
    .Y(_2103_));
 sg13g2_xnor2_1 _5548_ (.Y(_2104_),
    .A(\main.adder.s4_exponent_adjust[1] ),
    .B(\main.adder.s4_exponent[1] ));
 sg13g2_xor2_1 _5549_ (.B(_2104_),
    .A(_2096_),
    .X(_2105_));
 sg13g2_and2_1 _5550_ (.A(_2101_),
    .B(_2105_),
    .X(_2106_));
 sg13g2_nand2_1 _5551_ (.Y(_2107_),
    .A(net1313),
    .B(net1558));
 sg13g2_o21ai_1 _5552_ (.B1(net1387),
    .Y(_2108_),
    .A1(_2101_),
    .A2(_2105_));
 sg13g2_o21ai_1 _5553_ (.B1(_2107_),
    .Y(_0391_),
    .A1(_2106_),
    .A2(_2108_));
 sg13g2_xor2_1 _5554_ (.B(\main.adder.s4_exponent[2] ),
    .A(net1282),
    .X(_2109_));
 sg13g2_a21oi_1 _5555_ (.A1(_2096_),
    .A2(_2104_),
    .Y(_2110_),
    .B1(_2103_));
 sg13g2_nor2_1 _5556_ (.A(_2109_),
    .B(_2110_),
    .Y(_2111_));
 sg13g2_xor2_1 _5557_ (.B(_2110_),
    .A(_2109_),
    .X(_2112_));
 sg13g2_nand2_1 _5558_ (.Y(_2113_),
    .A(_2106_),
    .B(_2112_));
 sg13g2_xnor2_1 _5559_ (.Y(_2114_),
    .A(_2106_),
    .B(_2112_));
 sg13g2_nor2_1 _5560_ (.A(net1386),
    .B(net910),
    .Y(_2115_));
 sg13g2_a21oi_1 _5561_ (.A1(net1386),
    .A2(_2114_),
    .Y(_0392_),
    .B1(_2115_));
 sg13g2_nor2b_1 _5562_ (.A(net1387),
    .B_N(net1605),
    .Y(_2116_));
 sg13g2_xor2_1 _5563_ (.B(\main.adder.s4_exponent[3] ),
    .A(net1281),
    .X(_2117_));
 sg13g2_a21oi_1 _5564_ (.A1(_0715_),
    .A2(\main.adder.s4_exponent[2] ),
    .Y(_2118_),
    .B1(_2111_));
 sg13g2_nor2_1 _5565_ (.A(_2117_),
    .B(_2118_),
    .Y(_2119_));
 sg13g2_xnor2_1 _5566_ (.Y(_2120_),
    .A(_2117_),
    .B(_2118_));
 sg13g2_or2_1 _5567_ (.X(_2121_),
    .B(_2120_),
    .A(_2113_));
 sg13g2_a21oi_1 _5568_ (.A1(_2113_),
    .A2(_2120_),
    .Y(_2122_),
    .B1(net1313));
 sg13g2_a21o_1 _5569_ (.A2(_2122_),
    .A1(_2121_),
    .B1(_2116_),
    .X(_0393_));
 sg13g2_nand2b_1 _5570_ (.Y(_2123_),
    .B(\main.adder.s4_exponent[4] ),
    .A_N(net1277));
 sg13g2_xor2_1 _5571_ (.B(\main.adder.s4_exponent[4] ),
    .A(net1277),
    .X(_2124_));
 sg13g2_a21oi_1 _5572_ (.A1(_0716_),
    .A2(\main.adder.s4_exponent[3] ),
    .Y(_2125_),
    .B1(_2119_));
 sg13g2_xnor2_1 _5573_ (.Y(_2126_),
    .A(_2124_),
    .B(_2125_));
 sg13g2_or2_1 _5574_ (.X(_2127_),
    .B(_2126_),
    .A(_2121_));
 sg13g2_nor2b_1 _5575_ (.A(net1386),
    .B_N(net1609),
    .Y(_2128_));
 sg13g2_a21oi_1 _5576_ (.A1(_2121_),
    .A2(_2126_),
    .Y(_2129_),
    .B1(net1313));
 sg13g2_a21o_1 _5577_ (.A2(_2129_),
    .A1(_2127_),
    .B1(_2128_),
    .X(_0394_));
 sg13g2_nor2_1 _5578_ (.A(net1386),
    .B(_0711_),
    .Y(_2130_));
 sg13g2_o21ai_1 _5579_ (.B1(_2123_),
    .Y(_2131_),
    .A1(_2124_),
    .A2(_2125_));
 sg13g2_nor2b_1 _5580_ (.A(\main.adder.s4_exponent_adjust[5] ),
    .B_N(\main.adder.s4_exponent[5] ),
    .Y(_2132_));
 sg13g2_xnor2_1 _5581_ (.Y(_2133_),
    .A(\main.adder.s4_exponent_adjust[5] ),
    .B(\main.adder.s4_exponent[5] ));
 sg13g2_xnor2_1 _5582_ (.Y(_2134_),
    .A(_2131_),
    .B(_2133_));
 sg13g2_or2_1 _5583_ (.X(_2135_),
    .B(_2134_),
    .A(_2127_));
 sg13g2_a21oi_1 _5584_ (.A1(_2127_),
    .A2(_2134_),
    .Y(_2136_),
    .B1(net1315));
 sg13g2_a21o_1 _5585_ (.A2(_2136_),
    .A1(_2135_),
    .B1(_2130_),
    .X(_0395_));
 sg13g2_nand2_1 _5586_ (.Y(_2137_),
    .A(net1315),
    .B(net934));
 sg13g2_xor2_1 _5587_ (.B(\main.adder.s4_exponent[6] ),
    .A(\main.adder.s4_exponent_adjust[6] ),
    .X(_2138_));
 sg13g2_a21oi_2 _5588_ (.B1(_2132_),
    .Y(_2139_),
    .A2(_2133_),
    .A1(_2131_));
 sg13g2_nor2_1 _5589_ (.A(_2138_),
    .B(_2139_),
    .Y(_2140_));
 sg13g2_xnor2_1 _5590_ (.Y(_2141_),
    .A(_2138_),
    .B(_2139_));
 sg13g2_nor2_2 _5591_ (.A(_2135_),
    .B(_2141_),
    .Y(_2142_));
 sg13g2_a21o_1 _5592_ (.A2(_2141_),
    .A1(_2135_),
    .B1(net1315),
    .X(_2143_));
 sg13g2_o21ai_1 _5593_ (.B1(_2137_),
    .Y(_0396_),
    .A1(_2142_),
    .A2(_2143_));
 sg13g2_a21oi_1 _5594_ (.A1(_0714_),
    .A2(\main.adder.s4_exponent[6] ),
    .Y(_2144_),
    .B1(_2140_));
 sg13g2_inv_1 _5595_ (.Y(_2145_),
    .A(_2144_));
 sg13g2_nor2b_1 _5596_ (.A(\main.adder.s4_exponent_adjust[7] ),
    .B_N(\main.adder.s4_exponent[7] ),
    .Y(_2146_));
 sg13g2_xnor2_1 _5597_ (.Y(_2147_),
    .A(\main.adder.s4_exponent_adjust[7] ),
    .B(\main.adder.s4_exponent[7] ));
 sg13g2_xnor2_1 _5598_ (.Y(_2148_),
    .A(_2144_),
    .B(_2147_));
 sg13g2_xnor2_1 _5599_ (.Y(_2149_),
    .A(_2142_),
    .B(_2148_));
 sg13g2_nor2_1 _5600_ (.A(net1386),
    .B(net903),
    .Y(_2150_));
 sg13g2_a21oi_1 _5601_ (.A1(net1386),
    .A2(_2149_),
    .Y(_0397_),
    .B1(_2150_));
 sg13g2_a21oi_1 _5602_ (.A1(_2145_),
    .A2(_2147_),
    .Y(_2151_),
    .B1(_2146_));
 sg13g2_xnor2_1 _5603_ (.Y(_2152_),
    .A(_0073_),
    .B(_2151_));
 sg13g2_nand3_1 _5604_ (.B(_2148_),
    .C(_2152_),
    .A(_2142_),
    .Y(_2153_));
 sg13g2_a21o_1 _5605_ (.A2(_2148_),
    .A1(_2142_),
    .B1(_2152_),
    .X(_2154_));
 sg13g2_a21oi_1 _5606_ (.A1(_2153_),
    .A2(_2154_),
    .Y(_2155_),
    .B1(net1315));
 sg13g2_a21oi_1 _5607_ (.A1(net1315),
    .A2(_0712_),
    .Y(_0398_),
    .B1(_2155_));
 sg13g2_nor2_1 _5608_ (.A(\main.adder.s4_exponent_adjust[8] ),
    .B(_2151_),
    .Y(_2156_));
 sg13g2_xnor2_1 _5609_ (.Y(_2157_),
    .A(\main.adder.s4_exponent_adjust[9] ),
    .B(_2156_));
 sg13g2_xnor2_1 _5610_ (.Y(_2158_),
    .A(_2153_),
    .B(_2157_));
 sg13g2_mux2_1 _5611_ (.A0(net1520),
    .A1(_2158_),
    .S(net1392),
    .X(_0399_));
 sg13g2_and2_1 _5612_ (.A(net1338),
    .B(net580),
    .X(_0400_));
 sg13g2_mux2_1 _5613_ (.A0(net718),
    .A1(\main.adder.s3_flipped ),
    .S(net1354),
    .X(_0401_));
 sg13g2_mux2_1 _5614_ (.A0(net658),
    .A1(net829),
    .S(net1379),
    .X(_0402_));
 sg13g2_mux2_1 _5615_ (.A0(net780),
    .A1(\main.adder.s3_nan ),
    .S(net1388),
    .X(_0403_));
 sg13g2_mux2_1 _5616_ (.A0(net793),
    .A1(net779),
    .S(net1388),
    .X(_0404_));
 sg13g2_nor2_1 _5617_ (.A(net1390),
    .B(net609),
    .Y(_2159_));
 sg13g2_a21oi_1 _5618_ (.A1(net1390),
    .A2(_1293_),
    .Y(_0405_),
    .B1(_2159_));
 sg13g2_nor2_1 _5619_ (.A(net1390),
    .B(net635),
    .Y(_2160_));
 sg13g2_a21oi_1 _5620_ (.A1(net1390),
    .A2(_1285_),
    .Y(_0406_),
    .B1(_2160_));
 sg13g2_nor2_1 _5621_ (.A(net1390),
    .B(net613),
    .Y(_2161_));
 sg13g2_a21oi_1 _5622_ (.A1(net1390),
    .A2(_1276_),
    .Y(_0407_),
    .B1(_2161_));
 sg13g2_mux2_1 _5623_ (.A0(net666),
    .A1(_1261_),
    .S(net1359),
    .X(_0408_));
 sg13g2_nor2_1 _5624_ (.A(net1390),
    .B(net605),
    .Y(_2162_));
 sg13g2_a21oi_1 _5625_ (.A1(net1366),
    .A2(_1265_),
    .Y(_0409_),
    .B1(_2162_));
 sg13g2_nor2_1 _5626_ (.A(net1368),
    .B(net597),
    .Y(_2163_));
 sg13g2_a21oi_1 _5627_ (.A1(net1368),
    .A2(_1253_),
    .Y(_0410_),
    .B1(_2163_));
 sg13g2_mux2_1 _5628_ (.A0(net662),
    .A1(_1249_),
    .S(net1368),
    .X(_0411_));
 sg13g2_nor2_1 _5629_ (.A(net1366),
    .B(net586),
    .Y(_2164_));
 sg13g2_a21oi_1 _5630_ (.A1(net1366),
    .A2(_1240_),
    .Y(_0412_),
    .B1(_2164_));
 sg13g2_nor2_1 _5631_ (.A(net1366),
    .B(net593),
    .Y(_2165_));
 sg13g2_a21oi_1 _5632_ (.A1(net1366),
    .A2(_1218_),
    .Y(_0413_),
    .B1(_2165_));
 sg13g2_nor2_1 _5633_ (.A(net1366),
    .B(net595),
    .Y(_2166_));
 sg13g2_a21oi_1 _5634_ (.A1(net1366),
    .A2(_1211_),
    .Y(_0414_),
    .B1(_2166_));
 sg13g2_nor2_1 _5635_ (.A(net1367),
    .B(net621),
    .Y(_2167_));
 sg13g2_a21oi_1 _5636_ (.A1(net1366),
    .A2(_1224_),
    .Y(_0415_),
    .B1(_2167_));
 sg13g2_nor2_1 _5637_ (.A(net1367),
    .B(net592),
    .Y(_2168_));
 sg13g2_a21oi_1 _5638_ (.A1(net1367),
    .A2(_1235_),
    .Y(_0416_),
    .B1(_2168_));
 sg13g2_nor2_1 _5639_ (.A(net1367),
    .B(net611),
    .Y(_2169_));
 sg13g2_a21oi_1 _5640_ (.A1(net1367),
    .A2(_1231_),
    .Y(_0417_),
    .B1(_2169_));
 sg13g2_mux2_1 _5641_ (.A0(net624),
    .A1(_1204_),
    .S(net1367),
    .X(_0418_));
 sg13g2_mux2_1 _5642_ (.A0(net625),
    .A1(_1199_),
    .S(net1367),
    .X(_0419_));
 sg13g2_nor2_1 _5643_ (.A(net1363),
    .B(net603),
    .Y(_2170_));
 sg13g2_a21oi_1 _5644_ (.A1(net1363),
    .A2(_1158_),
    .Y(_0420_),
    .B1(_2170_));
 sg13g2_nor2_1 _5645_ (.A(net1370),
    .B(net590),
    .Y(_2171_));
 sg13g2_a21oi_1 _5646_ (.A1(net1370),
    .A2(_1189_),
    .Y(_0421_),
    .B1(_2171_));
 sg13g2_nor2_1 _5647_ (.A(net1376),
    .B(net599),
    .Y(_2172_));
 sg13g2_a21oi_1 _5648_ (.A1(net1376),
    .A2(_1183_),
    .Y(_0422_),
    .B1(_2172_));
 sg13g2_nor2_1 _5649_ (.A(net1376),
    .B(net607),
    .Y(_2173_));
 sg13g2_a21oi_1 _5650_ (.A1(net1376),
    .A2(_1164_),
    .Y(_0423_),
    .B1(_2173_));
 sg13g2_nor2_1 _5651_ (.A(net1376),
    .B(net617),
    .Y(_2174_));
 sg13g2_a21oi_1 _5652_ (.A1(net1376),
    .A2(_1174_),
    .Y(_0424_),
    .B1(_2174_));
 sg13g2_nor2_1 _5653_ (.A(net1375),
    .B(net799),
    .Y(_2175_));
 sg13g2_a21oi_1 _5654_ (.A1(net1375),
    .A2(_1186_),
    .Y(_0425_),
    .B1(_2175_));
 sg13g2_nor2_1 _5655_ (.A(net1372),
    .B(net1540),
    .Y(_2176_));
 sg13g2_a21oi_1 _5656_ (.A1(net1372),
    .A2(_1145_),
    .Y(_0426_),
    .B1(_2176_));
 sg13g2_nor2_1 _5657_ (.A(net1374),
    .B(net1499),
    .Y(_2177_));
 sg13g2_a21oi_1 _5658_ (.A1(net1374),
    .A2(_1161_),
    .Y(_0427_),
    .B1(_2177_));
 sg13g2_nor2_1 _5659_ (.A(net1371),
    .B(net1562),
    .Y(_2178_));
 sg13g2_a21oi_1 _5660_ (.A1(net1371),
    .A2(_1153_),
    .Y(_0428_),
    .B1(_2178_));
 sg13g2_nor2_1 _5661_ (.A(net1372),
    .B(net1564),
    .Y(_2179_));
 sg13g2_a21oi_1 _5662_ (.A1(net1372),
    .A2(_1167_),
    .Y(_0429_),
    .B1(_2179_));
 sg13g2_nor2_1 _5663_ (.A(net1371),
    .B(net1517),
    .Y(_2180_));
 sg13g2_a21oi_1 _5664_ (.A1(net1371),
    .A2(_1171_),
    .Y(_0430_),
    .B1(_2180_));
 sg13g2_nor2_1 _5665_ (.A(net1372),
    .B(net1467),
    .Y(_2181_));
 sg13g2_a21oi_1 _5666_ (.A1(net1372),
    .A2(_1181_),
    .Y(_0431_),
    .B1(_2181_));
 sg13g2_nor2_1 _5667_ (.A(net1363),
    .B(net1509),
    .Y(_2182_));
 sg13g2_a21oi_1 _5668_ (.A1(net1364),
    .A2(_1169_),
    .Y(_0432_),
    .B1(_2182_));
 sg13g2_nor2_1 _5669_ (.A(net1371),
    .B(net1444),
    .Y(_2183_));
 sg13g2_a21oi_1 _5670_ (.A1(net1371),
    .A2(_1177_),
    .Y(_0433_),
    .B1(_2183_));
 sg13g2_nor2_1 _5671_ (.A(net1371),
    .B(net824),
    .Y(_2184_));
 sg13g2_a21oi_1 _5672_ (.A1(net1373),
    .A2(_1151_),
    .Y(_0434_),
    .B1(_2184_));
 sg13g2_nor2_1 _5673_ (.A(net1373),
    .B(net1464),
    .Y(_2185_));
 sg13g2_a21oi_1 _5674_ (.A1(net1373),
    .A2(_1156_),
    .Y(_0435_),
    .B1(_2185_));
 sg13g2_nor2_1 _5675_ (.A(net1364),
    .B(net935),
    .Y(_2186_));
 sg13g2_a21oi_1 _5676_ (.A1(net1363),
    .A2(_1121_),
    .Y(_0436_),
    .B1(_2186_));
 sg13g2_nor2_1 _5677_ (.A(net1373),
    .B(net1403),
    .Y(_2187_));
 sg13g2_a21oi_1 _5678_ (.A1(net1373),
    .A2(_1117_),
    .Y(_0437_),
    .B1(_2187_));
 sg13g2_nor2_1 _5679_ (.A(net1372),
    .B(net850),
    .Y(_2188_));
 sg13g2_a21oi_1 _5680_ (.A1(net1372),
    .A2(_1130_),
    .Y(_0438_),
    .B1(_2188_));
 sg13g2_nor2_1 _5681_ (.A(net1374),
    .B(net945),
    .Y(_2189_));
 sg13g2_a21oi_1 _5682_ (.A1(net1374),
    .A2(_1125_),
    .Y(_0439_),
    .B1(_2189_));
 sg13g2_nor2_1 _5683_ (.A(net1375),
    .B(net649),
    .Y(_2190_));
 sg13g2_a21oi_1 _5684_ (.A1(net1374),
    .A2(_1104_),
    .Y(_0440_),
    .B1(_2190_));
 sg13g2_nor2_1 _5685_ (.A(net1374),
    .B(net1046),
    .Y(_2191_));
 sg13g2_a21oi_1 _5686_ (.A1(net1375),
    .A2(_1119_),
    .Y(_0441_),
    .B1(_2191_));
 sg13g2_nor2_1 _5687_ (.A(net1375),
    .B(net637),
    .Y(_2192_));
 sg13g2_a21oi_1 _5688_ (.A1(net1374),
    .A2(_1128_),
    .Y(_0442_),
    .B1(_2192_));
 sg13g2_mux2_1 _5689_ (.A0(net1407),
    .A1(_1110_),
    .S(net1374),
    .X(_0443_));
 sg13g2_nor2_1 _5690_ (.A(net1371),
    .B(net1496),
    .Y(_2193_));
 sg13g2_a21oi_1 _5691_ (.A1(net1370),
    .A2(_1123_),
    .Y(_0444_),
    .B1(_2193_));
 sg13g2_nor2_1 _5692_ (.A(net1369),
    .B(net1485),
    .Y(_2194_));
 sg13g2_a21oi_1 _5693_ (.A1(net1370),
    .A2(_1127_),
    .Y(_0445_),
    .B1(_2194_));
 sg13g2_nor2_1 _5694_ (.A(net1370),
    .B(net938),
    .Y(_2195_));
 sg13g2_a21oi_1 _5695_ (.A1(net1370),
    .A2(_1106_),
    .Y(_0446_),
    .B1(_2195_));
 sg13g2_nor2_1 _5696_ (.A(net1369),
    .B(net1523),
    .Y(_2196_));
 sg13g2_a21oi_1 _5697_ (.A1(net1369),
    .A2(_1100_),
    .Y(_0447_),
    .B1(_2196_));
 sg13g2_nor2_1 _5698_ (.A(net1369),
    .B(net954),
    .Y(_2197_));
 sg13g2_a21oi_1 _5699_ (.A1(net1369),
    .A2(_1105_),
    .Y(_0448_),
    .B1(_2197_));
 sg13g2_nor2_1 _5700_ (.A(net1369),
    .B(net1472),
    .Y(_2198_));
 sg13g2_a21oi_1 _5701_ (.A1(net1369),
    .A2(_1112_),
    .Y(_0449_),
    .B1(_2198_));
 sg13g2_nor2_1 _5702_ (.A(net1376),
    .B(net1415),
    .Y(_2199_));
 sg13g2_a21oi_1 _5703_ (.A1(net1367),
    .A2(_1114_),
    .Y(_0450_),
    .B1(_2199_));
 sg13g2_nor2_1 _5704_ (.A(net1369),
    .B(net980),
    .Y(_2200_));
 sg13g2_a21oi_1 _5705_ (.A1(net1377),
    .A2(_1095_),
    .Y(_0451_),
    .B1(_2200_));
 sg13g2_mux2_1 _5706_ (.A0(net633),
    .A1(\main.adder.s3_sum[0] ),
    .S(net1383),
    .X(_0452_));
 sg13g2_nor2_1 _5707_ (.A(net1358),
    .B(net660),
    .Y(_2201_));
 sg13g2_a21oi_1 _5708_ (.A1(_0687_),
    .A2(net1357),
    .Y(_0453_),
    .B1(_2201_));
 sg13g2_and2_1 _5709_ (.A(net1338),
    .B(net585),
    .X(_0454_));
 sg13g2_mux2_1 _5710_ (.A0(\main.adder.s3_nan ),
    .A1(net782),
    .S(net1388),
    .X(_0455_));
 sg13g2_mux2_1 _5711_ (.A0(net779),
    .A1(net756),
    .S(net1388),
    .X(_0456_));
 sg13g2_mux2_1 _5712_ (.A0(net778),
    .A1(net1258),
    .S(net1354),
    .X(_0457_));
 sg13g2_mux2_1 _5713_ (.A0(\main.adder.s3_shared_sign ),
    .A1(net726),
    .S(net1354),
    .X(_0458_));
 sg13g2_mux2_1 _5714_ (.A0(net866),
    .A1(net714),
    .S(net1358),
    .X(_0459_));
 sg13g2_mux2_1 _5715_ (.A0(net877),
    .A1(net694),
    .S(net1357),
    .X(_0460_));
 sg13g2_mux2_1 _5716_ (.A0(net919),
    .A1(net697),
    .S(net1358),
    .X(_0461_));
 sg13g2_nor2_1 _5717_ (.A(net929),
    .B(net1359),
    .Y(_2202_));
 sg13g2_a21oi_1 _5718_ (.A1(net1357),
    .A2(_0760_),
    .Y(_0462_),
    .B1(_2202_));
 sg13g2_mux2_1 _5719_ (.A0(net831),
    .A1(net777),
    .S(net1357),
    .X(_0463_));
 sg13g2_mux2_1 _5720_ (.A0(net814),
    .A1(net768),
    .S(net1359),
    .X(_0464_));
 sg13g2_mux2_1 _5721_ (.A0(\main.adder.s3_sum[6] ),
    .A1(net730),
    .S(net1354),
    .X(_0465_));
 sg13g2_nor2_1 _5722_ (.A(net707),
    .B(net1356),
    .Y(_2203_));
 sg13g2_a21oi_1 _5723_ (.A1(net1356),
    .A2(_0761_),
    .Y(_0466_),
    .B1(_2203_));
 sg13g2_nor2_1 _5724_ (.A(net751),
    .B(net1355),
    .Y(_2204_));
 sg13g2_a21oi_1 _5725_ (.A1(net1355),
    .A2(_0762_),
    .Y(_0467_),
    .B1(_2204_));
 sg13g2_nor2_1 _5726_ (.A(net795),
    .B(net1356),
    .Y(_2205_));
 sg13g2_a21oi_1 _5727_ (.A1(net1355),
    .A2(_0763_),
    .Y(_0468_),
    .B1(_2205_));
 sg13g2_mux2_1 _5728_ (.A0(net924),
    .A1(net743),
    .S(net1353),
    .X(_0469_));
 sg13g2_mux2_1 _5729_ (.A0(\main.adder.s3_sum[11] ),
    .A1(net1396),
    .S(net1355),
    .X(_0470_));
 sg13g2_nand2_1 _5730_ (.Y(_2206_),
    .A(net1352),
    .B(net705));
 sg13g2_o21ai_1 _5731_ (.B1(_2206_),
    .Y(_0471_),
    .A1(_0682_),
    .A2(net1355));
 sg13g2_mux2_1 _5732_ (.A0(\main.adder.s3_sum[13] ),
    .A1(net883),
    .S(net1356),
    .X(_0472_));
 sg13g2_mux2_1 _5733_ (.A0(\main.adder.s3_sum[14] ),
    .A1(net864),
    .S(net1356),
    .X(_0473_));
 sg13g2_nand2_1 _5734_ (.Y(_2207_),
    .A(net1362),
    .B(net927));
 sg13g2_o21ai_1 _5735_ (.B1(_2207_),
    .Y(_0474_),
    .A1(_0681_),
    .A2(net1361));
 sg13g2_mux2_1 _5736_ (.A0(\main.adder.s3_sum[16] ),
    .A1(net906),
    .S(net1350),
    .X(_0475_));
 sg13g2_mux2_1 _5737_ (.A0(\main.adder.s3_sum[17] ),
    .A1(net1020),
    .S(net1350),
    .X(_0476_));
 sg13g2_mux2_1 _5738_ (.A0(\main.adder.s3_sum[18] ),
    .A1(net982),
    .S(net1350),
    .X(_0477_));
 sg13g2_nor2_1 _5739_ (.A(net716),
    .B(net1349),
    .Y(_2208_));
 sg13g2_a21oi_1 _5740_ (.A1(net1349),
    .A2(_0757_),
    .Y(_0478_),
    .B1(_2208_));
 sg13g2_mux2_1 _5741_ (.A0(\main.adder.s3_sum[20] ),
    .A1(net1566),
    .S(net1363),
    .X(_0479_));
 sg13g2_nor2_1 _5742_ (.A(net1497),
    .B(net1363),
    .Y(_2209_));
 sg13g2_a21oi_1 _5743_ (.A1(net1363),
    .A2(_0758_),
    .Y(_0480_),
    .B1(_2209_));
 sg13g2_nor2_1 _5744_ (.A(net689),
    .B(net1364),
    .Y(_2210_));
 sg13g2_a21oi_1 _5745_ (.A1(net1364),
    .A2(_0759_),
    .Y(_0481_),
    .B1(_2210_));
 sg13g2_and2_1 _5746_ (.A(\main.adder.s2_smaler[23] ),
    .B(\main.adder.s2_larger[23] ),
    .X(_2211_));
 sg13g2_xor2_1 _5747_ (.B(\main.adder.s2_larger[23] ),
    .A(\main.adder.s2_smaler[23] ),
    .X(_2212_));
 sg13g2_mux2_1 _5748_ (.A0(net904),
    .A1(_2212_),
    .S(net1362),
    .X(_0482_));
 sg13g2_nor2_1 _5749_ (.A(net776),
    .B(net1362),
    .Y(_2213_));
 sg13g2_nor2_1 _5750_ (.A(net1256),
    .B(_0099_),
    .Y(_2214_));
 sg13g2_nor2_1 _5751_ (.A(\main.adder.s2_larger[23] ),
    .B(\main.adder.s2_larger[24] ),
    .Y(_2215_));
 sg13g2_xor2_1 _5752_ (.B(\main.adder.s2_larger[24] ),
    .A(\main.adder.s2_larger[23] ),
    .X(_2216_));
 sg13g2_a21oi_2 _5753_ (.B1(_2214_),
    .Y(_2217_),
    .A2(_2216_),
    .A1(net1256));
 sg13g2_nor2b_1 _5754_ (.A(_2217_),
    .B_N(\main.adder.s2_smaler[24] ),
    .Y(_2218_));
 sg13g2_xnor2_1 _5755_ (.Y(_2219_),
    .A(\main.adder.s2_smaler[24] ),
    .B(_2217_));
 sg13g2_xnor2_1 _5756_ (.Y(_2220_),
    .A(_2211_),
    .B(_2219_));
 sg13g2_a21oi_1 _5757_ (.A1(net1362),
    .A2(_2220_),
    .Y(_0483_),
    .B1(_2213_));
 sg13g2_a21oi_1 _5758_ (.A1(_2211_),
    .A2(_2219_),
    .Y(_2221_),
    .B1(_2218_));
 sg13g2_nor2_1 _5759_ (.A(net1256),
    .B(_0101_),
    .Y(_2222_));
 sg13g2_xnor2_1 _5760_ (.Y(_2223_),
    .A(\main.adder.s2_larger[25] ),
    .B(_2215_));
 sg13g2_a21o_1 _5761_ (.A2(_2223_),
    .A1(net1256),
    .B1(_2222_),
    .X(_2224_));
 sg13g2_nand2_1 _5762_ (.Y(_2225_),
    .A(\main.adder.s2_smaler[25] ),
    .B(_2224_));
 sg13g2_xnor2_1 _5763_ (.Y(_2226_),
    .A(\main.adder.s2_smaler[25] ),
    .B(_2224_));
 sg13g2_xnor2_1 _5764_ (.Y(_2227_),
    .A(_2221_),
    .B(_2226_));
 sg13g2_nor2_1 _5765_ (.A(net963),
    .B(net1362),
    .Y(_2228_));
 sg13g2_a21oi_1 _5766_ (.A1(net1362),
    .A2(_2227_),
    .Y(_0484_),
    .B1(_2228_));
 sg13g2_o21ai_1 _5767_ (.B1(_2225_),
    .Y(_2229_),
    .A1(_2221_),
    .A2(_2226_));
 sg13g2_nor2_1 _5768_ (.A(\main.adder.s2_larger[24] ),
    .B(\main.adder.s2_larger[25] ),
    .Y(_2230_));
 sg13g2_nand2_1 _5769_ (.Y(_2231_),
    .A(_0103_),
    .B(_2230_));
 sg13g2_xnor2_1 _5770_ (.Y(_2232_),
    .A(\main.adder.s2_larger[26] ),
    .B(_2231_));
 sg13g2_mux2_1 _5771_ (.A0(_0102_),
    .A1(_2232_),
    .S(net1258),
    .X(_2233_));
 sg13g2_nor2b_1 _5772_ (.A(_2233_),
    .B_N(\main.adder.s2_smaler[26] ),
    .Y(_2234_));
 sg13g2_nand2b_1 _5773_ (.Y(_2235_),
    .B(_2233_),
    .A_N(\main.adder.s2_smaler[26] ));
 sg13g2_nand2b_1 _5774_ (.Y(_2236_),
    .B(_2235_),
    .A_N(_2234_));
 sg13g2_xnor2_1 _5775_ (.Y(_2237_),
    .A(_2229_),
    .B(_2236_));
 sg13g2_mux2_1 _5776_ (.A0(net1587),
    .A1(_2237_),
    .S(net1363),
    .X(_0485_));
 sg13g2_a21oi_1 _5777_ (.A1(_2229_),
    .A2(_2235_),
    .Y(_2238_),
    .B1(_2234_));
 sg13g2_o21ai_1 _5778_ (.B1(\main.adder.s2_larger[27] ),
    .Y(_2239_),
    .A1(\main.adder.s2_larger[26] ),
    .A2(_2231_));
 sg13g2_nand4_1 _5779_ (.B(_0103_),
    .C(_0748_),
    .A(_0747_),
    .Y(_2240_),
    .D(_2230_));
 sg13g2_nand3_1 _5780_ (.B(_2239_),
    .C(_2240_),
    .A(net1256),
    .Y(_2241_));
 sg13g2_o21ai_1 _5781_ (.B1(_2241_),
    .Y(_2242_),
    .A1(net1256),
    .A2(_0104_));
 sg13g2_nand2_1 _5782_ (.Y(_2243_),
    .A(\main.adder.s2_smaler[27] ),
    .B(_2242_));
 sg13g2_nor2_1 _5783_ (.A(\main.adder.s2_smaler[27] ),
    .B(_2242_),
    .Y(_2244_));
 sg13g2_xnor2_1 _5784_ (.Y(_2245_),
    .A(\main.adder.s2_smaler[27] ),
    .B(_2242_));
 sg13g2_xnor2_1 _5785_ (.Y(_2246_),
    .A(_2238_),
    .B(_2245_));
 sg13g2_nor2_1 _5786_ (.A(net1547),
    .B(net1365),
    .Y(_2247_));
 sg13g2_a21oi_1 _5787_ (.A1(net1365),
    .A2(_2246_),
    .Y(_0486_),
    .B1(_2247_));
 sg13g2_o21ai_1 _5788_ (.B1(_2243_),
    .Y(_2248_),
    .A1(_2238_),
    .A2(_2244_));
 sg13g2_nand2_1 _5789_ (.Y(_2249_),
    .A(\main.adder.s2_larger[28] ),
    .B(_2240_));
 sg13g2_or2_2 _5790_ (.X(_2250_),
    .B(_2240_),
    .A(\main.adder.s2_larger[28] ));
 sg13g2_nand3_1 _5791_ (.B(_2249_),
    .C(_2250_),
    .A(net1254),
    .Y(_2251_));
 sg13g2_o21ai_1 _5792_ (.B1(_2251_),
    .Y(_2252_),
    .A1(net1254),
    .A2(_0105_));
 sg13g2_and2_1 _5793_ (.A(\main.adder.s2_smaler[28] ),
    .B(_2252_),
    .X(_2253_));
 sg13g2_xnor2_1 _5794_ (.Y(_2254_),
    .A(\main.adder.s2_smaler[28] ),
    .B(_2252_));
 sg13g2_inv_1 _5795_ (.Y(_2255_),
    .A(_2254_));
 sg13g2_xnor2_1 _5796_ (.Y(_2256_),
    .A(_2248_),
    .B(_2255_));
 sg13g2_nor2_1 _5797_ (.A(net1533),
    .B(net1365),
    .Y(_2257_));
 sg13g2_a21oi_1 _5798_ (.A1(net1365),
    .A2(_2256_),
    .Y(_0487_),
    .B1(_2257_));
 sg13g2_nor2_1 _5799_ (.A(net1530),
    .B(net1365),
    .Y(_2258_));
 sg13g2_a21oi_1 _5800_ (.A1(_2248_),
    .A2(_2255_),
    .Y(_2259_),
    .B1(_2253_));
 sg13g2_xnor2_1 _5801_ (.Y(_2260_),
    .A(\main.adder.s2_larger[29] ),
    .B(_2250_));
 sg13g2_nor2b_1 _5802_ (.A(net1254),
    .B_N(_0106_),
    .Y(_2261_));
 sg13g2_a21oi_2 _5803_ (.B1(_2261_),
    .Y(_2262_),
    .A2(_2260_),
    .A1(net1254));
 sg13g2_nor2_1 _5804_ (.A(\main.adder.s2_smaler[29] ),
    .B(_2262_),
    .Y(_2263_));
 sg13g2_xnor2_1 _5805_ (.Y(_2264_),
    .A(\main.adder.s2_smaler[29] ),
    .B(_2262_));
 sg13g2_xnor2_1 _5806_ (.Y(_2265_),
    .A(_2259_),
    .B(_2264_));
 sg13g2_a21oi_1 _5807_ (.A1(net1365),
    .A2(_2265_),
    .Y(_0488_),
    .B1(_2258_));
 sg13g2_o21ai_1 _5808_ (.B1(\main.adder.s2_larger[30] ),
    .Y(_2266_),
    .A1(\main.adder.s2_larger[29] ),
    .A2(_2250_));
 sg13g2_nor3_2 _5809_ (.A(\main.adder.s2_larger[29] ),
    .B(\main.adder.s2_larger[30] ),
    .C(_2250_),
    .Y(_2267_));
 sg13g2_nand3b_1 _5810_ (.B(net1254),
    .C(_2266_),
    .Y(_2268_),
    .A_N(_2267_));
 sg13g2_o21ai_1 _5811_ (.B1(_2268_),
    .Y(_2269_),
    .A1(net1254),
    .A2(_0107_));
 sg13g2_nand2_1 _5812_ (.Y(_2270_),
    .A(\main.adder.s2_smaler[30] ),
    .B(_2269_));
 sg13g2_xnor2_1 _5813_ (.Y(_2271_),
    .A(\main.adder.s2_smaler[30] ),
    .B(_2269_));
 sg13g2_a221oi_1 _5814_ (.B2(\main.adder.s2_smaler[29] ),
    .C1(_2253_),
    .B1(_2262_),
    .A1(_2248_),
    .Y(_2272_),
    .A2(_2255_));
 sg13g2_or3_1 _5815_ (.A(_2263_),
    .B(_2271_),
    .C(_2272_),
    .X(_2273_));
 sg13g2_o21ai_1 _5816_ (.B1(_2271_),
    .Y(_2274_),
    .A1(_2263_),
    .A2(_2272_));
 sg13g2_and2_1 _5817_ (.A(net1347),
    .B(_2274_),
    .X(_2275_));
 sg13g2_a22oi_1 _5818_ (.Y(_2276_),
    .B1(_2273_),
    .B2(_2275_),
    .A2(net1308),
    .A1(net1424));
 sg13g2_inv_1 _5819_ (.Y(_0489_),
    .A(_2276_));
 sg13g2_nor2_1 _5820_ (.A(net1252),
    .B(_0108_),
    .Y(_2277_));
 sg13g2_nand2b_2 _5821_ (.Y(_2278_),
    .B(_2267_),
    .A_N(\main.adder.s2_larger[31] ));
 sg13g2_xnor2_1 _5822_ (.Y(_2279_),
    .A(\main.adder.s2_larger[31] ),
    .B(_2267_));
 sg13g2_a21oi_2 _5823_ (.B1(_2277_),
    .Y(_2280_),
    .A2(_2279_),
    .A1(net1252));
 sg13g2_nand2b_1 _5824_ (.Y(_2281_),
    .B(\main.adder.s2_smaler[31] ),
    .A_N(_2280_));
 sg13g2_xor2_1 _5825_ (.B(_2280_),
    .A(\main.adder.s2_smaler[31] ),
    .X(_2282_));
 sg13g2_a21o_1 _5826_ (.A2(_2273_),
    .A1(_2270_),
    .B1(_2282_),
    .X(_2283_));
 sg13g2_nand3_1 _5827_ (.B(_2273_),
    .C(_2282_),
    .A(_2270_),
    .Y(_2284_));
 sg13g2_nand3_1 _5828_ (.B(_2283_),
    .C(_2284_),
    .A(net1349),
    .Y(_2285_));
 sg13g2_o21ai_1 _5829_ (.B1(_2285_),
    .Y(_0490_),
    .A1(_0684_),
    .A2(net1361));
 sg13g2_nor2_1 _5830_ (.A(net1578),
    .B(net1361),
    .Y(_2286_));
 sg13g2_nor2_1 _5831_ (.A(net1253),
    .B(_0109_),
    .Y(_2287_));
 sg13g2_xor2_1 _5832_ (.B(_2278_),
    .A(\main.adder.s2_larger[32] ),
    .X(_2288_));
 sg13g2_a21oi_2 _5833_ (.B1(_2287_),
    .Y(_2289_),
    .A2(_2288_),
    .A1(net1253));
 sg13g2_nand2b_1 _5834_ (.Y(_2290_),
    .B(\main.adder.s2_smaler[32] ),
    .A_N(_2289_));
 sg13g2_xor2_1 _5835_ (.B(_2289_),
    .A(\main.adder.s2_smaler[32] ),
    .X(_2291_));
 sg13g2_a21o_1 _5836_ (.A2(_2283_),
    .A1(_2281_),
    .B1(_2291_),
    .X(_2292_));
 sg13g2_nand3_1 _5837_ (.B(_2283_),
    .C(_2291_),
    .A(_2281_),
    .Y(_2293_));
 sg13g2_nand2_1 _5838_ (.Y(_2294_),
    .A(_2292_),
    .B(_2293_));
 sg13g2_a21oi_1 _5839_ (.A1(net1361),
    .A2(_2294_),
    .Y(_0491_),
    .B1(_2286_));
 sg13g2_nor2_1 _5840_ (.A(net1253),
    .B(_0110_),
    .Y(_2295_));
 sg13g2_nor3_2 _5841_ (.A(\main.adder.s2_larger[32] ),
    .B(\main.adder.s2_larger[33] ),
    .C(_2278_),
    .Y(_2296_));
 sg13g2_o21ai_1 _5842_ (.B1(\main.adder.s2_larger[33] ),
    .Y(_2297_),
    .A1(\main.adder.s2_larger[32] ),
    .A2(_2278_));
 sg13g2_nor2b_1 _5843_ (.A(_2296_),
    .B_N(_2297_),
    .Y(_2298_));
 sg13g2_a21oi_2 _5844_ (.B1(_2295_),
    .Y(_2299_),
    .A2(_2298_),
    .A1(net1253));
 sg13g2_nand2b_1 _5845_ (.Y(_2300_),
    .B(_2299_),
    .A_N(\main.adder.s2_smaler[33] ));
 sg13g2_nand2b_1 _5846_ (.Y(_2301_),
    .B(\main.adder.s2_smaler[33] ),
    .A_N(_2299_));
 sg13g2_a22oi_1 _5847_ (.Y(_2302_),
    .B1(_2300_),
    .B2(_2301_),
    .A2(_2292_),
    .A1(_2290_));
 sg13g2_and4_1 _5848_ (.A(_2290_),
    .B(_2292_),
    .C(_2300_),
    .D(_2301_),
    .X(_2303_));
 sg13g2_o21ai_1 _5849_ (.B1(net1349),
    .Y(_2304_),
    .A1(_2302_),
    .A2(_2303_));
 sg13g2_o21ai_1 _5850_ (.B1(_2304_),
    .Y(_0492_),
    .A1(_0694_),
    .A2(net1361));
 sg13g2_nor2_1 _5851_ (.A(net1252),
    .B(_0111_),
    .Y(_2305_));
 sg13g2_nand2b_2 _5852_ (.Y(_2306_),
    .B(_2296_),
    .A_N(\main.adder.s2_larger[34] ));
 sg13g2_xnor2_1 _5853_ (.Y(_2307_),
    .A(\main.adder.s2_larger[34] ),
    .B(_2296_));
 sg13g2_a21oi_2 _5854_ (.B1(_2305_),
    .Y(_2308_),
    .A2(_2307_),
    .A1(net1252));
 sg13g2_nand2b_1 _5855_ (.Y(_2309_),
    .B(net1516),
    .A_N(_2308_));
 sg13g2_xnor2_1 _5856_ (.Y(_2310_),
    .A(\main.adder.s2_smaler[34] ),
    .B(_2308_));
 sg13g2_nand3_1 _5857_ (.B(_2292_),
    .C(_2301_),
    .A(_2290_),
    .Y(_2311_));
 sg13g2_nand3_1 _5858_ (.B(_2310_),
    .C(_2311_),
    .A(_2300_),
    .Y(_2312_));
 sg13g2_a21o_1 _5859_ (.A2(_2311_),
    .A1(_2300_),
    .B1(_2310_),
    .X(_2313_));
 sg13g2_nand3_1 _5860_ (.B(_2312_),
    .C(_2313_),
    .A(net1349),
    .Y(_2314_));
 sg13g2_o21ai_1 _5861_ (.B1(_2314_),
    .Y(_0493_),
    .A1(_0693_),
    .A2(net1361));
 sg13g2_nor2_1 _5862_ (.A(net1252),
    .B(_0112_),
    .Y(_2315_));
 sg13g2_xor2_1 _5863_ (.B(_2306_),
    .A(\main.adder.s2_larger[35] ),
    .X(_2316_));
 sg13g2_a21oi_2 _5864_ (.B1(_2315_),
    .Y(_2317_),
    .A2(_2316_),
    .A1(net1252));
 sg13g2_nand2b_1 _5865_ (.Y(_2318_),
    .B(net1041),
    .A_N(_2317_));
 sg13g2_xnor2_1 _5866_ (.Y(_2319_),
    .A(_0749_),
    .B(_2317_));
 sg13g2_a21o_1 _5867_ (.A2(_2312_),
    .A1(_2309_),
    .B1(_2319_),
    .X(_2320_));
 sg13g2_nand3_1 _5868_ (.B(_2312_),
    .C(_2319_),
    .A(_2309_),
    .Y(_2321_));
 sg13g2_a21oi_1 _5869_ (.A1(_2320_),
    .A2(_2321_),
    .Y(_2322_),
    .B1(net1308));
 sg13g2_a21oi_1 _5870_ (.A1(_0692_),
    .A2(net1310),
    .Y(_0494_),
    .B1(_2322_));
 sg13g2_nor2_1 _5871_ (.A(net1252),
    .B(_0113_),
    .Y(_2323_));
 sg13g2_nor3_2 _5872_ (.A(\main.adder.s2_larger[35] ),
    .B(\main.adder.s2_larger[36] ),
    .C(_2306_),
    .Y(_2324_));
 sg13g2_o21ai_1 _5873_ (.B1(\main.adder.s2_larger[36] ),
    .Y(_2325_),
    .A1(\main.adder.s2_larger[35] ),
    .A2(_2306_));
 sg13g2_nor2b_1 _5874_ (.A(_2324_),
    .B_N(_2325_),
    .Y(_2326_));
 sg13g2_a21oi_2 _5875_ (.B1(_2323_),
    .Y(_2327_),
    .A2(_2326_),
    .A1(net1252));
 sg13g2_nor2b_1 _5876_ (.A(_2327_),
    .B_N(\main.adder.s2_smaler[36] ),
    .Y(_2328_));
 sg13g2_xor2_1 _5877_ (.B(_2327_),
    .A(\main.adder.s2_smaler[36] ),
    .X(_2329_));
 sg13g2_a21o_1 _5878_ (.A2(_2320_),
    .A1(_2318_),
    .B1(_2329_),
    .X(_2330_));
 sg13g2_nand3_1 _5879_ (.B(_2320_),
    .C(_2329_),
    .A(_2318_),
    .Y(_2331_));
 sg13g2_a21oi_1 _5880_ (.A1(_2330_),
    .A2(_2331_),
    .Y(_2332_),
    .B1(net1308));
 sg13g2_a21oi_1 _5881_ (.A1(_0691_),
    .A2(net1310),
    .Y(_0495_),
    .B1(_2332_));
 sg13g2_nor2_1 _5882_ (.A(net1254),
    .B(_0114_),
    .Y(_2333_));
 sg13g2_nand2b_2 _5883_ (.Y(_2334_),
    .B(_2324_),
    .A_N(\main.adder.s2_larger[37] ));
 sg13g2_xnor2_1 _5884_ (.Y(_2335_),
    .A(\main.adder.s2_larger[37] ),
    .B(_2324_));
 sg13g2_a21oi_2 _5885_ (.B1(_2333_),
    .Y(_2336_),
    .A2(_2335_),
    .A1(net1254));
 sg13g2_nor2_1 _5886_ (.A(_0750_),
    .B(_2336_),
    .Y(_2337_));
 sg13g2_xnor2_1 _5887_ (.Y(_2338_),
    .A(\main.adder.s2_smaler[37] ),
    .B(_2336_));
 sg13g2_nor2b_1 _5888_ (.A(_2328_),
    .B_N(_2330_),
    .Y(_2339_));
 sg13g2_xnor2_1 _5889_ (.Y(_2340_),
    .A(_2338_),
    .B(_2339_));
 sg13g2_mux2_1 _5890_ (.A0(net1549),
    .A1(_2340_),
    .S(net1361),
    .X(_0496_));
 sg13g2_nor2_1 _5891_ (.A(net1255),
    .B(_0115_),
    .Y(_2341_));
 sg13g2_xor2_1 _5892_ (.B(_2334_),
    .A(\main.adder.s2_larger[38] ),
    .X(_2342_));
 sg13g2_a21oi_2 _5893_ (.B1(_2341_),
    .Y(_2343_),
    .A2(_2342_),
    .A1(net1255));
 sg13g2_nand2b_1 _5894_ (.Y(_2344_),
    .B(\main.adder.s2_smaler[38] ),
    .A_N(_2343_));
 sg13g2_inv_1 _5895_ (.Y(_2345_),
    .A(_2344_));
 sg13g2_xnor2_1 _5896_ (.Y(_2346_),
    .A(\main.adder.s2_smaler[38] ),
    .B(_2343_));
 sg13g2_nor2_1 _5897_ (.A(_2328_),
    .B(_2337_),
    .Y(_2347_));
 sg13g2_a22oi_1 _5898_ (.Y(_2348_),
    .B1(_2347_),
    .B2(_2330_),
    .A2(_2336_),
    .A1(_0750_));
 sg13g2_o21ai_1 _5899_ (.B1(net1347),
    .Y(_2349_),
    .A1(_2346_),
    .A2(_2348_));
 sg13g2_a21oi_1 _5900_ (.A1(_2346_),
    .A2(_2348_),
    .Y(_2350_),
    .B1(_2349_));
 sg13g2_a21o_1 _5901_ (.A2(net1308),
    .A1(net1519),
    .B1(_2350_),
    .X(_0497_));
 sg13g2_nor2_1 _5902_ (.A(net1255),
    .B(_0116_),
    .Y(_2351_));
 sg13g2_nor3_2 _5903_ (.A(\main.adder.s2_larger[38] ),
    .B(\main.adder.s2_larger[39] ),
    .C(_2334_),
    .Y(_2352_));
 sg13g2_o21ai_1 _5904_ (.B1(\main.adder.s2_larger[39] ),
    .Y(_2353_),
    .A1(\main.adder.s2_larger[38] ),
    .A2(_2334_));
 sg13g2_nor2b_1 _5905_ (.A(_2352_),
    .B_N(_2353_),
    .Y(_2354_));
 sg13g2_a21oi_2 _5906_ (.B1(_2351_),
    .Y(_2355_),
    .A2(_2354_),
    .A1(net1255));
 sg13g2_nand2b_1 _5907_ (.Y(_2356_),
    .B(\main.adder.s2_smaler[39] ),
    .A_N(_2355_));
 sg13g2_nor2b_1 _5908_ (.A(\main.adder.s2_smaler[39] ),
    .B_N(_2355_),
    .Y(_2357_));
 sg13g2_xnor2_1 _5909_ (.Y(_2358_),
    .A(\main.adder.s2_smaler[39] ),
    .B(_2355_));
 sg13g2_a21oi_1 _5910_ (.A1(_2346_),
    .A2(_2348_),
    .Y(_2359_),
    .B1(_2345_));
 sg13g2_xor2_1 _5911_ (.B(_2359_),
    .A(_2358_),
    .X(_2360_));
 sg13g2_nor2_1 _5912_ (.A(net1476),
    .B(net1349),
    .Y(_2361_));
 sg13g2_a21oi_1 _5913_ (.A1(net1349),
    .A2(_2360_),
    .Y(_0498_),
    .B1(_2361_));
 sg13g2_nand2b_2 _5914_ (.Y(_2362_),
    .B(_2352_),
    .A_N(\main.adder.s2_larger[40] ));
 sg13g2_nand2b_1 _5915_ (.Y(_2363_),
    .B(\main.adder.s2_larger[40] ),
    .A_N(_2352_));
 sg13g2_nand3_1 _5916_ (.B(_2362_),
    .C(_2363_),
    .A(net1257),
    .Y(_2364_));
 sg13g2_o21ai_1 _5917_ (.B1(_2364_),
    .Y(_2365_),
    .A1(net1257),
    .A2(_0117_));
 sg13g2_nand2_1 _5918_ (.Y(_2366_),
    .A(\main.adder.s2_smaler[40] ),
    .B(_2365_));
 sg13g2_xor2_1 _5919_ (.B(_2365_),
    .A(\main.adder.s2_smaler[40] ),
    .X(_2367_));
 sg13g2_o21ai_1 _5920_ (.B1(_2356_),
    .Y(_2368_),
    .A1(_2344_),
    .A2(_2357_));
 sg13g2_nand2_1 _5921_ (.Y(_2369_),
    .A(_2346_),
    .B(_2358_));
 sg13g2_a221oi_1 _5922_ (.B2(_2330_),
    .C1(_2369_),
    .B1(_2347_),
    .A1(_0750_),
    .Y(_2370_),
    .A2(_2336_));
 sg13g2_o21ai_1 _5923_ (.B1(_2367_),
    .Y(_2371_),
    .A1(_2368_),
    .A2(_2370_));
 sg13g2_or3_1 _5924_ (.A(_2367_),
    .B(_2368_),
    .C(_2370_),
    .X(_2372_));
 sg13g2_a21oi_1 _5925_ (.A1(_2371_),
    .A2(_2372_),
    .Y(_2373_),
    .B1(net1307));
 sg13g2_a21oi_1 _5926_ (.A1(_0690_),
    .A2(net1310),
    .Y(_0499_),
    .B1(_2373_));
 sg13g2_nor2_1 _5927_ (.A(net1257),
    .B(_0118_),
    .Y(_2374_));
 sg13g2_xor2_1 _5928_ (.B(_2362_),
    .A(\main.adder.s2_larger[41] ),
    .X(_2375_));
 sg13g2_a21oi_1 _5929_ (.A1(net1257),
    .A2(_2375_),
    .Y(_2376_),
    .B1(_2374_));
 sg13g2_nand2b_1 _5930_ (.Y(_2377_),
    .B(_2376_),
    .A_N(\main.adder.s2_smaler[41] ));
 sg13g2_nand2b_1 _5931_ (.Y(_2378_),
    .B(\main.adder.s2_smaler[41] ),
    .A_N(_2376_));
 sg13g2_and2_1 _5932_ (.A(_2377_),
    .B(_2378_),
    .X(_2379_));
 sg13g2_nand2_1 _5933_ (.Y(_2380_),
    .A(_2366_),
    .B(_2371_));
 sg13g2_o21ai_1 _5934_ (.B1(net1347),
    .Y(_2381_),
    .A1(_2379_),
    .A2(_2380_));
 sg13g2_a21oi_1 _5935_ (.A1(_2379_),
    .A2(_2380_),
    .Y(_2382_),
    .B1(_2381_));
 sg13g2_a21o_1 _5936_ (.A2(net1310),
    .A1(net1582),
    .B1(_2382_),
    .X(_0500_));
 sg13g2_nor2_1 _5937_ (.A(net1257),
    .B(_0119_),
    .Y(_2383_));
 sg13g2_nor3_2 _5938_ (.A(\main.adder.s2_larger[41] ),
    .B(\main.adder.s2_larger[42] ),
    .C(_2362_),
    .Y(_2384_));
 sg13g2_o21ai_1 _5939_ (.B1(\main.adder.s2_larger[42] ),
    .Y(_2385_),
    .A1(\main.adder.s2_larger[41] ),
    .A2(_2362_));
 sg13g2_nor2b_1 _5940_ (.A(_2384_),
    .B_N(_2385_),
    .Y(_2386_));
 sg13g2_a21oi_1 _5941_ (.A1(net1257),
    .A2(_2386_),
    .Y(_2387_),
    .B1(_2383_));
 sg13g2_nand2b_1 _5942_ (.Y(_2388_),
    .B(\main.adder.s2_smaler[42] ),
    .A_N(_2387_));
 sg13g2_xnor2_1 _5943_ (.Y(_2389_),
    .A(\main.adder.s2_smaler[42] ),
    .B(_2387_));
 sg13g2_nand2b_1 _5944_ (.Y(_2390_),
    .B(_2377_),
    .A_N(_2366_));
 sg13g2_and2_1 _5945_ (.A(_2367_),
    .B(_2379_),
    .X(_2391_));
 sg13g2_o21ai_1 _5946_ (.B1(_2391_),
    .Y(_2392_),
    .A1(_2368_),
    .A2(_2370_));
 sg13g2_nand3_1 _5947_ (.B(_2390_),
    .C(_2392_),
    .A(_2378_),
    .Y(_2393_));
 sg13g2_nand2_1 _5948_ (.Y(_2394_),
    .A(_2389_),
    .B(_2393_));
 sg13g2_o21ai_1 _5949_ (.B1(net1347),
    .Y(_2395_),
    .A1(_2389_),
    .A2(_2393_));
 sg13g2_nand2b_1 _5950_ (.Y(_2396_),
    .B(_2394_),
    .A_N(_2395_));
 sg13g2_o21ai_1 _5951_ (.B1(_2396_),
    .Y(_0501_),
    .A1(_0689_),
    .A2(net1361));
 sg13g2_nand2b_2 _5952_ (.Y(_2397_),
    .B(_2384_),
    .A_N(\main.adder.s2_larger[43] ));
 sg13g2_xor2_1 _5953_ (.B(_2384_),
    .A(\main.adder.s2_larger[43] ),
    .X(_2398_));
 sg13g2_nand2_1 _5954_ (.Y(_2399_),
    .A(net1257),
    .B(_2398_));
 sg13g2_nand2b_1 _5955_ (.Y(_2400_),
    .B(_0120_),
    .A_N(net1257));
 sg13g2_a21o_1 _5956_ (.A2(_2400_),
    .A1(_2399_),
    .B1(\main.adder.s2_smaler[43] ),
    .X(_2401_));
 sg13g2_inv_1 _5957_ (.Y(_2402_),
    .A(_2401_));
 sg13g2_nand3_1 _5958_ (.B(_2399_),
    .C(_2400_),
    .A(\main.adder.s2_smaler[43] ),
    .Y(_2403_));
 sg13g2_and2_1 _5959_ (.A(_2401_),
    .B(_2403_),
    .X(_2404_));
 sg13g2_nand2_1 _5960_ (.Y(_2405_),
    .A(_2388_),
    .B(_2394_));
 sg13g2_o21ai_1 _5961_ (.B1(net1347),
    .Y(_2406_),
    .A1(_2404_),
    .A2(_2405_));
 sg13g2_a21oi_1 _5962_ (.A1(_2404_),
    .A2(_2405_),
    .Y(_2407_),
    .B1(_2406_));
 sg13g2_a21o_1 _5963_ (.A2(net1310),
    .A1(net1560),
    .B1(_2407_),
    .X(_0502_));
 sg13g2_nor2_1 _5964_ (.A(net1259),
    .B(_0121_),
    .Y(_2408_));
 sg13g2_xor2_1 _5965_ (.B(_2397_),
    .A(\main.adder.s2_larger[44] ),
    .X(_2409_));
 sg13g2_a21oi_1 _5966_ (.A1(net1259),
    .A2(_2409_),
    .Y(_2410_),
    .B1(_2408_));
 sg13g2_nor2_1 _5967_ (.A(_0753_),
    .B(_2410_),
    .Y(_2411_));
 sg13g2_xnor2_1 _5968_ (.Y(_2412_),
    .A(\main.adder.s2_smaler[44] ),
    .B(_2410_));
 sg13g2_o21ai_1 _5969_ (.B1(_2403_),
    .Y(_2413_),
    .A1(_2388_),
    .A2(_2402_));
 sg13g2_and2_1 _5970_ (.A(_2389_),
    .B(_2404_),
    .X(_2414_));
 sg13g2_a21o_2 _5971_ (.A2(_2414_),
    .A1(_2393_),
    .B1(_2413_),
    .X(_2415_));
 sg13g2_xnor2_1 _5972_ (.Y(_2416_),
    .A(_2412_),
    .B(_2415_));
 sg13g2_nor2_1 _5973_ (.A(net1588),
    .B(net1352),
    .Y(_2417_));
 sg13g2_a21oi_1 _5974_ (.A1(net1352),
    .A2(_2416_),
    .Y(_0503_),
    .B1(_2417_));
 sg13g2_a21oi_1 _5975_ (.A1(_2412_),
    .A2(_2415_),
    .Y(_2418_),
    .B1(_2411_));
 sg13g2_or2_1 _5976_ (.X(_2419_),
    .B(_0122_),
    .A(net1258));
 sg13g2_nor3_2 _5977_ (.A(\main.adder.s2_larger[44] ),
    .B(\main.adder.s2_larger[45] ),
    .C(_2397_),
    .Y(_2420_));
 sg13g2_o21ai_1 _5978_ (.B1(\main.adder.s2_larger[45] ),
    .Y(_2421_),
    .A1(\main.adder.s2_larger[44] ),
    .A2(_2397_));
 sg13g2_nand2_1 _5979_ (.Y(_2422_),
    .A(net1258),
    .B(_2421_));
 sg13g2_o21ai_1 _5980_ (.B1(_2419_),
    .Y(_2423_),
    .A1(_2420_),
    .A2(_2422_));
 sg13g2_nor2_1 _5981_ (.A(\main.adder.s2_smaler[45] ),
    .B(_2423_),
    .Y(_2424_));
 sg13g2_xnor2_1 _5982_ (.Y(_2425_),
    .A(net1001),
    .B(_2423_));
 sg13g2_xnor2_1 _5983_ (.Y(_2426_),
    .A(_2418_),
    .B(_2425_));
 sg13g2_nand2_1 _5984_ (.Y(_2427_),
    .A(net1490),
    .B(net1309));
 sg13g2_o21ai_1 _5985_ (.B1(_2427_),
    .Y(_0504_),
    .A1(net1309),
    .A2(_2426_));
 sg13g2_nor2_1 _5986_ (.A(net1258),
    .B(_0123_),
    .Y(_2428_));
 sg13g2_xnor2_1 _5987_ (.Y(_2429_),
    .A(\main.adder.s2_larger[46] ),
    .B(_2420_));
 sg13g2_a21oi_1 _5988_ (.A1(net1258),
    .A2(_2429_),
    .Y(_2430_),
    .B1(_2428_));
 sg13g2_nor2_1 _5989_ (.A(_0756_),
    .B(_2430_),
    .Y(_2431_));
 sg13g2_xnor2_1 _5990_ (.Y(_2432_),
    .A(_0756_),
    .B(_2430_));
 sg13g2_a221oi_1 _5991_ (.B2(\main.adder.s2_smaler[45] ),
    .C1(_2411_),
    .B1(_2423_),
    .A1(_2412_),
    .Y(_2433_),
    .A2(_2415_));
 sg13g2_nor3_2 _5992_ (.A(_2424_),
    .B(_2432_),
    .C(_2433_),
    .Y(_2434_));
 sg13g2_o21ai_1 _5993_ (.B1(_2432_),
    .Y(_2435_),
    .A1(_2424_),
    .A2(_2433_));
 sg13g2_nand2_1 _5994_ (.Y(_2436_),
    .A(net1534),
    .B(net1309));
 sg13g2_nand2_1 _5995_ (.Y(_2437_),
    .A(net1353),
    .B(_2435_));
 sg13g2_o21ai_1 _5996_ (.B1(_2436_),
    .Y(_0505_),
    .A1(_2434_),
    .A2(_2437_));
 sg13g2_a21o_1 _5997_ (.A2(_2420_),
    .A1(_0755_),
    .B1(net1603),
    .X(_2438_));
 sg13g2_o21ai_1 _5998_ (.B1(_2438_),
    .Y(_2439_),
    .A1(_2431_),
    .A2(_2434_));
 sg13g2_nor3_1 _5999_ (.A(_2431_),
    .B(_2434_),
    .C(_2438_),
    .Y(_2440_));
 sg13g2_nor2_1 _6000_ (.A(net1309),
    .B(_2440_),
    .Y(_2441_));
 sg13g2_a22oi_1 _6001_ (.Y(_0506_),
    .B1(_2439_),
    .B2(_2441_),
    .A2(net1310),
    .A1(_0688_));
 sg13g2_a21oi_1 _6002_ (.A1(_0687_),
    .A2(net1310),
    .Y(_0507_),
    .B1(_2441_));
 sg13g2_and2_1 _6003_ (.A(net1340),
    .B(net584),
    .X(_0508_));
 sg13g2_nor2_1 _6004_ (.A(net1333),
    .B(net1258),
    .Y(_2442_));
 sg13g2_xnor2_1 _6005_ (.Y(_2443_),
    .A(net760),
    .B(net813));
 sg13g2_a21oi_1 _6006_ (.A1(net1333),
    .A2(_2443_),
    .Y(_0509_),
    .B1(_2442_));
 sg13g2_mux2_1 _6007_ (.A0(\main.adder.s2_nan ),
    .A1(net720),
    .S(net1345),
    .X(_0510_));
 sg13g2_mux2_1 _6008_ (.A0(net756),
    .A1(\main.adder.s1_inf ),
    .S(net1345),
    .X(_0511_));
 sg13g2_nand2_1 _6009_ (.Y(_2444_),
    .A(net1307),
    .B(net944));
 sg13g2_o21ai_1 _6010_ (.B1(_2444_),
    .Y(_0512_),
    .A1(_1854_),
    .A2(net1130));
 sg13g2_mux2_1 _6011_ (.A0(net726),
    .A1(net760),
    .S(net1333),
    .X(_0513_));
 sg13g2_mux2_1 _6012_ (.A0(net771),
    .A1(\main.adder.s1_larger[23] ),
    .S(net1383),
    .X(_0514_));
 sg13g2_mux2_1 _6013_ (.A0(net737),
    .A1(net742),
    .S(net1383),
    .X(_0515_));
 sg13g2_mux2_1 _6014_ (.A0(net765),
    .A1(\main.adder.s1_larger[25] ),
    .S(net1380),
    .X(_0516_));
 sg13g2_mux2_1 _6015_ (.A0(net601),
    .A1(net711),
    .S(net1383),
    .X(_0517_));
 sg13g2_mux2_1 _6016_ (.A0(net822),
    .A1(\main.adder.s1_larger[27] ),
    .S(net1380),
    .X(_0518_));
 sg13g2_mux2_1 _6017_ (.A0(net922),
    .A1(\main.adder.s1_larger[28] ),
    .S(net1379),
    .X(_0519_));
 sg13g2_mux2_1 _6018_ (.A0(net788),
    .A1(net844),
    .S(net1380),
    .X(_0520_));
 sg13g2_mux2_1 _6019_ (.A0(net819),
    .A1(\main.adder.s1_larger[30] ),
    .S(net1380),
    .X(_0521_));
 sg13g2_nand2_1 _6020_ (.Y(_2445_),
    .A(\main.spi.state[0] ),
    .B(\main.spi.SPI_not_chip_select_sampled ));
 sg13g2_o21ai_1 _6021_ (.B1(net1345),
    .Y(_2446_),
    .A1(\main.spi.state[0] ),
    .A2(\main.spi.SPI_not_chip_select_sampled ));
 sg13g2_a21oi_1 _6022_ (.A1(net577),
    .A2(_2445_),
    .Y(_0522_),
    .B1(_2446_));
 sg13g2_mux4_1 _6023_ (.S0(net1232),
    .A0(\main.float_registers[0][15] ),
    .A1(\main.float_registers[1][15] ),
    .A2(\main.float_registers[2][15] ),
    .A3(\main.float_registers[3][15] ),
    .S1(net1227),
    .X(_2447_));
 sg13g2_mux4_1 _6024_ (.S0(net1233),
    .A0(\main.float_registers[0][0] ),
    .A1(\main.float_registers[1][0] ),
    .A2(\main.float_registers[2][0] ),
    .A3(\main.float_registers[3][0] ),
    .S1(net1228),
    .X(_2448_));
 sg13g2_mux4_1 _6025_ (.S0(net1232),
    .A0(\main.float_registers[0][11] ),
    .A1(\main.float_registers[1][11] ),
    .A2(\main.float_registers[2][11] ),
    .A3(\main.float_registers[3][11] ),
    .S1(net1227),
    .X(_2449_));
 sg13g2_mux4_1 _6026_ (.S0(net1231),
    .A0(\main.float_registers[0][17] ),
    .A1(\main.float_registers[1][17] ),
    .A2(\main.float_registers[2][17] ),
    .A3(\main.float_registers[3][17] ),
    .S1(net1226),
    .X(_2450_));
 sg13g2_mux4_1 _6027_ (.S0(net1233),
    .A0(\main.float_registers[0][19] ),
    .A1(\main.float_registers[1][19] ),
    .A2(\main.float_registers[2][19] ),
    .A3(\main.float_registers[3][19] ),
    .S1(net1228),
    .X(_2451_));
 sg13g2_mux4_1 _6028_ (.S0(net1235),
    .A0(\main.float_registers[0][3] ),
    .A1(\main.float_registers[1][3] ),
    .A2(\main.float_registers[2][3] ),
    .A3(\main.float_registers[3][3] ),
    .S1(net1230),
    .X(_2452_));
 sg13g2_mux4_1 _6029_ (.S0(net1235),
    .A0(\main.float_registers[0][6] ),
    .A1(\main.float_registers[1][6] ),
    .A2(\main.float_registers[2][6] ),
    .A3(\main.float_registers[3][6] ),
    .S1(net1230),
    .X(_2453_));
 sg13g2_mux4_1 _6030_ (.S0(net1232),
    .A0(\main.float_registers[0][13] ),
    .A1(\main.float_registers[1][13] ),
    .A2(\main.float_registers[2][13] ),
    .A3(\main.float_registers[3][13] ),
    .S1(net1227),
    .X(_2454_));
 sg13g2_mux4_1 _6031_ (.S0(net1232),
    .A0(\main.float_registers[0][8] ),
    .A1(\main.float_registers[1][8] ),
    .A2(\main.float_registers[2][8] ),
    .A3(\main.float_registers[3][8] ),
    .S1(net1227),
    .X(_2455_));
 sg13g2_mux4_1 _6032_ (.S0(net1231),
    .A0(\main.float_registers[0][20] ),
    .A1(\main.float_registers[1][20] ),
    .A2(\main.float_registers[2][20] ),
    .A3(\main.float_registers[3][20] ),
    .S1(net1226),
    .X(_2456_));
 sg13g2_mux4_1 _6033_ (.S0(net1233),
    .A0(\main.float_registers[0][4] ),
    .A1(\main.float_registers[1][4] ),
    .A2(\main.float_registers[2][4] ),
    .A3(\main.float_registers[3][4] ),
    .S1(net1228),
    .X(_2457_));
 sg13g2_mux4_1 _6034_ (.S0(net1231),
    .A0(\main.float_registers[0][22] ),
    .A1(\main.float_registers[1][22] ),
    .A2(\main.float_registers[2][22] ),
    .A3(\main.float_registers[3][22] ),
    .S1(net1226),
    .X(_2458_));
 sg13g2_mux4_1 _6035_ (.S0(net1232),
    .A0(\main.float_registers[0][9] ),
    .A1(\main.float_registers[1][9] ),
    .A2(\main.float_registers[2][9] ),
    .A3(\main.float_registers[3][9] ),
    .S1(net1227),
    .X(_2459_));
 sg13g2_mux4_1 _6036_ (.S0(net1231),
    .A0(\main.float_registers[0][18] ),
    .A1(\main.float_registers[1][18] ),
    .A2(\main.float_registers[2][18] ),
    .A3(\main.float_registers[3][18] ),
    .S1(net1226),
    .X(_2460_));
 sg13g2_mux4_1 _6037_ (.S0(net1231),
    .A0(\main.float_registers[0][1] ),
    .A1(\main.float_registers[1][1] ),
    .A2(\main.float_registers[2][1] ),
    .A3(\main.float_registers[3][1] ),
    .S1(net1226),
    .X(_2461_));
 sg13g2_mux4_1 _6038_ (.S0(net1235),
    .A0(\main.float_registers[0][2] ),
    .A1(\main.float_registers[1][2] ),
    .A2(\main.float_registers[2][2] ),
    .A3(\main.float_registers[3][2] ),
    .S1(net1230),
    .X(_2462_));
 sg13g2_mux4_1 _6039_ (.S0(net1231),
    .A0(\main.float_registers[0][21] ),
    .A1(\main.float_registers[1][21] ),
    .A2(\main.float_registers[2][21] ),
    .A3(\main.float_registers[3][21] ),
    .S1(net1226),
    .X(_2463_));
 sg13g2_mux4_1 _6040_ (.S0(net1231),
    .A0(\main.float_registers[0][16] ),
    .A1(\main.float_registers[1][16] ),
    .A2(\main.float_registers[2][16] ),
    .A3(\main.float_registers[3][16] ),
    .S1(net1226),
    .X(_2464_));
 sg13g2_mux4_1 _6041_ (.S0(net1232),
    .A0(\main.float_registers[0][12] ),
    .A1(\main.float_registers[1][12] ),
    .A2(\main.float_registers[2][12] ),
    .A3(\main.float_registers[3][12] ),
    .S1(net1227),
    .X(_2465_));
 sg13g2_mux4_1 _6042_ (.S0(net1235),
    .A0(\main.float_registers[0][5] ),
    .A1(\main.float_registers[1][5] ),
    .A2(\main.float_registers[2][5] ),
    .A3(\main.float_registers[3][5] ),
    .S1(net1230),
    .X(_2466_));
 sg13g2_mux4_1 _6043_ (.S0(net1231),
    .A0(\main.float_registers[0][14] ),
    .A1(\main.float_registers[1][14] ),
    .A2(\main.float_registers[2][14] ),
    .A3(\main.float_registers[3][14] ),
    .S1(net1226),
    .X(_2467_));
 sg13g2_mux4_1 _6044_ (.S0(net1234),
    .A0(\main.float_registers[0][7] ),
    .A1(\main.float_registers[1][7] ),
    .A2(\main.float_registers[2][7] ),
    .A3(\main.float_registers[3][7] ),
    .S1(net1229),
    .X(_2468_));
 sg13g2_mux4_1 _6045_ (.S0(net1232),
    .A0(\main.float_registers[0][10] ),
    .A1(\main.float_registers[1][10] ),
    .A2(\main.float_registers[2][10] ),
    .A3(\main.float_registers[3][10] ),
    .S1(net1227),
    .X(_2469_));
 sg13g2_nor4_1 _6046_ (.A(_2448_),
    .B(_2453_),
    .C(_2454_),
    .D(_2459_),
    .Y(_2470_));
 sg13g2_nor4_1 _6047_ (.A(_2447_),
    .B(_2464_),
    .C(_2466_),
    .D(_2467_),
    .Y(_2471_));
 sg13g2_nor4_2 _6048_ (.A(_2451_),
    .B(_2452_),
    .C(_2462_),
    .Y(_2472_),
    .D(_2468_));
 sg13g2_nor4_1 _6049_ (.A(_2450_),
    .B(_2455_),
    .C(_2457_),
    .D(_2465_),
    .Y(_2473_));
 sg13g2_nand2_1 _6050_ (.Y(_2474_),
    .A(_2472_),
    .B(_2473_));
 sg13g2_nor4_1 _6051_ (.A(_2449_),
    .B(_2460_),
    .C(_2461_),
    .D(_2474_),
    .Y(_2475_));
 sg13g2_nor4_1 _6052_ (.A(_2456_),
    .B(_2458_),
    .C(_2463_),
    .D(_2469_),
    .Y(_2476_));
 sg13g2_and4_2 _6053_ (.A(_2470_),
    .B(_2471_),
    .C(_2475_),
    .D(_2476_),
    .X(_2477_));
 sg13g2_mux4_1 _6054_ (.S0(net1234),
    .A0(\main.float_registers[0][25] ),
    .A1(\main.float_registers[1][25] ),
    .A2(\main.float_registers[2][25] ),
    .A3(\main.float_registers[3][25] ),
    .S1(net1229),
    .X(_2478_));
 sg13g2_mux4_1 _6055_ (.S0(net1234),
    .A0(\main.float_registers[0][29] ),
    .A1(\main.float_registers[1][29] ),
    .A2(\main.float_registers[2][29] ),
    .A3(\main.float_registers[3][29] ),
    .S1(net1229),
    .X(_2479_));
 sg13g2_mux4_1 _6056_ (.S0(net1235),
    .A0(\main.float_registers[0][27] ),
    .A1(\main.float_registers[1][27] ),
    .A2(\main.float_registers[2][27] ),
    .A3(\main.float_registers[3][27] ),
    .S1(net1230),
    .X(_2480_));
 sg13g2_mux4_1 _6057_ (.S0(net1234),
    .A0(\main.float_registers[0][30] ),
    .A1(\main.float_registers[1][30] ),
    .A2(\main.float_registers[2][30] ),
    .A3(\main.float_registers[3][30] ),
    .S1(net1229),
    .X(_2481_));
 sg13g2_mux4_1 _6058_ (.S0(net1234),
    .A0(\main.float_registers[0][28] ),
    .A1(\main.float_registers[1][28] ),
    .A2(\main.float_registers[2][28] ),
    .A3(\main.float_registers[3][28] ),
    .S1(net1229),
    .X(_2482_));
 sg13g2_mux4_1 _6059_ (.S0(net1234),
    .A0(\main.float_registers[0][24] ),
    .A1(\main.float_registers[1][24] ),
    .A2(\main.float_registers[2][24] ),
    .A3(\main.float_registers[3][24] ),
    .S1(net1229),
    .X(_2483_));
 sg13g2_inv_1 _6060_ (.Y(_2484_),
    .A(_2483_));
 sg13g2_mux4_1 _6061_ (.S0(net1232),
    .A0(\main.float_registers[0][23] ),
    .A1(\main.float_registers[1][23] ),
    .A2(\main.float_registers[2][23] ),
    .A3(\main.float_registers[3][23] ),
    .S1(net1227),
    .X(_2485_));
 sg13g2_mux4_1 _6062_ (.S0(net1234),
    .A0(\main.float_registers[0][26] ),
    .A1(\main.float_registers[1][26] ),
    .A2(\main.float_registers[2][26] ),
    .A3(\main.float_registers[3][26] ),
    .S1(net1229),
    .X(_2486_));
 sg13g2_mux4_1 _6063_ (.S0(net1244),
    .A0(\main.float_registers[0][28] ),
    .A1(\main.float_registers[1][28] ),
    .A2(\main.float_registers[2][28] ),
    .A3(\main.float_registers[3][28] ),
    .S1(net1239),
    .X(_2487_));
 sg13g2_mux4_1 _6064_ (.S0(net1244),
    .A0(\main.float_registers[0][26] ),
    .A1(\main.float_registers[1][26] ),
    .A2(\main.float_registers[2][26] ),
    .A3(\main.float_registers[3][26] ),
    .S1(net1239),
    .X(_2488_));
 sg13g2_mux4_1 _6065_ (.S0(net1244),
    .A0(\main.float_registers[0][24] ),
    .A1(\main.float_registers[1][24] ),
    .A2(\main.float_registers[2][24] ),
    .A3(\main.float_registers[3][24] ),
    .S1(net1239),
    .X(_2489_));
 sg13g2_mux4_1 _6066_ (.S0(net1245),
    .A0(\main.float_registers[0][30] ),
    .A1(\main.float_registers[1][30] ),
    .A2(\main.float_registers[2][30] ),
    .A3(\main.float_registers[3][30] ),
    .S1(net1240),
    .X(_2490_));
 sg13g2_mux4_1 _6067_ (.S0(net1244),
    .A0(\main.float_registers[0][29] ),
    .A1(\main.float_registers[1][29] ),
    .A2(\main.float_registers[2][29] ),
    .A3(\main.float_registers[3][29] ),
    .S1(net1239),
    .X(_2491_));
 sg13g2_mux4_1 _6068_ (.S0(net1244),
    .A0(\main.float_registers[0][27] ),
    .A1(\main.float_registers[1][27] ),
    .A2(\main.float_registers[2][27] ),
    .A3(\main.float_registers[3][27] ),
    .S1(net1239),
    .X(_2492_));
 sg13g2_mux4_1 _6069_ (.S0(net1243),
    .A0(\main.float_registers[0][23] ),
    .A1(\main.float_registers[1][23] ),
    .A2(\main.float_registers[2][23] ),
    .A3(\main.float_registers[3][23] ),
    .S1(net1238),
    .X(_2493_));
 sg13g2_mux4_1 _6070_ (.S0(net1244),
    .A0(\main.float_registers[0][25] ),
    .A1(\main.float_registers[1][25] ),
    .A2(\main.float_registers[2][25] ),
    .A3(\main.float_registers[3][25] ),
    .S1(net1239),
    .X(_2494_));
 sg13g2_nand4_1 _6071_ (.B(_2488_),
    .C(_2493_),
    .A(_2487_),
    .Y(_2495_),
    .D(_2494_));
 sg13g2_nand4_1 _6072_ (.B(_2490_),
    .C(_2491_),
    .A(_2489_),
    .Y(_2496_),
    .D(_2492_));
 sg13g2_nor2_1 _6073_ (.A(_2495_),
    .B(_2496_),
    .Y(_2497_));
 sg13g2_mux4_1 _6074_ (.S0(net1242),
    .A0(\main.float_registers[0][19] ),
    .A1(\main.float_registers[1][19] ),
    .A2(\main.float_registers[2][19] ),
    .A3(\main.float_registers[3][19] ),
    .S1(net1237),
    .X(_2498_));
 sg13g2_mux4_1 _6075_ (.S0(_0002_),
    .A0(\main.float_registers[0][13] ),
    .A1(\main.float_registers[1][13] ),
    .A2(\main.float_registers[2][13] ),
    .A3(\main.float_registers[3][13] ),
    .S1(_0003_),
    .X(_2499_));
 sg13g2_mux4_1 _6076_ (.S0(net1241),
    .A0(\main.float_registers[0][22] ),
    .A1(\main.float_registers[1][22] ),
    .A2(\main.float_registers[2][22] ),
    .A3(\main.float_registers[3][22] ),
    .S1(net1236),
    .X(_2500_));
 sg13g2_mux4_1 _6077_ (.S0(net1245),
    .A0(\main.float_registers[0][2] ),
    .A1(\main.float_registers[1][2] ),
    .A2(\main.float_registers[2][2] ),
    .A3(\main.float_registers[3][2] ),
    .S1(net1240),
    .X(_2501_));
 sg13g2_mux4_1 _6078_ (.S0(net1241),
    .A0(\main.float_registers[0][0] ),
    .A1(\main.float_registers[1][0] ),
    .A2(\main.float_registers[2][0] ),
    .A3(\main.float_registers[3][0] ),
    .S1(net1236),
    .X(_2502_));
 sg13g2_mux4_1 _6079_ (.S0(net1242),
    .A0(\main.float_registers[0][4] ),
    .A1(\main.float_registers[1][4] ),
    .A2(\main.float_registers[2][4] ),
    .A3(\main.float_registers[3][4] ),
    .S1(net1237),
    .X(_2503_));
 sg13g2_mux4_1 _6080_ (.S0(net1242),
    .A0(\main.float_registers[0][14] ),
    .A1(\main.float_registers[1][14] ),
    .A2(\main.float_registers[2][14] ),
    .A3(\main.float_registers[3][14] ),
    .S1(net1237),
    .X(_2504_));
 sg13g2_mux4_1 _6081_ (.S0(net1241),
    .A0(\main.float_registers[0][8] ),
    .A1(\main.float_registers[1][8] ),
    .A2(\main.float_registers[2][8] ),
    .A3(\main.float_registers[3][8] ),
    .S1(net1236),
    .X(_2505_));
 sg13g2_mux4_1 _6082_ (.S0(net1241),
    .A0(\main.float_registers[0][16] ),
    .A1(\main.float_registers[1][16] ),
    .A2(\main.float_registers[2][16] ),
    .A3(\main.float_registers[3][16] ),
    .S1(net1236),
    .X(_2506_));
 sg13g2_mux4_1 _6083_ (.S0(net1241),
    .A0(\main.float_registers[0][18] ),
    .A1(\main.float_registers[1][18] ),
    .A2(\main.float_registers[2][18] ),
    .A3(\main.float_registers[3][18] ),
    .S1(net1236),
    .X(_2507_));
 sg13g2_mux4_1 _6084_ (.S0(net1242),
    .A0(\main.float_registers[0][1] ),
    .A1(\main.float_registers[1][1] ),
    .A2(\main.float_registers[2][1] ),
    .A3(\main.float_registers[3][1] ),
    .S1(net1237),
    .X(_2508_));
 sg13g2_mux4_1 _6085_ (.S0(net1241),
    .A0(\main.float_registers[0][17] ),
    .A1(\main.float_registers[1][17] ),
    .A2(\main.float_registers[2][17] ),
    .A3(\main.float_registers[3][17] ),
    .S1(net1236),
    .X(_2509_));
 sg13g2_mux4_1 _6086_ (.S0(net1243),
    .A0(\main.float_registers[0][10] ),
    .A1(\main.float_registers[1][10] ),
    .A2(\main.float_registers[2][10] ),
    .A3(\main.float_registers[3][10] ),
    .S1(net1238),
    .X(_2510_));
 sg13g2_mux4_1 _6087_ (.S0(net1245),
    .A0(\main.float_registers[0][3] ),
    .A1(\main.float_registers[1][3] ),
    .A2(\main.float_registers[2][3] ),
    .A3(\main.float_registers[3][3] ),
    .S1(net1240),
    .X(_2511_));
 sg13g2_mux4_1 _6088_ (.S0(net1241),
    .A0(\main.float_registers[0][21] ),
    .A1(\main.float_registers[1][21] ),
    .A2(\main.float_registers[2][21] ),
    .A3(\main.float_registers[3][21] ),
    .S1(net1236),
    .X(_2512_));
 sg13g2_mux4_1 _6089_ (.S0(net1243),
    .A0(\main.float_registers[0][11] ),
    .A1(\main.float_registers[1][11] ),
    .A2(\main.float_registers[2][11] ),
    .A3(\main.float_registers[3][11] ),
    .S1(net1238),
    .X(_2513_));
 sg13g2_mux4_1 _6090_ (.S0(net1243),
    .A0(\main.float_registers[0][15] ),
    .A1(\main.float_registers[1][15] ),
    .A2(\main.float_registers[2][15] ),
    .A3(\main.float_registers[3][15] ),
    .S1(net1238),
    .X(_2514_));
 sg13g2_mux4_1 _6091_ (.S0(net1245),
    .A0(\main.float_registers[0][6] ),
    .A1(\main.float_registers[1][6] ),
    .A2(\main.float_registers[2][6] ),
    .A3(\main.float_registers[3][6] ),
    .S1(net1240),
    .X(_2515_));
 sg13g2_mux4_1 _6092_ (.S0(net1243),
    .A0(\main.float_registers[0][9] ),
    .A1(\main.float_registers[1][9] ),
    .A2(\main.float_registers[2][9] ),
    .A3(\main.float_registers[3][9] ),
    .S1(net1238),
    .X(_2516_));
 sg13g2_mux4_1 _6093_ (.S0(net1245),
    .A0(\main.float_registers[0][5] ),
    .A1(\main.float_registers[1][5] ),
    .A2(\main.float_registers[2][5] ),
    .A3(\main.float_registers[3][5] ),
    .S1(net1240),
    .X(_2517_));
 sg13g2_mux4_1 _6094_ (.S0(net1241),
    .A0(\main.float_registers[0][20] ),
    .A1(\main.float_registers[1][20] ),
    .A2(\main.float_registers[2][20] ),
    .A3(\main.float_registers[3][20] ),
    .S1(net1236),
    .X(_2518_));
 sg13g2_mux4_1 _6095_ (.S0(net1243),
    .A0(\main.float_registers[0][12] ),
    .A1(\main.float_registers[1][12] ),
    .A2(\main.float_registers[2][12] ),
    .A3(\main.float_registers[3][12] ),
    .S1(net1238),
    .X(_2519_));
 sg13g2_mux4_1 _6096_ (.S0(net1244),
    .A0(\main.float_registers[0][7] ),
    .A1(\main.float_registers[1][7] ),
    .A2(\main.float_registers[2][7] ),
    .A3(\main.float_registers[3][7] ),
    .S1(net1239),
    .X(_2520_));
 sg13g2_nor4_1 _6097_ (.A(_2500_),
    .B(_2501_),
    .C(_2511_),
    .D(_2512_),
    .Y(_2521_));
 sg13g2_nor4_1 _6098_ (.A(_2510_),
    .B(_2515_),
    .C(_2519_),
    .D(_2520_),
    .Y(_2522_));
 sg13g2_nor4_1 _6099_ (.A(_2503_),
    .B(_2513_),
    .C(_2514_),
    .D(_2516_),
    .Y(_2523_));
 sg13g2_nor4_1 _6100_ (.A(_2498_),
    .B(_2499_),
    .C(_2504_),
    .D(_2507_),
    .Y(_2524_));
 sg13g2_nand2_1 _6101_ (.Y(_2525_),
    .A(_2523_),
    .B(_2524_));
 sg13g2_nor4_1 _6102_ (.A(_2502_),
    .B(_2506_),
    .C(_2508_),
    .D(_2525_),
    .Y(_2526_));
 sg13g2_nor4_1 _6103_ (.A(_2505_),
    .B(_2509_),
    .C(_2517_),
    .D(_2518_),
    .Y(_2527_));
 sg13g2_and4_2 _6104_ (.A(_2521_),
    .B(_2522_),
    .C(_2526_),
    .D(_2527_),
    .X(_2528_));
 sg13g2_nand2b_1 _6105_ (.Y(_2529_),
    .B(_2497_),
    .A_N(_2528_));
 sg13g2_nand4_1 _6106_ (.B(_2479_),
    .C(_2480_),
    .A(_2478_),
    .Y(_2530_),
    .D(_2485_));
 sg13g2_nand4_1 _6107_ (.B(_2482_),
    .C(_2483_),
    .A(_2481_),
    .Y(_2531_),
    .D(_2486_));
 sg13g2_nor2_1 _6108_ (.A(_2530_),
    .B(_2531_),
    .Y(_2532_));
 sg13g2_nand2b_1 _6109_ (.Y(_2533_),
    .B(_2532_),
    .A_N(_2477_));
 sg13g2_mux4_1 _6110_ (.S0(net1244),
    .A0(\main.float_registers[0][31] ),
    .A1(\main.float_registers[1][31] ),
    .A2(\main.float_registers[2][31] ),
    .A3(\main.float_registers[3][31] ),
    .S1(net1239),
    .X(_2534_));
 sg13g2_mux4_1 _6111_ (.S0(net1234),
    .A0(\main.float_registers[0][31] ),
    .A1(\main.float_registers[1][31] ),
    .A2(\main.float_registers[2][31] ),
    .A3(\main.float_registers[3][31] ),
    .S1(net1229),
    .X(_2535_));
 sg13g2_xnor2_1 _6112_ (.Y(_2536_),
    .A(_2534_),
    .B(_2535_));
 sg13g2_and2_1 _6113_ (.A(_2497_),
    .B(_2528_),
    .X(_2537_));
 sg13g2_nand3_1 _6114_ (.B(_2532_),
    .C(_2537_),
    .A(_2477_),
    .Y(_2538_));
 sg13g2_or2_1 _6115_ (.X(_2539_),
    .B(_2538_),
    .A(_2536_));
 sg13g2_nand4_1 _6116_ (.B(_2529_),
    .C(_2533_),
    .A(net1342),
    .Y(_2540_),
    .D(_2539_));
 sg13g2_o21ai_1 _6117_ (.B1(_2540_),
    .Y(_2541_),
    .A1(net1345),
    .A2(net720));
 sg13g2_inv_1 _6118_ (.Y(_0524_),
    .A(_2541_));
 sg13g2_nand2_1 _6119_ (.Y(_2542_),
    .A(net1304),
    .B(net1505));
 sg13g2_a21o_1 _6120_ (.A2(_2532_),
    .A1(_2477_),
    .B1(_2537_),
    .X(_2543_));
 sg13g2_a22oi_1 _6121_ (.Y(_2544_),
    .B1(_2538_),
    .B2(_2543_),
    .A2(_2535_),
    .A1(_2534_));
 sg13g2_a21o_1 _6122_ (.A2(_2538_),
    .A1(_2536_),
    .B1(net1304),
    .X(_2545_));
 sg13g2_o21ai_1 _6123_ (.B1(_2542_),
    .Y(_0525_),
    .A1(_2544_),
    .A2(_2545_));
 sg13g2_nand2b_1 _6124_ (.Y(_2546_),
    .B(_2491_),
    .A_N(_2479_));
 sg13g2_xnor2_1 _6125_ (.Y(_2547_),
    .A(_2479_),
    .B(_2491_));
 sg13g2_nor2b_1 _6126_ (.A(_2482_),
    .B_N(_2487_),
    .Y(_2548_));
 sg13g2_nand2b_1 _6127_ (.Y(_2549_),
    .B(_2482_),
    .A_N(_2487_));
 sg13g2_nand2b_1 _6128_ (.Y(_2550_),
    .B(_2492_),
    .A_N(_2480_));
 sg13g2_xor2_1 _6129_ (.B(_2492_),
    .A(_2480_),
    .X(_2551_));
 sg13g2_nor2b_1 _6130_ (.A(_2486_),
    .B_N(_2488_),
    .Y(_2552_));
 sg13g2_nand2b_1 _6131_ (.Y(_2553_),
    .B(_2486_),
    .A_N(_2488_));
 sg13g2_nand2b_1 _6132_ (.Y(_2554_),
    .B(_2494_),
    .A_N(_2478_));
 sg13g2_xnor2_1 _6133_ (.Y(_2555_),
    .A(_2478_),
    .B(_2494_));
 sg13g2_inv_1 _6134_ (.Y(_2556_),
    .A(_2555_));
 sg13g2_xnor2_1 _6135_ (.Y(_2557_),
    .A(_2483_),
    .B(_2489_));
 sg13g2_nor3_1 _6136_ (.A(_2488_),
    .B(_2489_),
    .C(_2491_),
    .Y(_2558_));
 sg13g2_nor4_1 _6137_ (.A(_2487_),
    .B(_2490_),
    .C(_2492_),
    .D(_2494_),
    .Y(_2559_));
 sg13g2_a21oi_1 _6138_ (.A1(_2558_),
    .A2(_2559_),
    .Y(_2560_),
    .B1(_2493_));
 sg13g2_nor3_1 _6139_ (.A(_2479_),
    .B(_2483_),
    .C(_2486_),
    .Y(_2561_));
 sg13g2_nor4_1 _6140_ (.A(_2478_),
    .B(_2480_),
    .C(_2481_),
    .D(_2482_),
    .Y(_2562_));
 sg13g2_a21oi_1 _6141_ (.A1(_2561_),
    .A2(_2562_),
    .Y(_2563_),
    .B1(_2485_));
 sg13g2_nor2b_1 _6142_ (.A(_2563_),
    .B_N(_2560_),
    .Y(_2564_));
 sg13g2_nor2b_1 _6143_ (.A(_2564_),
    .B_N(_2557_),
    .Y(_2565_));
 sg13g2_a21oi_1 _6144_ (.A1(_2484_),
    .A2(_2489_),
    .Y(_2566_),
    .B1(_2565_));
 sg13g2_o21ai_1 _6145_ (.B1(_2554_),
    .Y(_2567_),
    .A1(_2556_),
    .A2(_2566_));
 sg13g2_o21ai_1 _6146_ (.B1(_2553_),
    .Y(_2568_),
    .A1(_2552_),
    .A2(_2567_));
 sg13g2_o21ai_1 _6147_ (.B1(_2550_),
    .Y(_2569_),
    .A1(_2551_),
    .A2(_2568_));
 sg13g2_o21ai_1 _6148_ (.B1(_2549_),
    .Y(_2570_),
    .A1(_2548_),
    .A2(_2569_));
 sg13g2_nand2b_1 _6149_ (.Y(_2571_),
    .B(_2547_),
    .A_N(_2570_));
 sg13g2_nand2_1 _6150_ (.Y(_2572_),
    .A(_2546_),
    .B(_2571_));
 sg13g2_nor2_1 _6151_ (.A(_2481_),
    .B(_2490_),
    .Y(_2573_));
 sg13g2_and2_1 _6152_ (.A(_2481_),
    .B(_2490_),
    .X(_2574_));
 sg13g2_nor2_1 _6153_ (.A(_2573_),
    .B(_2574_),
    .Y(_2575_));
 sg13g2_a21oi_1 _6154_ (.A1(_2546_),
    .A2(_2571_),
    .Y(_2576_),
    .B1(_2575_));
 sg13g2_nor2b_1 _6155_ (.A(_2481_),
    .B_N(_2490_),
    .Y(_2577_));
 sg13g2_nor2_1 _6156_ (.A(_2576_),
    .B(_2577_),
    .Y(_2578_));
 sg13g2_mux2_1 _6157_ (.A0(_2448_),
    .A1(_2502_),
    .S(net1063),
    .X(_2579_));
 sg13g2_mux2_1 _6158_ (.A0(net1048),
    .A1(_2579_),
    .S(net1335),
    .X(_0526_));
 sg13g2_mux2_1 _6159_ (.A0(_2461_),
    .A1(_2508_),
    .S(net1061),
    .X(_2580_));
 sg13g2_mux2_1 _6160_ (.A0(net685),
    .A1(_2580_),
    .S(net1336),
    .X(_0527_));
 sg13g2_mux2_1 _6161_ (.A0(_2462_),
    .A1(_2501_),
    .S(net1064),
    .X(_2581_));
 sg13g2_mux2_1 _6162_ (.A0(net641),
    .A1(_2581_),
    .S(net1336),
    .X(_0528_));
 sg13g2_mux2_1 _6163_ (.A0(_2452_),
    .A1(_2511_),
    .S(net1064),
    .X(_2582_));
 sg13g2_mux2_1 _6164_ (.A0(net647),
    .A1(_2582_),
    .S(net1336),
    .X(_0529_));
 sg13g2_mux2_1 _6165_ (.A0(_2457_),
    .A1(_2503_),
    .S(net1061),
    .X(_2583_));
 sg13g2_mux2_1 _6166_ (.A0(net644),
    .A1(_2583_),
    .S(net1328),
    .X(_0530_));
 sg13g2_mux2_1 _6167_ (.A0(_2466_),
    .A1(_2517_),
    .S(net1062),
    .X(_2584_));
 sg13g2_mux2_1 _6168_ (.A0(net664),
    .A1(_2584_),
    .S(net1336),
    .X(_0531_));
 sg13g2_mux2_1 _6169_ (.A0(_2453_),
    .A1(_2515_),
    .S(net1062),
    .X(_2585_));
 sg13g2_mux2_1 _6170_ (.A0(net655),
    .A1(_2585_),
    .S(net1336),
    .X(_0532_));
 sg13g2_mux2_1 _6171_ (.A0(_2468_),
    .A1(_2520_),
    .S(net1062),
    .X(_2586_));
 sg13g2_mux2_1 _6172_ (.A0(net650),
    .A1(_2586_),
    .S(net1336),
    .X(_0533_));
 sg13g2_mux2_1 _6173_ (.A0(_2455_),
    .A1(_2505_),
    .S(net1058),
    .X(_2587_));
 sg13g2_mux2_1 _6174_ (.A0(net651),
    .A1(_2587_),
    .S(net1328),
    .X(_0534_));
 sg13g2_mux2_1 _6175_ (.A0(_2459_),
    .A1(_2516_),
    .S(net1058),
    .X(_2588_));
 sg13g2_mux2_1 _6176_ (.A0(net645),
    .A1(_2588_),
    .S(net1323),
    .X(_0535_));
 sg13g2_mux2_1 _6177_ (.A0(_2469_),
    .A1(_2510_),
    .S(net1058),
    .X(_2589_));
 sg13g2_mux2_1 _6178_ (.A0(net619),
    .A1(_2589_),
    .S(net1328),
    .X(_0536_));
 sg13g2_mux2_1 _6179_ (.A0(_2449_),
    .A1(_2513_),
    .S(net1058),
    .X(_2590_));
 sg13g2_mux2_1 _6180_ (.A0(net620),
    .A1(_2590_),
    .S(net1325),
    .X(_0537_));
 sg13g2_mux2_1 _6181_ (.A0(_2465_),
    .A1(_2519_),
    .S(net1061),
    .X(_2591_));
 sg13g2_mux2_1 _6182_ (.A0(net652),
    .A1(_2591_),
    .S(net1325),
    .X(_0538_));
 sg13g2_mux2_1 _6183_ (.A0(_2454_),
    .A1(_2499_),
    .S(net1059),
    .X(_2592_));
 sg13g2_mux2_1 _6184_ (.A0(net643),
    .A1(_2592_),
    .S(net1325),
    .X(_0539_));
 sg13g2_mux2_1 _6185_ (.A0(_2467_),
    .A1(_2504_),
    .S(net1059),
    .X(_2593_));
 sg13g2_mux2_1 _6186_ (.A0(net638),
    .A1(_2593_),
    .S(net1325),
    .X(_0540_));
 sg13g2_mux2_1 _6187_ (.A0(_2447_),
    .A1(_2514_),
    .S(net1060),
    .X(_2594_));
 sg13g2_mux2_1 _6188_ (.A0(net646),
    .A1(_2594_),
    .S(net1323),
    .X(_0541_));
 sg13g2_mux2_1 _6189_ (.A0(_2464_),
    .A1(_2506_),
    .S(net1062),
    .X(_2595_));
 sg13g2_mux2_1 _6190_ (.A0(net668),
    .A1(_2595_),
    .S(net1325),
    .X(_0542_));
 sg13g2_mux2_1 _6191_ (.A0(_2450_),
    .A1(_2509_),
    .S(net1060),
    .X(_2596_));
 sg13g2_mux2_1 _6192_ (.A0(net642),
    .A1(_2596_),
    .S(net1323),
    .X(_0543_));
 sg13g2_mux2_1 _6193_ (.A0(_2460_),
    .A1(_2507_),
    .S(net1060),
    .X(_2597_));
 sg13g2_mux2_1 _6194_ (.A0(net623),
    .A1(_2597_),
    .S(net1323),
    .X(_0544_));
 sg13g2_mux2_1 _6195_ (.A0(_2451_),
    .A1(_2498_),
    .S(net1063),
    .X(_2598_));
 sg13g2_mux2_1 _6196_ (.A0(net648),
    .A1(_2598_),
    .S(net1336),
    .X(_0545_));
 sg13g2_mux2_1 _6197_ (.A0(_2456_),
    .A1(_2518_),
    .S(net1060),
    .X(_2599_));
 sg13g2_mux2_1 _6198_ (.A0(net629),
    .A1(_2599_),
    .S(net1328),
    .X(_0546_));
 sg13g2_mux2_1 _6199_ (.A0(_2463_),
    .A1(_2512_),
    .S(net1069),
    .X(_2600_));
 sg13g2_mux2_1 _6200_ (.A0(net682),
    .A1(_2600_),
    .S(net1336),
    .X(_0547_));
 sg13g2_mux2_1 _6201_ (.A0(_2458_),
    .A1(_2500_),
    .S(net1064),
    .X(_2601_));
 sg13g2_mux2_1 _6202_ (.A0(net630),
    .A1(_2601_),
    .S(net1334),
    .X(_0548_));
 sg13g2_mux2_1 _6203_ (.A0(_2485_),
    .A1(_2493_),
    .S(net1066),
    .X(_2602_));
 sg13g2_mux2_1 _6204_ (.A0(net733),
    .A1(_2602_),
    .S(net1381),
    .X(_0549_));
 sg13g2_mux2_1 _6205_ (.A0(_2483_),
    .A1(_2489_),
    .S(net1066),
    .X(_2603_));
 sg13g2_mux2_1 _6206_ (.A0(net767),
    .A1(_2603_),
    .S(net1343),
    .X(_0550_));
 sg13g2_mux2_1 _6207_ (.A0(_2478_),
    .A1(_2494_),
    .S(net1066),
    .X(_2604_));
 sg13g2_mux2_1 _6208_ (.A0(net722),
    .A1(_2604_),
    .S(net1381),
    .X(_0551_));
 sg13g2_mux2_1 _6209_ (.A0(_2486_),
    .A1(_2488_),
    .S(net1066),
    .X(_2605_));
 sg13g2_mux2_1 _6210_ (.A0(net769),
    .A1(_2605_),
    .S(net1379),
    .X(_0552_));
 sg13g2_mux2_1 _6211_ (.A0(_2480_),
    .A1(_2492_),
    .S(net1067),
    .X(_2606_));
 sg13g2_mux2_1 _6212_ (.A0(net900),
    .A1(_2606_),
    .S(net1342),
    .X(_0553_));
 sg13g2_mux2_1 _6213_ (.A0(_2482_),
    .A1(_2487_),
    .S(net1066),
    .X(_2607_));
 sg13g2_mux2_1 _6214_ (.A0(net856),
    .A1(_2607_),
    .S(net1342),
    .X(_0554_));
 sg13g2_mux2_1 _6215_ (.A0(_2479_),
    .A1(_2491_),
    .S(net1067),
    .X(_2608_));
 sg13g2_mux2_1 _6216_ (.A0(net911),
    .A1(_2608_),
    .S(net1343),
    .X(_0555_));
 sg13g2_mux2_1 _6217_ (.A0(net836),
    .A1(_2574_),
    .S(net1343),
    .X(_0556_));
 sg13g2_mux2_1 _6218_ (.A0(_2535_),
    .A1(_2534_),
    .S(net1065),
    .X(_2609_));
 sg13g2_mux2_1 _6219_ (.A0(net813),
    .A1(_2609_),
    .S(net1334),
    .X(_0557_));
 sg13g2_mux2_1 _6220_ (.A0(_2502_),
    .A1(_2448_),
    .S(net1061),
    .X(_2610_));
 sg13g2_mux2_1 _6221_ (.A0(net728),
    .A1(_2610_),
    .S(net1326),
    .X(_0558_));
 sg13g2_mux2_1 _6222_ (.A0(_2508_),
    .A1(_2461_),
    .S(net1061),
    .X(_2611_));
 sg13g2_mux2_1 _6223_ (.A0(net868),
    .A1(_2611_),
    .S(net1326),
    .X(_0559_));
 sg13g2_mux2_1 _6224_ (.A0(_2501_),
    .A1(_2462_),
    .S(net1064),
    .X(_2612_));
 sg13g2_mux2_1 _6225_ (.A0(net752),
    .A1(_2612_),
    .S(net1332),
    .X(_0560_));
 sg13g2_mux2_1 _6226_ (.A0(_2511_),
    .A1(_2452_),
    .S(net1064),
    .X(_2613_));
 sg13g2_mux2_1 _6227_ (.A0(net639),
    .A1(_2613_),
    .S(net1332),
    .X(_0561_));
 sg13g2_mux2_1 _6228_ (.A0(_2503_),
    .A1(_2457_),
    .S(net1061),
    .X(_2614_));
 sg13g2_mux2_1 _6229_ (.A0(net753),
    .A1(_2614_),
    .S(net1326),
    .X(_0562_));
 sg13g2_mux2_1 _6230_ (.A0(_2517_),
    .A1(_2466_),
    .S(net1062),
    .X(_2615_));
 sg13g2_mux2_1 _6231_ (.A0(net926),
    .A1(_2615_),
    .S(net1326),
    .X(_0563_));
 sg13g2_mux2_2 _6232_ (.A0(_2515_),
    .A1(_2453_),
    .S(net1062),
    .X(_2616_));
 sg13g2_mux2_1 _6233_ (.A0(net770),
    .A1(_2616_),
    .S(net1329),
    .X(_0564_));
 sg13g2_mux2_1 _6234_ (.A0(_2520_),
    .A1(_2468_),
    .S(net1062),
    .X(_2617_));
 sg13g2_mux2_1 _6235_ (.A0(net784),
    .A1(_2617_),
    .S(net1329),
    .X(_0565_));
 sg13g2_mux2_1 _6236_ (.A0(_2505_),
    .A1(_2455_),
    .S(net1060),
    .X(_2618_));
 sg13g2_mux2_1 _6237_ (.A0(net914),
    .A1(_2618_),
    .S(net1328),
    .X(_0566_));
 sg13g2_mux2_1 _6238_ (.A0(_2516_),
    .A1(_2459_),
    .S(net1060),
    .X(_2619_));
 sg13g2_mux2_1 _6239_ (.A0(net857),
    .A1(_2619_),
    .S(net1323),
    .X(_0567_));
 sg13g2_mux2_1 _6240_ (.A0(_2510_),
    .A1(_2469_),
    .S(net1058),
    .X(_2620_));
 sg13g2_mux2_1 _6241_ (.A0(net794),
    .A1(_2620_),
    .S(net1325),
    .X(_0568_));
 sg13g2_mux2_1 _6242_ (.A0(_2513_),
    .A1(_2449_),
    .S(net1058),
    .X(_2621_));
 sg13g2_mux2_1 _6243_ (.A0(net843),
    .A1(_2621_),
    .S(net1323),
    .X(_0569_));
 sg13g2_mux2_1 _6244_ (.A0(_2519_),
    .A1(_2465_),
    .S(net1061),
    .X(_2622_));
 sg13g2_mux2_1 _6245_ (.A0(net798),
    .A1(_2622_),
    .S(net1327),
    .X(_0570_));
 sg13g2_mux2_1 _6246_ (.A0(_2499_),
    .A1(_2454_),
    .S(net1059),
    .X(_2623_));
 sg13g2_mux2_1 _6247_ (.A0(net891),
    .A1(_2623_),
    .S(net1324),
    .X(_0571_));
 sg13g2_mux2_1 _6248_ (.A0(_2504_),
    .A1(_2467_),
    .S(net1059),
    .X(_2624_));
 sg13g2_mux2_1 _6249_ (.A0(net698),
    .A1(_2624_),
    .S(net1324),
    .X(_0572_));
 sg13g2_mux2_1 _6250_ (.A0(_2514_),
    .A1(_2447_),
    .S(net1058),
    .X(_2625_));
 sg13g2_mux2_1 _6251_ (.A0(net859),
    .A1(_2625_),
    .S(net1324),
    .X(_0573_));
 sg13g2_mux2_2 _6252_ (.A0(_2506_),
    .A1(_2464_),
    .S(net1061),
    .X(_2626_));
 sg13g2_mux2_1 _6253_ (.A0(net746),
    .A1(_2626_),
    .S(net1324),
    .X(_0574_));
 sg13g2_mux2_1 _6254_ (.A0(_2509_),
    .A1(_2450_),
    .S(net1060),
    .X(_2627_));
 sg13g2_mux2_1 _6255_ (.A0(net1529),
    .A1(_2627_),
    .S(net1323),
    .X(_0575_));
 sg13g2_mux2_1 _6256_ (.A0(_2507_),
    .A1(_2460_),
    .S(net1058),
    .X(_2628_));
 sg13g2_mux2_1 _6257_ (.A0(net901),
    .A1(_2628_),
    .S(net1324),
    .X(_0576_));
 sg13g2_mux2_2 _6258_ (.A0(_2498_),
    .A1(_2451_),
    .S(net1064),
    .X(_2629_));
 sg13g2_mux2_1 _6259_ (.A0(net739),
    .A1(_2629_),
    .S(net1330),
    .X(_0577_));
 sg13g2_mux2_1 _6260_ (.A0(_2518_),
    .A1(_2456_),
    .S(net1060),
    .X(_2630_));
 sg13g2_mux2_1 _6261_ (.A0(net1542),
    .A1(_2630_),
    .S(net1323),
    .X(_0578_));
 sg13g2_mux2_1 _6262_ (.A0(_2512_),
    .A1(_2463_),
    .S(net1064),
    .X(_2631_));
 sg13g2_mux2_1 _6263_ (.A0(net723),
    .A1(_2631_),
    .S(net1333),
    .X(_0579_));
 sg13g2_mux2_1 _6264_ (.A0(_2500_),
    .A1(_2458_),
    .S(net1064),
    .X(_2632_));
 sg13g2_mux2_1 _6265_ (.A0(net847),
    .A1(_2632_),
    .S(net1334),
    .X(_0580_));
 sg13g2_mux2_1 _6266_ (.A0(_2493_),
    .A1(_2485_),
    .S(net1066),
    .X(_2633_));
 sg13g2_mux2_1 _6267_ (.A0(net1493),
    .A1(_2633_),
    .S(net1382),
    .X(_0581_));
 sg13g2_o21ai_1 _6268_ (.B1(net1342),
    .Y(_2634_),
    .A1(_2489_),
    .A2(net1068));
 sg13g2_a21oi_1 _6269_ (.A1(_2484_),
    .A2(net1068),
    .Y(_2635_),
    .B1(_2634_));
 sg13g2_a21o_1 _6270_ (.A2(net742),
    .A1(net1314),
    .B1(_2635_),
    .X(_0582_));
 sg13g2_mux2_1 _6271_ (.A0(_2494_),
    .A1(_2478_),
    .S(net1067),
    .X(_2636_));
 sg13g2_mux2_1 _6272_ (.A0(net1038),
    .A1(_2636_),
    .S(net1380),
    .X(_0583_));
 sg13g2_mux2_1 _6273_ (.A0(_2488_),
    .A1(_2486_),
    .S(net1065),
    .X(_2637_));
 sg13g2_mux2_1 _6274_ (.A0(net711),
    .A1(_2637_),
    .S(net1382),
    .X(_0584_));
 sg13g2_mux2_1 _6275_ (.A0(_2492_),
    .A1(_2480_),
    .S(net1066),
    .X(_2638_));
 sg13g2_mux2_1 _6276_ (.A0(net876),
    .A1(_2638_),
    .S(net1381),
    .X(_0585_));
 sg13g2_mux2_1 _6277_ (.A0(_2487_),
    .A1(_2482_),
    .S(net1066),
    .X(_2639_));
 sg13g2_mux2_1 _6278_ (.A0(net1436),
    .A1(_2639_),
    .S(net1379),
    .X(_0586_));
 sg13g2_mux2_1 _6279_ (.A0(_2491_),
    .A1(_2479_),
    .S(net1067),
    .X(_2640_));
 sg13g2_mux2_1 _6280_ (.A0(net844),
    .A1(_2640_),
    .S(net1381),
    .X(_0587_));
 sg13g2_nor2_1 _6281_ (.A(net1380),
    .B(net943),
    .Y(_2641_));
 sg13g2_a21oi_1 _6282_ (.A1(net1380),
    .A2(_2573_),
    .Y(_0588_),
    .B1(_2641_));
 sg13g2_mux2_1 _6283_ (.A0(_2534_),
    .A1(_2535_),
    .S(net1065),
    .X(_2642_));
 sg13g2_mux2_1 _6284_ (.A0(net760),
    .A1(_2642_),
    .S(net1334),
    .X(_0589_));
 sg13g2_nor2b_1 _6285_ (.A(net1392),
    .B_N(net964),
    .Y(_0590_));
 sg13g2_nor2_1 _6286_ (.A(net1334),
    .B(net1471),
    .Y(_2643_));
 sg13g2_xnor2_1 _6287_ (.Y(_2644_),
    .A(_2560_),
    .B(_2563_));
 sg13g2_a21oi_1 _6288_ (.A1(net1334),
    .A2(_2644_),
    .Y(_0591_),
    .B1(_2643_));
 sg13g2_nand2b_1 _6289_ (.Y(_2645_),
    .B(net1065),
    .A_N(_2644_));
 sg13g2_xnor2_1 _6290_ (.Y(_2646_),
    .A(_2557_),
    .B(_2564_));
 sg13g2_o21ai_1 _6291_ (.B1(net1342),
    .Y(_2647_),
    .A1(_2645_),
    .A2(_2646_));
 sg13g2_a21oi_1 _6292_ (.A1(_2645_),
    .A2(_2646_),
    .Y(_2648_),
    .B1(_2647_));
 sg13g2_a21oi_1 _6293_ (.A1(net1298),
    .A2(_0746_),
    .Y(_0592_),
    .B1(_2648_));
 sg13g2_nand2_1 _6294_ (.Y(_2649_),
    .A(_2557_),
    .B(_2644_));
 sg13g2_nand2_1 _6295_ (.Y(_2650_),
    .A(net1065),
    .B(_2649_));
 sg13g2_xnor2_1 _6296_ (.Y(_2651_),
    .A(_2555_),
    .B(_2566_));
 sg13g2_xnor2_1 _6297_ (.Y(_2652_),
    .A(_2650_),
    .B(_2651_));
 sg13g2_mux2_1 _6298_ (.A0(net1409),
    .A1(_2652_),
    .S(net1335),
    .X(_0593_));
 sg13g2_nor2_1 _6299_ (.A(net1342),
    .B(net861),
    .Y(_2653_));
 sg13g2_nor2_1 _6300_ (.A(_2556_),
    .B(_2649_),
    .Y(_2654_));
 sg13g2_nor3_1 _6301_ (.A(_2576_),
    .B(_2577_),
    .C(_2654_),
    .Y(_2655_));
 sg13g2_nor2b_1 _6302_ (.A(_2552_),
    .B_N(_2553_),
    .Y(_2656_));
 sg13g2_xor2_1 _6303_ (.B(_2656_),
    .A(_2567_),
    .X(_2657_));
 sg13g2_xnor2_1 _6304_ (.Y(_2658_),
    .A(_2655_),
    .B(_2657_));
 sg13g2_a21oi_1 _6305_ (.A1(net1342),
    .A2(_2658_),
    .Y(_0594_),
    .B1(_2653_));
 sg13g2_nand2_1 _6306_ (.Y(_2659_),
    .A(_2654_),
    .B(_2656_));
 sg13g2_nand2_1 _6307_ (.Y(_2660_),
    .A(net1065),
    .B(_2659_));
 sg13g2_xnor2_1 _6308_ (.Y(_2661_),
    .A(_2551_),
    .B(_2568_));
 sg13g2_xnor2_1 _6309_ (.Y(_2662_),
    .A(_2660_),
    .B(_2661_));
 sg13g2_nor2_1 _6310_ (.A(net1379),
    .B(net678),
    .Y(_2663_));
 sg13g2_a21oi_1 _6311_ (.A1(net1379),
    .A2(_2662_),
    .Y(_0595_),
    .B1(_2663_));
 sg13g2_nor2_1 _6312_ (.A(net1379),
    .B(net761),
    .Y(_2664_));
 sg13g2_nor2_1 _6313_ (.A(_2551_),
    .B(_2659_),
    .Y(_2665_));
 sg13g2_nor3_1 _6314_ (.A(_2576_),
    .B(_2577_),
    .C(_2665_),
    .Y(_2666_));
 sg13g2_nor2b_1 _6315_ (.A(_2548_),
    .B_N(_2549_),
    .Y(_2667_));
 sg13g2_xor2_1 _6316_ (.B(_2667_),
    .A(_2569_),
    .X(_2668_));
 sg13g2_xnor2_1 _6317_ (.Y(_2669_),
    .A(_2666_),
    .B(_2668_));
 sg13g2_a21oi_1 _6318_ (.A1(net1379),
    .A2(_2669_),
    .Y(_0596_),
    .B1(_2664_));
 sg13g2_xnor2_1 _6319_ (.Y(_2670_),
    .A(_2547_),
    .B(_2570_));
 sg13g2_nand2_1 _6320_ (.Y(_2671_),
    .A(_2665_),
    .B(_2667_));
 sg13g2_nand2_1 _6321_ (.Y(_2672_),
    .A(net1065),
    .B(_2671_));
 sg13g2_o21ai_1 _6322_ (.B1(net1342),
    .Y(_2673_),
    .A1(_2670_),
    .A2(_2672_));
 sg13g2_a21oi_1 _6323_ (.A1(_2670_),
    .A2(_2672_),
    .Y(_2674_),
    .B1(_2673_));
 sg13g2_a21oi_1 _6324_ (.A1(net1298),
    .A2(_0713_),
    .Y(_0597_),
    .B1(_2674_));
 sg13g2_nor2_1 _6325_ (.A(net1334),
    .B(net997),
    .Y(_2675_));
 sg13g2_xor2_1 _6326_ (.B(_2575_),
    .A(_2572_),
    .X(_2676_));
 sg13g2_o21ai_1 _6327_ (.B1(net1065),
    .Y(_2677_),
    .A1(_2670_),
    .A2(_2671_));
 sg13g2_xnor2_1 _6328_ (.Y(_2678_),
    .A(_2676_),
    .B(_2677_));
 sg13g2_a21oi_1 _6329_ (.A1(net1335),
    .A2(_2678_),
    .Y(_0598_),
    .B1(_2675_));
 sg13g2_nor2b_1 _6330_ (.A(net1333),
    .B_N(net717),
    .Y(_0599_));
 sg13g2_nor2b_1 _6331_ (.A(net1333),
    .B_N(net687),
    .Y(_0600_));
 sg13g2_o21ai_1 _6332_ (.B1(net1340),
    .Y(_2679_),
    .A1(net669),
    .A2(_1371_));
 sg13g2_a21oi_1 _6333_ (.A1(_0680_),
    .A2(_1371_),
    .Y(_0601_),
    .B1(net670));
 sg13g2_nand3_1 _6334_ (.B(\main.spi.state[0] ),
    .C(net1220),
    .A(\main.spi.out_bit_counter[0] ),
    .Y(_2680_));
 sg13g2_or2_1 _6335_ (.X(_2681_),
    .B(_2680_),
    .A(_0679_));
 sg13g2_nand2_1 _6336_ (.Y(_2682_),
    .A(net1339),
    .B(_2681_));
 sg13g2_a21oi_1 _6337_ (.A1(_0679_),
    .A2(_2680_),
    .Y(_0602_),
    .B1(_2682_));
 sg13g2_nand2_1 _6338_ (.Y(_2683_),
    .A(net1429),
    .B(\main.spi.out_bit_counter[1] ));
 sg13g2_o21ai_1 _6339_ (.B1(net1339),
    .Y(_2684_),
    .A1(_2680_),
    .A2(_2683_));
 sg13g2_a21oi_1 _6340_ (.A1(_0678_),
    .A2(_2681_),
    .Y(_0603_),
    .B1(_2684_));
 sg13g2_nand3_1 _6341_ (.B(\main.state[6] ),
    .C(_0767_),
    .A(\main.SPI_output_data_ready ),
    .Y(_2685_));
 sg13g2_nor2b_2 _6342_ (.A(\main.spi.SPI_clock_sampler.sample_register[0] ),
    .B_N(\main.spi.SPI_clock_sampled ),
    .Y(_2686_));
 sg13g2_and4_1 _6343_ (.A(net1429),
    .B(net1592),
    .C(\main.spi.out_bit_counter[0] ),
    .D(_2686_),
    .X(_2687_));
 sg13g2_o21ai_1 _6344_ (.B1(net1128),
    .Y(_2688_),
    .A1(net1596),
    .A2(_2687_));
 sg13g2_nand2_1 _6345_ (.Y(_0604_),
    .A(net1338),
    .B(_2688_));
 sg13g2_nor2_2 _6346_ (.A(_0031_),
    .B(net1128),
    .Y(_2689_));
 sg13g2_mux4_1 _6347_ (.S0(net1268),
    .A0(\main.float_registers[0][16] ),
    .A1(\main.float_registers[1][16] ),
    .A2(\main.float_registers[2][16] ),
    .A3(\main.float_registers[3][16] ),
    .S1(net1263),
    .X(_2690_));
 sg13g2_mux4_1 _6348_ (.S0(net1271),
    .A0(\main.float_registers[0][24] ),
    .A1(\main.float_registers[1][24] ),
    .A2(\main.float_registers[2][24] ),
    .A3(\main.float_registers[3][24] ),
    .S1(net1266),
    .X(_2691_));
 sg13g2_a22oi_1 _6349_ (.Y(_2692_),
    .B1(_2691_),
    .B2(net1224),
    .A2(_2690_),
    .A1(net1223));
 sg13g2_mux4_1 _6350_ (.S0(net1269),
    .A0(\main.float_registers[0][0] ),
    .A1(\main.float_registers[1][0] ),
    .A2(\main.float_registers[2][0] ),
    .A3(\main.float_registers[3][0] ),
    .S1(net1264),
    .X(_2693_));
 sg13g2_mux4_1 _6351_ (.S0(net1269),
    .A0(\main.float_registers[0][8] ),
    .A1(\main.float_registers[1][8] ),
    .A2(\main.float_registers[2][8] ),
    .A3(\main.float_registers[3][8] ),
    .S1(net1264),
    .X(_2694_));
 sg13g2_a22oi_1 _6352_ (.Y(_2695_),
    .B1(_2694_),
    .B2(net1221),
    .A2(_2693_),
    .A1(net1222));
 sg13g2_nand2_1 _6353_ (.Y(_2696_),
    .A(_2692_),
    .B(_2695_));
 sg13g2_a22oi_1 _6354_ (.Y(_2697_),
    .B1(_2689_),
    .B2(_2696_),
    .A2(_2685_),
    .A1(net897));
 sg13g2_nor2_1 _6355_ (.A(net1299),
    .B(net898),
    .Y(_0605_));
 sg13g2_mux4_1 _6356_ (.S0(net1268),
    .A0(\main.float_registers[0][17] ),
    .A1(\main.float_registers[1][17] ),
    .A2(\main.float_registers[2][17] ),
    .A3(\main.float_registers[3][17] ),
    .S1(net1263),
    .X(_2698_));
 sg13g2_mux4_1 _6357_ (.S0(net1268),
    .A0(\main.float_registers[0][1] ),
    .A1(\main.float_registers[1][1] ),
    .A2(\main.float_registers[2][1] ),
    .A3(\main.float_registers[3][1] ),
    .S1(net1263),
    .X(_2699_));
 sg13g2_a22oi_1 _6358_ (.Y(_2700_),
    .B1(_2699_),
    .B2(net1222),
    .A2(_2698_),
    .A1(net1223));
 sg13g2_mux4_1 _6359_ (.S0(net1271),
    .A0(\main.float_registers[0][25] ),
    .A1(\main.float_registers[1][25] ),
    .A2(\main.float_registers[2][25] ),
    .A3(\main.float_registers[3][25] ),
    .S1(net1266),
    .X(_2701_));
 sg13g2_mux4_1 _6360_ (.S0(net1269),
    .A0(\main.float_registers[0][9] ),
    .A1(\main.float_registers[1][9] ),
    .A2(\main.float_registers[2][9] ),
    .A3(\main.float_registers[3][9] ),
    .S1(net1264),
    .X(_2702_));
 sg13g2_a22oi_1 _6361_ (.Y(_2703_),
    .B1(_2702_),
    .B2(_0793_),
    .A2(_2701_),
    .A1(net1224));
 sg13g2_nand2_1 _6362_ (.Y(_2704_),
    .A(_2700_),
    .B(_2703_));
 sg13g2_a22oi_1 _6363_ (.Y(_2705_),
    .B1(_2689_),
    .B2(_2704_),
    .A2(_2685_),
    .A1(net786));
 sg13g2_nor2_1 _6364_ (.A(net1299),
    .B(net787),
    .Y(_0606_));
 sg13g2_mux4_1 _6365_ (.S0(net1268),
    .A0(\main.float_registers[0][18] ),
    .A1(\main.float_registers[1][18] ),
    .A2(\main.float_registers[2][18] ),
    .A3(\main.float_registers[3][18] ),
    .S1(net1263),
    .X(_2706_));
 sg13g2_mux4_1 _6366_ (.S0(net1272),
    .A0(\main.float_registers[0][2] ),
    .A1(\main.float_registers[1][2] ),
    .A2(\main.float_registers[2][2] ),
    .A3(\main.float_registers[3][2] ),
    .S1(net1267),
    .X(_2707_));
 sg13g2_a22oi_1 _6367_ (.Y(_2708_),
    .B1(_2707_),
    .B2(net1222),
    .A2(_2706_),
    .A1(net1223));
 sg13g2_mux4_1 _6368_ (.S0(net1271),
    .A0(\main.float_registers[0][26] ),
    .A1(\main.float_registers[1][26] ),
    .A2(\main.float_registers[2][26] ),
    .A3(\main.float_registers[3][26] ),
    .S1(net1266),
    .X(_2709_));
 sg13g2_mux4_1 _6369_ (.S0(net1269),
    .A0(\main.float_registers[0][10] ),
    .A1(\main.float_registers[1][10] ),
    .A2(\main.float_registers[2][10] ),
    .A3(\main.float_registers[3][10] ),
    .S1(net1264),
    .X(_2710_));
 sg13g2_a22oi_1 _6370_ (.Y(_2711_),
    .B1(_2710_),
    .B2(net1221),
    .A2(_2709_),
    .A1(net1224));
 sg13g2_nand2_1 _6371_ (.Y(_2712_),
    .A(_2708_),
    .B(_2711_));
 sg13g2_a22oi_1 _6372_ (.Y(_2713_),
    .B1(_2689_),
    .B2(_2712_),
    .A2(net1128),
    .A1(net888));
 sg13g2_nor2_1 _6373_ (.A(net1299),
    .B(net889),
    .Y(_0607_));
 sg13g2_mux4_1 _6374_ (.S0(net1270),
    .A0(\main.float_registers[0][19] ),
    .A1(\main.float_registers[1][19] ),
    .A2(\main.float_registers[2][19] ),
    .A3(\main.float_registers[3][19] ),
    .S1(net1265),
    .X(_2714_));
 sg13g2_mux4_1 _6375_ (.S0(net1272),
    .A0(\main.float_registers[0][3] ),
    .A1(\main.float_registers[1][3] ),
    .A2(\main.float_registers[2][3] ),
    .A3(\main.float_registers[3][3] ),
    .S1(net1267),
    .X(_2715_));
 sg13g2_a22oi_1 _6376_ (.Y(_2716_),
    .B1(_2715_),
    .B2(net1222),
    .A2(_2714_),
    .A1(net1223));
 sg13g2_mux4_1 _6377_ (.S0(net1272),
    .A0(\main.float_registers[0][27] ),
    .A1(\main.float_registers[1][27] ),
    .A2(\main.float_registers[2][27] ),
    .A3(\main.float_registers[3][27] ),
    .S1(net1267),
    .X(_2717_));
 sg13g2_mux4_1 _6378_ (.S0(net1269),
    .A0(\main.float_registers[0][11] ),
    .A1(\main.float_registers[1][11] ),
    .A2(\main.float_registers[2][11] ),
    .A3(\main.float_registers[3][11] ),
    .S1(net1264),
    .X(_2718_));
 sg13g2_a22oi_1 _6379_ (.Y(_2719_),
    .B1(_2718_),
    .B2(net1221),
    .A2(_2717_),
    .A1(net1224));
 sg13g2_nand2_1 _6380_ (.Y(_2720_),
    .A(_2716_),
    .B(_2719_));
 sg13g2_a22oi_1 _6381_ (.Y(_2721_),
    .B1(_2689_),
    .B2(_2720_),
    .A2(net1128),
    .A1(net680));
 sg13g2_nor2_1 _6382_ (.A(net1299),
    .B(net681),
    .Y(_0608_));
 sg13g2_mux4_1 _6383_ (.S0(net1268),
    .A0(\main.float_registers[0][20] ),
    .A1(\main.float_registers[1][20] ),
    .A2(\main.float_registers[2][20] ),
    .A3(\main.float_registers[3][20] ),
    .S1(net1263),
    .X(_2722_));
 sg13g2_mux4_1 _6384_ (.S0(net1268),
    .A0(\main.float_registers[0][4] ),
    .A1(\main.float_registers[1][4] ),
    .A2(\main.float_registers[2][4] ),
    .A3(\main.float_registers[3][4] ),
    .S1(net1263),
    .X(_2723_));
 sg13g2_a22oi_1 _6385_ (.Y(_2724_),
    .B1(_2723_),
    .B2(net1222),
    .A2(_2722_),
    .A1(net1223));
 sg13g2_mux4_1 _6386_ (.S0(net1271),
    .A0(\main.float_registers[0][28] ),
    .A1(\main.float_registers[1][28] ),
    .A2(\main.float_registers[2][28] ),
    .A3(\main.float_registers[3][28] ),
    .S1(net1266),
    .X(_2725_));
 sg13g2_mux4_1 _6387_ (.S0(net1269),
    .A0(\main.float_registers[0][12] ),
    .A1(\main.float_registers[1][12] ),
    .A2(\main.float_registers[2][12] ),
    .A3(\main.float_registers[3][12] ),
    .S1(net1264),
    .X(_2726_));
 sg13g2_a22oi_1 _6388_ (.Y(_2727_),
    .B1(_2726_),
    .B2(net1221),
    .A2(_2725_),
    .A1(net1224));
 sg13g2_nand2_1 _6389_ (.Y(_2728_),
    .A(_2724_),
    .B(_2727_));
 sg13g2_a22oi_1 _6390_ (.Y(_2729_),
    .B1(_2689_),
    .B2(_2728_),
    .A2(net1128),
    .A1(net744));
 sg13g2_nor2_1 _6391_ (.A(net1299),
    .B(net745),
    .Y(_0609_));
 sg13g2_mux4_1 _6392_ (.S0(net1268),
    .A0(\main.float_registers[0][21] ),
    .A1(\main.float_registers[1][21] ),
    .A2(\main.float_registers[2][21] ),
    .A3(\main.float_registers[3][21] ),
    .S1(net1263),
    .X(_2730_));
 sg13g2_mux4_1 _6393_ (.S0(net1272),
    .A0(\main.float_registers[0][5] ),
    .A1(\main.float_registers[1][5] ),
    .A2(\main.float_registers[2][5] ),
    .A3(\main.float_registers[3][5] ),
    .S1(net1267),
    .X(_2731_));
 sg13g2_a22oi_1 _6394_ (.Y(_2732_),
    .B1(_2731_),
    .B2(net1222),
    .A2(_2730_),
    .A1(net1223));
 sg13g2_mux4_1 _6395_ (.S0(net1271),
    .A0(\main.float_registers[0][29] ),
    .A1(\main.float_registers[1][29] ),
    .A2(\main.float_registers[2][29] ),
    .A3(\main.float_registers[3][29] ),
    .S1(net1266),
    .X(_2733_));
 sg13g2_mux4_1 _6396_ (.S0(net1269),
    .A0(\main.float_registers[0][13] ),
    .A1(\main.float_registers[1][13] ),
    .A2(\main.float_registers[2][13] ),
    .A3(\main.float_registers[3][13] ),
    .S1(net1264),
    .X(_2734_));
 sg13g2_a22oi_1 _6397_ (.Y(_2735_),
    .B1(_2734_),
    .B2(net1221),
    .A2(_2733_),
    .A1(net1224));
 sg13g2_nand2_1 _6398_ (.Y(_2736_),
    .A(_2732_),
    .B(_2735_));
 sg13g2_a22oi_1 _6399_ (.Y(_2737_),
    .B1(_2689_),
    .B2(_2736_),
    .A2(net1128),
    .A1(net740));
 sg13g2_nor2_1 _6400_ (.A(net1299),
    .B(net741),
    .Y(_0610_));
 sg13g2_mux4_1 _6401_ (.S0(net1268),
    .A0(\main.float_registers[0][22] ),
    .A1(\main.float_registers[1][22] ),
    .A2(\main.float_registers[2][22] ),
    .A3(\main.float_registers[3][22] ),
    .S1(net1263),
    .X(_2738_));
 sg13g2_mux4_1 _6402_ (.S0(net1272),
    .A0(\main.float_registers[0][6] ),
    .A1(\main.float_registers[1][6] ),
    .A2(\main.float_registers[2][6] ),
    .A3(\main.float_registers[3][6] ),
    .S1(net1267),
    .X(_2739_));
 sg13g2_a22oi_1 _6403_ (.Y(_2740_),
    .B1(_2739_),
    .B2(net1222),
    .A2(_2738_),
    .A1(net1223));
 sg13g2_mux4_1 _6404_ (.S0(net1271),
    .A0(\main.float_registers[0][30] ),
    .A1(\main.float_registers[1][30] ),
    .A2(\main.float_registers[2][30] ),
    .A3(\main.float_registers[3][30] ),
    .S1(net1266),
    .X(_2741_));
 sg13g2_mux4_1 _6405_ (.S0(net1270),
    .A0(\main.float_registers[0][14] ),
    .A1(\main.float_registers[1][14] ),
    .A2(\main.float_registers[2][14] ),
    .A3(\main.float_registers[3][14] ),
    .S1(net1265),
    .X(_2742_));
 sg13g2_a22oi_1 _6406_ (.Y(_2743_),
    .B1(_2742_),
    .B2(net1221),
    .A2(_2741_),
    .A1(net1224));
 sg13g2_nand2_1 _6407_ (.Y(_2744_),
    .A(_2740_),
    .B(_2743_));
 sg13g2_a22oi_1 _6408_ (.Y(_2745_),
    .B1(_2689_),
    .B2(_2744_),
    .A2(net1128),
    .A1(net834));
 sg13g2_nor2_1 _6409_ (.A(net1299),
    .B(net835),
    .Y(_0611_));
 sg13g2_mux4_1 _6410_ (.S0(net1270),
    .A0(\main.float_registers[0][23] ),
    .A1(\main.float_registers[1][23] ),
    .A2(\main.float_registers[2][23] ),
    .A3(\main.float_registers[3][23] ),
    .S1(net1265),
    .X(_2746_));
 sg13g2_mux4_1 _6411_ (.S0(net1271),
    .A0(\main.float_registers[0][7] ),
    .A1(\main.float_registers[1][7] ),
    .A2(\main.float_registers[2][7] ),
    .A3(\main.float_registers[3][7] ),
    .S1(net1266),
    .X(_2747_));
 sg13g2_a22oi_1 _6412_ (.Y(_2748_),
    .B1(_2747_),
    .B2(net1222),
    .A2(_2746_),
    .A1(net1223));
 sg13g2_mux4_1 _6413_ (.S0(net1271),
    .A0(\main.float_registers[0][31] ),
    .A1(\main.float_registers[1][31] ),
    .A2(\main.float_registers[2][31] ),
    .A3(\main.float_registers[3][31] ),
    .S1(net1266),
    .X(_2749_));
 sg13g2_mux4_1 _6414_ (.S0(net1269),
    .A0(\main.float_registers[0][15] ),
    .A1(\main.float_registers[1][15] ),
    .A2(\main.float_registers[2][15] ),
    .A3(\main.float_registers[3][15] ),
    .S1(net1264),
    .X(_2750_));
 sg13g2_a22oi_1 _6415_ (.Y(_2751_),
    .B1(_2750_),
    .B2(net1221),
    .A2(_2749_),
    .A1(net1224));
 sg13g2_nand2_1 _6416_ (.Y(_2752_),
    .A(_2748_),
    .B(_2751_));
 sg13g2_a22oi_1 _6417_ (.Y(_2753_),
    .B1(_2689_),
    .B2(_2752_),
    .A2(net1128),
    .A1(net762));
 sg13g2_nor2_1 _6418_ (.A(net1299),
    .B(net763),
    .Y(_0612_));
 sg13g2_mux4_1 _6419_ (.S0(\main.spi.out_bit_counter[0] ),
    .A0(\main.spi.out_data_r[7] ),
    .A1(\main.spi.out_data_r[6] ),
    .A2(\main.spi.out_data_r[5] ),
    .A3(\main.spi.out_data_r[4] ),
    .S1(\main.spi.out_bit_counter[1] ),
    .X(_2754_));
 sg13g2_a21o_1 _6420_ (.A2(_0680_),
    .A1(\main.spi.out_data_r[1] ),
    .B1(_0679_),
    .X(_2755_));
 sg13g2_a21oi_1 _6421_ (.A1(\main.spi.out_data_r[0] ),
    .A2(\main.spi.out_bit_counter[0] ),
    .Y(_2756_),
    .B1(_2755_));
 sg13g2_mux2_1 _6422_ (.A0(\main.spi.out_data_r[3] ),
    .A1(\main.spi.out_data_r[2] ),
    .S(\main.spi.out_bit_counter[0] ),
    .X(_2757_));
 sg13g2_o21ai_1 _6423_ (.B1(\main.spi.out_bit_counter[2] ),
    .Y(_2758_),
    .A1(\main.spi.out_bit_counter[1] ),
    .A2(_2757_));
 sg13g2_o21ai_1 _6424_ (.B1(_2686_),
    .Y(_2759_),
    .A1(_2756_),
    .A2(_2758_));
 sg13g2_a21oi_1 _6425_ (.A1(_0678_),
    .A2(_2754_),
    .Y(_2760_),
    .B1(_2759_));
 sg13g2_nor2_1 _6426_ (.A(net790),
    .B(_2686_),
    .Y(_2761_));
 sg13g2_nor2_1 _6427_ (.A(_2760_),
    .B(net791),
    .Y(_0613_));
 sg13g2_nand2_1 _6428_ (.Y(_2762_),
    .A(\main.spi.state[0] ),
    .B(_2686_));
 sg13g2_a21oi_1 _6429_ (.A1(\main.spi.in_bit_counter[0] ),
    .A2(_2762_),
    .Y(_2763_),
    .B1(net1304));
 sg13g2_o21ai_1 _6430_ (.B1(_2763_),
    .Y(_0614_),
    .A1(_0677_),
    .A2(_2762_));
 sg13g2_nand3_1 _6431_ (.B(\main.spi.state[0] ),
    .C(_2686_),
    .A(net1612),
    .Y(_2764_));
 sg13g2_nand4_1 _6432_ (.B(net1612),
    .C(\main.spi.state[0] ),
    .A(net1477),
    .Y(_2765_),
    .D(_2686_));
 sg13g2_nand2b_1 _6433_ (.Y(_2766_),
    .B(_2764_),
    .A_N(net1477));
 sg13g2_a21o_1 _6434_ (.A2(_2766_),
    .A1(_2765_),
    .B1(net1300),
    .X(_0615_));
 sg13g2_a21oi_1 _6435_ (.A1(net700),
    .A2(_2765_),
    .Y(_2767_),
    .B1(net1300));
 sg13g2_o21ai_1 _6436_ (.B1(_2767_),
    .Y(_0616_),
    .A1(net700),
    .A2(_2765_));
 sg13g2_o21ai_1 _6437_ (.B1(net1344),
    .Y(_2768_),
    .A1(net1246),
    .A2(net1219));
 sg13g2_a21oi_1 _6438_ (.A1(_0676_),
    .A2(net1219),
    .Y(_0617_),
    .B1(_2768_));
 sg13g2_o21ai_1 _6439_ (.B1(net1339),
    .Y(_2769_),
    .A1(net702),
    .A2(net1220));
 sg13g2_a21oi_1 _6440_ (.A1(_0666_),
    .A2(net1220),
    .Y(_0618_),
    .B1(_2769_));
 sg13g2_o21ai_1 _6441_ (.B1(net1344),
    .Y(_2770_),
    .A1(net1544),
    .A2(net1220));
 sg13g2_a21oi_1 _6442_ (.A1(_0664_),
    .A2(net1220),
    .Y(_0619_),
    .B1(_2770_));
 sg13g2_o21ai_1 _6443_ (.B1(net1344),
    .Y(_2771_),
    .A1(net1537),
    .A2(net1218));
 sg13g2_a21oi_1 _6444_ (.A1(_0675_),
    .A2(net1218),
    .Y(_0620_),
    .B1(_2771_));
 sg13g2_o21ai_1 _6445_ (.B1(net1344),
    .Y(_2772_),
    .A1(\main.SPI_input_data[4] ),
    .A2(net1219));
 sg13g2_a21oi_1 _6446_ (.A1(_0674_),
    .A2(net1219),
    .Y(_0621_),
    .B1(_2772_));
 sg13g2_o21ai_1 _6447_ (.B1(net1344),
    .Y(_2773_),
    .A1(net1531),
    .A2(net1218));
 sg13g2_a21oi_1 _6448_ (.A1(_0673_),
    .A2(net1218),
    .Y(_0622_),
    .B1(_2773_));
 sg13g2_o21ai_1 _6449_ (.B1(net1344),
    .Y(_2774_),
    .A1(\main.SPI_input_data[6] ),
    .A2(net1218));
 sg13g2_a21oi_1 _6450_ (.A1(_0672_),
    .A2(net1218),
    .Y(_0623_),
    .B1(_2774_));
 sg13g2_o21ai_1 _6451_ (.B1(net1344),
    .Y(_2775_),
    .A1(\main.SPI_input_data[7] ),
    .A2(net1218));
 sg13g2_a21oi_1 _6452_ (.A1(_0671_),
    .A2(net1218),
    .Y(_0624_),
    .B1(_2775_));
 sg13g2_nand3_1 _6453_ (.B(_0764_),
    .C(_0792_),
    .A(net1274),
    .Y(_2776_));
 sg13g2_o21ai_1 _6454_ (.B1(net1338),
    .Y(_2777_),
    .A1(net1246),
    .A2(_2776_));
 sg13g2_a21oi_1 _6455_ (.A1(_0668_),
    .A2(_2776_),
    .Y(_0625_),
    .B1(_2777_));
 sg13g2_o21ai_1 _6456_ (.B1(net1338),
    .Y(_2778_),
    .A1(net702),
    .A2(_2776_));
 sg13g2_a21oi_1 _6457_ (.A1(_0667_),
    .A2(_2776_),
    .Y(_0626_),
    .B1(_2778_));
 sg13g2_nand3_1 _6458_ (.B(_0764_),
    .C(net1221),
    .A(net1274),
    .Y(_2779_));
 sg13g2_o21ai_1 _6459_ (.B1(net1338),
    .Y(_2780_),
    .A1(net1246),
    .A2(_2779_));
 sg13g2_a21oi_1 _6460_ (.A1(_0670_),
    .A2(_2779_),
    .Y(_0627_),
    .B1(_2780_));
 sg13g2_o21ai_1 _6461_ (.B1(net1338),
    .Y(_2781_),
    .A1(net702),
    .A2(_2779_));
 sg13g2_a21oi_1 _6462_ (.A1(_0669_),
    .A2(_2779_),
    .Y(_0628_),
    .B1(_2781_));
 sg13g2_a21oi_1 _6463_ (.A1(_0698_),
    .A2(_0781_),
    .Y(_0633_),
    .B1(_0782_));
 sg13g2_a21oi_1 _6464_ (.A1(_0699_),
    .A2(_0781_),
    .Y(_0634_),
    .B1(_0784_));
 sg13g2_nor2_1 _6465_ (.A(net1358),
    .B(net714),
    .Y(_2782_));
 sg13g2_a22oi_1 _6466_ (.Y(_2783_),
    .B1(_2004_),
    .B2(net1247),
    .A2(_1900_),
    .A1(_1819_));
 sg13g2_a21oi_1 _6467_ (.A1(net1358),
    .A2(_2783_),
    .Y(_0635_),
    .B1(_2782_));
 sg13g2_nor2_1 _6468_ (.A(net1357),
    .B(net694),
    .Y(_2784_));
 sg13g2_a22oi_1 _6469_ (.Y(_2785_),
    .B1(_2006_),
    .B2(net1247),
    .A2(_1919_),
    .A1(_1819_));
 sg13g2_a21oi_1 _6470_ (.A1(net1357),
    .A2(_2785_),
    .Y(_0636_),
    .B1(_2784_));
 sg13g2_nor2_1 _6471_ (.A(net1357),
    .B(net697),
    .Y(_2786_));
 sg13g2_a22oi_1 _6472_ (.Y(_2787_),
    .B1(_2008_),
    .B2(net1247),
    .A2(_1937_),
    .A1(_1819_));
 sg13g2_a21oi_1 _6473_ (.A1(net1357),
    .A2(_2787_),
    .Y(_0637_),
    .B1(_2786_));
 sg13g2_nand3_1 _6474_ (.B(net1136),
    .C(_1941_),
    .A(net1248),
    .Y(_2788_));
 sg13g2_a21oi_1 _6475_ (.A1(_1819_),
    .A2(_1945_),
    .Y(_2789_),
    .B1(net1306));
 sg13g2_a22oi_1 _6476_ (.Y(_0638_),
    .B1(_2788_),
    .B2(_2789_),
    .A2(_0760_),
    .A1(net1305));
 sg13g2_nand3b_1 _6477_ (.B(net1136),
    .C(net1248),
    .Y(_2790_),
    .A_N(_1950_));
 sg13g2_o21ai_1 _6478_ (.B1(_2790_),
    .Y(_2791_),
    .A1(_1820_),
    .A2(_1955_));
 sg13g2_mux2_1 _6479_ (.A0(net777),
    .A1(_2791_),
    .S(net1354),
    .X(_0639_));
 sg13g2_nand3_1 _6480_ (.B(net1136),
    .C(_1960_),
    .A(net1248),
    .Y(_2792_));
 sg13g2_o21ai_1 _6481_ (.B1(_2792_),
    .Y(_2793_),
    .A1(_1820_),
    .A2(_1965_));
 sg13g2_mux2_1 _6482_ (.A0(net768),
    .A1(_2793_),
    .S(net1355),
    .X(_0640_));
 sg13g2_nand3_1 _6483_ (.B(net1136),
    .C(_1970_),
    .A(net1248),
    .Y(_2794_));
 sg13g2_o21ai_1 _6484_ (.B1(_2794_),
    .Y(_2795_),
    .A1(_1820_),
    .A2(_1973_));
 sg13g2_mux2_1 _6485_ (.A0(net730),
    .A1(_2795_),
    .S(net1354),
    .X(_0641_));
 sg13g2_a221oi_1 _6486_ (.B2(_1816_),
    .C1(net1305),
    .B1(_2015_),
    .A1(_1819_),
    .Y(_2796_),
    .A2(_1978_));
 sg13g2_a21oi_1 _6487_ (.A1(net1308),
    .A2(_0761_),
    .Y(_0642_),
    .B1(_2796_));
 sg13g2_o21ai_1 _6488_ (.B1(_1818_),
    .Y(_2797_),
    .A1(_1885_),
    .A2(_1980_));
 sg13g2_nand2b_1 _6489_ (.Y(_2798_),
    .B(_1898_),
    .A_N(_1866_));
 sg13g2_o21ai_1 _6490_ (.B1(_2798_),
    .Y(_2799_),
    .A1(net1135),
    .A2(_1983_));
 sg13g2_o21ai_1 _6491_ (.B1(_2797_),
    .Y(_2800_),
    .A1(_1816_),
    .A2(_2799_));
 sg13g2_o21ai_1 _6492_ (.B1(_2800_),
    .Y(_0643_),
    .A1(net1353),
    .A2(_0762_));
 sg13g2_o21ai_1 _6493_ (.B1(_1818_),
    .Y(_2801_),
    .A1(_1885_),
    .A2(_1984_));
 sg13g2_nor2_1 _6494_ (.A(net1134),
    .B(_1985_),
    .Y(_2802_));
 sg13g2_o21ai_1 _6495_ (.B1(_1815_),
    .Y(_2803_),
    .A1(_1866_),
    .A2(_1917_));
 sg13g2_o21ai_1 _6496_ (.B1(_2801_),
    .Y(_2804_),
    .A1(_2802_),
    .A2(_2803_));
 sg13g2_o21ai_1 _6497_ (.B1(_2804_),
    .Y(_0644_),
    .A1(net1355),
    .A2(_0763_));
 sg13g2_nand2_1 _6498_ (.Y(_2805_),
    .A(net1309),
    .B(net743));
 sg13g2_a21oi_1 _6499_ (.A1(_1884_),
    .A2(_1988_),
    .Y(_2806_),
    .B1(net1131));
 sg13g2_nor2_1 _6500_ (.A(net1135),
    .B(_1990_),
    .Y(_2807_));
 sg13g2_nor3_1 _6501_ (.A(net1155),
    .B(_1866_),
    .C(_1935_),
    .Y(_2808_));
 sg13g2_nor3_1 _6502_ (.A(_1816_),
    .B(_2807_),
    .C(_2808_),
    .Y(_2809_));
 sg13g2_o21ai_1 _6503_ (.B1(_2805_),
    .Y(_0645_),
    .A1(_2806_),
    .A2(_2809_));
 sg13g2_nor2_1 _6504_ (.A(net1134),
    .B(_1991_),
    .Y(_2810_));
 sg13g2_nor2_1 _6505_ (.A(_1866_),
    .B(_1944_),
    .Y(_2811_));
 sg13g2_o21ai_1 _6506_ (.B1(_1815_),
    .Y(_2812_),
    .A1(_2810_),
    .A2(_2811_));
 sg13g2_nand3_1 _6507_ (.B(net1134),
    .C(_1992_),
    .A(net1247),
    .Y(_2813_));
 sg13g2_nand3_1 _6508_ (.B(_2812_),
    .C(_2813_),
    .A(net1348),
    .Y(_2814_));
 sg13g2_o21ai_1 _6509_ (.B1(_2814_),
    .Y(_2815_),
    .A1(net1352),
    .A2(net1396));
 sg13g2_inv_1 _6510_ (.Y(_0646_),
    .A(_2815_));
 sg13g2_or2_1 _6511_ (.X(_2816_),
    .B(_1953_),
    .A(_1866_));
 sg13g2_o21ai_1 _6512_ (.B1(_2816_),
    .Y(_2817_),
    .A1(net1135),
    .A2(_1995_));
 sg13g2_nand4_1 _6513_ (.B(net1247),
    .C(net1135),
    .A(net1352),
    .Y(_2818_),
    .D(_1996_));
 sg13g2_a22oi_1 _6514_ (.Y(_2819_),
    .B1(net1131),
    .B2(_2817_),
    .A2(net705),
    .A1(net1298));
 sg13g2_nand2_1 _6515_ (.Y(_0647_),
    .A(_2818_),
    .B(_2819_));
 sg13g2_nand2b_1 _6516_ (.Y(_2820_),
    .B(_1962_),
    .A_N(_1866_));
 sg13g2_o21ai_1 _6517_ (.B1(_2820_),
    .Y(_2821_),
    .A1(net1134),
    .A2(_1998_));
 sg13g2_nand2_1 _6518_ (.Y(_2822_),
    .A(_1815_),
    .B(_2821_));
 sg13g2_nand3_1 _6519_ (.B(net1134),
    .C(_1999_),
    .A(net1247),
    .Y(_2823_));
 sg13g2_nand3_1 _6520_ (.B(_2822_),
    .C(_2823_),
    .A(net1348),
    .Y(_2824_));
 sg13g2_o21ai_1 _6521_ (.B1(_2824_),
    .Y(_2825_),
    .A1(net1350),
    .A2(net883));
 sg13g2_inv_1 _6522_ (.Y(_0648_),
    .A(_2825_));
 sg13g2_nor2_1 _6523_ (.A(net1137),
    .B(_2001_),
    .Y(_2826_));
 sg13g2_nor2_1 _6524_ (.A(_1866_),
    .B(_1971_),
    .Y(_2827_));
 sg13g2_o21ai_1 _6525_ (.B1(_1815_),
    .Y(_2828_),
    .A1(_2826_),
    .A2(_2827_));
 sg13g2_nand3_1 _6526_ (.B(net1136),
    .C(_2002_),
    .A(net1248),
    .Y(_2829_));
 sg13g2_nand3_1 _6527_ (.B(_2828_),
    .C(_2829_),
    .A(net1353),
    .Y(_2830_));
 sg13g2_o21ai_1 _6528_ (.B1(_2830_),
    .Y(_2831_),
    .A1(net1355),
    .A2(net864));
 sg13g2_inv_1 _6529_ (.Y(_0649_),
    .A(_2831_));
 sg13g2_nor2_1 _6530_ (.A(net1453),
    .B(net1104),
    .Y(_2832_));
 sg13g2_a21oi_1 _6531_ (.A1(net1104),
    .A2(_0846_),
    .Y(_0650_),
    .B1(_2832_));
 sg13g2_nor2_1 _6532_ (.A(net1481),
    .B(net1101),
    .Y(_2833_));
 sg13g2_a21oi_1 _6533_ (.A1(net1101),
    .A2(_0940_),
    .Y(_0651_),
    .B1(_2833_));
 sg13g2_nor2_1 _6534_ (.A(net1463),
    .B(net1090),
    .Y(_2834_));
 sg13g2_a21oi_1 _6535_ (.A1(_0930_),
    .A2(net1090),
    .Y(_0652_),
    .B1(_2834_));
 sg13g2_nor2_1 _6536_ (.A(net989),
    .B(net1101),
    .Y(_2835_));
 sg13g2_a21oi_1 _6537_ (.A1(net1101),
    .A2(_0895_),
    .Y(_0653_),
    .B1(_2835_));
 sg13g2_nor2_1 _6538_ (.A(net979),
    .B(net1101),
    .Y(_2836_));
 sg13g2_a21oi_1 _6539_ (.A1(net1101),
    .A2(_0870_),
    .Y(_0654_),
    .B1(_2836_));
 sg13g2_nand2_1 _6540_ (.Y(_2837_),
    .A(net937),
    .B(net1093));
 sg13g2_o21ai_1 _6541_ (.B1(_2837_),
    .Y(_0655_),
    .A1(net1093),
    .A2(_1003_));
 sg13g2_nor2_1 _6542_ (.A(net1009),
    .B(net1110),
    .Y(_2838_));
 sg13g2_a21oi_1 _6543_ (.A1(_0930_),
    .A2(net1110),
    .Y(_0656_),
    .B1(_2838_));
 sg13g2_nor2_1 _6544_ (.A(net1425),
    .B(net1076),
    .Y(_2839_));
 sg13g2_a21oi_1 _6545_ (.A1(_0953_),
    .A2(net1076),
    .Y(_0657_),
    .B1(_2839_));
 sg13g2_nor2_1 _6546_ (.A(net1034),
    .B(net1076),
    .Y(_2840_));
 sg13g2_a21oi_1 _6547_ (.A1(_0949_),
    .A2(net1076),
    .Y(_0660_),
    .B1(_2840_));
 sg13g2_nor2_1 _6548_ (.A(net1506),
    .B(net1105),
    .Y(_2841_));
 sg13g2_a21oi_1 _6549_ (.A1(net1105),
    .A2(_0966_),
    .Y(_0661_),
    .B1(_2841_));
 sg13g2_nor2_1 _6550_ (.A(net1450),
    .B(net1077),
    .Y(_2842_));
 sg13g2_a21oi_1 _6551_ (.A1(_0945_),
    .A2(net1077),
    .Y(_0662_),
    .B1(_2842_));
 sg13g2_nor2_1 _6552_ (.A(net1454),
    .B(net1077),
    .Y(_2843_));
 sg13g2_a21oi_1 _6553_ (.A1(_1003_),
    .A2(net1077),
    .Y(_0663_),
    .B1(_2843_));
 sg13g2_a21oi_1 _6554_ (.A1(_0668_),
    .A2(_2776_),
    .Y(_0629_),
    .B1(_2777_));
 sg13g2_a21oi_1 _6555_ (.A1(_0667_),
    .A2(_2776_),
    .Y(_0630_),
    .B1(_2778_));
 sg13g2_a21oi_1 _6556_ (.A1(_0666_),
    .A2(_2032_),
    .Y(_0631_),
    .B1(_2033_));
 sg13g2_a21oi_1 _6557_ (.A1(_0664_),
    .A2(_2032_),
    .Y(_0632_),
    .B1(_2034_));
 sg13g2_a21oi_1 _6558_ (.A1(_0670_),
    .A2(_2779_),
    .Y(_0658_),
    .B1(_2780_));
 sg13g2_a21oi_1 _6559_ (.A1(_0669_),
    .A2(_2779_),
    .Y(_0659_),
    .B1(_2781_));
 sg13g2_dfrbp_1 _6560_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net142),
    .D(_0126_),
    .Q_N(_0064_),
    .Q(\main.byte_counter[1] ));
 sg13g2_dfrbp_1 _6561_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net322),
    .D(_0127_),
    .Q_N(_3270_),
    .Q(\main.byte_counter[0] ));
 sg13g2_dfrbp_1 _6562_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net320),
    .D(net1487),
    .Q_N(_3269_),
    .Q(\main.float_registers[2][30] ));
 sg13g2_dfrbp_1 _6563_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net318),
    .D(_0129_),
    .Q_N(_3268_),
    .Q(\main.float_registers[3][3] ));
 sg13g2_dfrbp_1 _6564_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net317),
    .D(_0130_),
    .Q_N(_3267_),
    .Q(\main.float_registers[3][4] ));
 sg13g2_dfrbp_1 _6565_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net316),
    .D(_0131_),
    .Q_N(_3266_),
    .Q(\main.float_registers[3][8] ));
 sg13g2_dfrbp_1 _6566_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net315),
    .D(_0132_),
    .Q_N(_3265_),
    .Q(\main.float_registers[0][7] ));
 sg13g2_dfrbp_1 _6567_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net313),
    .D(_0133_),
    .Q_N(_3264_),
    .Q(\main.float_registers[0][6] ));
 sg13g2_dfrbp_1 _6568_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net311),
    .D(_0134_),
    .Q_N(_3263_),
    .Q(\main.float_registers[0][16] ));
 sg13g2_dfrbp_1 _6569_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net309),
    .D(_0135_),
    .Q_N(_3262_),
    .Q(\main.float_registers[0][5] ));
 sg13g2_dfrbp_1 _6570_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net307),
    .D(_0136_),
    .Q_N(_3261_),
    .Q(\main.float_registers[0][4] ));
 sg13g2_dfrbp_1 _6571_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net305),
    .D(_0137_),
    .Q_N(_3260_),
    .Q(\main.float_registers[0][15] ));
 sg13g2_dfrbp_1 _6572_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net303),
    .D(_0138_),
    .Q_N(_3259_),
    .Q(\main.float_registers[0][3] ));
 sg13g2_dfrbp_1 _6573_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net301),
    .D(net863),
    .Q_N(_3258_),
    .Q(\main.float_registers[0][9] ));
 sg13g2_dfrbp_1 _6574_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net299),
    .D(_0140_),
    .Q_N(_3257_),
    .Q(\main.float_registers[0][8] ));
 sg13g2_dfrbp_1 _6575_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net297),
    .D(_0141_),
    .Q_N(_3256_),
    .Q(\main.float_registers[0][23] ));
 sg13g2_dfrbp_1 _6576_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net295),
    .D(_0142_),
    .Q_N(_3255_),
    .Q(\main.float_registers[0][22] ));
 sg13g2_dfrbp_1 _6577_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net293),
    .D(_0143_),
    .Q_N(_3254_),
    .Q(\main.float_registers[0][12] ));
 sg13g2_dfrbp_1 _6578_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net291),
    .D(_0144_),
    .Q_N(_3253_),
    .Q(\main.float_registers[0][11] ));
 sg13g2_dfrbp_1 _6579_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net289),
    .D(net913),
    .Q_N(_3252_),
    .Q(\main.float_registers[0][10] ));
 sg13g2_dfrbp_1 _6580_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net287),
    .D(_0146_),
    .Q_N(_3251_),
    .Q(\main.float_registers[0][21] ));
 sg13g2_dfrbp_1 _6581_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net285),
    .D(_0147_),
    .Q_N(_3250_),
    .Q(\main.float_registers[0][20] ));
 sg13g2_dfrbp_1 _6582_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net283),
    .D(_0148_),
    .Q_N(_3249_),
    .Q(\main.float_registers[0][19] ));
 sg13g2_dfrbp_1 _6583_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net281),
    .D(_0149_),
    .Q_N(_3248_),
    .Q(\main.float_registers[0][18] ));
 sg13g2_dfrbp_1 _6584_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net279),
    .D(_0150_),
    .Q_N(_3247_),
    .Q(\main.float_registers[0][17] ));
 sg13g2_dfrbp_1 _6585_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net277),
    .D(_0151_),
    .Q_N(_3246_),
    .Q(\main.float_registers[0][2] ));
 sg13g2_dfrbp_1 _6586_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net275),
    .D(_0152_),
    .Q_N(_3245_),
    .Q(\main.float_registers[0][0] ));
 sg13g2_dfrbp_1 _6587_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net273),
    .D(_0153_),
    .Q_N(_3244_),
    .Q(\main.float_registers[0][13] ));
 sg13g2_dfrbp_1 _6588_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net271),
    .D(net818),
    .Q_N(_3243_),
    .Q(\main.float_registers[0][14] ));
 sg13g2_dfrbp_1 _6589_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net269),
    .D(net881),
    .Q_N(_3242_),
    .Q(\main.float_registers[0][25] ));
 sg13g2_dfrbp_1 _6590_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net267),
    .D(_0156_),
    .Q_N(_3241_),
    .Q(\main.float_registers[0][26] ));
 sg13g2_dfrbp_1 _6591_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net265),
    .D(net896),
    .Q_N(_3240_),
    .Q(\main.float_registers[0][27] ));
 sg13g2_dfrbp_1 _6592_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net263),
    .D(net804),
    .Q_N(_3239_),
    .Q(\main.float_registers[0][28] ));
 sg13g2_dfrbp_1 _6593_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net261),
    .D(net949),
    .Q_N(_3238_),
    .Q(\main.float_registers[0][29] ));
 sg13g2_dfrbp_1 _6594_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net259),
    .D(_0160_),
    .Q_N(_3237_),
    .Q(\main.float_registers[0][30] ));
 sg13g2_dfrbp_1 _6595_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net257),
    .D(net872),
    .Q_N(_3236_),
    .Q(\main.float_registers[0][31] ));
 sg13g2_dfrbp_1 _6596_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net255),
    .D(_0162_),
    .Q_N(_3235_),
    .Q(\main.float_registers[0][1] ));
 sg13g2_dfrbp_1 _6597_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net253),
    .D(_0163_),
    .Q_N(_3234_),
    .Q(\main.float_registers[1][1] ));
 sg13g2_dfrbp_1 _6598_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net251),
    .D(_0164_),
    .Q_N(_3233_),
    .Q(\main.float_registers[1][2] ));
 sg13g2_dfrbp_1 _6599_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net249),
    .D(_0165_),
    .Q_N(_3232_),
    .Q(\main.float_registers[1][3] ));
 sg13g2_dfrbp_1 _6600_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net247),
    .D(_0166_),
    .Q_N(_3231_),
    .Q(\main.float_registers[1][4] ));
 sg13g2_dfrbp_1 _6601_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net245),
    .D(_0167_),
    .Q_N(_3230_),
    .Q(\main.float_registers[1][5] ));
 sg13g2_dfrbp_1 _6602_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net243),
    .D(_0168_),
    .Q_N(_3229_),
    .Q(\main.float_registers[1][6] ));
 sg13g2_dfrbp_1 _6603_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net241),
    .D(_0169_),
    .Q_N(_3228_),
    .Q(\main.float_registers[1][7] ));
 sg13g2_dfrbp_1 _6604_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net239),
    .D(_0170_),
    .Q_N(_3227_),
    .Q(\main.float_registers[1][8] ));
 sg13g2_dfrbp_1 _6605_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net237),
    .D(net1495),
    .Q_N(_3226_),
    .Q(\main.float_registers[1][9] ));
 sg13g2_dfrbp_1 _6606_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net235),
    .D(net1414),
    .Q_N(_3225_),
    .Q(\main.float_registers[1][10] ));
 sg13g2_dfrbp_1 _6607_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net233),
    .D(_0173_),
    .Q_N(_3224_),
    .Q(\main.float_registers[1][11] ));
 sg13g2_dfrbp_1 _6608_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net231),
    .D(_0174_),
    .Q_N(_3223_),
    .Q(\main.float_registers[1][12] ));
 sg13g2_dfrbp_1 _6609_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net229),
    .D(_0175_),
    .Q_N(_3222_),
    .Q(\main.float_registers[1][13] ));
 sg13g2_dfrbp_1 _6610_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net227),
    .D(net1512),
    .Q_N(_3221_),
    .Q(\main.float_registers[1][14] ));
 sg13g2_dfrbp_1 _6611_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net225),
    .D(net1033),
    .Q_N(_3220_),
    .Q(\main.float_registers[1][15] ));
 sg13g2_dfrbp_1 _6612_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net223),
    .D(_0178_),
    .Q_N(_3219_),
    .Q(\main.float_registers[1][16] ));
 sg13g2_dfrbp_1 _6613_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net221),
    .D(_0179_),
    .Q_N(_3218_),
    .Q(\main.float_registers[1][17] ));
 sg13g2_dfrbp_1 _6614_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net219),
    .D(_0180_),
    .Q_N(_3217_),
    .Q(\main.float_registers[1][18] ));
 sg13g2_dfrbp_1 _6615_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net217),
    .D(_0181_),
    .Q_N(_3216_),
    .Q(\main.float_registers[1][19] ));
 sg13g2_dfrbp_1 _6616_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net215),
    .D(_0182_),
    .Q_N(_3215_),
    .Q(\main.float_registers[1][20] ));
 sg13g2_dfrbp_1 _6617_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net213),
    .D(_0183_),
    .Q_N(_3214_),
    .Q(\main.float_registers[1][21] ));
 sg13g2_dfrbp_1 _6618_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net211),
    .D(_0184_),
    .Q_N(_3213_),
    .Q(\main.float_registers[1][22] ));
 sg13g2_dfrbp_1 _6619_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net209),
    .D(_0185_),
    .Q_N(_3212_),
    .Q(\main.float_registers[1][23] ));
 sg13g2_dfrbp_1 _6620_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net207),
    .D(_0186_),
    .Q_N(_3211_),
    .Q(\main.float_registers[1][24] ));
 sg13g2_dfrbp_1 _6621_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net205),
    .D(net1428),
    .Q_N(_3210_),
    .Q(\main.float_registers[1][25] ));
 sg13g2_dfrbp_1 _6622_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net203),
    .D(_0188_),
    .Q_N(_3209_),
    .Q(\main.float_registers[1][26] ));
 sg13g2_dfrbp_1 _6623_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net201),
    .D(_0189_),
    .Q_N(_3208_),
    .Q(\main.float_registers[1][27] ));
 sg13g2_dfrbp_1 _6624_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net199),
    .D(net1037),
    .Q_N(_3207_),
    .Q(\main.float_registers[1][28] ));
 sg13g2_dfrbp_1 _6625_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net197),
    .D(net974),
    .Q_N(_3206_),
    .Q(\main.float_registers[1][29] ));
 sg13g2_dfrbp_1 _6626_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net195),
    .D(_0192_),
    .Q_N(_3205_),
    .Q(\main.float_registers[1][30] ));
 sg13g2_dfrbp_1 _6627_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net193),
    .D(net1014),
    .Q_N(_3204_),
    .Q(\main.float_registers[1][31] ));
 sg13g2_dfrbp_1 _6628_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net191),
    .D(_0194_),
    .Q_N(_3203_),
    .Q(\main.float_registers[2][1] ));
 sg13g2_dfrbp_1 _6629_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net189),
    .D(_0195_),
    .Q_N(_3202_),
    .Q(\main.float_registers[2][2] ));
 sg13g2_dfrbp_1 _6630_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net187),
    .D(_0196_),
    .Q_N(_3201_),
    .Q(\main.float_registers[2][3] ));
 sg13g2_dfrbp_1 _6631_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net185),
    .D(_0197_),
    .Q_N(_3200_),
    .Q(\main.float_registers[2][4] ));
 sg13g2_dfrbp_1 _6632_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net183),
    .D(_0198_),
    .Q_N(_3199_),
    .Q(\main.float_registers[2][5] ));
 sg13g2_dfrbp_1 _6633_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net181),
    .D(_0199_),
    .Q_N(_3198_),
    .Q(\main.float_registers[2][6] ));
 sg13g2_dfrbp_1 _6634_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net179),
    .D(_0200_),
    .Q_N(_3197_),
    .Q(\main.float_registers[2][7] ));
 sg13g2_dfrbp_1 _6635_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net177),
    .D(_0201_),
    .Q_N(_3196_),
    .Q(\main.float_registers[2][8] ));
 sg13g2_dfrbp_1 _6636_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net175),
    .D(net1525),
    .Q_N(_3195_),
    .Q(\main.float_registers[2][9] ));
 sg13g2_dfrbp_1 _6637_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net173),
    .D(net1418),
    .Q_N(_3194_),
    .Q(\main.float_registers[2][10] ));
 sg13g2_dfrbp_1 _6638_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net171),
    .D(_0204_),
    .Q_N(_3193_),
    .Q(\main.float_registers[2][11] ));
 sg13g2_dfrbp_1 _6639_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net169),
    .D(_0205_),
    .Q_N(_3192_),
    .Q(\main.float_registers[2][12] ));
 sg13g2_dfrbp_1 _6640_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net167),
    .D(_0206_),
    .Q_N(_3191_),
    .Q(\main.float_registers[2][13] ));
 sg13g2_dfrbp_1 _6641_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net165),
    .D(net1492),
    .Q_N(_3190_),
    .Q(\main.float_registers[2][14] ));
 sg13g2_dfrbp_1 _6642_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net163),
    .D(_0208_),
    .Q_N(_3189_),
    .Q(\main.float_registers[2][15] ));
 sg13g2_dfrbp_1 _6643_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net161),
    .D(_0209_),
    .Q_N(_3188_),
    .Q(\main.float_registers[2][16] ));
 sg13g2_dfrbp_1 _6644_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net159),
    .D(_0210_),
    .Q_N(_3187_),
    .Q(\main.float_registers[2][17] ));
 sg13g2_dfrbp_1 _6645_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net157),
    .D(_0211_),
    .Q_N(_3186_),
    .Q(\main.float_registers[2][18] ));
 sg13g2_dfrbp_1 _6646_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net155),
    .D(_0212_),
    .Q_N(_3185_),
    .Q(\main.float_registers[2][19] ));
 sg13g2_dfrbp_1 _6647_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net153),
    .D(_0213_),
    .Q_N(_3184_),
    .Q(\main.float_registers[2][20] ));
 sg13g2_dfrbp_1 _6648_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net151),
    .D(_0214_),
    .Q_N(_3183_),
    .Q(\main.float_registers[2][21] ));
 sg13g2_dfrbp_1 _6649_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net149),
    .D(_0215_),
    .Q_N(_3182_),
    .Q(\main.float_registers[2][22] ));
 sg13g2_dfrbp_1 _6650_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net141),
    .D(_0216_),
    .Q_N(_3181_),
    .Q(\main.float_registers[2][23] ));
 sg13g2_dfrbp_1 _6651_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net139),
    .D(_0217_),
    .Q_N(_3180_),
    .Q(\main.float_registers[2][24] ));
 sg13g2_dfrbp_1 _6652_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net137),
    .D(net1003),
    .Q_N(_3179_),
    .Q(\main.float_registers[2][25] ));
 sg13g2_dfrbp_1 _6653_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net135),
    .D(_0219_),
    .Q_N(_3178_),
    .Q(\main.float_registers[2][26] ));
 sg13g2_dfrbp_1 _6654_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net133),
    .D(_0220_),
    .Q_N(_3177_),
    .Q(\main.float_registers[2][27] ));
 sg13g2_dfrbp_1 _6655_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(net1011),
    .Q_N(_3176_),
    .Q(\main.float_registers[2][28] ));
 sg13g2_dfrbp_1 _6656_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net129),
    .D(net1459),
    .Q_N(_3175_),
    .Q(\main.float_registers[2][29] ));
 sg13g2_dfrbp_1 _6657_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net127),
    .D(net1443),
    .Q_N(_3174_),
    .Q(\main.float_registers[3][31] ));
 sg13g2_dfrbp_1 _6658_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net126),
    .D(net1016),
    .Q_N(_3173_),
    .Q(\main.float_registers[3][30] ));
 sg13g2_dfrbp_1 _6659_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net125),
    .D(net1551),
    .Q_N(_3172_),
    .Q(\main.adder.s4_exponent_adjust[0] ));
 sg13g2_dfrbp_1 _6660_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net124),
    .D(_0226_),
    .Q_N(_3171_),
    .Q(\main.adder.s4_exponent_adjust[1] ));
 sg13g2_dfrbp_1 _6661_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net123),
    .D(_0227_),
    .Q_N(_3170_),
    .Q(\main.adder.s4_exponent_adjust[2] ));
 sg13g2_dfrbp_1 _6662_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net122),
    .D(_0228_),
    .Q_N(_3169_),
    .Q(\main.adder.s4_exponent_adjust[3] ));
 sg13g2_dfrbp_1 _6663_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net121),
    .D(_0229_),
    .Q_N(_3168_),
    .Q(\main.adder.s4_exponent_adjust[4] ));
 sg13g2_dfrbp_1 _6664_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net120),
    .D(_0230_),
    .Q_N(_3167_),
    .Q(\main.adder.s4_exponent_adjust[5] ));
 sg13g2_dfrbp_1 _6665_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net119),
    .D(net1522),
    .Q_N(_3166_),
    .Q(\main.adder.s4_exponent_adjust[6] ));
 sg13g2_dfrbp_1 _6666_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net118),
    .D(_0232_),
    .Q_N(_3165_),
    .Q(\main.adder.s4_exponent_adjust[7] ));
 sg13g2_dfrbp_1 _6667_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net117),
    .D(_0233_),
    .Q_N(_0073_),
    .Q(\main.adder.s4_exponent_adjust[8] ));
 sg13g2_dfrbp_1 _6668_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net116),
    .D(_0234_),
    .Q_N(_3164_),
    .Q(\main.float_registers[3][17] ));
 sg13g2_dfrbp_1 _6669_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net115),
    .D(_0235_),
    .Q_N(_3163_),
    .Q(\main.float_registers[3][16] ));
 sg13g2_dfrbp_1 _6670_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net114),
    .D(_0236_),
    .Q_N(_3162_),
    .Q(\main.float_registers[3][22] ));
 sg13g2_dfrbp_1 _6671_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net113),
    .D(_0237_),
    .Q_N(_3161_),
    .Q(\main.float_registers[3][23] ));
 sg13g2_dfrbp_1 _6672_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net112),
    .D(net985),
    .Q_N(_3160_),
    .Q(\main.float_registers[3][9] ));
 sg13g2_dfrbp_1 _6673_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net111),
    .D(net1420),
    .Q_N(_3159_),
    .Q(\main.float_registers[3][29] ));
 sg13g2_dfrbp_1 _6674_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net143),
    .D(_0240_),
    .Q_N(_3271_),
    .Q(\main.float_registers[3][0] ));
 sg13g2_dfrbp_1 _6675_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net144),
    .D(_0006_),
    .Q_N(_3272_),
    .Q(\main.state[0] ));
 sg13g2_dfrbp_1 _6676_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net145),
    .D(_0007_),
    .Q_N(_3273_),
    .Q(\main.state[1] ));
 sg13g2_dfrbp_1 _6677_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net146),
    .D(net750),
    .Q_N(_3274_),
    .Q(\main.state[2] ));
 sg13g2_dfrbp_1 _6678_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net147),
    .D(net589),
    .Q_N(_3275_),
    .Q(\main.state[4] ));
 sg13g2_dfrbp_1 _6679_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net524),
    .D(net710),
    .Q_N(_3276_),
    .Q(\main.adder.in_valid ));
 sg13g2_dfrbp_1 _6680_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net110),
    .D(net852),
    .Q_N(_0031_),
    .Q(\main.state[6] ));
 sg13g2_dfrbp_1 _6681_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net109),
    .D(net1479),
    .Q_N(_0032_),
    .Q(\main.SPI_input_data_valid ));
 sg13g2_dfrbp_1 _6682_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net108),
    .D(_0242_),
    .Q_N(_3158_),
    .Q(\main.float_registers[3][5] ));
 sg13g2_dfrbp_1 _6683_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net107),
    .D(_0243_),
    .Q_N(_3157_),
    .Q(\main.float_registers[3][2] ));
 sg13g2_dfrbp_1 _6684_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net106),
    .D(_0244_),
    .Q_N(_3156_),
    .Q(\main.float_registers[3][21] ));
 sg13g2_dfrbp_1 _6685_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net105),
    .D(_0245_),
    .Q_N(_0076_),
    .Q(\main.adder.s3_exponent[0] ));
 sg13g2_dfrbp_1 _6686_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net104),
    .D(net738),
    .Q_N(_0075_),
    .Q(\main.adder.s3_exponent[1] ));
 sg13g2_dfrbp_1 _6687_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net103),
    .D(_0247_),
    .Q_N(_3155_),
    .Q(\main.adder.s3_exponent[2] ));
 sg13g2_dfrbp_1 _6688_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net102),
    .D(net602),
    .Q_N(_3154_),
    .Q(\main.adder.s3_exponent[3] ));
 sg13g2_dfrbp_1 _6689_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net101),
    .D(_0249_),
    .Q_N(_3153_),
    .Q(\main.adder.s3_exponent[4] ));
 sg13g2_dfrbp_1 _6690_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net100),
    .D(_0250_),
    .Q_N(_3152_),
    .Q(\main.adder.s3_exponent[5] ));
 sg13g2_dfrbp_1 _6691_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net99),
    .D(net789),
    .Q_N(_3151_),
    .Q(\main.adder.s3_exponent[6] ));
 sg13g2_dfrbp_1 _6692_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net98),
    .D(_0252_),
    .Q_N(_0074_),
    .Q(\main.adder.s3_exponent[7] ));
 sg13g2_dfrbp_1 _6693_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net97),
    .D(_0253_),
    .Q_N(_3150_),
    .Q(\main.adder.s4_exponent[0] ));
 sg13g2_dfrbp_1 _6694_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net96),
    .D(net995),
    .Q_N(_3149_),
    .Q(\main.adder.s4_exponent[1] ));
 sg13g2_dfrbp_1 _6695_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net95),
    .D(_0255_),
    .Q_N(_3148_),
    .Q(\main.adder.s4_exponent[2] ));
 sg13g2_dfrbp_1 _6696_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net94),
    .D(net810),
    .Q_N(_3147_),
    .Q(\main.adder.s4_exponent[3] ));
 sg13g2_dfrbp_1 _6697_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net93),
    .D(_0257_),
    .Q_N(_3146_),
    .Q(\main.adder.s4_exponent[4] ));
 sg13g2_dfrbp_1 _6698_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net92),
    .D(_0258_),
    .Q_N(_3145_),
    .Q(\main.adder.s4_exponent[5] ));
 sg13g2_dfrbp_1 _6699_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net91),
    .D(net952),
    .Q_N(_3144_),
    .Q(\main.adder.s4_exponent[6] ));
 sg13g2_dfrbp_1 _6700_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net90),
    .D(net1007),
    .Q_N(_3143_),
    .Q(\main.adder.s4_exponent[7] ));
 sg13g2_dfrbp_1 _6701_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net89),
    .D(net966),
    .Q_N(_3142_),
    .Q(\main.adder.out[1] ));
 sg13g2_dfrbp_1 _6702_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net87),
    .D(net909),
    .Q_N(_3141_),
    .Q(\main.adder.out[2] ));
 sg13g2_dfrbp_1 _6703_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net85),
    .D(net999),
    .Q_N(_3140_),
    .Q(\main.adder.out[3] ));
 sg13g2_dfrbp_1 _6704_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net83),
    .D(net1504),
    .Q_N(_3139_),
    .Q(\main.adder.out[4] ));
 sg13g2_dfrbp_1 _6705_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net81),
    .D(net921),
    .Q_N(_3138_),
    .Q(\main.adder.out[5] ));
 sg13g2_dfrbp_1 _6706_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net79),
    .D(net736),
    .Q_N(_3137_),
    .Q(\main.adder.out[6] ));
 sg13g2_dfrbp_1 _6707_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net77),
    .D(net704),
    .Q_N(_3136_),
    .Q(\main.adder.out[7] ));
 sg13g2_dfrbp_1 _6708_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net75),
    .D(net673),
    .Q_N(_3135_),
    .Q(\main.adder.out[8] ));
 sg13g2_dfrbp_1 _6709_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net73),
    .D(net775),
    .Q_N(_3134_),
    .Q(\main.adder.out[9] ));
 sg13g2_dfrbp_1 _6710_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net71),
    .D(net797),
    .Q_N(_3133_),
    .Q(\main.adder.out[10] ));
 sg13g2_dfrbp_1 _6711_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net69),
    .D(net894),
    .Q_N(_3132_),
    .Q(\main.adder.out[11] ));
 sg13g2_dfrbp_1 _6712_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net67),
    .D(net842),
    .Q_N(_3131_),
    .Q(\main.adder.out[12] ));
 sg13g2_dfrbp_1 _6713_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net65),
    .D(net838),
    .Q_N(_3130_),
    .Q(\main.adder.out[13] ));
 sg13g2_dfrbp_1 _6714_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net63),
    .D(net942),
    .Q_N(_3129_),
    .Q(\main.adder.out[14] ));
 sg13g2_dfrbp_1 _6715_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net61),
    .D(net755),
    .Q_N(_3128_),
    .Q(\main.adder.out[15] ));
 sg13g2_dfrbp_1 _6716_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net59),
    .D(net691),
    .Q_N(_3127_),
    .Q(\main.adder.out[16] ));
 sg13g2_dfrbp_1 _6717_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net57),
    .D(net684),
    .Q_N(_3126_),
    .Q(\main.adder.out[17] ));
 sg13g2_dfrbp_1 _6718_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net55),
    .D(net657),
    .Q_N(_3125_),
    .Q(\main.adder.out[18] ));
 sg13g2_dfrbp_1 _6719_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net53),
    .D(net654),
    .Q_N(_3124_),
    .Q(\main.adder.out[19] ));
 sg13g2_dfrbp_1 _6720_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net51),
    .D(net677),
    .Q_N(_3123_),
    .Q(\main.adder.out[20] ));
 sg13g2_dfrbp_1 _6721_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net49),
    .D(net675),
    .Q_N(_3122_),
    .Q(\main.adder.out[21] ));
 sg13g2_dfrbp_1 _6722_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net47),
    .D(net696),
    .Q_N(_3121_),
    .Q(\main.adder.out[22] ));
 sg13g2_dfrbp_1 _6723_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net45),
    .D(_0283_),
    .Q_N(_3120_),
    .Q(\main.adder.s5_mant[8] ));
 sg13g2_dfrbp_1 _6724_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net44),
    .D(_0284_),
    .Q_N(_3119_),
    .Q(\main.adder.s5_mant[9] ));
 sg13g2_dfrbp_1 _6725_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net43),
    .D(_0285_),
    .Q_N(_3118_),
    .Q(\main.adder.s5_mant[10] ));
 sg13g2_dfrbp_1 _6726_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net42),
    .D(_0286_),
    .Q_N(_3117_),
    .Q(\main.adder.s5_mant[11] ));
 sg13g2_dfrbp_1 _6727_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net41),
    .D(_0287_),
    .Q_N(_3116_),
    .Q(\main.adder.s5_mant[12] ));
 sg13g2_dfrbp_1 _6728_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net40),
    .D(_0288_),
    .Q_N(_3115_),
    .Q(\main.adder.s5_mant[13] ));
 sg13g2_dfrbp_1 _6729_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net39),
    .D(_0289_),
    .Q_N(_3114_),
    .Q(\main.adder.s5_mant[14] ));
 sg13g2_dfrbp_1 _6730_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net38),
    .D(_0290_),
    .Q_N(_3113_),
    .Q(\main.adder.s5_mant[15] ));
 sg13g2_dfrbp_1 _6731_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net37),
    .D(_0291_),
    .Q_N(_3112_),
    .Q(\main.adder.s5_mant[16] ));
 sg13g2_dfrbp_1 _6732_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net36),
    .D(_0292_),
    .Q_N(_3111_),
    .Q(\main.adder.s5_mant[17] ));
 sg13g2_dfrbp_1 _6733_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net35),
    .D(_0293_),
    .Q_N(_3110_),
    .Q(\main.adder.s5_mant[18] ));
 sg13g2_dfrbp_1 _6734_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net34),
    .D(_0294_),
    .Q_N(_3109_),
    .Q(\main.adder.s5_mant[19] ));
 sg13g2_dfrbp_1 _6735_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net33),
    .D(_0295_),
    .Q_N(_3108_),
    .Q(\main.adder.s5_mant[20] ));
 sg13g2_dfrbp_1 _6736_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net32),
    .D(_0296_),
    .Q_N(_3107_),
    .Q(\main.adder.s5_mant[21] ));
 sg13g2_dfrbp_1 _6737_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net31),
    .D(_0297_),
    .Q_N(_3106_),
    .Q(\main.adder.s5_mant[22] ));
 sg13g2_dfrbp_1 _6738_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net30),
    .D(_0298_),
    .Q_N(_3105_),
    .Q(\main.adder.s5_mant[23] ));
 sg13g2_dfrbp_1 _6739_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net29),
    .D(net729),
    .Q_N(_0103_),
    .Q(\main.adder.s2_larger[23] ));
 sg13g2_dfrbp_1 _6740_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net28),
    .D(net869),
    .Q_N(_0099_),
    .Q(\main.adder.s2_larger[24] ));
 sg13g2_dfrbp_1 _6741_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net27),
    .D(_0301_),
    .Q_N(_0101_),
    .Q(\main.adder.s2_larger[25] ));
 sg13g2_dfrbp_1 _6742_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net576),
    .D(net640),
    .Q_N(_0102_),
    .Q(\main.adder.s2_larger[26] ));
 sg13g2_dfrbp_1 _6743_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net575),
    .D(_0303_),
    .Q_N(_0104_),
    .Q(\main.adder.s2_larger[27] ));
 sg13g2_dfrbp_1 _6744_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net574),
    .D(net874),
    .Q_N(_0105_),
    .Q(\main.adder.s2_larger[28] ));
 sg13g2_dfrbp_1 _6745_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net573),
    .D(_0305_),
    .Q_N(_0106_),
    .Q(\main.adder.s2_larger[29] ));
 sg13g2_dfrbp_1 _6746_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net572),
    .D(net785),
    .Q_N(_0107_),
    .Q(\main.adder.s2_larger[30] ));
 sg13g2_dfrbp_1 _6747_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net571),
    .D(_0307_),
    .Q_N(_0108_),
    .Q(\main.adder.s2_larger[31] ));
 sg13g2_dfrbp_1 _6748_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net570),
    .D(_0308_),
    .Q_N(_0109_),
    .Q(\main.adder.s2_larger[32] ));
 sg13g2_dfrbp_1 _6749_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net569),
    .D(_0309_),
    .Q_N(_0110_),
    .Q(\main.adder.s2_larger[33] ));
 sg13g2_dfrbp_1 _6750_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net568),
    .D(_0310_),
    .Q_N(_0111_),
    .Q(\main.adder.s2_larger[34] ));
 sg13g2_dfrbp_1 _6751_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net567),
    .D(_0311_),
    .Q_N(_0112_),
    .Q(\main.adder.s2_larger[35] ));
 sg13g2_dfrbp_1 _6752_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net566),
    .D(_0312_),
    .Q_N(_0113_),
    .Q(\main.adder.s2_larger[36] ));
 sg13g2_dfrbp_1 _6753_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net565),
    .D(net699),
    .Q_N(_0114_),
    .Q(\main.adder.s2_larger[37] ));
 sg13g2_dfrbp_1 _6754_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net564),
    .D(net860),
    .Q_N(_0115_),
    .Q(\main.adder.s2_larger[38] ));
 sg13g2_dfrbp_1 _6755_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net563),
    .D(net747),
    .Q_N(_0116_),
    .Q(\main.adder.s2_larger[39] ));
 sg13g2_dfrbp_1 _6756_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net562),
    .D(net1423),
    .Q_N(_0117_),
    .Q(\main.adder.s2_larger[40] ));
 sg13g2_dfrbp_1 _6757_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net561),
    .D(net902),
    .Q_N(_0118_),
    .Q(\main.adder.s2_larger[41] ));
 sg13g2_dfrbp_1 _6758_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net560),
    .D(_0318_),
    .Q_N(_0119_),
    .Q(\main.adder.s2_larger[42] ));
 sg13g2_dfrbp_1 _6759_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net559),
    .D(net976),
    .Q_N(_0120_),
    .Q(\main.adder.s2_larger[43] ));
 sg13g2_dfrbp_1 _6760_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net558),
    .D(net724),
    .Q_N(_0121_),
    .Q(\main.adder.s2_larger[44] ));
 sg13g2_dfrbp_1 _6761_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net557),
    .D(_0321_),
    .Q_N(_0122_),
    .Q(\main.adder.s2_larger[45] ));
 sg13g2_dfrbp_1 _6762_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net556),
    .D(_0322_),
    .Q_N(_0123_),
    .Q(\main.adder.s2_larger[46] ));
 sg13g2_dfrbp_1 _6763_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net555),
    .D(_0323_),
    .Q_N(_3104_),
    .Q(\main.adder.s2_smaler[15] ));
 sg13g2_dfrbp_1 _6764_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net553),
    .D(_0324_),
    .Q_N(_3103_),
    .Q(\main.adder.s2_smaler[16] ));
 sg13g2_dfrbp_1 _6765_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net551),
    .D(_0325_),
    .Q_N(_3102_),
    .Q(\main.adder.s2_smaler[17] ));
 sg13g2_dfrbp_1 _6766_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net549),
    .D(_0326_),
    .Q_N(_3101_),
    .Q(\main.adder.s2_smaler[18] ));
 sg13g2_dfrbp_1 _6767_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net547),
    .D(_0327_),
    .Q_N(_3100_),
    .Q(\main.adder.s2_smaler[19] ));
 sg13g2_dfrbp_1 _6768_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net545),
    .D(_0328_),
    .Q_N(_3099_),
    .Q(\main.adder.s2_smaler[20] ));
 sg13g2_dfrbp_1 _6769_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net543),
    .D(_0329_),
    .Q_N(_3098_),
    .Q(\main.adder.s2_smaler[21] ));
 sg13g2_dfrbp_1 _6770_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net541),
    .D(_0330_),
    .Q_N(_3097_),
    .Q(\main.adder.s2_smaler[22] ));
 sg13g2_dfrbp_1 _6771_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net539),
    .D(_0331_),
    .Q_N(_3096_),
    .Q(\main.adder.s2_smaler[23] ));
 sg13g2_dfrbp_1 _6772_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net537),
    .D(_0332_),
    .Q_N(_3095_),
    .Q(\main.adder.s2_smaler[24] ));
 sg13g2_dfrbp_1 _6773_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net535),
    .D(_0333_),
    .Q_N(_3094_),
    .Q(\main.adder.s2_smaler[25] ));
 sg13g2_dfrbp_1 _6774_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net533),
    .D(_0334_),
    .Q_N(_3093_),
    .Q(\main.adder.s2_smaler[26] ));
 sg13g2_dfrbp_1 _6775_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net531),
    .D(_0335_),
    .Q_N(_3092_),
    .Q(\main.adder.s2_smaler[27] ));
 sg13g2_dfrbp_1 _6776_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net523),
    .D(_0336_),
    .Q_N(_3091_),
    .Q(\main.adder.s2_smaler[28] ));
 sg13g2_dfrbp_1 _6777_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net521),
    .D(_0337_),
    .Q_N(_3090_),
    .Q(\main.adder.s2_smaler[29] ));
 sg13g2_dfrbp_1 _6778_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net519),
    .D(_0338_),
    .Q_N(_3089_),
    .Q(\main.adder.s2_smaler[30] ));
 sg13g2_dfrbp_1 _6779_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net517),
    .D(_0339_),
    .Q_N(_3088_),
    .Q(\main.adder.s2_smaler[32] ));
 sg13g2_dfrbp_1 _6780_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net515),
    .D(_0340_),
    .Q_N(_3087_),
    .Q(\main.adder.s2_smaler[33] ));
 sg13g2_dfrbp_1 _6781_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net513),
    .D(_0341_),
    .Q_N(_3086_),
    .Q(\main.adder.s2_smaler[34] ));
 sg13g2_dfrbp_1 _6782_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net511),
    .D(_0342_),
    .Q_N(_3085_),
    .Q(\main.adder.s2_smaler[35] ));
 sg13g2_dfrbp_1 _6783_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net509),
    .D(_0343_),
    .Q_N(_3084_),
    .Q(\main.adder.s2_smaler[36] ));
 sg13g2_dfrbp_1 _6784_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net507),
    .D(_0344_),
    .Q_N(_3083_),
    .Q(\main.adder.s2_smaler[37] ));
 sg13g2_dfrbp_1 _6785_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net505),
    .D(_0345_),
    .Q_N(_3082_),
    .Q(\main.adder.s2_smaler[38] ));
 sg13g2_dfrbp_1 _6786_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net503),
    .D(_0346_),
    .Q_N(_3081_),
    .Q(\main.adder.s2_smaler[39] ));
 sg13g2_dfrbp_1 _6787_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net501),
    .D(_0347_),
    .Q_N(_3080_),
    .Q(\main.adder.s2_smaler[40] ));
 sg13g2_dfrbp_1 _6788_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net499),
    .D(_0348_),
    .Q_N(_3079_),
    .Q(\main.adder.s2_smaler[41] ));
 sg13g2_dfrbp_1 _6789_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net497),
    .D(_0349_),
    .Q_N(_3078_),
    .Q(\main.adder.s2_smaler[42] ));
 sg13g2_dfrbp_1 _6790_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net495),
    .D(_0350_),
    .Q_N(_3077_),
    .Q(\main.adder.s2_smaler[43] ));
 sg13g2_dfrbp_1 _6791_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net493),
    .D(_0351_),
    .Q_N(_3076_),
    .Q(\main.adder.s2_smaler[44] ));
 sg13g2_dfrbp_1 _6792_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net491),
    .D(_0352_),
    .Q_N(_3075_),
    .Q(\main.adder.s2_smaler[45] ));
 sg13g2_dfrbp_1 _6793_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net489),
    .D(net960),
    .Q_N(_3074_),
    .Q(\main.adder.s2_smaler[46] ));
 sg13g2_dfrbp_1 _6794_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net487),
    .D(_0354_),
    .Q_N(_3073_),
    .Q(\main.float_registers[3][19] ));
 sg13g2_dfrbp_1 _6795_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net486),
    .D(_0355_),
    .Q_N(_3072_),
    .Q(\main.float_registers[3][28] ));
 sg13g2_dfrbp_1 _6796_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net485),
    .D(_0356_),
    .Q_N(_3071_),
    .Q(\main.float_registers[3][1] ));
 sg13g2_dfrbp_1 _6797_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net484),
    .D(_0357_),
    .Q_N(_3070_),
    .Q(\main.float_registers[3][20] ));
 sg13g2_dfrbp_1 _6798_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net483),
    .D(_0358_),
    .Q_N(_3069_),
    .Q(\main.float_registers[3][12] ));
 sg13g2_dfrbp_1 _6799_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net482),
    .D(_0359_),
    .Q_N(_3068_),
    .Q(\main.float_registers[3][18] ));
 sg13g2_dfrbp_1 _6800_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net481),
    .D(_0360_),
    .Q_N(_3067_),
    .Q(\main.float_registers[3][13] ));
 sg13g2_dfrbp_1 _6801_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net480),
    .D(_0361_),
    .Q_N(_3066_),
    .Q(_0004_));
 sg13g2_dfrbp_1 _6802_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net479),
    .D(_0362_),
    .Q_N(_3065_),
    .Q(_0005_));
 sg13g2_dfrbp_1 _6803_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net478),
    .D(net1470),
    .Q_N(_3064_),
    .Q(\main.float_registers[3][10] ));
 sg13g2_dfrbp_1 _6804_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net477),
    .D(_0364_),
    .Q_N(_3063_),
    .Q(\main.float_registers[3][6] ));
 sg13g2_dfrbp_1 _6805_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net476),
    .D(_0365_),
    .Q_N(_3062_),
    .Q(\main.adder.out_valid ));
 sg13g2_dfrbp_1 _6806_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net475),
    .D(_0366_),
    .Q_N(_3061_),
    .Q(\main.adder.out[0] ));
 sg13g2_dfrbp_1 _6807_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net473),
    .D(net947),
    .Q_N(_3060_),
    .Q(\main.adder.out[23] ));
 sg13g2_dfrbp_1 _6808_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net471),
    .D(net887),
    .Q_N(_3059_),
    .Q(\main.adder.out[24] ));
 sg13g2_dfrbp_1 _6809_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net469),
    .D(net759),
    .Q_N(_3058_),
    .Q(\main.adder.out[25] ));
 sg13g2_dfrbp_1 _6810_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net467),
    .D(net1023),
    .Q_N(_3057_),
    .Q(\main.adder.out[26] ));
 sg13g2_dfrbp_1 _6811_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net465),
    .D(net1005),
    .Q_N(_3056_),
    .Q(\main.adder.out[27] ));
 sg13g2_dfrbp_1 _6812_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net463),
    .D(net917),
    .Q_N(_3055_),
    .Q(\main.adder.out[28] ));
 sg13g2_dfrbp_1 _6813_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net461),
    .D(net1399),
    .Q_N(_3054_),
    .Q(\main.adder.out[29] ));
 sg13g2_dfrbp_1 _6814_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net459),
    .D(net969),
    .Q_N(_3053_),
    .Q(\main.adder.out[30] ));
 sg13g2_dfrbp_1 _6815_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net457),
    .D(net632),
    .Q_N(_3052_),
    .Q(\main.adder.out[31] ));
 sg13g2_dfrbp_1 _6816_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net456),
    .D(_0376_),
    .Q_N(_3051_),
    .Q(\main.adder.s5_valid ));
 sg13g2_dfrbp_1 _6817_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net455),
    .D(_0377_),
    .Q_N(_3050_),
    .Q(\main.adder.s5_mant[0] ));
 sg13g2_dfrbp_1 _6818_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net453),
    .D(_0378_),
    .Q_N(_3049_),
    .Q(\main.adder.s5_mant[1] ));
 sg13g2_dfrbp_1 _6819_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net451),
    .D(_0379_),
    .Q_N(_3048_),
    .Q(\main.adder.s5_mant[2] ));
 sg13g2_dfrbp_1 _6820_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net449),
    .D(_0380_),
    .Q_N(_3047_),
    .Q(\main.adder.s5_mant[3] ));
 sg13g2_dfrbp_1 _6821_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net447),
    .D(_0381_),
    .Q_N(_3046_),
    .Q(\main.adder.s5_mant[4] ));
 sg13g2_dfrbp_1 _6822_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net445),
    .D(_0382_),
    .Q_N(_3045_),
    .Q(\main.adder.s5_mant[5] ));
 sg13g2_dfrbp_1 _6823_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net443),
    .D(_0383_),
    .Q_N(_3044_),
    .Q(\main.adder.s5_mant[6] ));
 sg13g2_dfrbp_1 _6824_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net441),
    .D(_0384_),
    .Q_N(_3043_),
    .Q(\main.adder.s5_mant[7] ));
 sg13g2_dfrbp_1 _6825_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net439),
    .D(_0385_),
    .Q_N(_0033_),
    .Q(\main.adder.s5_R ));
 sg13g2_dfrbp_1 _6826_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net437),
    .D(_0386_),
    .Q_N(_3042_),
    .Q(\main.adder.s5_sign ));
 sg13g2_dfrbp_1 _6827_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net436),
    .D(_0387_),
    .Q_N(_3041_),
    .Q(\main.adder.s5_S ));
 sg13g2_dfrbp_1 _6828_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net435),
    .D(_0388_),
    .Q_N(_3040_),
    .Q(\main.adder.s5_nan ));
 sg13g2_dfrbp_1 _6829_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net434),
    .D(_0389_),
    .Q_N(_3039_),
    .Q(\main.adder.s5_inf ));
 sg13g2_dfrbp_1 _6830_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net433),
    .D(_0390_),
    .Q_N(_0034_),
    .Q(\main.adder.s5_exponent[0] ));
 sg13g2_dfrbp_1 _6831_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net432),
    .D(_0391_),
    .Q_N(_0035_),
    .Q(\main.adder.s5_exponent[1] ));
 sg13g2_dfrbp_1 _6832_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net431),
    .D(_0392_),
    .Q_N(_0036_),
    .Q(\main.adder.s5_exponent[2] ));
 sg13g2_dfrbp_1 _6833_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net430),
    .D(_0393_),
    .Q_N(_0037_),
    .Q(\main.adder.s5_exponent[3] ));
 sg13g2_dfrbp_1 _6834_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net429),
    .D(_0394_),
    .Q_N(_0038_),
    .Q(\main.adder.s5_exponent[4] ));
 sg13g2_dfrbp_1 _6835_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net428),
    .D(_0395_),
    .Q_N(_0039_),
    .Q(\main.adder.s5_exponent[5] ));
 sg13g2_dfrbp_1 _6836_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net427),
    .D(_0396_),
    .Q_N(_0040_),
    .Q(\main.adder.s5_exponent[6] ));
 sg13g2_dfrbp_1 _6837_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net426),
    .D(_0397_),
    .Q_N(_0041_),
    .Q(\main.adder.s5_exponent[7] ));
 sg13g2_dfrbp_1 _6838_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net425),
    .D(net1402),
    .Q_N(_3038_),
    .Q(\main.adder.s5_exponent[8] ));
 sg13g2_dfrbp_1 _6839_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net424),
    .D(_0399_),
    .Q_N(_3037_),
    .Q(\main.adder.s5_exponent[9] ));
 sg13g2_dfrbp_1 _6840_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net423),
    .D(_0400_),
    .Q_N(_3036_),
    .Q(\main.adder.s4_valid ));
 sg13g2_dfrbp_1 _6841_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net422),
    .D(net719),
    .Q_N(_3035_),
    .Q(\main.adder.s4_flipped ));
 sg13g2_dfrbp_1 _6842_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net421),
    .D(_0402_),
    .Q_N(_3034_),
    .Q(\main.adder.s4_shared_sign ));
 sg13g2_dfrbp_1 _6843_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net420),
    .D(net781),
    .Q_N(_3033_),
    .Q(\main.adder.s4_nan ));
 sg13g2_dfrbp_1 _6844_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net419),
    .D(_0404_),
    .Q_N(_3032_),
    .Q(\main.adder.s4_inf ));
 sg13g2_dfrbp_1 _6845_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net418),
    .D(net610),
    .Q_N(_0043_),
    .Q(\main.adder.s4_mant[1] ));
 sg13g2_dfrbp_1 _6846_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net417),
    .D(net636),
    .Q_N(_0044_),
    .Q(\main.adder.s4_mant[2] ));
 sg13g2_dfrbp_1 _6847_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net416),
    .D(net614),
    .Q_N(_0045_),
    .Q(\main.adder.s4_mant[3] ));
 sg13g2_dfrbp_1 _6848_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net415),
    .D(net667),
    .Q_N(_0046_),
    .Q(\main.adder.s4_mant[4] ));
 sg13g2_dfrbp_1 _6849_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net414),
    .D(net606),
    .Q_N(_0047_),
    .Q(\main.adder.s4_mant[5] ));
 sg13g2_dfrbp_1 _6850_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net413),
    .D(net598),
    .Q_N(_0048_),
    .Q(\main.adder.s4_mant[6] ));
 sg13g2_dfrbp_1 _6851_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net412),
    .D(net663),
    .Q_N(_0049_),
    .Q(\main.adder.s4_mant[7] ));
 sg13g2_dfrbp_1 _6852_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net411),
    .D(net587),
    .Q_N(_0050_),
    .Q(\main.adder.s4_mant[8] ));
 sg13g2_dfrbp_1 _6853_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net410),
    .D(net594),
    .Q_N(_0051_),
    .Q(\main.adder.s4_mant[9] ));
 sg13g2_dfrbp_1 _6854_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net409),
    .D(net596),
    .Q_N(_0052_),
    .Q(\main.adder.s4_mant[10] ));
 sg13g2_dfrbp_1 _6855_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net408),
    .D(net622),
    .Q_N(_0053_),
    .Q(\main.adder.s4_mant[11] ));
 sg13g2_dfrbp_1 _6856_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net407),
    .D(_0416_),
    .Q_N(_0054_),
    .Q(\main.adder.s4_mant[12] ));
 sg13g2_dfrbp_1 _6857_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net406),
    .D(net612),
    .Q_N(_0055_),
    .Q(\main.adder.s4_mant[13] ));
 sg13g2_dfrbp_1 _6858_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net405),
    .D(_0418_),
    .Q_N(_0056_),
    .Q(\main.adder.s4_mant[14] ));
 sg13g2_dfrbp_1 _6859_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net404),
    .D(net626),
    .Q_N(_0057_),
    .Q(\main.adder.s4_mant[15] ));
 sg13g2_dfrbp_1 _6860_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net403),
    .D(net604),
    .Q_N(_0058_),
    .Q(\main.adder.s4_mant[16] ));
 sg13g2_dfrbp_1 _6861_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net402),
    .D(net591),
    .Q_N(_0059_),
    .Q(\main.adder.s4_mant[17] ));
 sg13g2_dfrbp_1 _6862_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net401),
    .D(net600),
    .Q_N(_0060_),
    .Q(\main.adder.s4_mant[18] ));
 sg13g2_dfrbp_1 _6863_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net400),
    .D(net608),
    .Q_N(_0061_),
    .Q(\main.adder.s4_mant[19] ));
 sg13g2_dfrbp_1 _6864_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net399),
    .D(net618),
    .Q_N(_0062_),
    .Q(\main.adder.s4_mant[20] ));
 sg13g2_dfrbp_1 _6865_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net398),
    .D(net800),
    .Q_N(_0063_),
    .Q(\main.adder.s4_mant[21] ));
 sg13g2_dfrbp_1 _6866_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net397),
    .D(net1541),
    .Q_N(_3031_),
    .Q(\main.adder.s4_mant[22] ));
 sg13g2_dfrbp_1 _6867_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net396),
    .D(net1500),
    .Q_N(_3030_),
    .Q(\main.adder.s4_mant[23] ));
 sg13g2_dfrbp_1 _6868_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net395),
    .D(net1563),
    .Q_N(_3029_),
    .Q(\main.adder.s4_mant[24] ));
 sg13g2_dfrbp_1 _6869_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net394),
    .D(net1565),
    .Q_N(_3028_),
    .Q(\main.adder.s4_mant[25] ));
 sg13g2_dfrbp_1 _6870_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net393),
    .D(net1518),
    .Q_N(_3027_),
    .Q(\main.adder.s4_mant[26] ));
 sg13g2_dfrbp_1 _6871_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net392),
    .D(net1468),
    .Q_N(_3026_),
    .Q(\main.adder.s4_mant[27] ));
 sg13g2_dfrbp_1 _6872_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net391),
    .D(net1510),
    .Q_N(_3025_),
    .Q(\main.adder.s4_mant[28] ));
 sg13g2_dfrbp_1 _6873_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net390),
    .D(net1445),
    .Q_N(_3024_),
    .Q(\main.adder.s4_mant[29] ));
 sg13g2_dfrbp_1 _6874_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net389),
    .D(net825),
    .Q_N(_3023_),
    .Q(\main.adder.s4_mant[30] ));
 sg13g2_dfrbp_1 _6875_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net388),
    .D(net1465),
    .Q_N(_3022_),
    .Q(\main.adder.s4_mant[31] ));
 sg13g2_dfrbp_1 _6876_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net387),
    .D(net936),
    .Q_N(_3021_),
    .Q(\main.adder.s4_mant[32] ));
 sg13g2_dfrbp_1 _6877_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net386),
    .D(net1404),
    .Q_N(_3020_),
    .Q(\main.adder.s4_mant[33] ));
 sg13g2_dfrbp_1 _6878_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net385),
    .D(_0438_),
    .Q_N(_3019_),
    .Q(\main.adder.s4_mant[34] ));
 sg13g2_dfrbp_1 _6879_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net384),
    .D(_0439_),
    .Q_N(_3018_),
    .Q(\main.adder.s4_mant[35] ));
 sg13g2_dfrbp_1 _6880_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net383),
    .D(_0440_),
    .Q_N(_3017_),
    .Q(\main.adder.s4_mant[36] ));
 sg13g2_dfrbp_1 _6881_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net382),
    .D(_0441_),
    .Q_N(_3016_),
    .Q(\main.adder.s4_mant[37] ));
 sg13g2_dfrbp_1 _6882_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net381),
    .D(_0442_),
    .Q_N(_3015_),
    .Q(\main.adder.s4_mant[38] ));
 sg13g2_dfrbp_1 _6883_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net380),
    .D(_0443_),
    .Q_N(_3014_),
    .Q(\main.adder.s4_mant[39] ));
 sg13g2_dfrbp_1 _6884_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net379),
    .D(_0444_),
    .Q_N(_3013_),
    .Q(\main.adder.s4_mant[40] ));
 sg13g2_dfrbp_1 _6885_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net378),
    .D(_0445_),
    .Q_N(_3012_),
    .Q(\main.adder.s4_mant[41] ));
 sg13g2_dfrbp_1 _6886_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net377),
    .D(net939),
    .Q_N(_3011_),
    .Q(\main.adder.s4_mant[42] ));
 sg13g2_dfrbp_1 _6887_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net376),
    .D(_0447_),
    .Q_N(_3010_),
    .Q(\main.adder.s4_mant[43] ));
 sg13g2_dfrbp_1 _6888_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net375),
    .D(net955),
    .Q_N(_3009_),
    .Q(\main.adder.s4_mant[44] ));
 sg13g2_dfrbp_1 _6889_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net374),
    .D(net1473),
    .Q_N(_3008_),
    .Q(\main.adder.s4_mant[45] ));
 sg13g2_dfrbp_1 _6890_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net373),
    .D(net1416),
    .Q_N(_3007_),
    .Q(\main.adder.s4_mant[46] ));
 sg13g2_dfrbp_1 _6891_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net372),
    .D(net981),
    .Q_N(_3006_),
    .Q(\main.adder.s4_mant[47] ));
 sg13g2_dfrbp_1 _6892_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net371),
    .D(net634),
    .Q_N(_0042_),
    .Q(\main.adder.s4_mant[0] ));
 sg13g2_dfrbp_1 _6893_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net370),
    .D(net661),
    .Q_N(_3005_),
    .Q(\main.adder.s4_sum[48] ));
 sg13g2_dfrbp_1 _6894_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net369),
    .D(_0454_),
    .Q_N(_3004_),
    .Q(\main.adder.s3_valid ));
 sg13g2_dfrbp_1 _6895_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net368),
    .D(net783),
    .Q_N(_3003_),
    .Q(\main.adder.s3_nan ));
 sg13g2_dfrbp_1 _6896_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net367),
    .D(_0456_),
    .Q_N(_3002_),
    .Q(\main.adder.s3_inf ));
 sg13g2_dfrbp_1 _6897_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net366),
    .D(_0457_),
    .Q_N(_3001_),
    .Q(\main.adder.s3_flipped ));
 sg13g2_dfrbp_1 _6898_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net365),
    .D(net727),
    .Q_N(_3000_),
    .Q(\main.adder.s3_shared_sign ));
 sg13g2_dfrbp_1 _6899_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net364),
    .D(_0459_),
    .Q_N(_2999_),
    .Q(\main.adder.s3_sum[0] ));
 sg13g2_dfrbp_1 _6900_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net363),
    .D(_0460_),
    .Q_N(_0065_),
    .Q(\main.adder.s3_sum[1] ));
 sg13g2_dfrbp_1 _6901_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net362),
    .D(_0461_),
    .Q_N(_2998_),
    .Q(\main.adder.s3_sum[2] ));
 sg13g2_dfrbp_1 _6902_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net361),
    .D(net930),
    .Q_N(_0066_),
    .Q(\main.adder.s3_sum[3] ));
 sg13g2_dfrbp_1 _6903_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net360),
    .D(_0463_),
    .Q_N(_2997_),
    .Q(\main.adder.s3_sum[4] ));
 sg13g2_dfrbp_1 _6904_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net359),
    .D(_0464_),
    .Q_N(_0067_),
    .Q(\main.adder.s3_sum[5] ));
 sg13g2_dfrbp_1 _6905_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net358),
    .D(net731),
    .Q_N(_2996_),
    .Q(\main.adder.s3_sum[6] ));
 sg13g2_dfrbp_1 _6906_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net357),
    .D(net708),
    .Q_N(_0068_),
    .Q(\main.adder.s3_sum[7] ));
 sg13g2_dfrbp_1 _6907_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net356),
    .D(_0467_),
    .Q_N(_2995_),
    .Q(\main.adder.s3_sum[8] ));
 sg13g2_dfrbp_1 _6908_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net355),
    .D(_0468_),
    .Q_N(_0069_),
    .Q(\main.adder.s3_sum[9] ));
 sg13g2_dfrbp_1 _6909_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net354),
    .D(_0469_),
    .Q_N(_2994_),
    .Q(\main.adder.s3_sum[10] ));
 sg13g2_dfrbp_1 _6910_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net353),
    .D(net1397),
    .Q_N(_0070_),
    .Q(\main.adder.s3_sum[11] ));
 sg13g2_dfrbp_1 _6911_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net352),
    .D(net706),
    .Q_N(_2993_),
    .Q(\main.adder.s3_sum[12] ));
 sg13g2_dfrbp_1 _6912_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net351),
    .D(net884),
    .Q_N(_0071_),
    .Q(\main.adder.s3_sum[13] ));
 sg13g2_dfrbp_1 _6913_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net350),
    .D(net865),
    .Q_N(_2992_),
    .Q(\main.adder.s3_sum[14] ));
 sg13g2_dfrbp_1 _6914_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net349),
    .D(net928),
    .Q_N(_0072_),
    .Q(\main.adder.s3_sum[15] ));
 sg13g2_dfrbp_1 _6915_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net348),
    .D(net907),
    .Q_N(_2991_),
    .Q(\main.adder.s3_sum[16] ));
 sg13g2_dfrbp_1 _6916_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net347),
    .D(net1021),
    .Q_N(_0016_),
    .Q(\main.adder.s3_sum[17] ));
 sg13g2_dfrbp_1 _6917_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net346),
    .D(net983),
    .Q_N(_0017_),
    .Q(\main.adder.s3_sum[18] ));
 sg13g2_dfrbp_1 _6918_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net345),
    .D(_0478_),
    .Q_N(_0018_),
    .Q(\main.adder.s3_sum[19] ));
 sg13g2_dfrbp_1 _6919_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net344),
    .D(net1567),
    .Q_N(_0019_),
    .Q(\main.adder.s3_sum[20] ));
 sg13g2_dfrbp_1 _6920_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net343),
    .D(_0480_),
    .Q_N(_0020_),
    .Q(\main.adder.s3_sum[21] ));
 sg13g2_dfrbp_1 _6921_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net342),
    .D(_0481_),
    .Q_N(_0021_),
    .Q(\main.adder.s3_sum[22] ));
 sg13g2_dfrbp_1 _6922_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net341),
    .D(net905),
    .Q_N(_0022_),
    .Q(\main.adder.s3_sum[23] ));
 sg13g2_dfrbp_1 _6923_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net340),
    .D(_0483_),
    .Q_N(_0023_),
    .Q(\main.adder.s3_sum[24] ));
 sg13g2_dfrbp_1 _6924_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net339),
    .D(_0484_),
    .Q_N(_0024_),
    .Q(\main.adder.s3_sum[25] ));
 sg13g2_dfrbp_1 _6925_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net338),
    .D(_0485_),
    .Q_N(_0025_),
    .Q(\main.adder.s3_sum[26] ));
 sg13g2_dfrbp_1 _6926_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net337),
    .D(_0486_),
    .Q_N(_0026_),
    .Q(\main.adder.s3_sum[27] ));
 sg13g2_dfrbp_1 _6927_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net336),
    .D(_0487_),
    .Q_N(_0027_),
    .Q(\main.adder.s3_sum[28] ));
 sg13g2_dfrbp_1 _6928_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net335),
    .D(_0488_),
    .Q_N(_0028_),
    .Q(\main.adder.s3_sum[29] ));
 sg13g2_dfrbp_1 _6929_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net334),
    .D(_0489_),
    .Q_N(_0029_),
    .Q(\main.adder.s3_sum[30] ));
 sg13g2_dfrbp_1 _6930_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net333),
    .D(_0490_),
    .Q_N(_0030_),
    .Q(\main.adder.s3_sum[31] ));
 sg13g2_dfrbp_1 _6931_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net332),
    .D(net1579),
    .Q_N(_2990_),
    .Q(\main.adder.s3_sum[32] ));
 sg13g2_dfrbp_1 _6932_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net331),
    .D(_0492_),
    .Q_N(_2989_),
    .Q(\main.adder.s3_sum[33] ));
 sg13g2_dfrbp_1 _6933_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net330),
    .D(_0493_),
    .Q_N(_2988_),
    .Q(\main.adder.s3_sum[34] ));
 sg13g2_dfrbp_1 _6934_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net329),
    .D(_0494_),
    .Q_N(_2987_),
    .Q(\main.adder.s3_sum[35] ));
 sg13g2_dfrbp_1 _6935_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net328),
    .D(_0495_),
    .Q_N(_2986_),
    .Q(\main.adder.s3_sum[36] ));
 sg13g2_dfrbp_1 _6936_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net327),
    .D(_0496_),
    .Q_N(_2985_),
    .Q(\main.adder.s3_sum[37] ));
 sg13g2_dfrbp_1 _6937_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net326),
    .D(_0497_),
    .Q_N(_2984_),
    .Q(\main.adder.s3_sum[38] ));
 sg13g2_dfrbp_1 _6938_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net325),
    .D(_0498_),
    .Q_N(_2983_),
    .Q(\main.adder.s3_sum[39] ));
 sg13g2_dfrbp_1 _6939_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net324),
    .D(_0499_),
    .Q_N(_2982_),
    .Q(\main.adder.s3_sum[40] ));
 sg13g2_dfrbp_1 _6940_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net323),
    .D(_0500_),
    .Q_N(_2981_),
    .Q(\main.adder.s3_sum[41] ));
 sg13g2_dfrbp_1 _6941_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net321),
    .D(_0501_),
    .Q_N(_2980_),
    .Q(\main.adder.s3_sum[42] ));
 sg13g2_dfrbp_1 _6942_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net319),
    .D(_0502_),
    .Q_N(_2979_),
    .Q(\main.adder.s3_sum[43] ));
 sg13g2_dfrbp_1 _6943_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net314),
    .D(net1589),
    .Q_N(_2978_),
    .Q(\main.adder.s3_sum[44] ));
 sg13g2_dfrbp_1 _6944_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net312),
    .D(_0504_),
    .Q_N(_2977_),
    .Q(\main.adder.s3_sum[45] ));
 sg13g2_dfrbp_1 _6945_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net310),
    .D(net1535),
    .Q_N(_2976_),
    .Q(\main.adder.s3_sum[46] ));
 sg13g2_dfrbp_1 _6946_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net308),
    .D(net1604),
    .Q_N(_2975_),
    .Q(\main.adder.s3_sum[47] ));
 sg13g2_dfrbp_1 _6947_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net306),
    .D(_0507_),
    .Q_N(_0015_),
    .Q(\main.adder.s3_sum[48] ));
 sg13g2_dfrbp_1 _6948_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net304),
    .D(_0508_),
    .Q_N(_2974_),
    .Q(\main.adder.s2_valid ));
 sg13g2_dfrbp_1 _6949_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net302),
    .D(_0509_),
    .Q_N(_0100_),
    .Q(\main.adder.s2_flip_sign ));
 sg13g2_dfrbp_1 _6950_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net300),
    .D(net721),
    .Q_N(_2973_),
    .Q(\main.adder.s2_nan ));
 sg13g2_dfrbp_1 _6951_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net298),
    .D(net757),
    .Q_N(_2972_),
    .Q(\main.adder.s2_inf ));
 sg13g2_dfrbp_1 _6952_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net296),
    .D(_0512_),
    .Q_N(_2971_),
    .Q(\main.adder.s2_smaler[31] ));
 sg13g2_dfrbp_1 _6953_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net292),
    .D(_0513_),
    .Q_N(_2970_),
    .Q(\main.adder.s2_shared_sign ));
 sg13g2_dfrbp_1 _6954_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net290),
    .D(net772),
    .Q_N(_2969_),
    .Q(\main.adder.s2_exponent[0] ));
 sg13g2_dfrbp_1 _6955_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net288),
    .D(_0515_),
    .Q_N(_2968_),
    .Q(\main.adder.s2_exponent[1] ));
 sg13g2_dfrbp_1 _6956_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net286),
    .D(net766),
    .Q_N(_2967_),
    .Q(\main.adder.s2_exponent[2] ));
 sg13g2_dfrbp_1 _6957_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net284),
    .D(_0517_),
    .Q_N(_2966_),
    .Q(\main.adder.s2_exponent[3] ));
 sg13g2_dfrbp_1 _6958_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net282),
    .D(net823),
    .Q_N(_2965_),
    .Q(\main.adder.s2_exponent[4] ));
 sg13g2_dfrbp_1 _6959_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net280),
    .D(net923),
    .Q_N(_2964_),
    .Q(\main.adder.s2_exponent[5] ));
 sg13g2_dfrbp_1 _6960_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net278),
    .D(_0520_),
    .Q_N(_2963_),
    .Q(\main.adder.s2_exponent[6] ));
 sg13g2_dfrbp_1 _6961_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net276),
    .D(net820),
    .Q_N(_2962_),
    .Q(\main.adder.s2_exponent[7] ));
 sg13g2_dfrbp_1 _6962_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net274),
    .D(net578),
    .Q_N(_2961_),
    .Q(\main.spi.state[0] ));
 sg13g2_dfrbp_1 _6963_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net270),
    .D(_0523_),
    .Q_N(_2960_),
    .Q(\main.adder.s1_valid ));
 sg13g2_dfrbp_1 _6964_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net268),
    .D(_0524_),
    .Q_N(_2959_),
    .Q(\main.adder.s1_nan ));
 sg13g2_dfrbp_1 _6965_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net266),
    .D(_0525_),
    .Q_N(_2958_),
    .Q(\main.adder.s1_inf ));
 sg13g2_dfrbp_1 _6966_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net264),
    .D(_0526_),
    .Q_N(_2957_),
    .Q(\main.adder.s1_rs.levels[0][23] ));
 sg13g2_dfrbp_1 _6967_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net262),
    .D(_0527_),
    .Q_N(_0078_),
    .Q(\main.adder.s1_rs.levels[0][24] ));
 sg13g2_dfrbp_1 _6968_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net260),
    .D(_0528_),
    .Q_N(_0077_),
    .Q(\main.adder.s1_rs.levels[0][25] ));
 sg13g2_dfrbp_1 _6969_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net258),
    .D(_0529_),
    .Q_N(_0080_),
    .Q(\main.adder.s1_rs.levels[0][26] ));
 sg13g2_dfrbp_1 _6970_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net256),
    .D(_0530_),
    .Q_N(_0079_),
    .Q(\main.adder.s1_rs.levels[0][27] ));
 sg13g2_dfrbp_1 _6971_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net254),
    .D(_0531_),
    .Q_N(_0082_),
    .Q(\main.adder.s1_rs.levels[0][28] ));
 sg13g2_dfrbp_1 _6972_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net252),
    .D(_0532_),
    .Q_N(_0081_),
    .Q(\main.adder.s1_rs.levels[0][29] ));
 sg13g2_dfrbp_1 _6973_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net250),
    .D(_0533_),
    .Q_N(_0084_),
    .Q(\main.adder.s1_rs.levels[0][30] ));
 sg13g2_dfrbp_1 _6974_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net248),
    .D(_0534_),
    .Q_N(_0083_),
    .Q(\main.adder.s1_rs.levels[0][31] ));
 sg13g2_dfrbp_1 _6975_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net246),
    .D(_0535_),
    .Q_N(_0086_),
    .Q(\main.adder.s1_rs.levels[0][32] ));
 sg13g2_dfrbp_1 _6976_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net244),
    .D(_0536_),
    .Q_N(_0085_),
    .Q(\main.adder.s1_rs.levels[0][33] ));
 sg13g2_dfrbp_1 _6977_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net242),
    .D(_0537_),
    .Q_N(_0088_),
    .Q(\main.adder.s1_rs.levels[0][34] ));
 sg13g2_dfrbp_1 _6978_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net240),
    .D(_0538_),
    .Q_N(_0087_),
    .Q(\main.adder.s1_rs.levels[0][35] ));
 sg13g2_dfrbp_1 _6979_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net238),
    .D(_0539_),
    .Q_N(_0090_),
    .Q(\main.adder.s1_rs.levels[0][36] ));
 sg13g2_dfrbp_1 _6980_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net236),
    .D(_0540_),
    .Q_N(_0089_),
    .Q(\main.adder.s1_rs.levels[0][37] ));
 sg13g2_dfrbp_1 _6981_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net234),
    .D(_0541_),
    .Q_N(_0092_),
    .Q(\main.adder.s1_rs.levels[0][38] ));
 sg13g2_dfrbp_1 _6982_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net232),
    .D(_0542_),
    .Q_N(_0091_),
    .Q(\main.adder.s1_rs.levels[0][39] ));
 sg13g2_dfrbp_1 _6983_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net230),
    .D(_0543_),
    .Q_N(_0094_),
    .Q(\main.adder.s1_rs.levels[0][40] ));
 sg13g2_dfrbp_1 _6984_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net228),
    .D(_0544_),
    .Q_N(_0093_),
    .Q(\main.adder.s1_rs.levels[0][41] ));
 sg13g2_dfrbp_1 _6985_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net226),
    .D(_0545_),
    .Q_N(_0096_),
    .Q(\main.adder.s1_rs.levels[0][42] ));
 sg13g2_dfrbp_1 _6986_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net224),
    .D(_0546_),
    .Q_N(_0095_),
    .Q(\main.adder.s1_rs.levels[0][43] ));
 sg13g2_dfrbp_1 _6987_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net222),
    .D(_0547_),
    .Q_N(_0098_),
    .Q(\main.adder.s1_rs.levels[0][44] ));
 sg13g2_dfrbp_1 _6988_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net220),
    .D(_0548_),
    .Q_N(_0097_),
    .Q(\main.adder.s1_rs.levels[0][45] ));
 sg13g2_dfrbp_1 _6989_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net218),
    .D(_0549_),
    .Q_N(_2956_),
    .Q(\main.adder.s1_smaler[23] ));
 sg13g2_dfrbp_1 _6990_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net216),
    .D(_0550_),
    .Q_N(_2955_),
    .Q(\main.adder.s1_smaler[24] ));
 sg13g2_dfrbp_1 _6991_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net214),
    .D(_0551_),
    .Q_N(_2954_),
    .Q(\main.adder.s1_smaler[25] ));
 sg13g2_dfrbp_1 _6992_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net212),
    .D(_0552_),
    .Q_N(_2953_),
    .Q(\main.adder.s1_smaler[26] ));
 sg13g2_dfrbp_1 _6993_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net210),
    .D(_0553_),
    .Q_N(_2952_),
    .Q(\main.adder.s1_smaler[27] ));
 sg13g2_dfrbp_1 _6994_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net208),
    .D(_0554_),
    .Q_N(_2951_),
    .Q(\main.adder.s1_smaler[28] ));
 sg13g2_dfrbp_1 _6995_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net206),
    .D(_0555_),
    .Q_N(_2950_),
    .Q(\main.adder.s1_smaler[29] ));
 sg13g2_dfrbp_1 _6996_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net204),
    .D(_0556_),
    .Q_N(_2949_),
    .Q(\main.adder.s1_smaler[30] ));
 sg13g2_dfrbp_1 _6997_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net202),
    .D(_0557_),
    .Q_N(_2948_),
    .Q(\main.adder.s1_smaler[31] ));
 sg13g2_dfrbp_1 _6998_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net200),
    .D(_0558_),
    .Q_N(_2947_),
    .Q(\main.adder.s1_larger[0] ));
 sg13g2_dfrbp_1 _6999_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net198),
    .D(_0559_),
    .Q_N(_2946_),
    .Q(\main.adder.s1_larger[1] ));
 sg13g2_dfrbp_1 _7000_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net196),
    .D(_0560_),
    .Q_N(_2945_),
    .Q(\main.adder.s1_larger[2] ));
 sg13g2_dfrbp_1 _7001_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net194),
    .D(_0561_),
    .Q_N(_2944_),
    .Q(\main.adder.s1_larger[3] ));
 sg13g2_dfrbp_1 _7002_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net192),
    .D(_0562_),
    .Q_N(_2943_),
    .Q(\main.adder.s1_larger[4] ));
 sg13g2_dfrbp_1 _7003_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net190),
    .D(_0563_),
    .Q_N(_2942_),
    .Q(\main.adder.s1_larger[5] ));
 sg13g2_dfrbp_1 _7004_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net188),
    .D(_0564_),
    .Q_N(_2941_),
    .Q(\main.adder.s1_larger[6] ));
 sg13g2_dfrbp_1 _7005_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net186),
    .D(_0565_),
    .Q_N(_2940_),
    .Q(\main.adder.s1_larger[7] ));
 sg13g2_dfrbp_1 _7006_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net184),
    .D(_0566_),
    .Q_N(_2939_),
    .Q(\main.adder.s1_larger[8] ));
 sg13g2_dfrbp_1 _7007_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net182),
    .D(_0567_),
    .Q_N(_2938_),
    .Q(\main.adder.s1_larger[9] ));
 sg13g2_dfrbp_1 _7008_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net180),
    .D(_0568_),
    .Q_N(_2937_),
    .Q(\main.adder.s1_larger[10] ));
 sg13g2_dfrbp_1 _7009_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net178),
    .D(_0569_),
    .Q_N(_2936_),
    .Q(\main.adder.s1_larger[11] ));
 sg13g2_dfrbp_1 _7010_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net176),
    .D(_0570_),
    .Q_N(_2935_),
    .Q(\main.adder.s1_larger[12] ));
 sg13g2_dfrbp_1 _7011_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net174),
    .D(_0571_),
    .Q_N(_2934_),
    .Q(\main.adder.s1_larger[13] ));
 sg13g2_dfrbp_1 _7012_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net172),
    .D(_0572_),
    .Q_N(_2933_),
    .Q(\main.adder.s1_larger[14] ));
 sg13g2_dfrbp_1 _7013_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net170),
    .D(_0573_),
    .Q_N(_2932_),
    .Q(\main.adder.s1_larger[15] ));
 sg13g2_dfrbp_1 _7014_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net168),
    .D(_0574_),
    .Q_N(_2931_),
    .Q(\main.adder.s1_larger[16] ));
 sg13g2_dfrbp_1 _7015_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net166),
    .D(_0575_),
    .Q_N(_2930_),
    .Q(\main.adder.s1_larger[17] ));
 sg13g2_dfrbp_1 _7016_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net164),
    .D(_0576_),
    .Q_N(_2929_),
    .Q(\main.adder.s1_larger[18] ));
 sg13g2_dfrbp_1 _7017_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net162),
    .D(_0577_),
    .Q_N(_2928_),
    .Q(\main.adder.s1_larger[19] ));
 sg13g2_dfrbp_1 _7018_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net160),
    .D(_0578_),
    .Q_N(_2927_),
    .Q(\main.adder.s1_larger[20] ));
 sg13g2_dfrbp_1 _7019_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net158),
    .D(_0579_),
    .Q_N(_2926_),
    .Q(\main.adder.s1_larger[21] ));
 sg13g2_dfrbp_1 _7020_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net156),
    .D(_0580_),
    .Q_N(_2925_),
    .Q(\main.adder.s1_larger[22] ));
 sg13g2_dfrbp_1 _7021_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net154),
    .D(_0581_),
    .Q_N(_2924_),
    .Q(\main.adder.s1_larger[23] ));
 sg13g2_dfrbp_1 _7022_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net152),
    .D(_0582_),
    .Q_N(_2923_),
    .Q(\main.adder.s1_larger[24] ));
 sg13g2_dfrbp_1 _7023_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net150),
    .D(_0583_),
    .Q_N(_2922_),
    .Q(\main.adder.s1_larger[25] ));
 sg13g2_dfrbp_1 _7024_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net148),
    .D(_0584_),
    .Q_N(_2921_),
    .Q(\main.adder.s1_larger[26] ));
 sg13g2_dfrbp_1 _7025_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net140),
    .D(_0585_),
    .Q_N(_2920_),
    .Q(\main.adder.s1_larger[27] ));
 sg13g2_dfrbp_1 _7026_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net138),
    .D(_0586_),
    .Q_N(_2919_),
    .Q(\main.adder.s1_larger[28] ));
 sg13g2_dfrbp_1 _7027_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net136),
    .D(_0587_),
    .Q_N(_2918_),
    .Q(\main.adder.s1_larger[29] ));
 sg13g2_dfrbp_1 _7028_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net134),
    .D(_0588_),
    .Q_N(_2917_),
    .Q(\main.adder.s1_larger[30] ));
 sg13g2_dfrbp_1 _7029_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net132),
    .D(_0589_),
    .Q_N(_2916_),
    .Q(\main.adder.s1_larger[31] ));
 sg13g2_dfrbp_1 _7030_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net130),
    .D(_0590_),
    .Q_N(_2915_),
    .Q(\main.adder.s4_exponent_adjust[9] ));
 sg13g2_dfrbp_1 _7031_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net88),
    .D(_0591_),
    .Q_N(_2914_),
    .Q(\main.adder.s1_exp_diff[0] ));
 sg13g2_dfrbp_1 _7032_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net86),
    .D(_0592_),
    .Q_N(_2913_),
    .Q(\main.adder.s1_exp_diff[1] ));
 sg13g2_dfrbp_1 _7033_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net84),
    .D(_0593_),
    .Q_N(_2912_),
    .Q(\main.adder.s1_exp_diff[2] ));
 sg13g2_dfrbp_1 _7034_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net82),
    .D(_0594_),
    .Q_N(_2911_),
    .Q(\main.adder.s1_exp_diff[3] ));
 sg13g2_dfrbp_1 _7035_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net80),
    .D(_0595_),
    .Q_N(_2910_),
    .Q(\main.adder.s1_exp_diff[4] ));
 sg13g2_dfrbp_1 _7036_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net78),
    .D(_0596_),
    .Q_N(_2909_),
    .Q(\main.adder.s1_exp_diff[5] ));
 sg13g2_dfrbp_1 _7037_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net76),
    .D(_0597_),
    .Q_N(_2908_),
    .Q(\main.adder.s1_exp_diff[6] ));
 sg13g2_dfrbp_1 _7038_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net74),
    .D(_0598_),
    .Q_N(_2907_),
    .Q(\main.adder.s1_exp_diff[7] ));
 sg13g2_dfrbp_1 _7039_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net72),
    .D(_0599_),
    .Q_N(_2906_),
    .Q(\main.adder.s1_exp_diff[8] ));
 sg13g2_dfrbp_1 _7040_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net70),
    .D(_0600_),
    .Q_N(_2905_),
    .Q(\main.adder.s1_exp_diff[9] ));
 sg13g2_dfrbp_1 _7041_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net68),
    .D(net671),
    .Q_N(_0125_),
    .Q(\main.spi.out_bit_counter[0] ));
 sg13g2_dfrbp_1 _7042_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net64),
    .D(net1593),
    .Q_N(_2904_),
    .Q(\main.spi.out_bit_counter[1] ));
 sg13g2_dfrbp_1 _7043_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net60),
    .D(net1430),
    .Q_N(_2903_),
    .Q(\main.spi.out_bit_counter[2] ));
 sg13g2_dfrbp_1 _7044_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net56),
    .D(_0604_),
    .Q_N(_2902_),
    .Q(\main.SPI_output_data_ready ));
 sg13g2_dfrbp_1 _7045_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net52),
    .D(_0605_),
    .Q_N(_2901_),
    .Q(\main.spi.out_data_r[0] ));
 sg13g2_dfrbp_1 _7046_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net48),
    .D(_0606_),
    .Q_N(_2900_),
    .Q(\main.spi.out_data_r[1] ));
 sg13g2_dfrbp_1 _7047_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net554),
    .D(_0607_),
    .Q_N(_2899_),
    .Q(\main.spi.out_data_r[2] ));
 sg13g2_dfrbp_1 _7048_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net550),
    .D(_0608_),
    .Q_N(_2898_),
    .Q(\main.spi.out_data_r[3] ));
 sg13g2_dfrbp_1 _7049_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net546),
    .D(_0609_),
    .Q_N(_2897_),
    .Q(\main.spi.out_data_r[4] ));
 sg13g2_dfrbp_1 _7050_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net542),
    .D(_0610_),
    .Q_N(_2896_),
    .Q(\main.spi.out_data_r[5] ));
 sg13g2_dfrbp_1 _7051_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net538),
    .D(_0611_),
    .Q_N(_2895_),
    .Q(\main.spi.out_data_r[6] ));
 sg13g2_dfrbp_1 _7052_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net534),
    .D(_0612_),
    .Q_N(_2894_),
    .Q(\main.spi.out_data_r[7] ));
 sg13g2_dfrbp_1 _7053_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net530),
    .D(net792),
    .Q_N(_2893_),
    .Q(\main.SPI_out ));
 sg13g2_dfrbp_1 _7054_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net522),
    .D(net583),
    .Q_N(_0124_),
    .Q(\main.spi.in_bit_counter[0] ));
 sg13g2_dfrbp_1 _7055_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net518),
    .D(_0615_),
    .Q_N(_2892_),
    .Q(\main.spi.in_bit_counter[1] ));
 sg13g2_dfrbp_1 _7056_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net525),
    .D(net701),
    .Q_N(_3277_),
    .Q(\main.spi.in_bit_counter[2] ));
 sg13g2_dfrbp_1 _7057_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net526),
    .D(net1),
    .Q_N(_3278_),
    .Q(\main.spi.SPI_clock_sampler.sample_register[0] ));
 sg13g2_dfrbp_1 _7058_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net527),
    .D(_0012_),
    .Q_N(_3279_),
    .Q(\main.spi.SPI_clock_sampled ));
 sg13g2_dfrbp_1 _7059_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net528),
    .D(net2),
    .Q_N(_3280_),
    .Q(\main.spi.SPI_not_chip_select_sampler.sample_register[0] ));
 sg13g2_dfrbp_1 _7060_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net529),
    .D(_0014_),
    .Q_N(_3281_),
    .Q(\main.spi.SPI_not_chip_select_sampled ));
 sg13g2_dfrbp_1 _7061_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net500),
    .D(net3),
    .Q_N(_3282_),
    .Q(\main.spi.SPI_in_sampler.sample_register[0] ));
 sg13g2_dfrbp_1 _7062_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net514),
    .D(_0013_),
    .Q_N(_2891_),
    .Q(\main.spi.SPI_in_sampled ));
 sg13g2_dfrbp_1 _7063_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net510),
    .D(net616),
    .Q_N(_2890_),
    .Q(\main.SPI_input_data[0] ));
 sg13g2_dfrbp_1 _7064_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net506),
    .D(_0618_),
    .Q_N(_2889_),
    .Q(\main.SPI_input_data[1] ));
 sg13g2_dfrbp_1 _7065_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net502),
    .D(_0619_),
    .Q_N(_2888_),
    .Q(\main.SPI_input_data[2] ));
 sg13g2_dfrbp_1 _7066_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net498),
    .D(_0620_),
    .Q_N(_2887_),
    .Q(\main.SPI_input_data[3] ));
 sg13g2_dfrbp_1 _7067_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net494),
    .D(net1538),
    .Q_N(_2886_),
    .Q(\main.SPI_input_data[4] ));
 sg13g2_dfrbp_1 _7068_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net490),
    .D(_0622_),
    .Q_N(_2885_),
    .Q(\main.SPI_input_data[5] ));
 sg13g2_dfrbp_1 _7069_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net474),
    .D(net1532),
    .Q_N(_2884_),
    .Q(\main.SPI_input_data[6] ));
 sg13g2_dfrbp_1 _7070_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net470),
    .D(net1556),
    .Q_N(_2883_),
    .Q(\main.SPI_input_data[7] ));
 sg13g2_dfrbp_1 _7071_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net466),
    .D(_0625_),
    .Q_N(_2882_),
    .Q(_0002_));
 sg13g2_dfrbp_1 _7072_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net464),
    .D(_0626_),
    .Q_N(_2881_),
    .Q(_0003_));
 sg13g2_dfrbp_1 _7073_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net462),
    .D(_0627_),
    .Q_N(_2880_),
    .Q(\main.register_id_input_b[0] ));
 sg13g2_dfrbp_1 _7074_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net458),
    .D(_0628_),
    .Q_N(_2879_),
    .Q(\main.register_id_input_b[1] ));
 sg13g2_dfrbp_1 _7075_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net452),
    .D(_0629_),
    .Q_N(_2878_),
    .Q(\main.register_id_input_a[0] ));
 sg13g2_dfrbp_1 _7076_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net448),
    .D(_0630_),
    .Q_N(_2877_),
    .Q(\main.register_id_input_a[1] ));
 sg13g2_dfrbp_1 _7077_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net444),
    .D(_0631_),
    .Q_N(_2876_),
    .Q(\main.register_id_result[0] ));
 sg13g2_dfrbp_1 _7078_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net440),
    .D(_0632_),
    .Q_N(_2875_),
    .Q(\main.register_id_result[1] ));
 sg13g2_dfrbp_1 _7079_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net294),
    .D(net1591),
    .Q_N(_2874_),
    .Q(\main.read_command[0] ));
 sg13g2_dfrbp_1 _7080_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net272),
    .D(net1528),
    .Q_N(_2873_),
    .Q(\main.read_command[1] ));
 sg13g2_dfrbp_1 _7081_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net128),
    .D(_0635_),
    .Q_N(_2872_),
    .Q(\main.adder.s2_smaler[0] ));
 sg13g2_dfrbp_1 _7082_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net66),
    .D(_0636_),
    .Q_N(_2871_),
    .Q(\main.adder.s2_smaler[1] ));
 sg13g2_dfrbp_1 _7083_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net62),
    .D(_0637_),
    .Q_N(_2870_),
    .Q(\main.adder.s2_smaler[2] ));
 sg13g2_dfrbp_1 _7084_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net58),
    .D(_0638_),
    .Q_N(_2869_),
    .Q(\main.adder.s2_smaler[3] ));
 sg13g2_dfrbp_1 _7085_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net54),
    .D(_0639_),
    .Q_N(_2868_),
    .Q(\main.adder.s2_smaler[4] ));
 sg13g2_dfrbp_1 _7086_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net50),
    .D(_0640_),
    .Q_N(_2867_),
    .Q(\main.adder.s2_smaler[5] ));
 sg13g2_dfrbp_1 _7087_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net46),
    .D(_0641_),
    .Q_N(_2866_),
    .Q(\main.adder.s2_smaler[6] ));
 sg13g2_dfrbp_1 _7088_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net552),
    .D(_0642_),
    .Q_N(_2865_),
    .Q(\main.adder.s2_smaler[7] ));
 sg13g2_dfrbp_1 _7089_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net548),
    .D(_0643_),
    .Q_N(_2864_),
    .Q(\main.adder.s2_smaler[8] ));
 sg13g2_dfrbp_1 _7090_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net544),
    .D(_0644_),
    .Q_N(_2863_),
    .Q(\main.adder.s2_smaler[9] ));
 sg13g2_dfrbp_1 _7091_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net540),
    .D(_0645_),
    .Q_N(_2862_),
    .Q(\main.adder.s2_smaler[10] ));
 sg13g2_dfrbp_1 _7092_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net536),
    .D(_0646_),
    .Q_N(_2861_),
    .Q(\main.adder.s2_smaler[11] ));
 sg13g2_dfrbp_1 _7093_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net532),
    .D(_0647_),
    .Q_N(_2860_),
    .Q(\main.adder.s2_smaler[12] ));
 sg13g2_dfrbp_1 _7094_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net520),
    .D(_0648_),
    .Q_N(_2859_),
    .Q(\main.adder.s2_smaler[13] ));
 sg13g2_dfrbp_1 _7095_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net516),
    .D(_0649_),
    .Q_N(_2858_),
    .Q(\main.adder.s2_smaler[14] ));
 sg13g2_dfrbp_1 _7096_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net512),
    .D(_0650_),
    .Q_N(_2857_),
    .Q(\main.float_registers[3][7] ));
 sg13g2_dfrbp_1 _7097_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net508),
    .D(net1482),
    .Q_N(_2856_),
    .Q(\main.float_registers[3][14] ));
 sg13g2_dfrbp_1 _7098_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net504),
    .D(_0652_),
    .Q_N(_2855_),
    .Q(\main.float_registers[1][0] ));
 sg13g2_dfrbp_1 _7099_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net496),
    .D(_0653_),
    .Q_N(_2854_),
    .Q(\main.float_registers[3][11] ));
 sg13g2_dfrbp_1 _7100_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net492),
    .D(_0654_),
    .Q_N(_2853_),
    .Q(\main.float_registers[3][15] ));
 sg13g2_dfrbp_1 _7101_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net488),
    .D(_0655_),
    .Q_N(_2852_),
    .Q(\main.float_registers[0][24] ));
 sg13g2_dfrbp_1 _7102_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net468),
    .D(_0656_),
    .Q_N(_2851_),
    .Q(\main.float_registers[2][0] ));
 sg13g2_dfrbp_1 _7103_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net454),
    .D(_0657_),
    .Q_N(_2850_),
    .Q(\main.float_registers[3][27] ));
 sg13g2_dfrbp_1 _7104_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net450),
    .D(net628),
    .Q_N(_2849_),
    .Q(_0000_));
 sg13g2_dfrbp_1 _7105_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net446),
    .D(net693),
    .Q_N(_2848_),
    .Q(_0001_));
 sg13g2_dfrbp_1 _7106_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net442),
    .D(_0660_),
    .Q_N(_2847_),
    .Q(\main.float_registers[3][26] ));
 sg13g2_dfrbp_1 _7107_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net438),
    .D(net1507),
    .Q_N(_2846_),
    .Q(\main.float_registers[2][31] ));
 sg13g2_dfrbp_1 _7108_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net472),
    .D(net1451),
    .Q_N(_2845_),
    .Q(\main.float_registers[3][25] ));
 sg13g2_dfrbp_1 _7109_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net460),
    .D(_0663_),
    .Q_N(_2844_),
    .Q(\main.float_registers[3][24] ));
 sg13g2_tiehi _6740__28 (.L_HI(net28));
 sg13g2_tiehi _6739__29 (.L_HI(net29));
 sg13g2_tiehi _6738__30 (.L_HI(net30));
 sg13g2_tiehi _6737__31 (.L_HI(net31));
 sg13g2_tiehi _6736__32 (.L_HI(net32));
 sg13g2_tiehi _6735__33 (.L_HI(net33));
 sg13g2_tiehi _6734__34 (.L_HI(net34));
 sg13g2_tiehi _6733__35 (.L_HI(net35));
 sg13g2_tiehi _6732__36 (.L_HI(net36));
 sg13g2_tiehi _6731__37 (.L_HI(net37));
 sg13g2_tiehi _6730__38 (.L_HI(net38));
 sg13g2_tiehi _6729__39 (.L_HI(net39));
 sg13g2_tiehi _6728__40 (.L_HI(net40));
 sg13g2_tiehi _6727__41 (.L_HI(net41));
 sg13g2_tiehi _6726__42 (.L_HI(net42));
 sg13g2_tiehi _6725__43 (.L_HI(net43));
 sg13g2_tiehi _6724__44 (.L_HI(net44));
 sg13g2_tiehi _6723__45 (.L_HI(net45));
 sg13g2_tiehi _7087__46 (.L_HI(net46));
 sg13g2_tiehi _6722__47 (.L_HI(net47));
 sg13g2_tiehi _7046__48 (.L_HI(net48));
 sg13g2_tiehi _6721__49 (.L_HI(net49));
 sg13g2_tiehi _7086__50 (.L_HI(net50));
 sg13g2_tiehi _6720__51 (.L_HI(net51));
 sg13g2_tiehi _7045__52 (.L_HI(net52));
 sg13g2_tiehi _6719__53 (.L_HI(net53));
 sg13g2_tiehi _7085__54 (.L_HI(net54));
 sg13g2_tiehi _6718__55 (.L_HI(net55));
 sg13g2_tiehi _7044__56 (.L_HI(net56));
 sg13g2_tiehi _6717__57 (.L_HI(net57));
 sg13g2_tiehi _7084__58 (.L_HI(net58));
 sg13g2_tiehi _6716__59 (.L_HI(net59));
 sg13g2_tiehi _7043__60 (.L_HI(net60));
 sg13g2_tiehi _6715__61 (.L_HI(net61));
 sg13g2_tiehi _7083__62 (.L_HI(net62));
 sg13g2_tiehi _6714__63 (.L_HI(net63));
 sg13g2_tiehi _7042__64 (.L_HI(net64));
 sg13g2_tiehi _6713__65 (.L_HI(net65));
 sg13g2_tiehi _7082__66 (.L_HI(net66));
 sg13g2_tiehi _6712__67 (.L_HI(net67));
 sg13g2_tiehi _7041__68 (.L_HI(net68));
 sg13g2_tiehi _6711__69 (.L_HI(net69));
 sg13g2_tiehi _7040__70 (.L_HI(net70));
 sg13g2_tiehi _6710__71 (.L_HI(net71));
 sg13g2_tiehi _7039__72 (.L_HI(net72));
 sg13g2_tiehi _6709__73 (.L_HI(net73));
 sg13g2_tiehi _7038__74 (.L_HI(net74));
 sg13g2_tiehi _6708__75 (.L_HI(net75));
 sg13g2_tiehi _7037__76 (.L_HI(net76));
 sg13g2_tiehi _6707__77 (.L_HI(net77));
 sg13g2_tiehi _7036__78 (.L_HI(net78));
 sg13g2_tiehi _6706__79 (.L_HI(net79));
 sg13g2_tiehi _7035__80 (.L_HI(net80));
 sg13g2_tiehi _6705__81 (.L_HI(net81));
 sg13g2_tiehi _7034__82 (.L_HI(net82));
 sg13g2_tiehi _6704__83 (.L_HI(net83));
 sg13g2_tiehi _7033__84 (.L_HI(net84));
 sg13g2_tiehi _6703__85 (.L_HI(net85));
 sg13g2_tiehi _7032__86 (.L_HI(net86));
 sg13g2_tiehi _6702__87 (.L_HI(net87));
 sg13g2_tiehi _7031__88 (.L_HI(net88));
 sg13g2_tiehi _6701__89 (.L_HI(net89));
 sg13g2_tiehi _6700__90 (.L_HI(net90));
 sg13g2_tiehi _6699__91 (.L_HI(net91));
 sg13g2_tiehi _6698__92 (.L_HI(net92));
 sg13g2_tiehi _6697__93 (.L_HI(net93));
 sg13g2_tiehi _6696__94 (.L_HI(net94));
 sg13g2_tiehi _6695__95 (.L_HI(net95));
 sg13g2_tiehi _6694__96 (.L_HI(net96));
 sg13g2_tiehi _6693__97 (.L_HI(net97));
 sg13g2_tiehi _6692__98 (.L_HI(net98));
 sg13g2_tiehi _6691__99 (.L_HI(net99));
 sg13g2_tiehi _6690__100 (.L_HI(net100));
 sg13g2_tiehi _6689__101 (.L_HI(net101));
 sg13g2_tiehi _6688__102 (.L_HI(net102));
 sg13g2_tiehi _6687__103 (.L_HI(net103));
 sg13g2_tiehi _6686__104 (.L_HI(net104));
 sg13g2_tiehi _6685__105 (.L_HI(net105));
 sg13g2_tiehi _6684__106 (.L_HI(net106));
 sg13g2_tiehi _6683__107 (.L_HI(net107));
 sg13g2_tiehi _6682__108 (.L_HI(net108));
 sg13g2_tiehi _6681__109 (.L_HI(net109));
 sg13g2_tiehi _6680__110 (.L_HI(net110));
 sg13g2_tiehi _6673__111 (.L_HI(net111));
 sg13g2_tiehi _6672__112 (.L_HI(net112));
 sg13g2_tiehi _6671__113 (.L_HI(net113));
 sg13g2_tiehi _6670__114 (.L_HI(net114));
 sg13g2_tiehi _6669__115 (.L_HI(net115));
 sg13g2_tiehi _6668__116 (.L_HI(net116));
 sg13g2_tiehi _6667__117 (.L_HI(net117));
 sg13g2_tiehi _6666__118 (.L_HI(net118));
 sg13g2_tiehi _6665__119 (.L_HI(net119));
 sg13g2_tiehi _6664__120 (.L_HI(net120));
 sg13g2_tiehi _6663__121 (.L_HI(net121));
 sg13g2_tiehi _6662__122 (.L_HI(net122));
 sg13g2_tiehi _6661__123 (.L_HI(net123));
 sg13g2_tiehi _6660__124 (.L_HI(net124));
 sg13g2_tiehi _6659__125 (.L_HI(net125));
 sg13g2_tiehi _6658__126 (.L_HI(net126));
 sg13g2_tiehi _6657__127 (.L_HI(net127));
 sg13g2_tiehi _7081__128 (.L_HI(net128));
 sg13g2_tiehi _6656__129 (.L_HI(net129));
 sg13g2_tiehi _7030__130 (.L_HI(net130));
 sg13g2_tiehi _6655__131 (.L_HI(net131));
 sg13g2_tiehi _7029__132 (.L_HI(net132));
 sg13g2_tiehi _6654__133 (.L_HI(net133));
 sg13g2_tiehi _7028__134 (.L_HI(net134));
 sg13g2_tiehi _6653__135 (.L_HI(net135));
 sg13g2_tiehi _7027__136 (.L_HI(net136));
 sg13g2_tiehi _6652__137 (.L_HI(net137));
 sg13g2_tiehi _7026__138 (.L_HI(net138));
 sg13g2_tiehi _6651__139 (.L_HI(net139));
 sg13g2_tiehi _7025__140 (.L_HI(net140));
 sg13g2_tiehi _6650__141 (.L_HI(net141));
 sg13g2_tiehi _6560__142 (.L_HI(net142));
 sg13g2_tiehi _6674__143 (.L_HI(net143));
 sg13g2_tiehi _6675__144 (.L_HI(net144));
 sg13g2_tiehi _6676__145 (.L_HI(net145));
 sg13g2_tiehi _6677__146 (.L_HI(net146));
 sg13g2_tiehi _6678__147 (.L_HI(net147));
 sg13g2_tiehi _7024__148 (.L_HI(net148));
 sg13g2_tiehi _6649__149 (.L_HI(net149));
 sg13g2_tiehi _7023__150 (.L_HI(net150));
 sg13g2_tiehi _6648__151 (.L_HI(net151));
 sg13g2_tiehi _7022__152 (.L_HI(net152));
 sg13g2_tiehi _6647__153 (.L_HI(net153));
 sg13g2_tiehi _7021__154 (.L_HI(net154));
 sg13g2_tiehi _6646__155 (.L_HI(net155));
 sg13g2_tiehi _7020__156 (.L_HI(net156));
 sg13g2_tiehi _6645__157 (.L_HI(net157));
 sg13g2_tiehi _7019__158 (.L_HI(net158));
 sg13g2_tiehi _6644__159 (.L_HI(net159));
 sg13g2_tiehi _7018__160 (.L_HI(net160));
 sg13g2_tiehi _6643__161 (.L_HI(net161));
 sg13g2_tiehi _7017__162 (.L_HI(net162));
 sg13g2_tiehi _6642__163 (.L_HI(net163));
 sg13g2_tiehi _7016__164 (.L_HI(net164));
 sg13g2_tiehi _6641__165 (.L_HI(net165));
 sg13g2_tiehi _7015__166 (.L_HI(net166));
 sg13g2_tiehi _6640__167 (.L_HI(net167));
 sg13g2_tiehi _7014__168 (.L_HI(net168));
 sg13g2_tiehi _6639__169 (.L_HI(net169));
 sg13g2_tiehi _7013__170 (.L_HI(net170));
 sg13g2_tiehi _6638__171 (.L_HI(net171));
 sg13g2_tiehi _7012__172 (.L_HI(net172));
 sg13g2_tiehi _6637__173 (.L_HI(net173));
 sg13g2_tiehi _7011__174 (.L_HI(net174));
 sg13g2_tiehi _6636__175 (.L_HI(net175));
 sg13g2_tiehi _7010__176 (.L_HI(net176));
 sg13g2_tiehi _6635__177 (.L_HI(net177));
 sg13g2_tiehi _7009__178 (.L_HI(net178));
 sg13g2_tiehi _6634__179 (.L_HI(net179));
 sg13g2_tiehi _7008__180 (.L_HI(net180));
 sg13g2_tiehi _6633__181 (.L_HI(net181));
 sg13g2_tiehi _7007__182 (.L_HI(net182));
 sg13g2_tiehi _6632__183 (.L_HI(net183));
 sg13g2_tiehi _7006__184 (.L_HI(net184));
 sg13g2_tiehi _6631__185 (.L_HI(net185));
 sg13g2_tiehi _7005__186 (.L_HI(net186));
 sg13g2_tiehi _6630__187 (.L_HI(net187));
 sg13g2_tiehi _7004__188 (.L_HI(net188));
 sg13g2_tiehi _6629__189 (.L_HI(net189));
 sg13g2_tiehi _7003__190 (.L_HI(net190));
 sg13g2_tiehi _6628__191 (.L_HI(net191));
 sg13g2_tiehi _7002__192 (.L_HI(net192));
 sg13g2_tiehi _6627__193 (.L_HI(net193));
 sg13g2_tiehi _7001__194 (.L_HI(net194));
 sg13g2_tiehi _6626__195 (.L_HI(net195));
 sg13g2_tiehi _7000__196 (.L_HI(net196));
 sg13g2_tiehi _6625__197 (.L_HI(net197));
 sg13g2_tiehi _6999__198 (.L_HI(net198));
 sg13g2_tiehi _6624__199 (.L_HI(net199));
 sg13g2_tiehi _6998__200 (.L_HI(net200));
 sg13g2_tiehi _6623__201 (.L_HI(net201));
 sg13g2_tiehi _6997__202 (.L_HI(net202));
 sg13g2_tiehi _6622__203 (.L_HI(net203));
 sg13g2_tiehi _6996__204 (.L_HI(net204));
 sg13g2_tiehi _6621__205 (.L_HI(net205));
 sg13g2_tiehi _6995__206 (.L_HI(net206));
 sg13g2_tiehi _6620__207 (.L_HI(net207));
 sg13g2_tiehi _6994__208 (.L_HI(net208));
 sg13g2_tiehi _6619__209 (.L_HI(net209));
 sg13g2_tiehi _6993__210 (.L_HI(net210));
 sg13g2_tiehi _6618__211 (.L_HI(net211));
 sg13g2_tiehi _6992__212 (.L_HI(net212));
 sg13g2_tiehi _6617__213 (.L_HI(net213));
 sg13g2_tiehi _6991__214 (.L_HI(net214));
 sg13g2_tiehi _6616__215 (.L_HI(net215));
 sg13g2_tiehi _6990__216 (.L_HI(net216));
 sg13g2_tiehi _6615__217 (.L_HI(net217));
 sg13g2_tiehi _6989__218 (.L_HI(net218));
 sg13g2_tiehi _6614__219 (.L_HI(net219));
 sg13g2_tiehi _6988__220 (.L_HI(net220));
 sg13g2_tiehi _6613__221 (.L_HI(net221));
 sg13g2_tiehi _6987__222 (.L_HI(net222));
 sg13g2_tiehi _6612__223 (.L_HI(net223));
 sg13g2_tiehi _6986__224 (.L_HI(net224));
 sg13g2_tiehi _6611__225 (.L_HI(net225));
 sg13g2_tiehi _6985__226 (.L_HI(net226));
 sg13g2_tiehi _6610__227 (.L_HI(net227));
 sg13g2_tiehi _6984__228 (.L_HI(net228));
 sg13g2_tiehi _6609__229 (.L_HI(net229));
 sg13g2_tiehi _6983__230 (.L_HI(net230));
 sg13g2_tiehi _6608__231 (.L_HI(net231));
 sg13g2_tiehi _6982__232 (.L_HI(net232));
 sg13g2_tiehi _6607__233 (.L_HI(net233));
 sg13g2_tiehi _6981__234 (.L_HI(net234));
 sg13g2_tiehi _6606__235 (.L_HI(net235));
 sg13g2_tiehi _6980__236 (.L_HI(net236));
 sg13g2_tiehi _6605__237 (.L_HI(net237));
 sg13g2_tiehi _6979__238 (.L_HI(net238));
 sg13g2_tiehi _6604__239 (.L_HI(net239));
 sg13g2_tiehi _6978__240 (.L_HI(net240));
 sg13g2_tiehi _6603__241 (.L_HI(net241));
 sg13g2_tiehi _6977__242 (.L_HI(net242));
 sg13g2_tiehi _6602__243 (.L_HI(net243));
 sg13g2_tiehi _6976__244 (.L_HI(net244));
 sg13g2_tiehi _6601__245 (.L_HI(net245));
 sg13g2_tiehi _6975__246 (.L_HI(net246));
 sg13g2_tiehi _6600__247 (.L_HI(net247));
 sg13g2_tiehi _6974__248 (.L_HI(net248));
 sg13g2_tiehi _6599__249 (.L_HI(net249));
 sg13g2_tiehi _6973__250 (.L_HI(net250));
 sg13g2_tiehi _6598__251 (.L_HI(net251));
 sg13g2_tiehi _6972__252 (.L_HI(net252));
 sg13g2_tiehi _6597__253 (.L_HI(net253));
 sg13g2_tiehi _6971__254 (.L_HI(net254));
 sg13g2_tiehi _6596__255 (.L_HI(net255));
 sg13g2_tiehi _6970__256 (.L_HI(net256));
 sg13g2_tiehi _6595__257 (.L_HI(net257));
 sg13g2_tiehi _6969__258 (.L_HI(net258));
 sg13g2_tiehi _6594__259 (.L_HI(net259));
 sg13g2_tiehi _6968__260 (.L_HI(net260));
 sg13g2_tiehi _6593__261 (.L_HI(net261));
 sg13g2_tiehi _6967__262 (.L_HI(net262));
 sg13g2_tiehi _6592__263 (.L_HI(net263));
 sg13g2_tiehi _6966__264 (.L_HI(net264));
 sg13g2_tiehi _6591__265 (.L_HI(net265));
 sg13g2_tiehi _6965__266 (.L_HI(net266));
 sg13g2_tiehi _6590__267 (.L_HI(net267));
 sg13g2_tiehi _6964__268 (.L_HI(net268));
 sg13g2_tiehi _6589__269 (.L_HI(net269));
 sg13g2_tiehi _6963__270 (.L_HI(net270));
 sg13g2_tiehi _6588__271 (.L_HI(net271));
 sg13g2_tiehi _7080__272 (.L_HI(net272));
 sg13g2_tiehi _6587__273 (.L_HI(net273));
 sg13g2_tiehi _6962__274 (.L_HI(net274));
 sg13g2_tiehi _6586__275 (.L_HI(net275));
 sg13g2_tiehi _6961__276 (.L_HI(net276));
 sg13g2_tiehi _6585__277 (.L_HI(net277));
 sg13g2_tiehi _6960__278 (.L_HI(net278));
 sg13g2_tiehi _6584__279 (.L_HI(net279));
 sg13g2_tiehi _6959__280 (.L_HI(net280));
 sg13g2_tiehi _6583__281 (.L_HI(net281));
 sg13g2_tiehi _6958__282 (.L_HI(net282));
 sg13g2_tiehi _6582__283 (.L_HI(net283));
 sg13g2_tiehi _6957__284 (.L_HI(net284));
 sg13g2_tiehi _6581__285 (.L_HI(net285));
 sg13g2_tiehi _6956__286 (.L_HI(net286));
 sg13g2_tiehi _6580__287 (.L_HI(net287));
 sg13g2_tiehi _6955__288 (.L_HI(net288));
 sg13g2_tiehi _6579__289 (.L_HI(net289));
 sg13g2_tiehi _6954__290 (.L_HI(net290));
 sg13g2_tiehi _6578__291 (.L_HI(net291));
 sg13g2_tiehi _6953__292 (.L_HI(net292));
 sg13g2_tiehi _6577__293 (.L_HI(net293));
 sg13g2_tiehi _7079__294 (.L_HI(net294));
 sg13g2_tiehi _6576__295 (.L_HI(net295));
 sg13g2_tiehi _6952__296 (.L_HI(net296));
 sg13g2_tiehi _6575__297 (.L_HI(net297));
 sg13g2_tiehi _6951__298 (.L_HI(net298));
 sg13g2_tiehi _6574__299 (.L_HI(net299));
 sg13g2_tiehi _6950__300 (.L_HI(net300));
 sg13g2_tiehi _6573__301 (.L_HI(net301));
 sg13g2_tiehi _6949__302 (.L_HI(net302));
 sg13g2_tiehi _6572__303 (.L_HI(net303));
 sg13g2_tiehi _6948__304 (.L_HI(net304));
 sg13g2_tiehi _6571__305 (.L_HI(net305));
 sg13g2_tiehi _6947__306 (.L_HI(net306));
 sg13g2_tiehi _6570__307 (.L_HI(net307));
 sg13g2_tiehi _6946__308 (.L_HI(net308));
 sg13g2_tiehi _6569__309 (.L_HI(net309));
 sg13g2_tiehi _6945__310 (.L_HI(net310));
 sg13g2_tiehi _6568__311 (.L_HI(net311));
 sg13g2_tiehi _6944__312 (.L_HI(net312));
 sg13g2_tiehi _6567__313 (.L_HI(net313));
 sg13g2_tiehi _6943__314 (.L_HI(net314));
 sg13g2_tiehi _6566__315 (.L_HI(net315));
 sg13g2_tiehi _6565__316 (.L_HI(net316));
 sg13g2_tiehi _6564__317 (.L_HI(net317));
 sg13g2_tiehi _6563__318 (.L_HI(net318));
 sg13g2_tiehi _6942__319 (.L_HI(net319));
 sg13g2_tiehi _6562__320 (.L_HI(net320));
 sg13g2_tiehi _6941__321 (.L_HI(net321));
 sg13g2_tiehi _6561__322 (.L_HI(net322));
 sg13g2_tiehi _6940__323 (.L_HI(net323));
 sg13g2_tiehi _6939__324 (.L_HI(net324));
 sg13g2_tiehi _6938__325 (.L_HI(net325));
 sg13g2_tiehi _6937__326 (.L_HI(net326));
 sg13g2_tiehi _6936__327 (.L_HI(net327));
 sg13g2_tiehi _6935__328 (.L_HI(net328));
 sg13g2_tiehi _6934__329 (.L_HI(net329));
 sg13g2_tiehi _6933__330 (.L_HI(net330));
 sg13g2_tiehi _6932__331 (.L_HI(net331));
 sg13g2_tiehi _6931__332 (.L_HI(net332));
 sg13g2_tiehi _6930__333 (.L_HI(net333));
 sg13g2_tiehi _6929__334 (.L_HI(net334));
 sg13g2_tiehi _6928__335 (.L_HI(net335));
 sg13g2_tiehi _6927__336 (.L_HI(net336));
 sg13g2_tiehi _6926__337 (.L_HI(net337));
 sg13g2_tiehi _6925__338 (.L_HI(net338));
 sg13g2_tiehi _6924__339 (.L_HI(net339));
 sg13g2_tiehi _6923__340 (.L_HI(net340));
 sg13g2_tiehi _6922__341 (.L_HI(net341));
 sg13g2_tiehi _6921__342 (.L_HI(net342));
 sg13g2_tiehi _6920__343 (.L_HI(net343));
 sg13g2_tiehi _6919__344 (.L_HI(net344));
 sg13g2_tiehi _6918__345 (.L_HI(net345));
 sg13g2_tiehi _6917__346 (.L_HI(net346));
 sg13g2_tiehi _6916__347 (.L_HI(net347));
 sg13g2_tiehi _6915__348 (.L_HI(net348));
 sg13g2_tiehi _6914__349 (.L_HI(net349));
 sg13g2_tiehi _6913__350 (.L_HI(net350));
 sg13g2_tiehi _6912__351 (.L_HI(net351));
 sg13g2_tiehi _6911__352 (.L_HI(net352));
 sg13g2_tiehi _6910__353 (.L_HI(net353));
 sg13g2_tiehi _6909__354 (.L_HI(net354));
 sg13g2_tiehi _6908__355 (.L_HI(net355));
 sg13g2_tiehi _6907__356 (.L_HI(net356));
 sg13g2_tiehi _6906__357 (.L_HI(net357));
 sg13g2_tiehi _6905__358 (.L_HI(net358));
 sg13g2_tiehi _6904__359 (.L_HI(net359));
 sg13g2_tiehi _6903__360 (.L_HI(net360));
 sg13g2_tiehi _6902__361 (.L_HI(net361));
 sg13g2_tiehi _6901__362 (.L_HI(net362));
 sg13g2_tiehi _6900__363 (.L_HI(net363));
 sg13g2_tiehi _6899__364 (.L_HI(net364));
 sg13g2_tiehi _6898__365 (.L_HI(net365));
 sg13g2_tiehi _6897__366 (.L_HI(net366));
 sg13g2_tiehi _6896__367 (.L_HI(net367));
 sg13g2_tiehi _6895__368 (.L_HI(net368));
 sg13g2_tiehi _6894__369 (.L_HI(net369));
 sg13g2_tiehi _6893__370 (.L_HI(net370));
 sg13g2_tiehi _6892__371 (.L_HI(net371));
 sg13g2_tiehi _6891__372 (.L_HI(net372));
 sg13g2_tiehi _6890__373 (.L_HI(net373));
 sg13g2_tiehi _6889__374 (.L_HI(net374));
 sg13g2_tiehi _6888__375 (.L_HI(net375));
 sg13g2_tiehi _6887__376 (.L_HI(net376));
 sg13g2_tiehi _6886__377 (.L_HI(net377));
 sg13g2_tiehi _6885__378 (.L_HI(net378));
 sg13g2_tiehi _6884__379 (.L_HI(net379));
 sg13g2_tiehi _6883__380 (.L_HI(net380));
 sg13g2_tiehi _6882__381 (.L_HI(net381));
 sg13g2_tiehi _6881__382 (.L_HI(net382));
 sg13g2_tiehi _6880__383 (.L_HI(net383));
 sg13g2_tiehi _6879__384 (.L_HI(net384));
 sg13g2_tiehi _6878__385 (.L_HI(net385));
 sg13g2_tiehi _6877__386 (.L_HI(net386));
 sg13g2_tiehi _6876__387 (.L_HI(net387));
 sg13g2_tiehi _6875__388 (.L_HI(net388));
 sg13g2_tiehi _6874__389 (.L_HI(net389));
 sg13g2_tiehi _6873__390 (.L_HI(net390));
 sg13g2_tiehi _6872__391 (.L_HI(net391));
 sg13g2_tiehi _6871__392 (.L_HI(net392));
 sg13g2_tiehi _6870__393 (.L_HI(net393));
 sg13g2_tiehi _6869__394 (.L_HI(net394));
 sg13g2_tiehi _6868__395 (.L_HI(net395));
 sg13g2_tiehi _6867__396 (.L_HI(net396));
 sg13g2_tiehi _6866__397 (.L_HI(net397));
 sg13g2_tiehi _6865__398 (.L_HI(net398));
 sg13g2_tiehi _6864__399 (.L_HI(net399));
 sg13g2_tiehi _6863__400 (.L_HI(net400));
 sg13g2_tiehi _6862__401 (.L_HI(net401));
 sg13g2_tiehi _6861__402 (.L_HI(net402));
 sg13g2_tiehi _6860__403 (.L_HI(net403));
 sg13g2_tiehi _6859__404 (.L_HI(net404));
 sg13g2_tiehi _6858__405 (.L_HI(net405));
 sg13g2_tiehi _6857__406 (.L_HI(net406));
 sg13g2_tiehi _6856__407 (.L_HI(net407));
 sg13g2_tiehi _6855__408 (.L_HI(net408));
 sg13g2_tiehi _6854__409 (.L_HI(net409));
 sg13g2_tiehi _6853__410 (.L_HI(net410));
 sg13g2_tiehi _6852__411 (.L_HI(net411));
 sg13g2_tiehi _6851__412 (.L_HI(net412));
 sg13g2_tiehi _6850__413 (.L_HI(net413));
 sg13g2_tiehi _6849__414 (.L_HI(net414));
 sg13g2_tiehi _6848__415 (.L_HI(net415));
 sg13g2_tiehi _6847__416 (.L_HI(net416));
 sg13g2_tiehi _6846__417 (.L_HI(net417));
 sg13g2_tiehi _6845__418 (.L_HI(net418));
 sg13g2_tiehi _6844__419 (.L_HI(net419));
 sg13g2_tiehi _6843__420 (.L_HI(net420));
 sg13g2_tiehi _6842__421 (.L_HI(net421));
 sg13g2_tiehi _6841__422 (.L_HI(net422));
 sg13g2_tiehi _6840__423 (.L_HI(net423));
 sg13g2_tiehi _6839__424 (.L_HI(net424));
 sg13g2_tiehi _6838__425 (.L_HI(net425));
 sg13g2_tiehi _6837__426 (.L_HI(net426));
 sg13g2_tiehi _6836__427 (.L_HI(net427));
 sg13g2_tiehi _6835__428 (.L_HI(net428));
 sg13g2_tiehi _6834__429 (.L_HI(net429));
 sg13g2_tiehi _6833__430 (.L_HI(net430));
 sg13g2_tiehi _6832__431 (.L_HI(net431));
 sg13g2_tiehi _6831__432 (.L_HI(net432));
 sg13g2_tiehi _6830__433 (.L_HI(net433));
 sg13g2_tiehi _6829__434 (.L_HI(net434));
 sg13g2_tiehi _6828__435 (.L_HI(net435));
 sg13g2_tiehi _6827__436 (.L_HI(net436));
 sg13g2_tiehi _6826__437 (.L_HI(net437));
 sg13g2_tiehi _7107__438 (.L_HI(net438));
 sg13g2_tiehi _6825__439 (.L_HI(net439));
 sg13g2_tiehi _7078__440 (.L_HI(net440));
 sg13g2_tiehi _6824__441 (.L_HI(net441));
 sg13g2_tiehi _7106__442 (.L_HI(net442));
 sg13g2_tiehi _6823__443 (.L_HI(net443));
 sg13g2_tiehi _7077__444 (.L_HI(net444));
 sg13g2_tiehi _6822__445 (.L_HI(net445));
 sg13g2_tiehi _7105__446 (.L_HI(net446));
 sg13g2_tiehi _6821__447 (.L_HI(net447));
 sg13g2_tiehi _7076__448 (.L_HI(net448));
 sg13g2_tiehi _6820__449 (.L_HI(net449));
 sg13g2_tiehi _7104__450 (.L_HI(net450));
 sg13g2_tiehi _6819__451 (.L_HI(net451));
 sg13g2_tiehi _7075__452 (.L_HI(net452));
 sg13g2_tiehi _6818__453 (.L_HI(net453));
 sg13g2_tiehi _7103__454 (.L_HI(net454));
 sg13g2_tiehi _6817__455 (.L_HI(net455));
 sg13g2_tiehi _6816__456 (.L_HI(net456));
 sg13g2_tiehi _6815__457 (.L_HI(net457));
 sg13g2_tiehi _7074__458 (.L_HI(net458));
 sg13g2_tiehi _6814__459 (.L_HI(net459));
 sg13g2_tiehi _7109__460 (.L_HI(net460));
 sg13g2_tiehi _6813__461 (.L_HI(net461));
 sg13g2_tiehi _7073__462 (.L_HI(net462));
 sg13g2_tiehi _6812__463 (.L_HI(net463));
 sg13g2_tiehi _7072__464 (.L_HI(net464));
 sg13g2_tiehi _6811__465 (.L_HI(net465));
 sg13g2_tiehi _7071__466 (.L_HI(net466));
 sg13g2_tiehi _6810__467 (.L_HI(net467));
 sg13g2_tiehi _7102__468 (.L_HI(net468));
 sg13g2_tiehi _6809__469 (.L_HI(net469));
 sg13g2_tiehi _7070__470 (.L_HI(net470));
 sg13g2_tiehi _6808__471 (.L_HI(net471));
 sg13g2_tiehi _7108__472 (.L_HI(net472));
 sg13g2_tiehi _6807__473 (.L_HI(net473));
 sg13g2_tiehi _7069__474 (.L_HI(net474));
 sg13g2_tiehi _6806__475 (.L_HI(net475));
 sg13g2_tiehi _6805__476 (.L_HI(net476));
 sg13g2_tiehi _6804__477 (.L_HI(net477));
 sg13g2_tiehi _6803__478 (.L_HI(net478));
 sg13g2_tiehi _6802__479 (.L_HI(net479));
 sg13g2_tiehi _6801__480 (.L_HI(net480));
 sg13g2_tiehi _6800__481 (.L_HI(net481));
 sg13g2_tiehi _6799__482 (.L_HI(net482));
 sg13g2_tiehi _6798__483 (.L_HI(net483));
 sg13g2_tiehi _6797__484 (.L_HI(net484));
 sg13g2_tiehi _6796__485 (.L_HI(net485));
 sg13g2_tiehi _6795__486 (.L_HI(net486));
 sg13g2_tiehi _6794__487 (.L_HI(net487));
 sg13g2_tiehi _7101__488 (.L_HI(net488));
 sg13g2_tiehi _6793__489 (.L_HI(net489));
 sg13g2_tiehi _7068__490 (.L_HI(net490));
 sg13g2_tiehi _6792__491 (.L_HI(net491));
 sg13g2_tiehi _7100__492 (.L_HI(net492));
 sg13g2_tiehi _6791__493 (.L_HI(net493));
 sg13g2_tiehi _7067__494 (.L_HI(net494));
 sg13g2_tiehi _6790__495 (.L_HI(net495));
 sg13g2_tiehi _7099__496 (.L_HI(net496));
 sg13g2_tiehi _6789__497 (.L_HI(net497));
 sg13g2_tiehi _7066__498 (.L_HI(net498));
 sg13g2_tiehi _6788__499 (.L_HI(net499));
 sg13g2_tiehi _7061__500 (.L_HI(net500));
 sg13g2_tiehi _6787__501 (.L_HI(net501));
 sg13g2_tiehi _7065__502 (.L_HI(net502));
 sg13g2_tiehi _6786__503 (.L_HI(net503));
 sg13g2_tiehi _7098__504 (.L_HI(net504));
 sg13g2_tiehi _6785__505 (.L_HI(net505));
 sg13g2_tiehi _7064__506 (.L_HI(net506));
 sg13g2_tiehi _6784__507 (.L_HI(net507));
 sg13g2_tiehi _7097__508 (.L_HI(net508));
 sg13g2_tiehi _6783__509 (.L_HI(net509));
 sg13g2_tiehi _7063__510 (.L_HI(net510));
 sg13g2_tiehi _6782__511 (.L_HI(net511));
 sg13g2_tiehi _7096__512 (.L_HI(net512));
 sg13g2_tiehi _6781__513 (.L_HI(net513));
 sg13g2_tiehi _7062__514 (.L_HI(net514));
 sg13g2_tiehi _6780__515 (.L_HI(net515));
 sg13g2_tiehi _7095__516 (.L_HI(net516));
 sg13g2_tiehi _6779__517 (.L_HI(net517));
 sg13g2_tiehi _7055__518 (.L_HI(net518));
 sg13g2_tiehi _6778__519 (.L_HI(net519));
 sg13g2_tiehi _7094__520 (.L_HI(net520));
 sg13g2_tiehi _6777__521 (.L_HI(net521));
 sg13g2_tiehi _7054__522 (.L_HI(net522));
 sg13g2_tiehi _6776__523 (.L_HI(net523));
 sg13g2_tiehi _6679__524 (.L_HI(net524));
 sg13g2_tiehi _7056__525 (.L_HI(net525));
 sg13g2_tiehi _7057__526 (.L_HI(net526));
 sg13g2_tiehi _7058__527 (.L_HI(net527));
 sg13g2_tiehi _7059__528 (.L_HI(net528));
 sg13g2_tiehi _7060__529 (.L_HI(net529));
 sg13g2_tiehi _7053__530 (.L_HI(net530));
 sg13g2_tiehi _6775__531 (.L_HI(net531));
 sg13g2_tiehi _7093__532 (.L_HI(net532));
 sg13g2_tiehi _6774__533 (.L_HI(net533));
 sg13g2_tiehi _7052__534 (.L_HI(net534));
 sg13g2_tiehi _6773__535 (.L_HI(net535));
 sg13g2_tiehi _7092__536 (.L_HI(net536));
 sg13g2_tiehi _6772__537 (.L_HI(net537));
 sg13g2_tiehi _7051__538 (.L_HI(net538));
 sg13g2_tiehi _6771__539 (.L_HI(net539));
 sg13g2_tiehi _7091__540 (.L_HI(net540));
 sg13g2_tiehi _6770__541 (.L_HI(net541));
 sg13g2_tiehi _7050__542 (.L_HI(net542));
 sg13g2_tiehi _6769__543 (.L_HI(net543));
 sg13g2_tiehi _7090__544 (.L_HI(net544));
 sg13g2_tiehi _6768__545 (.L_HI(net545));
 sg13g2_tiehi _7049__546 (.L_HI(net546));
 sg13g2_tiehi _6767__547 (.L_HI(net547));
 sg13g2_tiehi _7089__548 (.L_HI(net548));
 sg13g2_tiehi _6766__549 (.L_HI(net549));
 sg13g2_tiehi _7048__550 (.L_HI(net550));
 sg13g2_tiehi _6765__551 (.L_HI(net551));
 sg13g2_tiehi _7088__552 (.L_HI(net552));
 sg13g2_tiehi _6764__553 (.L_HI(net553));
 sg13g2_tiehi _7047__554 (.L_HI(net554));
 sg13g2_tiehi _6763__555 (.L_HI(net555));
 sg13g2_tiehi _6762__556 (.L_HI(net556));
 sg13g2_tiehi _6761__557 (.L_HI(net557));
 sg13g2_tiehi _6760__558 (.L_HI(net558));
 sg13g2_tiehi _6759__559 (.L_HI(net559));
 sg13g2_tiehi _6758__560 (.L_HI(net560));
 sg13g2_tiehi _6757__561 (.L_HI(net561));
 sg13g2_tiehi _6756__562 (.L_HI(net562));
 sg13g2_tiehi _6755__563 (.L_HI(net563));
 sg13g2_tiehi _6754__564 (.L_HI(net564));
 sg13g2_tiehi _6753__565 (.L_HI(net565));
 sg13g2_tiehi _6752__566 (.L_HI(net566));
 sg13g2_tiehi _6751__567 (.L_HI(net567));
 sg13g2_tiehi _6750__568 (.L_HI(net568));
 sg13g2_tiehi _6749__569 (.L_HI(net569));
 sg13g2_tiehi _6748__570 (.L_HI(net570));
 sg13g2_tiehi _6747__571 (.L_HI(net571));
 sg13g2_tiehi _6746__572 (.L_HI(net572));
 sg13g2_tiehi _6745__573 (.L_HI(net573));
 sg13g2_tiehi _6744__574 (.L_HI(net574));
 sg13g2_tiehi _6743__575 (.L_HI(net575));
 sg13g2_tiehi _6742__576 (.L_HI(net576));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_5 (.L_LO(net5));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_6 (.L_LO(net6));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_7 (.L_LO(net7));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_8 (.L_LO(net8));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_9 (.L_LO(net9));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_10 (.L_LO(net10));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_11 (.L_LO(net11));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_12 (.L_LO(net12));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_13 (.L_LO(net13));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_14 (.L_LO(net14));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_15 (.L_LO(net15));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_16 (.L_LO(net16));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_17 (.L_LO(net17));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_18 (.L_LO(net18));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_19 (.L_LO(net19));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_20 (.L_LO(net20));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_21 (.L_LO(net21));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_22 (.L_LO(net22));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_23 (.L_LO(net23));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_24 (.L_LO(net24));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_25 (.L_LO(net25));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_26 (.L_LO(net26));
 sg13g2_tiehi _6741__27 (.L_HI(net27));
 sg13g2_buf_1 _7683_ (.A(\main.SPI_out ),
    .X(uo_out[0]));
 sg13g2_buf_2 fanout1050 (.A(net1054),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(net1052),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(net1054),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(net1054),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(_1444_),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_1326_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(_1399_),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_1399_),
    .X(net1057));
 sg13g2_buf_4 fanout1058 (.X(net1058),
    .A(net1063));
 sg13g2_buf_1 fanout1059 (.A(net1063),
    .X(net1059));
 sg13g2_buf_4 fanout1060 (.X(net1060),
    .A(net1063));
 sg13g2_buf_4 fanout1061 (.X(net1061),
    .A(net1062));
 sg13g2_buf_4 fanout1062 (.X(net1062),
    .A(net1063));
 sg13g2_buf_2 fanout1063 (.A(net1069),
    .X(net1063));
 sg13g2_buf_4 fanout1064 (.X(net1064),
    .A(net1069));
 sg13g2_buf_2 fanout1065 (.A(net1068),
    .X(net1065));
 sg13g2_buf_4 fanout1066 (.X(net1066),
    .A(net1068));
 sg13g2_buf_2 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(net1069),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(_2578_),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(net1071),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(_1137_),
    .X(net1071));
 sg13g2_buf_2 fanout1072 (.A(_1136_),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(net1074),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(net1075),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(_1361_),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(net1077),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_1043_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(net1079),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(net1080),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(_1028_),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(_1019_),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(_1019_),
    .X(net1082));
 sg13g2_buf_2 fanout1083 (.A(net1084),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(_0999_),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(net1086),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(net1087),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_0990_),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(_0981_),
    .X(net1088));
 sg13g2_buf_2 fanout1089 (.A(_0981_),
    .X(net1089));
 sg13g2_buf_2 fanout1090 (.A(_0973_),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(_0973_),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(net1093),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(_0942_),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(_0866_),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(_0866_),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(net1097),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(net1098),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(_0854_),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(_0842_),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(_0842_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(_0835_),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(_0835_),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(_0823_),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(_0823_),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(net1106),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(_0815_),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(net1108),
    .X(net1107));
 sg13g2_buf_1 fanout1108 (.A(net1109),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(_1086_),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(_1011_),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(_1011_),
    .X(net1111));
 sg13g2_buf_4 fanout1112 (.X(net1112),
    .A(_1090_));
 sg13g2_buf_2 fanout1113 (.A(_1090_),
    .X(net1113));
 sg13g2_buf_4 fanout1114 (.X(net1114),
    .A(net1115));
 sg13g2_buf_2 fanout1115 (.A(_1089_),
    .X(net1115));
 sg13g2_buf_4 fanout1116 (.X(net1116),
    .A(net1117));
 sg13g2_buf_2 fanout1117 (.A(_1089_),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(net1119),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(_1088_),
    .X(net1119));
 sg13g2_buf_2 fanout1120 (.A(net1121),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(_1084_),
    .X(net1121));
 sg13g2_buf_4 fanout1122 (.X(net1122),
    .A(net1123));
 sg13g2_buf_4 fanout1123 (.X(net1123),
    .A(net1124));
 sg13g2_buf_4 fanout1124 (.X(net1124),
    .A(_0809_));
 sg13g2_buf_4 fanout1125 (.X(net1125),
    .A(net1126));
 sg13g2_buf_4 fanout1126 (.X(net1126),
    .A(_0809_));
 sg13g2_buf_4 fanout1127 (.X(net1127),
    .A(_1066_));
 sg13g2_buf_2 fanout1128 (.A(_2685_),
    .X(net1128));
 sg13g2_buf_2 fanout1129 (.A(_1887_),
    .X(net1129));
 sg13g2_buf_2 fanout1130 (.A(_1887_),
    .X(net1130));
 sg13g2_buf_2 fanout1131 (.A(_1817_),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(net1133),
    .X(net1132));
 sg13g2_buf_2 fanout1133 (.A(_1500_),
    .X(net1133));
 sg13g2_buf_2 fanout1134 (.A(net1137),
    .X(net1134));
 sg13g2_buf_1 fanout1135 (.A(net1137),
    .X(net1135));
 sg13g2_buf_2 fanout1136 (.A(net1137),
    .X(net1136));
 sg13g2_buf_1 fanout1137 (.A(_1864_),
    .X(net1137));
 sg13g2_buf_4 fanout1138 (.X(net1138),
    .A(net1139));
 sg13g2_buf_4 fanout1139 (.X(net1139),
    .A(net1140));
 sg13g2_buf_1 fanout1140 (.A(net1141),
    .X(net1140));
 sg13g2_buf_2 fanout1141 (.A(net1142),
    .X(net1141));
 sg13g2_buf_2 fanout1142 (.A(_1829_),
    .X(net1142));
 sg13g2_buf_2 fanout1143 (.A(net1144),
    .X(net1143));
 sg13g2_buf_2 fanout1144 (.A(net1145),
    .X(net1144));
 sg13g2_buf_2 fanout1145 (.A(_1828_),
    .X(net1145));
 sg13g2_buf_4 fanout1146 (.X(net1146),
    .A(net1149));
 sg13g2_buf_1 fanout1147 (.A(net1149),
    .X(net1147));
 sg13g2_buf_2 fanout1148 (.A(net1149),
    .X(net1148));
 sg13g2_buf_1 fanout1149 (.A(_1827_),
    .X(net1149));
 sg13g2_buf_2 fanout1150 (.A(net1152),
    .X(net1150));
 sg13g2_buf_4 fanout1151 (.X(net1151),
    .A(net1152));
 sg13g2_buf_2 fanout1152 (.A(_1826_),
    .X(net1152));
 sg13g2_buf_4 fanout1153 (.X(net1153),
    .A(net1154));
 sg13g2_buf_2 fanout1154 (.A(net1155),
    .X(net1154));
 sg13g2_buf_2 fanout1155 (.A(_1825_),
    .X(net1155));
 sg13g2_buf_2 fanout1156 (.A(net1157),
    .X(net1156));
 sg13g2_buf_2 fanout1157 (.A(_1824_),
    .X(net1157));
 sg13g2_buf_2 fanout1158 (.A(net1160),
    .X(net1158));
 sg13g2_buf_2 fanout1159 (.A(net1160),
    .X(net1159));
 sg13g2_buf_4 fanout1160 (.X(net1160),
    .A(_1823_));
 sg13g2_buf_2 fanout1161 (.A(net1162),
    .X(net1161));
 sg13g2_buf_2 fanout1162 (.A(_1518_),
    .X(net1162));
 sg13g2_buf_1 fanout1163 (.A(_1518_),
    .X(net1163));
 sg13g2_buf_2 fanout1164 (.A(net1165),
    .X(net1164));
 sg13g2_buf_1 fanout1165 (.A(net1170),
    .X(net1165));
 sg13g2_buf_2 fanout1166 (.A(net1170),
    .X(net1166));
 sg13g2_buf_2 fanout1167 (.A(net1168),
    .X(net1167));
 sg13g2_buf_2 fanout1168 (.A(net1169),
    .X(net1168));
 sg13g2_buf_2 fanout1169 (.A(net1170),
    .X(net1169));
 sg13g2_buf_1 fanout1170 (.A(_1517_),
    .X(net1170));
 sg13g2_buf_2 fanout1171 (.A(net1174),
    .X(net1171));
 sg13g2_buf_2 fanout1172 (.A(net1174),
    .X(net1172));
 sg13g2_buf_2 fanout1173 (.A(net1174),
    .X(net1173));
 sg13g2_buf_1 fanout1174 (.A(_1512_),
    .X(net1174));
 sg13g2_buf_4 fanout1175 (.X(net1175),
    .A(net1176));
 sg13g2_buf_2 fanout1176 (.A(net1181),
    .X(net1176));
 sg13g2_buf_4 fanout1177 (.X(net1177),
    .A(net1180));
 sg13g2_buf_2 fanout1178 (.A(net1179),
    .X(net1178));
 sg13g2_buf_2 fanout1179 (.A(net1180),
    .X(net1179));
 sg13g2_buf_1 fanout1180 (.A(net1181),
    .X(net1180));
 sg13g2_buf_2 fanout1181 (.A(_1511_),
    .X(net1181));
 sg13g2_buf_4 fanout1182 (.X(net1182),
    .A(net1183));
 sg13g2_buf_2 fanout1183 (.A(net1184),
    .X(net1183));
 sg13g2_buf_2 fanout1184 (.A(_1507_),
    .X(net1184));
 sg13g2_buf_4 fanout1185 (.X(net1185),
    .A(net1187));
 sg13g2_buf_1 fanout1186 (.A(net1187),
    .X(net1186));
 sg13g2_buf_4 fanout1187 (.X(net1187),
    .A(net1188));
 sg13g2_buf_4 fanout1188 (.X(net1188),
    .A(_1506_));
 sg13g2_buf_4 fanout1189 (.X(net1189),
    .A(net1190));
 sg13g2_buf_2 fanout1190 (.A(net1191),
    .X(net1190));
 sg13g2_buf_4 fanout1191 (.X(net1191),
    .A(_1506_));
 sg13g2_buf_2 fanout1192 (.A(net1193),
    .X(net1192));
 sg13g2_buf_2 fanout1193 (.A(_1505_),
    .X(net1193));
 sg13g2_buf_2 fanout1194 (.A(_1505_),
    .X(net1194));
 sg13g2_buf_2 fanout1195 (.A(_1505_),
    .X(net1195));
 sg13g2_buf_2 fanout1196 (.A(net1201),
    .X(net1196));
 sg13g2_buf_2 fanout1197 (.A(net1201),
    .X(net1197));
 sg13g2_buf_2 fanout1198 (.A(net1199),
    .X(net1198));
 sg13g2_buf_1 fanout1199 (.A(net1200),
    .X(net1199));
 sg13g2_buf_2 fanout1200 (.A(net1201),
    .X(net1200));
 sg13g2_buf_2 fanout1201 (.A(_1504_),
    .X(net1201));
 sg13g2_buf_2 fanout1202 (.A(net1203),
    .X(net1202));
 sg13g2_buf_2 fanout1203 (.A(net1206),
    .X(net1203));
 sg13g2_buf_2 fanout1204 (.A(net1206),
    .X(net1204));
 sg13g2_buf_1 fanout1205 (.A(net1206),
    .X(net1205));
 sg13g2_buf_1 fanout1206 (.A(_1502_),
    .X(net1206));
 sg13g2_buf_2 fanout1207 (.A(net1208),
    .X(net1207));
 sg13g2_buf_2 fanout1208 (.A(_1501_),
    .X(net1208));
 sg13g2_buf_2 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_2 fanout1210 (.A(_0807_),
    .X(net1210));
 sg13g2_buf_2 fanout1211 (.A(net1212),
    .X(net1211));
 sg13g2_buf_2 fanout1212 (.A(net1213),
    .X(net1212));
 sg13g2_buf_2 fanout1213 (.A(_0807_),
    .X(net1213));
 sg13g2_buf_2 fanout1214 (.A(net1216),
    .X(net1214));
 sg13g2_buf_2 fanout1215 (.A(net1216),
    .X(net1215));
 sg13g2_buf_2 fanout1216 (.A(_0807_),
    .X(net1216));
 sg13g2_buf_2 fanout1217 (.A(_0806_),
    .X(net1217));
 sg13g2_buf_2 fanout1218 (.A(net1220),
    .X(net1218));
 sg13g2_buf_1 fanout1219 (.A(net1220),
    .X(net1219));
 sg13g2_buf_2 fanout1220 (.A(_1370_),
    .X(net1220));
 sg13g2_buf_4 fanout1221 (.X(net1221),
    .A(_0793_));
 sg13g2_buf_4 fanout1222 (.X(net1222),
    .A(_0792_));
 sg13g2_buf_4 fanout1223 (.X(net1223),
    .A(_0777_));
 sg13g2_buf_2 fanout1224 (.A(_0770_),
    .X(net1224));
 sg13g2_buf_2 fanout1225 (.A(_0765_),
    .X(net1225));
 sg13g2_buf_4 fanout1226 (.X(net1226),
    .A(net1228));
 sg13g2_buf_4 fanout1227 (.X(net1227),
    .A(net1228));
 sg13g2_buf_2 fanout1228 (.A(_0001_),
    .X(net1228));
 sg13g2_buf_4 fanout1229 (.X(net1229),
    .A(net1230));
 sg13g2_buf_4 fanout1230 (.X(net1230),
    .A(_0001_));
 sg13g2_buf_8 fanout1231 (.A(net1233),
    .X(net1231));
 sg13g2_buf_8 fanout1232 (.A(net1233),
    .X(net1232));
 sg13g2_buf_4 fanout1233 (.X(net1233),
    .A(_0000_));
 sg13g2_buf_8 fanout1234 (.A(net1235),
    .X(net1234));
 sg13g2_buf_8 fanout1235 (.A(_0000_),
    .X(net1235));
 sg13g2_buf_4 fanout1236 (.X(net1236),
    .A(net1238));
 sg13g2_buf_2 fanout1237 (.A(net1238),
    .X(net1237));
 sg13g2_buf_4 fanout1238 (.X(net1238),
    .A(_0003_));
 sg13g2_buf_4 fanout1239 (.X(net1239),
    .A(net1240));
 sg13g2_buf_4 fanout1240 (.X(net1240),
    .A(_0003_));
 sg13g2_buf_8 fanout1241 (.A(net1243),
    .X(net1241));
 sg13g2_buf_4 fanout1242 (.X(net1242),
    .A(net1243));
 sg13g2_buf_8 fanout1243 (.A(_0002_),
    .X(net1243));
 sg13g2_buf_8 fanout1244 (.A(net1245),
    .X(net1244));
 sg13g2_buf_8 fanout1245 (.A(_0002_),
    .X(net1245));
 sg13g2_buf_4 fanout1246 (.X(net1246),
    .A(net665));
 sg13g2_buf_4 fanout1247 (.X(net1247),
    .A(net761));
 sg13g2_buf_1 fanout1248 (.A(net761),
    .X(net1248));
 sg13g2_buf_4 fanout1249 (.X(net1249),
    .A(net678));
 sg13g2_buf_2 fanout1250 (.A(net1251),
    .X(net1250));
 sg13g2_buf_1 fanout1251 (.A(net1455),
    .X(net1251));
 sg13g2_buf_2 fanout1252 (.A(net1259),
    .X(net1252));
 sg13g2_buf_1 fanout1253 (.A(net1259),
    .X(net1253));
 sg13g2_buf_2 fanout1254 (.A(net1256),
    .X(net1254));
 sg13g2_buf_1 fanout1255 (.A(net1256),
    .X(net1255));
 sg13g2_buf_2 fanout1256 (.A(net1259),
    .X(net1256));
 sg13g2_buf_2 fanout1257 (.A(net1258),
    .X(net1257));
 sg13g2_buf_4 fanout1258 (.X(net1258),
    .A(net1259));
 sg13g2_buf_4 fanout1259 (.X(net1259),
    .A(\main.adder.s2_flip_sign ));
 sg13g2_buf_2 fanout1260 (.A(net1262),
    .X(net1260));
 sg13g2_buf_1 fanout1261 (.A(net1262),
    .X(net1261));
 sg13g2_buf_2 fanout1262 (.A(_0015_),
    .X(net1262));
 sg13g2_buf_4 fanout1263 (.X(net1263),
    .A(net1265));
 sg13g2_buf_4 fanout1264 (.X(net1264),
    .A(net1265));
 sg13g2_buf_2 fanout1265 (.A(_0005_),
    .X(net1265));
 sg13g2_buf_4 fanout1266 (.X(net1266),
    .A(net1267));
 sg13g2_buf_4 fanout1267 (.X(net1267),
    .A(_0005_));
 sg13g2_buf_8 fanout1268 (.A(net1270),
    .X(net1268));
 sg13g2_buf_8 fanout1269 (.A(net1270),
    .X(net1269));
 sg13g2_buf_4 fanout1270 (.X(net1270),
    .A(_0004_));
 sg13g2_buf_8 fanout1271 (.A(net1272),
    .X(net1271));
 sg13g2_buf_8 fanout1272 (.A(_0004_),
    .X(net1272));
 sg13g2_buf_2 fanout1273 (.A(\main.SPI_input_data_valid ),
    .X(net1273));
 sg13g2_buf_2 fanout1274 (.A(net1577),
    .X(net1274));
 sg13g2_buf_2 fanout1275 (.A(net1277),
    .X(net1275));
 sg13g2_buf_1 fanout1276 (.A(net1277),
    .X(net1276));
 sg13g2_buf_2 fanout1277 (.A(net1595),
    .X(net1277));
 sg13g2_buf_2 fanout1278 (.A(net1279),
    .X(net1278));
 sg13g2_buf_2 fanout1279 (.A(net1280),
    .X(net1279));
 sg13g2_buf_1 fanout1280 (.A(net1281),
    .X(net1280));
 sg13g2_buf_2 fanout1281 (.A(net1610),
    .X(net1281));
 sg13g2_buf_4 fanout1282 (.X(net1282),
    .A(net1619));
 sg13g2_buf_2 fanout1283 (.A(net1284),
    .X(net1283));
 sg13g2_buf_1 fanout1284 (.A(\main.byte_counter[0] ),
    .X(net1284));
 sg13g2_buf_2 fanout1285 (.A(net1287),
    .X(net1285));
 sg13g2_buf_1 fanout1286 (.A(net1287),
    .X(net1286));
 sg13g2_buf_2 fanout1287 (.A(net1288),
    .X(net1287));
 sg13g2_buf_2 fanout1288 (.A(\main.byte_counter[0] ),
    .X(net1288));
 sg13g2_buf_2 fanout1289 (.A(net1290),
    .X(net1289));
 sg13g2_buf_2 fanout1290 (.A(net1291),
    .X(net1290));
 sg13g2_buf_1 fanout1291 (.A(net1606),
    .X(net1291));
 sg13g2_buf_2 fanout1292 (.A(net1296),
    .X(net1292));
 sg13g2_buf_2 fanout1293 (.A(net1294),
    .X(net1293));
 sg13g2_buf_1 fanout1294 (.A(net1295),
    .X(net1294));
 sg13g2_buf_1 fanout1295 (.A(net1296),
    .X(net1295));
 sg13g2_buf_1 fanout1296 (.A(\main.byte_counter[1] ),
    .X(net1296));
 sg13g2_buf_2 fanout1297 (.A(net1298),
    .X(net1297));
 sg13g2_buf_2 fanout1298 (.A(net1322),
    .X(net1298));
 sg13g2_buf_2 fanout1299 (.A(net1300),
    .X(net1299));
 sg13g2_buf_2 fanout1300 (.A(net1304),
    .X(net1300));
 sg13g2_buf_2 fanout1301 (.A(net1303),
    .X(net1301));
 sg13g2_buf_2 fanout1302 (.A(net1303),
    .X(net1302));
 sg13g2_buf_2 fanout1303 (.A(net1304),
    .X(net1303));
 sg13g2_buf_2 fanout1304 (.A(net1322),
    .X(net1304));
 sg13g2_buf_2 fanout1305 (.A(net1307),
    .X(net1305));
 sg13g2_buf_1 fanout1306 (.A(net1307),
    .X(net1306));
 sg13g2_buf_2 fanout1307 (.A(net1308),
    .X(net1307));
 sg13g2_buf_2 fanout1308 (.A(net1309),
    .X(net1308));
 sg13g2_buf_2 fanout1309 (.A(net1310),
    .X(net1309));
 sg13g2_buf_4 fanout1310 (.X(net1310),
    .A(net1322));
 sg13g2_buf_2 fanout1311 (.A(net1313),
    .X(net1311));
 sg13g2_buf_1 fanout1312 (.A(net1313),
    .X(net1312));
 sg13g2_buf_4 fanout1313 (.X(net1313),
    .A(net1314));
 sg13g2_buf_2 fanout1314 (.A(net1322),
    .X(net1314));
 sg13g2_buf_2 fanout1315 (.A(net1316),
    .X(net1315));
 sg13g2_buf_1 fanout1316 (.A(net1320),
    .X(net1316));
 sg13g2_buf_2 fanout1317 (.A(net1318),
    .X(net1317));
 sg13g2_buf_1 fanout1318 (.A(net1319),
    .X(net1318));
 sg13g2_buf_2 fanout1319 (.A(net1320),
    .X(net1319));
 sg13g2_buf_1 fanout1320 (.A(net1321),
    .X(net1320));
 sg13g2_buf_4 fanout1321 (.X(net1321),
    .A(net1322));
 sg13g2_buf_4 fanout1322 (.X(net1322),
    .A(_0700_));
 sg13g2_buf_4 fanout1323 (.X(net1323),
    .A(net1328));
 sg13g2_buf_4 fanout1324 (.X(net1324),
    .A(net1327));
 sg13g2_buf_4 fanout1325 (.X(net1325),
    .A(net1327));
 sg13g2_buf_2 fanout1326 (.A(net1327),
    .X(net1326));
 sg13g2_buf_2 fanout1327 (.A(net1328),
    .X(net1327));
 sg13g2_buf_4 fanout1328 (.X(net1328),
    .A(net1337));
 sg13g2_buf_4 fanout1329 (.X(net1329),
    .A(net1331));
 sg13g2_buf_2 fanout1330 (.A(net1331),
    .X(net1330));
 sg13g2_buf_2 fanout1331 (.A(net1332),
    .X(net1331));
 sg13g2_buf_2 fanout1332 (.A(net1337),
    .X(net1332));
 sg13g2_buf_4 fanout1333 (.X(net1333),
    .A(net1334));
 sg13g2_buf_4 fanout1334 (.X(net1334),
    .A(net1335));
 sg13g2_buf_2 fanout1335 (.A(net1337),
    .X(net1335));
 sg13g2_buf_4 fanout1336 (.X(net1336),
    .A(net1337));
 sg13g2_buf_2 fanout1337 (.A(net1346),
    .X(net1337));
 sg13g2_buf_2 fanout1338 (.A(net1340),
    .X(net1338));
 sg13g2_buf_2 fanout1339 (.A(net1340),
    .X(net1339));
 sg13g2_buf_2 fanout1340 (.A(net1341),
    .X(net1340));
 sg13g2_buf_2 fanout1341 (.A(net1346),
    .X(net1341));
 sg13g2_buf_4 fanout1342 (.X(net1342),
    .A(net1343));
 sg13g2_buf_2 fanout1343 (.A(net1346),
    .X(net1343));
 sg13g2_buf_2 fanout1344 (.A(net1345),
    .X(net1344));
 sg13g2_buf_4 fanout1345 (.X(net1345),
    .A(net1346));
 sg13g2_buf_4 fanout1346 (.X(net1346),
    .A(rst_n));
 sg13g2_buf_2 fanout1347 (.A(net1351),
    .X(net1347));
 sg13g2_buf_1 fanout1348 (.A(net1351),
    .X(net1348));
 sg13g2_buf_2 fanout1349 (.A(net1351),
    .X(net1349));
 sg13g2_buf_2 fanout1350 (.A(net1351),
    .X(net1350));
 sg13g2_buf_2 fanout1351 (.A(net1395),
    .X(net1351));
 sg13g2_buf_2 fanout1352 (.A(net1354),
    .X(net1352));
 sg13g2_buf_1 fanout1353 (.A(net1354),
    .X(net1353));
 sg13g2_buf_4 fanout1354 (.X(net1354),
    .A(net1360));
 sg13g2_buf_2 fanout1355 (.A(net1360),
    .X(net1355));
 sg13g2_buf_2 fanout1356 (.A(net1360),
    .X(net1356));
 sg13g2_buf_2 fanout1357 (.A(net1359),
    .X(net1357));
 sg13g2_buf_2 fanout1358 (.A(net1359),
    .X(net1358));
 sg13g2_buf_2 fanout1359 (.A(net1360),
    .X(net1359));
 sg13g2_buf_2 fanout1360 (.A(net1395),
    .X(net1360));
 sg13g2_buf_4 fanout1361 (.X(net1361),
    .A(net1378));
 sg13g2_buf_2 fanout1362 (.A(net1378),
    .X(net1362));
 sg13g2_buf_2 fanout1363 (.A(net1365),
    .X(net1363));
 sg13g2_buf_1 fanout1364 (.A(net1365),
    .X(net1364));
 sg13g2_buf_2 fanout1365 (.A(net1378),
    .X(net1365));
 sg13g2_buf_2 fanout1366 (.A(net1368),
    .X(net1366));
 sg13g2_buf_2 fanout1367 (.A(net1368),
    .X(net1367));
 sg13g2_buf_2 fanout1368 (.A(net1377),
    .X(net1368));
 sg13g2_buf_2 fanout1369 (.A(net1370),
    .X(net1369));
 sg13g2_buf_2 fanout1370 (.A(net1377),
    .X(net1370));
 sg13g2_buf_2 fanout1371 (.A(net1373),
    .X(net1371));
 sg13g2_buf_2 fanout1372 (.A(net1373),
    .X(net1372));
 sg13g2_buf_2 fanout1373 (.A(net1377),
    .X(net1373));
 sg13g2_buf_2 fanout1374 (.A(net1375),
    .X(net1374));
 sg13g2_buf_2 fanout1375 (.A(net1376),
    .X(net1375));
 sg13g2_buf_2 fanout1376 (.A(net1377),
    .X(net1376));
 sg13g2_buf_2 fanout1377 (.A(net1378),
    .X(net1377));
 sg13g2_buf_2 fanout1378 (.A(net1395),
    .X(net1378));
 sg13g2_buf_2 fanout1379 (.A(net1382),
    .X(net1379));
 sg13g2_buf_4 fanout1380 (.X(net1380),
    .A(net1381));
 sg13g2_buf_2 fanout1381 (.A(net1382),
    .X(net1381));
 sg13g2_buf_2 fanout1382 (.A(net1389),
    .X(net1382));
 sg13g2_buf_4 fanout1383 (.X(net1383),
    .A(net1385));
 sg13g2_buf_4 fanout1384 (.X(net1384),
    .A(net1385));
 sg13g2_buf_2 fanout1385 (.A(net1389),
    .X(net1385));
 sg13g2_buf_2 fanout1386 (.A(net1387),
    .X(net1386));
 sg13g2_buf_2 fanout1387 (.A(net1389),
    .X(net1387));
 sg13g2_buf_4 fanout1388 (.X(net1388),
    .A(net1389));
 sg13g2_buf_2 fanout1389 (.A(net1395),
    .X(net1389));
 sg13g2_buf_2 fanout1390 (.A(net1394),
    .X(net1390));
 sg13g2_buf_2 fanout1391 (.A(net1394),
    .X(net1391));
 sg13g2_buf_4 fanout1392 (.X(net1392),
    .A(net1394));
 sg13g2_buf_2 fanout1393 (.A(net1394),
    .X(net1393));
 sg13g2_buf_2 fanout1394 (.A(net1395),
    .X(net1394));
 sg13g2_buf_4 fanout1395 (.X(net1395),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_tielo tt_um_Qwendu_spi_fpu_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_3_0_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_4_4_0_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_4_5_0_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_4_8_0_clk));
 sg13g2_buf_1 clkload9 (.A(clknet_4_9_0_clk));
 sg13g2_buf_1 clkload10 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_11_0_clk));
 sg13g2_buf_1 clkload12 (.A(clknet_4_12_0_clk));
 sg13g2_buf_1 clkload13 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_0_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_5_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_11_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_68_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_14_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_20_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_9_clk));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_27_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_24_clk));
 sg13g2_inv_4 clkload24 (.A(clknet_leaf_61_clk));
 sg13g2_inv_8 clkload25 (.A(clknet_leaf_57_clk));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_58_clk));
 sg13g2_inv_2 clkload27 (.A(clknet_leaf_44_clk));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_52_clk));
 sg13g2_inv_2 clkload29 (.A(clknet_leaf_36_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_41_clk));
 sg13g2_inv_4 clkload31 (.A(clknet_leaf_42_clk));
 sg13g2_inv_1 clkload32 (.A(clknet_leaf_31_clk));
 sg13g2_inv_4 clkload33 (.A(clknet_leaf_37_clk));
 sg13g2_inv_4 clkload34 (.A(clknet_leaf_45_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\main.spi.SPI_not_chip_select_sampler.sample_register[0] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0522_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold3 (.A(\main.adder.s4_valid ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold4 (.A(\main.adder.s3_valid ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold5 (.A(\main.adder.s5_valid ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0124_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0614_),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold8 (.A(\main.adder.s1_valid ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold9 (.A(\main.adder.s2_valid ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold10 (.A(\main.adder.s4_mant[8] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0412_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold12 (.A(\main.state[0] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0009_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold14 (.A(\main.adder.s4_mant[17] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0421_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold16 (.A(\main.adder.s4_mant[12] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold17 (.A(\main.adder.s4_mant[9] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0413_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold19 (.A(\main.adder.s4_mant[10] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0414_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold21 (.A(\main.adder.s4_mant[6] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0410_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold23 (.A(\main.adder.s4_mant[18] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0422_),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold25 (.A(\main.adder.s2_exponent[3] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0248_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold27 (.A(\main.adder.s4_mant[16] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0420_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold29 (.A(\main.adder.s4_mant[5] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0409_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold31 (.A(\main.adder.s4_mant[19] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0423_),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold33 (.A(\main.adder.s4_mant[1] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0405_),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold35 (.A(\main.adder.s4_mant[13] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0417_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold37 (.A(\main.adder.s4_mant[3] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0407_),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold39 (.A(\main.spi.SPI_in_sampled ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0617_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold41 (.A(\main.adder.s4_mant[20] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0424_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold43 (.A(\main.adder.s1_rs.levels[0][33] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold44 (.A(\main.adder.s1_rs.levels[0][34] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold45 (.A(\main.adder.s4_mant[11] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0415_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold47 (.A(\main.adder.s1_rs.levels[0][41] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold48 (.A(\main.adder.s4_mant[14] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold49 (.A(\main.adder.s4_mant[15] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0419_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold51 (.A(\main.register_id_input_b[0] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0658_),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold53 (.A(\main.adder.s1_rs.levels[0][43] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold54 (.A(\main.adder.s1_rs.levels[0][45] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold55 (.A(\main.adder.s5_sign ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0375_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold57 (.A(\main.adder.s4_mant[0] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0452_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold59 (.A(\main.adder.s4_mant[2] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0406_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold61 (.A(\main.adder.s4_mant[38] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold62 (.A(\main.adder.s1_rs.levels[0][37] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold63 (.A(\main.adder.s1_larger[3] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0302_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold65 (.A(\main.adder.s1_rs.levels[0][25] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold66 (.A(\main.adder.s1_rs.levels[0][40] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold67 (.A(\main.adder.s1_rs.levels[0][36] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold68 (.A(\main.adder.s1_rs.levels[0][27] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold69 (.A(\main.adder.s1_rs.levels[0][32] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold70 (.A(\main.adder.s1_rs.levels[0][38] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold71 (.A(\main.adder.s1_rs.levels[0][26] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold72 (.A(\main.adder.s1_rs.levels[0][42] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold73 (.A(\main.adder.s4_mant[36] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold74 (.A(\main.adder.s1_rs.levels[0][30] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold75 (.A(\main.adder.s1_rs.levels[0][31] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold76 (.A(\main.adder.s1_rs.levels[0][35] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold77 (.A(\main.adder.out[19] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0279_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold79 (.A(\main.adder.s1_rs.levels[0][29] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold80 (.A(\main.adder.out[18] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0278_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold82 (.A(\main.adder.s4_shared_sign ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold83 (.A(_2084_),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold84 (.A(\main.adder.s4_sum[48] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0453_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold86 (.A(\main.adder.s4_mant[7] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0411_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold88 (.A(\main.adder.s1_rs.levels[0][28] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold89 (.A(\main.SPI_input_data[0] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold90 (.A(\main.adder.s4_mant[4] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0408_),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold92 (.A(\main.adder.s1_rs.levels[0][39] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0125_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold94 (.A(_2679_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0601_),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold96 (.A(\main.adder.out[8] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0268_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold98 (.A(\main.adder.out[21] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0281_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold100 (.A(\main.adder.out[20] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0280_),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold102 (.A(\main.adder.s1_exp_diff[4] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold103 (.A(\main.adder.s5_R ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold104 (.A(\main.spi.out_data_r[3] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold105 (.A(_2721_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold106 (.A(\main.adder.s1_rs.levels[0][44] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold107 (.A(\main.adder.out[17] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0277_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold109 (.A(\main.adder.s1_rs.levels[0][24] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold110 (.A(\main.adder.s2_smaler[22] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold111 (.A(\main.adder.s1_exp_diff[9] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold112 (.A(\main.adder.s2_smaler[19] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold113 (.A(\main.adder.s3_sum[22] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold114 (.A(\main.adder.out[16] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0276_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold116 (.A(\main.register_id_input_b[1] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0659_),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold118 (.A(\main.adder.s2_smaler[1] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold119 (.A(\main.adder.out[22] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0282_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold121 (.A(\main.adder.s2_smaler[2] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold122 (.A(\main.adder.s1_larger[14] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0313_),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold124 (.A(\main.spi.in_bit_counter[2] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0616_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold126 (.A(\main.SPI_input_data[1] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold127 (.A(\main.adder.out[7] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0267_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold129 (.A(\main.adder.s2_smaler[12] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0471_),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold131 (.A(\main.adder.s3_sum[7] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0466_),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold133 (.A(\main.adder.out_valid ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0010_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold135 (.A(\main.adder.s1_larger[26] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold136 (.A(\main.register_id_input_a[1] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold137 (.A(\main.register_id_input_a[0] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold138 (.A(\main.adder.s2_smaler[0] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold139 (.A(\main.adder.s2_smaler[8] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold140 (.A(\main.adder.s3_sum[19] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold141 (.A(\main.adder.s1_exp_diff[8] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold142 (.A(\main.adder.s4_flipped ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0401_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold144 (.A(\main.adder.s1_nan ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0510_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold146 (.A(\main.adder.s1_smaler[25] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold147 (.A(\main.adder.s1_larger[21] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0320_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold149 (.A(\main.adder.s2_smaler[41] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold150 (.A(\main.adder.s2_shared_sign ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0458_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold152 (.A(\main.adder.s1_larger[0] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0299_),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold154 (.A(\main.adder.s2_smaler[6] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0465_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold156 (.A(\main.adder.s2_smaler[9] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold157 (.A(\main.adder.s1_smaler[23] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold158 (.A(\main.float_registers[1][3] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold159 (.A(\main.adder.out[6] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0266_),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold161 (.A(\main.adder.s2_exponent[1] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0246_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold163 (.A(\main.adder.s1_larger[19] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold164 (.A(\main.spi.out_data_r[5] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold165 (.A(_2737_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold166 (.A(\main.adder.s1_larger[24] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold167 (.A(\main.adder.s2_smaler[10] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold168 (.A(\main.spi.out_data_r[4] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold169 (.A(_2729_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold170 (.A(\main.adder.s1_larger[16] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0315_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold172 (.A(\main.adder.s2_smaler[43] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold173 (.A(\main.state[2] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0008_),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold175 (.A(\main.adder.s3_sum[8] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold176 (.A(\main.adder.s1_larger[2] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold177 (.A(\main.adder.s1_larger[4] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold178 (.A(\main.adder.out[15] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0275_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold180 (.A(\main.adder.s2_inf ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0511_),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold182 (.A(\main.adder.out[25] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0369_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold184 (.A(\main.adder.s1_larger[31] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold185 (.A(\main.adder.s1_exp_diff[5] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold186 (.A(\main.spi.out_data_r[7] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold187 (.A(_2753_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold188 (.A(\main.spi.SPI_in_sampler.sample_register[0] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold189 (.A(\main.adder.s2_exponent[2] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0516_),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold191 (.A(\main.adder.s1_smaler[24] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold192 (.A(\main.adder.s2_smaler[5] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold193 (.A(\main.adder.s1_smaler[26] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold194 (.A(\main.adder.s1_larger[6] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold195 (.A(\main.adder.s2_exponent[0] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0514_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold197 (.A(\main.float_registers[1][21] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold198 (.A(\main.adder.out[9] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0269_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold200 (.A(\main.adder.s3_sum[24] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold201 (.A(\main.adder.s2_smaler[4] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold202 (.A(\main.adder.s3_flipped ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold203 (.A(\main.adder.s3_inf ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold204 (.A(\main.adder.s4_nan ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0403_),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold206 (.A(\main.adder.s2_nan ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0455_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold208 (.A(\main.adder.s1_larger[7] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0306_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold210 (.A(\main.spi.out_data_r[1] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold211 (.A(_2705_),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold212 (.A(\main.adder.s2_exponent[6] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0251_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold214 (.A(\main.SPI_out ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold215 (.A(_2761_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0613_),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold217 (.A(\main.adder.s4_inf ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold218 (.A(\main.adder.s1_larger[10] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold219 (.A(\main.adder.s3_sum[9] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold220 (.A(\main.adder.out[10] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0270_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold222 (.A(\main.adder.s1_larger[12] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold223 (.A(\main.adder.s4_mant[21] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0425_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold225 (.A(\main.adder.s2_larger[27] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold226 (.A(\main.adder.s2_larger[33] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold227 (.A(\main.float_registers[0][28] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0158_),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold229 (.A(\main.adder.s5_mant[18] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold230 (.A(\main.adder.s2_larger[42] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold231 (.A(\main.adder.s2_smaler[7] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold232 (.A(\main.adder.s3_exponent[2] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold233 (.A(\main.adder.s4_exponent[3] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0256_),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold235 (.A(\main.float_registers[0][20] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold236 (.A(\main.float_registers[0][12] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold237 (.A(\main.adder.s1_smaler[31] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold238 (.A(\main.adder.s3_sum[5] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold239 (.A(\main.float_registers[0][16] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold240 (.A(\main.adder.s2_larger[29] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold241 (.A(\main.float_registers[0][14] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0154_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold243 (.A(\main.adder.s2_exponent[7] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0521_),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold245 (.A(\main.float_registers[0][5] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold246 (.A(\main.adder.s2_exponent[4] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0518_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold248 (.A(\main.adder.s4_mant[30] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0434_),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold250 (.A(\main.adder.s3_exponent[0] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold251 (.A(\main.float_registers[0][13] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold252 (.A(\main.adder.s5_nan ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold253 (.A(\main.adder.s3_shared_sign ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold254 (.A(\main.adder.s2_larger[25] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold255 (.A(\main.adder.s3_sum[4] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold256 (.A(\main.float_registers[0][11] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold257 (.A(\main.adder.s5_inf ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold258 (.A(\main.spi.out_data_r[6] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold259 (.A(_2745_),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold260 (.A(\main.adder.s1_smaler[30] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold261 (.A(\main.adder.out[13] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0273_),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold263 (.A(\main.float_registers[0][7] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold264 (.A(\main.float_registers[0][22] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold265 (.A(\main.adder.out[12] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0272_),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold267 (.A(\main.adder.s1_larger[11] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold268 (.A(\main.adder.s1_larger[29] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold269 (.A(\main.float_registers[0][19] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold270 (.A(\main.float_registers[0][2] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold271 (.A(\main.adder.s1_larger[22] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold272 (.A(\main.float_registers[0][21] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold273 (.A(\main.float_registers[0][17] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold274 (.A(\main.adder.s4_mant[34] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold275 (.A(\main.state[6] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0011_),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold277 (.A(\main.float_registers[0][6] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold278 (.A(\main.float_registers[0][26] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold279 (.A(\main.float_registers[0][23] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold280 (.A(\main.adder.s1_smaler[28] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold281 (.A(\main.adder.s1_larger[9] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold282 (.A(\main.adder.s2_larger[35] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold283 (.A(\main.adder.s1_larger[15] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0314_),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold285 (.A(\main.adder.s1_exp_diff[3] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold286 (.A(\main.float_registers[0][9] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0139_),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold288 (.A(\main.adder.s2_smaler[14] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0473_),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold290 (.A(\main.adder.s3_sum[0] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold291 (.A(\main.adder.s3_exponent[4] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold292 (.A(\main.adder.s1_larger[1] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0300_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold294 (.A(\main.adder.s2_larger[32] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold295 (.A(\main.float_registers[0][31] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0161_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold297 (.A(\main.adder.s2_larger[28] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0304_),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold299 (.A(\main.adder.s2_smaler[40] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold300 (.A(\main.adder.s1_larger[27] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold301 (.A(\main.adder.s3_sum[1] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold302 (.A(\main.float_registers[0][15] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold303 (.A(\main.adder.in_valid ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold304 (.A(\main.float_registers[0][25] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0155_),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold306 (.A(\main.float_registers[0][0] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold307 (.A(\main.adder.s2_smaler[13] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0472_),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold309 (.A(\main.adder.s2_smaler[44] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold310 (.A(\main.adder.out[24] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0368_),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold312 (.A(\main.spi.out_data_r[2] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold313 (.A(_2713_),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold314 (.A(\main.float_registers[0][30] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold315 (.A(\main.adder.s1_larger[13] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold316 (.A(\main.float_registers[1][1] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold317 (.A(\main.adder.out[11] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0271_),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold319 (.A(\main.float_registers[0][27] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0157_),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold321 (.A(\main.spi.out_data_r[0] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold322 (.A(_2697_),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold323 (.A(\main.adder.s2_smaler[38] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold324 (.A(\main.adder.s1_smaler[27] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold325 (.A(\main.adder.s1_larger[18] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0317_),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold327 (.A(\main.adder.s5_exponent[7] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold328 (.A(\main.adder.s3_sum[23] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0482_),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold330 (.A(\main.adder.s2_smaler[16] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0475_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold332 (.A(\main.adder.out[2] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0262_),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold334 (.A(\main.adder.s5_exponent[2] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold335 (.A(\main.adder.s1_smaler[29] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold336 (.A(\main.float_registers[0][10] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0145_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold338 (.A(\main.adder.s1_larger[8] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold339 (.A(\main.float_registers[0][8] ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold340 (.A(\main.adder.out[28] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0372_),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold342 (.A(\main.adder.s2_larger[36] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold343 (.A(\main.adder.s3_sum[2] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold344 (.A(\main.adder.out[5] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0265_),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold346 (.A(\main.adder.s2_exponent[5] ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0519_),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold348 (.A(\main.adder.s3_sum[10] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold349 (.A(\main.float_registers[0][18] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold350 (.A(\main.adder.s1_larger[5] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold351 (.A(\main.adder.s2_smaler[15] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0474_),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold353 (.A(\main.adder.s3_sum[3] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0462_),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold355 (.A(\main.adder.s2_larger[34] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold356 (.A(\main.float_registers[0][3] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold357 (.A(\main.adder.s2_larger[45] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold358 (.A(\main.adder.s5_exponent[6] ),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold359 (.A(\main.adder.s4_mant[32] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0436_),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold361 (.A(\main.float_registers[0][24] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold362 (.A(\main.adder.s4_mant[42] ),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0446_),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold364 (.A(\main.adder.s5_mant[9] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold365 (.A(\main.adder.out[14] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0274_),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold367 (.A(\main.adder.s1_larger[30] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold368 (.A(\main.adder.s2_smaler[31] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold369 (.A(\main.adder.s4_mant[35] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold370 (.A(\main.adder.out[23] ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0367_),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold372 (.A(\main.float_registers[0][29] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0159_),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold374 (.A(\main.adder.s4_exponent[0] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold375 (.A(\main.adder.s4_exponent[6] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0259_),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold377 (.A(\main.adder.s3_sum[31] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold378 (.A(\main.adder.s4_mant[44] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0448_),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold380 (.A(\main.adder.s2_larger[31] ),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold381 (.A(\main.float_registers[1][11] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold382 (.A(\main.adder.s3_exponent[5] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold383 (.A(\main.adder.s2_smaler[46] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0353_),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold385 (.A(\main.adder.s4_exponent[5] ),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold386 (.A(\main.adder.s1_exp_diff[6] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold387 (.A(\main.adder.s3_sum[25] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold388 (.A(\main.adder.s4_exponent_adjust[9] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold389 (.A(\main.adder.out[1] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0261_),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold391 (.A(\main.adder.s4_exponent[4] ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold392 (.A(\main.adder.out[30] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0374_),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold394 (.A(\main.float_registers[0][4] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold395 (.A(\main.float_registers[2][2] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold396 (.A(\main.float_registers[1][18] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold397 (.A(\main.float_registers[1][29] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold398 (.A(_0191_),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold399 (.A(\main.adder.s2_larger[43] ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold400 (.A(_0319_),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold401 (.A(\main.float_registers[2][3] ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold402 (.A(\main.float_registers[1][5] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold403 (.A(\main.float_registers[3][15] ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold404 (.A(\main.adder.s4_mant[47] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0451_),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold406 (.A(\main.adder.s2_smaler[18] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0477_),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold408 (.A(\main.float_registers[3][9] ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0238_),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold410 (.A(\main.float_registers[1][20] ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold411 (.A(\main.float_registers[3][17] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold412 (.A(\main.float_registers[3][0] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold413 (.A(\main.float_registers[3][11] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold414 (.A(\main.float_registers[2][5] ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold415 (.A(\main.float_registers[1][6] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold416 (.A(\main.float_registers[1][2] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold417 (.A(\main.float_registers[3][21] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold418 (.A(\main.adder.s4_exponent[1] ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0254_),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold420 (.A(\main.float_registers[0][1] ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold421 (.A(\main.adder.s1_exp_diff[7] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold422 (.A(\main.adder.out[3] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0263_),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold424 (.A(\main.float_registers[3][2] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold425 (.A(\main.adder.s2_smaler[45] ),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold426 (.A(\main.float_registers[2][25] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0218_),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold428 (.A(\main.adder.out[27] ),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold429 (.A(_0371_),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold430 (.A(\main.adder.s4_exponent[7] ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold431 (.A(_0260_),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold432 (.A(\main.float_registers[1][13] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold433 (.A(\main.float_registers[2][0] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold434 (.A(\main.float_registers[2][28] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold435 (.A(_0221_),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold436 (.A(\main.float_registers[1][7] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold437 (.A(\main.float_registers[1][31] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold438 (.A(_0193_),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold439 (.A(\main.float_registers[3][30] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold440 (.A(_0224_),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold441 (.A(\main.float_registers[2][27] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold442 (.A(\main.float_registers[1][8] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold443 (.A(\main.float_registers[1][30] ),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold444 (.A(\main.adder.s2_smaler[17] ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold445 (.A(_0476_),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold446 (.A(\main.adder.out[26] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold447 (.A(_0370_),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold448 (.A(\main.float_registers[2][7] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold449 (.A(\main.float_registers[2][26] ),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold450 (.A(\main.float_registers[3][8] ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold451 (.A(\main.float_registers[2][11] ),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold452 (.A(\main.adder.s2_smaler[21] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold453 (.A(\main.adder.s4_exponent[2] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold454 (.A(\main.float_registers[3][6] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold455 (.A(\main.adder.s5_mant[23] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold456 (.A(\main.float_registers[1][15] ),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold457 (.A(_0177_),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold458 (.A(\main.float_registers[3][26] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold459 (.A(\main.float_registers[1][22] ),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold460 (.A(\main.float_registers[1][28] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0190_),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold462 (.A(\main.adder.s1_larger[25] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold463 (.A(\main.float_registers[2][12] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold464 (.A(\main.float_registers[2][22] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold465 (.A(\main.adder.s2_smaler[35] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold466 (.A(\main.float_registers[2][23] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold467 (.A(\main.float_registers[2][21] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold468 (.A(\main.float_registers[2][16] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold469 (.A(\main.float_registers[3][12] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold470 (.A(\main.adder.s4_mant[37] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold471 (.A(\main.float_registers[3][23] ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold472 (.A(\main.adder.s1_rs.levels[0][23] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold473 (.A(\main.float_registers[2][6] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold474 (.A(\main.adder.s2_smaler[11] ),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0470_),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold476 (.A(\main.adder.out[29] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold477 (.A(_0373_),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold478 (.A(\main.float_registers[3][1] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold479 (.A(\main.adder.s5_exponent[8] ),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0398_),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold481 (.A(\main.adder.s4_mant[33] ),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold482 (.A(_0437_),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold483 (.A(\main.adder.s3_exponent[7] ),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold484 (.A(\main.float_registers[3][5] ),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold485 (.A(\main.adder.s4_mant[39] ),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold486 (.A(\main.float_registers[1][17] ),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold487 (.A(\main.adder.s1_exp_diff[2] ),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold488 (.A(\main.float_registers[3][22] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold489 (.A(\main.float_registers[3][16] ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold490 (.A(\main.float_registers[3][18] ),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold491 (.A(\main.float_registers[1][10] ),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold492 (.A(_0172_),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold493 (.A(\main.adder.s4_mant[46] ),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold494 (.A(_0450_),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold495 (.A(\main.float_registers[2][10] ),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold496 (.A(_0203_),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold497 (.A(\main.float_registers[3][29] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold498 (.A(_0239_),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold499 (.A(\main.float_registers[1][16] ),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold500 (.A(\main.adder.s2_larger[40] ),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold501 (.A(_0316_),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold502 (.A(\main.adder.s3_sum[30] ),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold503 (.A(\main.float_registers[3][27] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold504 (.A(\main.adder.s2_smaler[39] ),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold505 (.A(\main.float_registers[1][25] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold506 (.A(_0187_),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold507 (.A(\main.spi.out_bit_counter[2] ),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold508 (.A(_0603_),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold509 (.A(\main.float_registers[2][8] ),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold510 (.A(\main.float_registers[2][20] ),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold511 (.A(\main.float_registers[1][4] ),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold512 (.A(\main.float_registers[1][19] ),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold513 (.A(\main.adder.s5_S ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold514 (.A(\main.adder.s1_larger[28] ),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold515 (.A(\main.float_registers[2][17] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold516 (.A(\main.float_registers[2][18] ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold517 (.A(\main.float_registers[1][24] ),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold518 (.A(\main.float_registers[2][15] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold519 (.A(\main.adder.s1_exp_diff[1] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold520 (.A(\main.float_registers[3][31] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold521 (.A(_0223_),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold522 (.A(\main.adder.s4_mant[29] ),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold523 (.A(_0433_),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold524 (.A(\main.float_registers[1][27] ),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold525 (.A(\main.float_registers[1][12] ),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold526 (.A(\main.float_registers[1][23] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold527 (.A(\main.float_registers[2][24] ),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold528 (.A(\main.float_registers[3][25] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold529 (.A(_0662_),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold530 (.A(\main.float_registers[3][19] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold531 (.A(\main.float_registers[3][7] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold532 (.A(\main.float_registers[3][24] ),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold533 (.A(\main.adder.s1_exp_diff[3] ),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold534 (.A(\main.adder.s2_smaler[33] ),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold535 (.A(\main.float_registers[2][13] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold536 (.A(\main.float_registers[2][29] ),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0222_),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold538 (.A(\main.float_registers[3][20] ),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold539 (.A(\main.adder.s5_mant[22] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold540 (.A(\main.float_registers[1][26] ),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold541 (.A(\main.float_registers[1][0] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold542 (.A(\main.adder.s4_mant[31] ),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold543 (.A(_0435_),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold544 (.A(\main.float_registers[2][4] ),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold545 (.A(\main.adder.s4_mant[27] ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold546 (.A(_0431_),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold547 (.A(\main.float_registers[3][10] ),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0363_),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold549 (.A(\main.adder.s1_exp_diff[0] ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold550 (.A(\main.adder.s4_mant[45] ),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold551 (.A(_0449_),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold552 (.A(\main.adder.s5_mant[10] ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold553 (.A(\main.adder.s5_exponent[0] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold554 (.A(\main.adder.s3_sum[39] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold555 (.A(\main.spi.in_bit_counter[1] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold556 (.A(_1372_),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold557 (.A(_0241_),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold558 (.A(\main.float_registers[3][28] ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold559 (.A(\main.float_registers[3][14] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold560 (.A(_0651_),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold561 (.A(\main.adder.s5_mant[0] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold562 (.A(\main.adder.s2_smaler[36] ),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold563 (.A(\main.adder.s4_mant[41] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold564 (.A(\main.float_registers[2][30] ),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold565 (.A(_0128_),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold566 (.A(\main.spi.SPI_clock_sampled ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold567 (.A(\main.float_registers[3][3] ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold568 (.A(\main.adder.s3_sum[45] ),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold569 (.A(\main.float_registers[2][14] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold570 (.A(_0207_),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold571 (.A(\main.adder.s1_larger[23] ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold572 (.A(\main.float_registers[1][9] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold573 (.A(_0171_),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold574 (.A(\main.adder.s4_mant[40] ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold575 (.A(\main.adder.s3_sum[21] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold576 (.A(\main.spi.SPI_clock_sampler.sample_register[0] ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold577 (.A(\main.adder.s4_mant[23] ),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold578 (.A(_0427_),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold579 (.A(\main.float_registers[2][19] ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold580 (.A(\main.float_registers[3][13] ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold581 (.A(\main.adder.out[4] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold582 (.A(_0264_),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold583 (.A(\main.adder.s1_inf ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold584 (.A(\main.float_registers[2][31] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold585 (.A(_0661_),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold586 (.A(\main.adder.s5_mant[19] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold587 (.A(\main.adder.s4_mant[28] ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold588 (.A(_0432_),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold589 (.A(\main.float_registers[1][14] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold590 (.A(_0176_),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold591 (.A(\main.adder.s5_mant[16] ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold592 (.A(\main.float_registers[3][4] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold593 (.A(\main.float_registers[2][1] ),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold594 (.A(\main.adder.s2_smaler[34] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold595 (.A(\main.adder.s4_mant[26] ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold596 (.A(_0430_),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold597 (.A(\main.adder.s3_sum[38] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold598 (.A(\main.adder.s5_exponent[9] ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold599 (.A(\main.adder.s4_exponent_adjust[6] ),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold600 (.A(_0231_),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold601 (.A(\main.adder.s4_mant[43] ),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold602 (.A(\main.float_registers[2][9] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold603 (.A(_0202_),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold604 (.A(\main.adder.s2_smaler[32] ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold605 (.A(\main.read_command[1] ),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold606 (.A(_0634_),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold607 (.A(\main.adder.s1_larger[17] ),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold608 (.A(\main.adder.s3_sum[29] ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold609 (.A(\main.SPI_input_data[5] ),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold610 (.A(_0623_),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold611 (.A(\main.adder.s3_sum[28] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold612 (.A(\main.adder.s3_sum[46] ),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold613 (.A(_0505_),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold614 (.A(\main.adder.s5_mant[1] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold615 (.A(\main.SPI_input_data[3] ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold616 (.A(_0621_),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold617 (.A(\main.adder.s2_smaler[26] ),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold618 (.A(\main.adder.s4_mant[22] ),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold619 (.A(_0426_),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold620 (.A(\main.adder.s1_larger[20] ),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold621 (.A(\main.adder.s3_sum[34] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold622 (.A(\main.SPI_input_data[2] ),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold623 (.A(\main.adder.s5_mant[8] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold624 (.A(\main.register_id_result[0] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold625 (.A(\main.adder.s3_sum[27] ),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold626 (.A(\main.adder.s3_sum[36] ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold627 (.A(\main.adder.s3_sum[37] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold628 (.A(_0076_),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold629 (.A(_0225_),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold630 (.A(\main.adder.s2_smaler[24] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold631 (.A(\main.adder.s2_smaler[30] ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold632 (.A(\main.adder.s2_smaler[3] ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold633 (.A(\main.SPI_input_data[6] ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold634 (.A(_0624_),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold635 (.A(\main.adder.s2_smaler[37] ),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold636 (.A(\main.adder.s5_exponent[1] ),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold637 (.A(\main.adder.s2_smaler[23] ),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold638 (.A(\main.adder.s3_sum[43] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold639 (.A(\main.adder.s5_mant[17] ),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold640 (.A(\main.adder.s4_mant[24] ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold641 (.A(_0428_),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold642 (.A(\main.adder.s4_mant[25] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold643 (.A(_0429_),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold644 (.A(\main.adder.s2_smaler[20] ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold645 (.A(_0479_),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold646 (.A(\main.adder.s3_sum[42] ),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold647 (.A(\main.adder.s5_mant[21] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold648 (.A(\main.adder.s2_smaler[28] ),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold649 (.A(\main.adder.s3_sum[35] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold650 (.A(\main.adder.s5_mant[13] ),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold651 (.A(\main.SPI_input_data[4] ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold652 (.A(\main.adder.out[0] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold653 (.A(\main.adder.s4_exponent_adjust[8] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold654 (.A(\main.adder.s2_smaler[25] ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold655 (.A(\main.state[1] ),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold656 (.A(\main.adder.s3_sum[32] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold657 (.A(_0491_),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold658 (.A(\main.adder.s3_sum[33] ),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold659 (.A(\main.adder.s2_larger[46] ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold660 (.A(\main.adder.s3_sum[41] ),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold661 (.A(\main.adder.s5_mant[7] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold662 (.A(\main.adder.s4_exponent_adjust[7] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold663 (.A(\main.adder.s2_smaler[29] ),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold664 (.A(\main.adder.s2_smaler[27] ),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold665 (.A(\main.adder.s3_sum[26] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold666 (.A(\main.adder.s3_sum[44] ),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold667 (.A(_0503_),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold668 (.A(\main.read_command[0] ),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold669 (.A(_0633_),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold670 (.A(\main.spi.out_bit_counter[1] ),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold671 (.A(_0602_),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold672 (.A(\main.register_id_result[1] ),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold673 (.A(\main.adder.s4_exponent_adjust[4] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold674 (.A(\main.SPI_output_data_ready ),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold675 (.A(\main.adder.s5_exponent[5] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold676 (.A(\main.adder.s5_mant[12] ),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold677 (.A(\main.adder.s5_mant[15] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold678 (.A(\main.adder.s3_sum[40] ),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold679 (.A(\main.adder.s2_smaler[42] ),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold680 (.A(\main.adder.s5_mant[20] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold681 (.A(_0100_),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold682 (.A(_0506_),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold683 (.A(\main.adder.s5_exponent[3] ),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold684 (.A(_0064_),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold685 (.A(_0798_),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold686 (.A(\main.adder.s4_exponent_adjust[5] ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold687 (.A(\main.adder.s5_exponent[4] ),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold688 (.A(\main.adder.s4_exponent_adjust[3] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold689 (.A(\main.adder.s5_mant[6] ),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold690 (.A(\main.spi.in_bit_counter[0] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold691 (.A(\main.adder.s4_exponent_adjust[1] ),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold692 (.A(\main.adder.s5_mant[4] ),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold693 (.A(\main.adder.s5_mant[3] ),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold694 (.A(\main.adder.s5_mant[2] ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold695 (.A(\main.adder.s5_mant[5] ),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold696 (.A(\main.adder.s3_sum[48] ),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold697 (.A(\main.adder.s4_exponent_adjust[2] ),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold698 (.A(\main.adder.s5_mant[14] ),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold699 (.A(\main.adder.s5_mant[11] ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold700 (.A(\main.state[6] ),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold701 (.A(\main.SPI_input_data[3] ),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold702 (.A(\main.SPI_input_data[5] ),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold703 (.A(\main.SPI_input_data[4] ),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold704 (.A(\main.adder.s3_sum[34] ),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold705 (.A(\main.SPI_input_data[2] ),
    .X(net1627));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_4 FILLER_16_280 ();
 sg13g2_fill_1 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_295 ();
 sg13g2_fill_2 FILLER_16_305 ();
 sg13g2_fill_1 FILLER_16_307 ();
 sg13g2_decap_8 FILLER_16_312 ();
 sg13g2_fill_1 FILLER_16_319 ();
 sg13g2_decap_8 FILLER_16_344 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_decap_8 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_decap_8 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_16_414 ();
 sg13g2_decap_8 FILLER_16_421 ();
 sg13g2_decap_8 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_16_435 ();
 sg13g2_decap_8 FILLER_16_442 ();
 sg13g2_decap_8 FILLER_16_449 ();
 sg13g2_decap_8 FILLER_16_456 ();
 sg13g2_decap_8 FILLER_16_463 ();
 sg13g2_decap_8 FILLER_16_470 ();
 sg13g2_decap_8 FILLER_16_477 ();
 sg13g2_decap_8 FILLER_16_484 ();
 sg13g2_decap_8 FILLER_16_491 ();
 sg13g2_decap_8 FILLER_16_498 ();
 sg13g2_decap_8 FILLER_16_505 ();
 sg13g2_decap_8 FILLER_16_512 ();
 sg13g2_decap_8 FILLER_16_519 ();
 sg13g2_decap_8 FILLER_16_526 ();
 sg13g2_decap_8 FILLER_16_533 ();
 sg13g2_decap_8 FILLER_16_540 ();
 sg13g2_decap_8 FILLER_16_547 ();
 sg13g2_decap_8 FILLER_16_554 ();
 sg13g2_decap_8 FILLER_16_561 ();
 sg13g2_decap_8 FILLER_16_568 ();
 sg13g2_decap_8 FILLER_16_575 ();
 sg13g2_decap_8 FILLER_16_582 ();
 sg13g2_decap_8 FILLER_16_589 ();
 sg13g2_decap_8 FILLER_16_596 ();
 sg13g2_decap_8 FILLER_16_603 ();
 sg13g2_decap_8 FILLER_16_610 ();
 sg13g2_decap_8 FILLER_16_617 ();
 sg13g2_decap_8 FILLER_16_624 ();
 sg13g2_decap_8 FILLER_16_631 ();
 sg13g2_decap_8 FILLER_16_638 ();
 sg13g2_decap_8 FILLER_16_645 ();
 sg13g2_decap_8 FILLER_16_652 ();
 sg13g2_decap_8 FILLER_16_659 ();
 sg13g2_decap_8 FILLER_16_666 ();
 sg13g2_decap_8 FILLER_16_673 ();
 sg13g2_decap_8 FILLER_16_680 ();
 sg13g2_decap_8 FILLER_16_687 ();
 sg13g2_decap_8 FILLER_16_694 ();
 sg13g2_decap_8 FILLER_16_701 ();
 sg13g2_decap_8 FILLER_16_708 ();
 sg13g2_decap_8 FILLER_16_715 ();
 sg13g2_decap_8 FILLER_16_722 ();
 sg13g2_decap_8 FILLER_16_729 ();
 sg13g2_decap_8 FILLER_16_736 ();
 sg13g2_decap_8 FILLER_16_743 ();
 sg13g2_decap_8 FILLER_16_750 ();
 sg13g2_decap_8 FILLER_16_757 ();
 sg13g2_decap_8 FILLER_16_764 ();
 sg13g2_decap_8 FILLER_16_771 ();
 sg13g2_decap_8 FILLER_16_778 ();
 sg13g2_decap_8 FILLER_16_785 ();
 sg13g2_decap_8 FILLER_16_792 ();
 sg13g2_decap_8 FILLER_16_799 ();
 sg13g2_decap_8 FILLER_16_806 ();
 sg13g2_decap_8 FILLER_16_813 ();
 sg13g2_decap_8 FILLER_16_820 ();
 sg13g2_decap_8 FILLER_16_827 ();
 sg13g2_decap_8 FILLER_16_834 ();
 sg13g2_decap_8 FILLER_16_841 ();
 sg13g2_decap_8 FILLER_16_848 ();
 sg13g2_decap_8 FILLER_16_855 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_191 ();
 sg13g2_fill_1 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_221 ();
 sg13g2_decap_8 FILLER_17_228 ();
 sg13g2_decap_8 FILLER_17_244 ();
 sg13g2_decap_8 FILLER_17_251 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_265 ();
 sg13g2_decap_8 FILLER_17_272 ();
 sg13g2_fill_2 FILLER_17_279 ();
 sg13g2_fill_1 FILLER_17_281 ();
 sg13g2_decap_4 FILLER_17_292 ();
 sg13g2_fill_1 FILLER_17_296 ();
 sg13g2_fill_2 FILLER_17_332 ();
 sg13g2_fill_1 FILLER_17_334 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_4 FILLER_17_350 ();
 sg13g2_fill_1 FILLER_17_354 ();
 sg13g2_decap_4 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_8 FILLER_17_403 ();
 sg13g2_decap_8 FILLER_17_410 ();
 sg13g2_decap_8 FILLER_17_417 ();
 sg13g2_decap_8 FILLER_17_424 ();
 sg13g2_fill_1 FILLER_17_431 ();
 sg13g2_fill_1 FILLER_17_471 ();
 sg13g2_decap_8 FILLER_17_475 ();
 sg13g2_decap_8 FILLER_17_482 ();
 sg13g2_fill_1 FILLER_17_489 ();
 sg13g2_decap_8 FILLER_17_516 ();
 sg13g2_decap_8 FILLER_17_523 ();
 sg13g2_decap_8 FILLER_17_530 ();
 sg13g2_decap_8 FILLER_17_537 ();
 sg13g2_decap_8 FILLER_17_544 ();
 sg13g2_decap_8 FILLER_17_551 ();
 sg13g2_decap_8 FILLER_17_558 ();
 sg13g2_decap_8 FILLER_17_565 ();
 sg13g2_decap_8 FILLER_17_572 ();
 sg13g2_decap_8 FILLER_17_579 ();
 sg13g2_decap_8 FILLER_17_586 ();
 sg13g2_decap_8 FILLER_17_593 ();
 sg13g2_decap_8 FILLER_17_600 ();
 sg13g2_decap_8 FILLER_17_607 ();
 sg13g2_decap_8 FILLER_17_614 ();
 sg13g2_decap_8 FILLER_17_621 ();
 sg13g2_decap_8 FILLER_17_628 ();
 sg13g2_decap_8 FILLER_17_635 ();
 sg13g2_decap_8 FILLER_17_642 ();
 sg13g2_decap_8 FILLER_17_649 ();
 sg13g2_decap_8 FILLER_17_656 ();
 sg13g2_decap_8 FILLER_17_663 ();
 sg13g2_decap_8 FILLER_17_670 ();
 sg13g2_decap_8 FILLER_17_677 ();
 sg13g2_decap_8 FILLER_17_684 ();
 sg13g2_decap_8 FILLER_17_691 ();
 sg13g2_decap_8 FILLER_17_698 ();
 sg13g2_decap_8 FILLER_17_705 ();
 sg13g2_decap_8 FILLER_17_712 ();
 sg13g2_decap_8 FILLER_17_719 ();
 sg13g2_decap_8 FILLER_17_726 ();
 sg13g2_decap_8 FILLER_17_733 ();
 sg13g2_decap_8 FILLER_17_740 ();
 sg13g2_decap_8 FILLER_17_747 ();
 sg13g2_decap_8 FILLER_17_754 ();
 sg13g2_decap_8 FILLER_17_761 ();
 sg13g2_decap_8 FILLER_17_768 ();
 sg13g2_decap_8 FILLER_17_775 ();
 sg13g2_decap_8 FILLER_17_782 ();
 sg13g2_decap_8 FILLER_17_789 ();
 sg13g2_decap_8 FILLER_17_796 ();
 sg13g2_decap_8 FILLER_17_803 ();
 sg13g2_decap_8 FILLER_17_810 ();
 sg13g2_decap_8 FILLER_17_817 ();
 sg13g2_decap_8 FILLER_17_824 ();
 sg13g2_decap_8 FILLER_17_831 ();
 sg13g2_decap_8 FILLER_17_838 ();
 sg13g2_decap_8 FILLER_17_845 ();
 sg13g2_decap_8 FILLER_17_852 ();
 sg13g2_fill_2 FILLER_17_859 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_fill_1 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_165 ();
 sg13g2_decap_4 FILLER_18_170 ();
 sg13g2_fill_2 FILLER_18_174 ();
 sg13g2_fill_2 FILLER_18_186 ();
 sg13g2_fill_2 FILLER_18_214 ();
 sg13g2_fill_1 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_233 ();
 sg13g2_decap_4 FILLER_18_240 ();
 sg13g2_fill_2 FILLER_18_244 ();
 sg13g2_fill_2 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_265 ();
 sg13g2_fill_1 FILLER_18_318 ();
 sg13g2_fill_2 FILLER_18_342 ();
 sg13g2_decap_8 FILLER_18_383 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_2 FILLER_18_408 ();
 sg13g2_decap_4 FILLER_18_415 ();
 sg13g2_fill_1 FILLER_18_419 ();
 sg13g2_decap_8 FILLER_18_424 ();
 sg13g2_fill_2 FILLER_18_431 ();
 sg13g2_decap_4 FILLER_18_437 ();
 sg13g2_fill_1 FILLER_18_441 ();
 sg13g2_fill_1 FILLER_18_464 ();
 sg13g2_fill_1 FILLER_18_487 ();
 sg13g2_fill_2 FILLER_18_498 ();
 sg13g2_fill_1 FILLER_18_500 ();
 sg13g2_decap_4 FILLER_18_505 ();
 sg13g2_fill_1 FILLER_18_509 ();
 sg13g2_decap_8 FILLER_18_530 ();
 sg13g2_decap_8 FILLER_18_537 ();
 sg13g2_fill_1 FILLER_18_544 ();
 sg13g2_decap_8 FILLER_18_552 ();
 sg13g2_decap_8 FILLER_18_559 ();
 sg13g2_decap_8 FILLER_18_566 ();
 sg13g2_decap_4 FILLER_18_573 ();
 sg13g2_fill_1 FILLER_18_577 ();
 sg13g2_decap_8 FILLER_18_587 ();
 sg13g2_fill_2 FILLER_18_594 ();
 sg13g2_decap_8 FILLER_18_605 ();
 sg13g2_decap_8 FILLER_18_612 ();
 sg13g2_decap_8 FILLER_18_619 ();
 sg13g2_decap_8 FILLER_18_626 ();
 sg13g2_decap_8 FILLER_18_633 ();
 sg13g2_decap_8 FILLER_18_640 ();
 sg13g2_decap_8 FILLER_18_647 ();
 sg13g2_decap_8 FILLER_18_654 ();
 sg13g2_decap_8 FILLER_18_661 ();
 sg13g2_decap_8 FILLER_18_668 ();
 sg13g2_decap_8 FILLER_18_675 ();
 sg13g2_decap_8 FILLER_18_682 ();
 sg13g2_decap_8 FILLER_18_689 ();
 sg13g2_decap_8 FILLER_18_696 ();
 sg13g2_decap_8 FILLER_18_703 ();
 sg13g2_decap_8 FILLER_18_710 ();
 sg13g2_decap_8 FILLER_18_717 ();
 sg13g2_decap_8 FILLER_18_724 ();
 sg13g2_decap_8 FILLER_18_731 ();
 sg13g2_decap_8 FILLER_18_738 ();
 sg13g2_decap_8 FILLER_18_745 ();
 sg13g2_decap_8 FILLER_18_752 ();
 sg13g2_decap_8 FILLER_18_759 ();
 sg13g2_decap_8 FILLER_18_766 ();
 sg13g2_decap_8 FILLER_18_773 ();
 sg13g2_decap_8 FILLER_18_780 ();
 sg13g2_decap_8 FILLER_18_787 ();
 sg13g2_decap_8 FILLER_18_794 ();
 sg13g2_decap_8 FILLER_18_801 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_8 FILLER_18_815 ();
 sg13g2_decap_8 FILLER_18_822 ();
 sg13g2_decap_8 FILLER_18_829 ();
 sg13g2_decap_8 FILLER_18_836 ();
 sg13g2_decap_8 FILLER_18_843 ();
 sg13g2_decap_8 FILLER_18_850 ();
 sg13g2_decap_4 FILLER_18_857 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_fill_2 FILLER_19_140 ();
 sg13g2_decap_4 FILLER_19_152 ();
 sg13g2_fill_2 FILLER_19_182 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_235 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_fill_2 FILLER_19_310 ();
 sg13g2_fill_1 FILLER_19_312 ();
 sg13g2_fill_2 FILLER_19_354 ();
 sg13g2_fill_1 FILLER_19_356 ();
 sg13g2_fill_2 FILLER_19_361 ();
 sg13g2_fill_1 FILLER_19_363 ();
 sg13g2_decap_4 FILLER_19_379 ();
 sg13g2_fill_1 FILLER_19_383 ();
 sg13g2_fill_2 FILLER_19_449 ();
 sg13g2_decap_8 FILLER_19_475 ();
 sg13g2_decap_4 FILLER_19_569 ();
 sg13g2_fill_1 FILLER_19_582 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_fill_1 FILLER_19_630 ();
 sg13g2_decap_4 FILLER_19_641 ();
 sg13g2_fill_1 FILLER_19_645 ();
 sg13g2_decap_8 FILLER_19_659 ();
 sg13g2_decap_8 FILLER_19_666 ();
 sg13g2_decap_8 FILLER_19_673 ();
 sg13g2_decap_8 FILLER_19_680 ();
 sg13g2_decap_8 FILLER_19_687 ();
 sg13g2_decap_8 FILLER_19_694 ();
 sg13g2_decap_8 FILLER_19_701 ();
 sg13g2_decap_8 FILLER_19_708 ();
 sg13g2_decap_8 FILLER_19_715 ();
 sg13g2_decap_8 FILLER_19_722 ();
 sg13g2_decap_8 FILLER_19_729 ();
 sg13g2_decap_8 FILLER_19_736 ();
 sg13g2_decap_8 FILLER_19_743 ();
 sg13g2_decap_8 FILLER_19_750 ();
 sg13g2_decap_8 FILLER_19_757 ();
 sg13g2_decap_8 FILLER_19_764 ();
 sg13g2_decap_8 FILLER_19_771 ();
 sg13g2_decap_8 FILLER_19_778 ();
 sg13g2_decap_8 FILLER_19_785 ();
 sg13g2_decap_8 FILLER_19_792 ();
 sg13g2_decap_8 FILLER_19_799 ();
 sg13g2_decap_8 FILLER_19_806 ();
 sg13g2_decap_8 FILLER_19_813 ();
 sg13g2_decap_8 FILLER_19_820 ();
 sg13g2_decap_8 FILLER_19_827 ();
 sg13g2_decap_8 FILLER_19_834 ();
 sg13g2_decap_8 FILLER_19_841 ();
 sg13g2_decap_8 FILLER_19_848 ();
 sg13g2_decap_8 FILLER_19_855 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_4 FILLER_20_126 ();
 sg13g2_fill_1 FILLER_20_130 ();
 sg13g2_fill_1 FILLER_20_206 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_fill_1 FILLER_20_268 ();
 sg13g2_fill_2 FILLER_20_278 ();
 sg13g2_fill_1 FILLER_20_280 ();
 sg13g2_decap_4 FILLER_20_327 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_fill_1 FILLER_20_390 ();
 sg13g2_fill_1 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_419 ();
 sg13g2_fill_1 FILLER_20_432 ();
 sg13g2_fill_2 FILLER_20_474 ();
 sg13g2_fill_1 FILLER_20_476 ();
 sg13g2_fill_2 FILLER_20_483 ();
 sg13g2_fill_1 FILLER_20_490 ();
 sg13g2_decap_4 FILLER_20_502 ();
 sg13g2_fill_2 FILLER_20_506 ();
 sg13g2_fill_2 FILLER_20_528 ();
 sg13g2_fill_1 FILLER_20_555 ();
 sg13g2_decap_4 FILLER_20_589 ();
 sg13g2_decap_8 FILLER_20_597 ();
 sg13g2_decap_8 FILLER_20_604 ();
 sg13g2_fill_2 FILLER_20_611 ();
 sg13g2_fill_1 FILLER_20_613 ();
 sg13g2_decap_4 FILLER_20_670 ();
 sg13g2_fill_1 FILLER_20_674 ();
 sg13g2_decap_8 FILLER_20_688 ();
 sg13g2_decap_8 FILLER_20_695 ();
 sg13g2_decap_8 FILLER_20_702 ();
 sg13g2_decap_8 FILLER_20_709 ();
 sg13g2_decap_8 FILLER_20_716 ();
 sg13g2_decap_8 FILLER_20_723 ();
 sg13g2_decap_8 FILLER_20_730 ();
 sg13g2_decap_8 FILLER_20_737 ();
 sg13g2_decap_8 FILLER_20_744 ();
 sg13g2_decap_8 FILLER_20_751 ();
 sg13g2_decap_8 FILLER_20_758 ();
 sg13g2_decap_8 FILLER_20_765 ();
 sg13g2_decap_8 FILLER_20_772 ();
 sg13g2_decap_8 FILLER_20_779 ();
 sg13g2_decap_8 FILLER_20_786 ();
 sg13g2_decap_8 FILLER_20_793 ();
 sg13g2_decap_8 FILLER_20_800 ();
 sg13g2_decap_8 FILLER_20_807 ();
 sg13g2_decap_8 FILLER_20_814 ();
 sg13g2_decap_8 FILLER_20_821 ();
 sg13g2_decap_8 FILLER_20_828 ();
 sg13g2_decap_8 FILLER_20_835 ();
 sg13g2_decap_8 FILLER_20_842 ();
 sg13g2_decap_8 FILLER_20_849 ();
 sg13g2_decap_4 FILLER_20_856 ();
 sg13g2_fill_2 FILLER_20_860 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_4 FILLER_21_133 ();
 sg13g2_fill_2 FILLER_21_137 ();
 sg13g2_decap_8 FILLER_21_153 ();
 sg13g2_decap_8 FILLER_21_160 ();
 sg13g2_fill_1 FILLER_21_167 ();
 sg13g2_fill_1 FILLER_21_173 ();
 sg13g2_fill_2 FILLER_21_184 ();
 sg13g2_fill_1 FILLER_21_186 ();
 sg13g2_fill_2 FILLER_21_213 ();
 sg13g2_fill_1 FILLER_21_215 ();
 sg13g2_fill_2 FILLER_21_236 ();
 sg13g2_fill_1 FILLER_21_264 ();
 sg13g2_fill_2 FILLER_21_296 ();
 sg13g2_fill_1 FILLER_21_298 ();
 sg13g2_fill_2 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_318 ();
 sg13g2_fill_2 FILLER_21_325 ();
 sg13g2_fill_1 FILLER_21_327 ();
 sg13g2_fill_1 FILLER_21_354 ();
 sg13g2_fill_2 FILLER_21_417 ();
 sg13g2_fill_1 FILLER_21_419 ();
 sg13g2_fill_2 FILLER_21_423 ();
 sg13g2_fill_1 FILLER_21_425 ();
 sg13g2_fill_1 FILLER_21_439 ();
 sg13g2_decap_8 FILLER_21_445 ();
 sg13g2_decap_4 FILLER_21_452 ();
 sg13g2_fill_1 FILLER_21_460 ();
 sg13g2_fill_1 FILLER_21_527 ();
 sg13g2_fill_2 FILLER_21_564 ();
 sg13g2_fill_2 FILLER_21_571 ();
 sg13g2_decap_8 FILLER_21_577 ();
 sg13g2_fill_1 FILLER_21_584 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_fill_1 FILLER_21_623 ();
 sg13g2_decap_4 FILLER_21_632 ();
 sg13g2_fill_2 FILLER_21_653 ();
 sg13g2_decap_8 FILLER_21_710 ();
 sg13g2_decap_8 FILLER_21_717 ();
 sg13g2_decap_8 FILLER_21_724 ();
 sg13g2_decap_8 FILLER_21_731 ();
 sg13g2_decap_8 FILLER_21_738 ();
 sg13g2_decap_8 FILLER_21_745 ();
 sg13g2_decap_8 FILLER_21_752 ();
 sg13g2_decap_8 FILLER_21_759 ();
 sg13g2_decap_8 FILLER_21_766 ();
 sg13g2_decap_8 FILLER_21_773 ();
 sg13g2_decap_8 FILLER_21_780 ();
 sg13g2_decap_8 FILLER_21_787 ();
 sg13g2_decap_8 FILLER_21_794 ();
 sg13g2_decap_8 FILLER_21_801 ();
 sg13g2_decap_8 FILLER_21_808 ();
 sg13g2_decap_8 FILLER_21_815 ();
 sg13g2_decap_8 FILLER_21_822 ();
 sg13g2_decap_8 FILLER_21_829 ();
 sg13g2_decap_8 FILLER_21_836 ();
 sg13g2_decap_8 FILLER_21_843 ();
 sg13g2_decap_8 FILLER_21_850 ();
 sg13g2_decap_4 FILLER_21_857 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_decap_4 FILLER_22_155 ();
 sg13g2_fill_1 FILLER_22_159 ();
 sg13g2_fill_2 FILLER_22_178 ();
 sg13g2_fill_2 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_208 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_4 FILLER_22_245 ();
 sg13g2_fill_2 FILLER_22_262 ();
 sg13g2_fill_2 FILLER_22_285 ();
 sg13g2_decap_8 FILLER_22_300 ();
 sg13g2_decap_4 FILLER_22_307 ();
 sg13g2_fill_2 FILLER_22_311 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_4 FILLER_22_329 ();
 sg13g2_fill_2 FILLER_22_333 ();
 sg13g2_fill_2 FILLER_22_371 ();
 sg13g2_fill_2 FILLER_22_385 ();
 sg13g2_fill_1 FILLER_22_387 ();
 sg13g2_fill_2 FILLER_22_416 ();
 sg13g2_fill_1 FILLER_22_418 ();
 sg13g2_decap_8 FILLER_22_457 ();
 sg13g2_fill_2 FILLER_22_491 ();
 sg13g2_fill_1 FILLER_22_493 ();
 sg13g2_decap_8 FILLER_22_502 ();
 sg13g2_fill_2 FILLER_22_509 ();
 sg13g2_fill_1 FILLER_22_511 ();
 sg13g2_fill_2 FILLER_22_538 ();
 sg13g2_fill_2 FILLER_22_548 ();
 sg13g2_fill_1 FILLER_22_550 ();
 sg13g2_decap_4 FILLER_22_568 ();
 sg13g2_fill_2 FILLER_22_572 ();
 sg13g2_fill_2 FILLER_22_597 ();
 sg13g2_fill_1 FILLER_22_599 ();
 sg13g2_fill_2 FILLER_22_639 ();
 sg13g2_fill_2 FILLER_22_653 ();
 sg13g2_fill_2 FILLER_22_672 ();
 sg13g2_decap_4 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_718 ();
 sg13g2_decap_8 FILLER_22_725 ();
 sg13g2_decap_8 FILLER_22_732 ();
 sg13g2_decap_8 FILLER_22_739 ();
 sg13g2_decap_8 FILLER_22_746 ();
 sg13g2_decap_8 FILLER_22_753 ();
 sg13g2_decap_8 FILLER_22_760 ();
 sg13g2_decap_8 FILLER_22_767 ();
 sg13g2_decap_8 FILLER_22_774 ();
 sg13g2_decap_8 FILLER_22_781 ();
 sg13g2_decap_8 FILLER_22_788 ();
 sg13g2_decap_8 FILLER_22_795 ();
 sg13g2_decap_8 FILLER_22_802 ();
 sg13g2_decap_8 FILLER_22_809 ();
 sg13g2_decap_8 FILLER_22_816 ();
 sg13g2_decap_8 FILLER_22_823 ();
 sg13g2_decap_8 FILLER_22_830 ();
 sg13g2_decap_8 FILLER_22_837 ();
 sg13g2_decap_8 FILLER_22_844 ();
 sg13g2_decap_8 FILLER_22_851 ();
 sg13g2_decap_4 FILLER_22_858 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_4 FILLER_23_105 ();
 sg13g2_fill_2 FILLER_23_132 ();
 sg13g2_fill_1 FILLER_23_160 ();
 sg13g2_fill_1 FILLER_23_210 ();
 sg13g2_fill_2 FILLER_23_227 ();
 sg13g2_decap_4 FILLER_23_297 ();
 sg13g2_fill_2 FILLER_23_301 ();
 sg13g2_fill_1 FILLER_23_337 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_fill_2 FILLER_23_366 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_450 ();
 sg13g2_decap_8 FILLER_23_463 ();
 sg13g2_fill_2 FILLER_23_470 ();
 sg13g2_fill_1 FILLER_23_482 ();
 sg13g2_fill_2 FILLER_23_571 ();
 sg13g2_decap_4 FILLER_23_604 ();
 sg13g2_decap_4 FILLER_23_617 ();
 sg13g2_fill_1 FILLER_23_621 ();
 sg13g2_fill_1 FILLER_23_635 ();
 sg13g2_fill_1 FILLER_23_653 ();
 sg13g2_decap_4 FILLER_23_670 ();
 sg13g2_fill_2 FILLER_23_674 ();
 sg13g2_decap_4 FILLER_23_729 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_4 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_88 ();
 sg13g2_fill_2 FILLER_24_187 ();
 sg13g2_fill_1 FILLER_24_189 ();
 sg13g2_decap_4 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_decap_4 FILLER_24_232 ();
 sg13g2_fill_2 FILLER_24_236 ();
 sg13g2_fill_2 FILLER_24_261 ();
 sg13g2_fill_1 FILLER_24_263 ();
 sg13g2_fill_1 FILLER_24_300 ();
 sg13g2_fill_2 FILLER_24_306 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_fill_1 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_388 ();
 sg13g2_fill_2 FILLER_24_415 ();
 sg13g2_fill_2 FILLER_24_434 ();
 sg13g2_fill_1 FILLER_24_436 ();
 sg13g2_fill_2 FILLER_24_470 ();
 sg13g2_fill_1 FILLER_24_472 ();
 sg13g2_decap_4 FILLER_24_493 ();
 sg13g2_fill_2 FILLER_24_523 ();
 sg13g2_decap_8 FILLER_24_566 ();
 sg13g2_decap_8 FILLER_24_573 ();
 sg13g2_fill_1 FILLER_24_580 ();
 sg13g2_fill_1 FILLER_24_624 ();
 sg13g2_fill_1 FILLER_24_634 ();
 sg13g2_fill_1 FILLER_24_672 ();
 sg13g2_fill_2 FILLER_24_697 ();
 sg13g2_fill_1 FILLER_24_711 ();
 sg13g2_fill_2 FILLER_24_773 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_8 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_847 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_4 FILLER_25_98 ();
 sg13g2_fill_1 FILLER_25_102 ();
 sg13g2_decap_8 FILLER_25_113 ();
 sg13g2_fill_2 FILLER_25_120 ();
 sg13g2_decap_8 FILLER_25_132 ();
 sg13g2_fill_1 FILLER_25_139 ();
 sg13g2_fill_2 FILLER_25_153 ();
 sg13g2_fill_2 FILLER_25_159 ();
 sg13g2_fill_1 FILLER_25_161 ();
 sg13g2_fill_2 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_207 ();
 sg13g2_fill_2 FILLER_25_222 ();
 sg13g2_fill_2 FILLER_25_236 ();
 sg13g2_fill_1 FILLER_25_238 ();
 sg13g2_fill_2 FILLER_25_275 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_fill_2 FILLER_25_300 ();
 sg13g2_fill_1 FILLER_25_302 ();
 sg13g2_fill_2 FILLER_25_307 ();
 sg13g2_fill_1 FILLER_25_309 ();
 sg13g2_fill_2 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_353 ();
 sg13g2_decap_4 FILLER_25_360 ();
 sg13g2_fill_2 FILLER_25_396 ();
 sg13g2_fill_2 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_415 ();
 sg13g2_decap_4 FILLER_25_422 ();
 sg13g2_fill_1 FILLER_25_426 ();
 sg13g2_decap_8 FILLER_25_432 ();
 sg13g2_fill_2 FILLER_25_444 ();
 sg13g2_fill_2 FILLER_25_449 ();
 sg13g2_fill_2 FILLER_25_468 ();
 sg13g2_fill_1 FILLER_25_470 ();
 sg13g2_decap_4 FILLER_25_475 ();
 sg13g2_fill_2 FILLER_25_483 ();
 sg13g2_fill_1 FILLER_25_485 ();
 sg13g2_decap_8 FILLER_25_491 ();
 sg13g2_fill_2 FILLER_25_498 ();
 sg13g2_fill_1 FILLER_25_500 ();
 sg13g2_fill_2 FILLER_25_512 ();
 sg13g2_fill_1 FILLER_25_514 ();
 sg13g2_decap_4 FILLER_25_533 ();
 sg13g2_fill_1 FILLER_25_537 ();
 sg13g2_decap_8 FILLER_25_543 ();
 sg13g2_decap_8 FILLER_25_550 ();
 sg13g2_decap_8 FILLER_25_557 ();
 sg13g2_fill_2 FILLER_25_564 ();
 sg13g2_fill_1 FILLER_25_566 ();
 sg13g2_fill_1 FILLER_25_599 ();
 sg13g2_fill_2 FILLER_25_631 ();
 sg13g2_decap_4 FILLER_25_636 ();
 sg13g2_fill_2 FILLER_25_640 ();
 sg13g2_fill_2 FILLER_25_647 ();
 sg13g2_fill_1 FILLER_25_649 ();
 sg13g2_decap_8 FILLER_25_666 ();
 sg13g2_decap_8 FILLER_25_673 ();
 sg13g2_fill_2 FILLER_25_680 ();
 sg13g2_fill_1 FILLER_25_696 ();
 sg13g2_fill_2 FILLER_25_710 ();
 sg13g2_fill_1 FILLER_25_730 ();
 sg13g2_decap_4 FILLER_25_738 ();
 sg13g2_fill_2 FILLER_25_742 ();
 sg13g2_fill_1 FILLER_25_754 ();
 sg13g2_decap_8 FILLER_25_786 ();
 sg13g2_decap_8 FILLER_25_793 ();
 sg13g2_decap_8 FILLER_25_800 ();
 sg13g2_decap_8 FILLER_25_807 ();
 sg13g2_decap_8 FILLER_25_814 ();
 sg13g2_decap_8 FILLER_25_821 ();
 sg13g2_decap_8 FILLER_25_828 ();
 sg13g2_decap_8 FILLER_25_835 ();
 sg13g2_decap_8 FILLER_25_842 ();
 sg13g2_decap_8 FILLER_25_849 ();
 sg13g2_decap_4 FILLER_25_856 ();
 sg13g2_fill_2 FILLER_25_860 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_4 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_102 ();
 sg13g2_fill_2 FILLER_26_155 ();
 sg13g2_fill_1 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_188 ();
 sg13g2_decap_4 FILLER_26_215 ();
 sg13g2_decap_8 FILLER_26_232 ();
 sg13g2_fill_1 FILLER_26_248 ();
 sg13g2_decap_8 FILLER_26_253 ();
 sg13g2_fill_1 FILLER_26_260 ();
 sg13g2_fill_2 FILLER_26_345 ();
 sg13g2_fill_1 FILLER_26_347 ();
 sg13g2_decap_4 FILLER_26_360 ();
 sg13g2_fill_2 FILLER_26_364 ();
 sg13g2_fill_1 FILLER_26_389 ();
 sg13g2_decap_4 FILLER_26_399 ();
 sg13g2_fill_1 FILLER_26_411 ();
 sg13g2_fill_1 FILLER_26_486 ();
 sg13g2_decap_4 FILLER_26_491 ();
 sg13g2_decap_4 FILLER_26_500 ();
 sg13g2_fill_1 FILLER_26_504 ();
 sg13g2_fill_2 FILLER_26_538 ();
 sg13g2_decap_4 FILLER_26_545 ();
 sg13g2_decap_8 FILLER_26_607 ();
 sg13g2_fill_1 FILLER_26_614 ();
 sg13g2_fill_2 FILLER_26_627 ();
 sg13g2_fill_1 FILLER_26_650 ();
 sg13g2_decap_8 FILLER_26_727 ();
 sg13g2_fill_1 FILLER_26_734 ();
 sg13g2_decap_8 FILLER_26_788 ();
 sg13g2_decap_8 FILLER_26_795 ();
 sg13g2_decap_8 FILLER_26_802 ();
 sg13g2_decap_8 FILLER_26_809 ();
 sg13g2_decap_8 FILLER_26_816 ();
 sg13g2_decap_8 FILLER_26_823 ();
 sg13g2_decap_8 FILLER_26_830 ();
 sg13g2_decap_8 FILLER_26_837 ();
 sg13g2_decap_8 FILLER_26_844 ();
 sg13g2_decap_8 FILLER_26_851 ();
 sg13g2_decap_4 FILLER_26_858 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_fill_1 FILLER_27_105 ();
 sg13g2_decap_4 FILLER_27_127 ();
 sg13g2_fill_1 FILLER_27_175 ();
 sg13g2_fill_1 FILLER_27_194 ();
 sg13g2_fill_2 FILLER_27_221 ();
 sg13g2_fill_1 FILLER_27_223 ();
 sg13g2_fill_1 FILLER_27_234 ();
 sg13g2_fill_1 FILLER_27_261 ();
 sg13g2_fill_1 FILLER_27_317 ();
 sg13g2_fill_2 FILLER_27_336 ();
 sg13g2_fill_1 FILLER_27_338 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_fill_2 FILLER_27_403 ();
 sg13g2_fill_1 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_27_414 ();
 sg13g2_decap_8 FILLER_27_421 ();
 sg13g2_decap_8 FILLER_27_436 ();
 sg13g2_fill_1 FILLER_27_443 ();
 sg13g2_decap_8 FILLER_27_449 ();
 sg13g2_decap_4 FILLER_27_473 ();
 sg13g2_decap_8 FILLER_27_515 ();
 sg13g2_fill_1 FILLER_27_522 ();
 sg13g2_fill_1 FILLER_27_527 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_fill_2 FILLER_27_539 ();
 sg13g2_decap_4 FILLER_27_663 ();
 sg13g2_fill_2 FILLER_27_667 ();
 sg13g2_decap_8 FILLER_27_674 ();
 sg13g2_decap_4 FILLER_27_681 ();
 sg13g2_fill_2 FILLER_27_705 ();
 sg13g2_decap_8 FILLER_27_725 ();
 sg13g2_fill_2 FILLER_27_732 ();
 sg13g2_decap_4 FILLER_27_759 ();
 sg13g2_fill_1 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_786 ();
 sg13g2_decap_8 FILLER_27_793 ();
 sg13g2_decap_8 FILLER_27_800 ();
 sg13g2_decap_8 FILLER_27_807 ();
 sg13g2_decap_8 FILLER_27_814 ();
 sg13g2_decap_8 FILLER_27_821 ();
 sg13g2_decap_8 FILLER_27_828 ();
 sg13g2_decap_8 FILLER_27_835 ();
 sg13g2_decap_8 FILLER_27_842 ();
 sg13g2_decap_8 FILLER_27_849 ();
 sg13g2_decap_4 FILLER_27_856 ();
 sg13g2_fill_2 FILLER_27_860 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_fill_2 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_164 ();
 sg13g2_fill_1 FILLER_28_201 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_decap_4 FILLER_28_261 ();
 sg13g2_fill_1 FILLER_28_265 ();
 sg13g2_decap_4 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_306 ();
 sg13g2_fill_1 FILLER_28_317 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_349 ();
 sg13g2_decap_4 FILLER_28_356 ();
 sg13g2_fill_2 FILLER_28_386 ();
 sg13g2_fill_1 FILLER_28_402 ();
 sg13g2_fill_2 FILLER_28_429 ();
 sg13g2_decap_4 FILLER_28_457 ();
 sg13g2_fill_2 FILLER_28_485 ();
 sg13g2_fill_2 FILLER_28_496 ();
 sg13g2_fill_1 FILLER_28_498 ();
 sg13g2_decap_4 FILLER_28_514 ();
 sg13g2_fill_1 FILLER_28_544 ();
 sg13g2_decap_4 FILLER_28_589 ();
 sg13g2_fill_2 FILLER_28_593 ();
 sg13g2_fill_1 FILLER_28_611 ();
 sg13g2_decap_4 FILLER_28_617 ();
 sg13g2_fill_1 FILLER_28_621 ();
 sg13g2_decap_8 FILLER_28_630 ();
 sg13g2_decap_4 FILLER_28_641 ();
 sg13g2_fill_1 FILLER_28_645 ();
 sg13g2_decap_8 FILLER_28_680 ();
 sg13g2_decap_4 FILLER_28_687 ();
 sg13g2_fill_2 FILLER_28_691 ();
 sg13g2_fill_1 FILLER_28_707 ();
 sg13g2_decap_4 FILLER_28_712 ();
 sg13g2_fill_2 FILLER_28_761 ();
 sg13g2_fill_2 FILLER_28_776 ();
 sg13g2_fill_1 FILLER_28_778 ();
 sg13g2_fill_2 FILLER_28_787 ();
 sg13g2_fill_2 FILLER_28_793 ();
 sg13g2_fill_1 FILLER_28_795 ();
 sg13g2_decap_8 FILLER_28_804 ();
 sg13g2_decap_8 FILLER_28_811 ();
 sg13g2_decap_8 FILLER_28_818 ();
 sg13g2_decap_8 FILLER_28_825 ();
 sg13g2_decap_8 FILLER_28_832 ();
 sg13g2_decap_8 FILLER_28_839 ();
 sg13g2_decap_8 FILLER_28_846 ();
 sg13g2_decap_8 FILLER_28_853 ();
 sg13g2_fill_2 FILLER_28_860 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_4 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_95 ();
 sg13g2_fill_2 FILLER_29_123 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_fill_2 FILLER_29_135 ();
 sg13g2_fill_1 FILLER_29_146 ();
 sg13g2_fill_2 FILLER_29_193 ();
 sg13g2_decap_8 FILLER_29_204 ();
 sg13g2_decap_4 FILLER_29_221 ();
 sg13g2_fill_1 FILLER_29_225 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_2 FILLER_29_273 ();
 sg13g2_fill_2 FILLER_29_280 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_decap_4 FILLER_29_307 ();
 sg13g2_fill_2 FILLER_29_311 ();
 sg13g2_decap_8 FILLER_29_340 ();
 sg13g2_decap_4 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_375 ();
 sg13g2_fill_1 FILLER_29_416 ();
 sg13g2_fill_2 FILLER_29_442 ();
 sg13g2_fill_1 FILLER_29_457 ();
 sg13g2_fill_1 FILLER_29_517 ();
 sg13g2_decap_4 FILLER_29_544 ();
 sg13g2_fill_2 FILLER_29_548 ();
 sg13g2_fill_1 FILLER_29_646 ();
 sg13g2_fill_2 FILLER_29_668 ();
 sg13g2_fill_1 FILLER_29_670 ();
 sg13g2_fill_2 FILLER_29_712 ();
 sg13g2_fill_1 FILLER_29_714 ();
 sg13g2_fill_2 FILLER_29_725 ();
 sg13g2_fill_1 FILLER_29_727 ();
 sg13g2_fill_2 FILLER_29_741 ();
 sg13g2_fill_1 FILLER_29_743 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_4 FILLER_29_756 ();
 sg13g2_fill_2 FILLER_29_760 ();
 sg13g2_fill_1 FILLER_29_783 ();
 sg13g2_decap_8 FILLER_29_822 ();
 sg13g2_decap_8 FILLER_29_829 ();
 sg13g2_decap_8 FILLER_29_836 ();
 sg13g2_decap_8 FILLER_29_843 ();
 sg13g2_decap_8 FILLER_29_850 ();
 sg13g2_decap_4 FILLER_29_857 ();
 sg13g2_fill_1 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_4 FILLER_30_77 ();
 sg13g2_fill_2 FILLER_30_81 ();
 sg13g2_fill_1 FILLER_30_116 ();
 sg13g2_fill_2 FILLER_30_153 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_fill_2 FILLER_30_208 ();
 sg13g2_fill_2 FILLER_30_225 ();
 sg13g2_fill_1 FILLER_30_252 ();
 sg13g2_fill_2 FILLER_30_257 ();
 sg13g2_fill_2 FILLER_30_283 ();
 sg13g2_fill_1 FILLER_30_285 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_decap_4 FILLER_30_307 ();
 sg13g2_fill_2 FILLER_30_311 ();
 sg13g2_fill_2 FILLER_30_323 ();
 sg13g2_decap_4 FILLER_30_351 ();
 sg13g2_fill_2 FILLER_30_375 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_fill_1 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_30_429 ();
 sg13g2_fill_2 FILLER_30_436 ();
 sg13g2_fill_1 FILLER_30_442 ();
 sg13g2_fill_2 FILLER_30_452 ();
 sg13g2_fill_2 FILLER_30_481 ();
 sg13g2_fill_2 FILLER_30_489 ();
 sg13g2_fill_2 FILLER_30_500 ();
 sg13g2_fill_1 FILLER_30_502 ();
 sg13g2_decap_8 FILLER_30_519 ();
 sg13g2_decap_4 FILLER_30_526 ();
 sg13g2_fill_2 FILLER_30_538 ();
 sg13g2_fill_1 FILLER_30_623 ();
 sg13g2_fill_2 FILLER_30_643 ();
 sg13g2_fill_2 FILLER_30_658 ();
 sg13g2_fill_1 FILLER_30_660 ();
 sg13g2_fill_2 FILLER_30_684 ();
 sg13g2_fill_1 FILLER_30_695 ();
 sg13g2_fill_2 FILLER_30_718 ();
 sg13g2_fill_1 FILLER_30_720 ();
 sg13g2_fill_2 FILLER_30_798 ();
 sg13g2_fill_2 FILLER_30_837 ();
 sg13g2_fill_1 FILLER_30_839 ();
 sg13g2_decap_8 FILLER_30_844 ();
 sg13g2_decap_8 FILLER_30_851 ();
 sg13g2_decap_4 FILLER_30_858 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_103 ();
 sg13g2_fill_1 FILLER_31_105 ();
 sg13g2_fill_2 FILLER_31_134 ();
 sg13g2_fill_1 FILLER_31_136 ();
 sg13g2_decap_4 FILLER_31_163 ();
 sg13g2_fill_1 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_191 ();
 sg13g2_decap_4 FILLER_31_228 ();
 sg13g2_decap_4 FILLER_31_253 ();
 sg13g2_fill_2 FILLER_31_257 ();
 sg13g2_fill_2 FILLER_31_285 ();
 sg13g2_fill_2 FILLER_31_295 ();
 sg13g2_decap_4 FILLER_31_307 ();
 sg13g2_decap_8 FILLER_31_326 ();
 sg13g2_decap_4 FILLER_31_333 ();
 sg13g2_fill_2 FILLER_31_363 ();
 sg13g2_fill_2 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_31_377 ();
 sg13g2_fill_1 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_2 FILLER_31_450 ();
 sg13g2_fill_1 FILLER_31_452 ();
 sg13g2_fill_2 FILLER_31_464 ();
 sg13g2_fill_2 FILLER_31_478 ();
 sg13g2_fill_1 FILLER_31_480 ();
 sg13g2_fill_2 FILLER_31_496 ();
 sg13g2_fill_2 FILLER_31_503 ();
 sg13g2_fill_1 FILLER_31_505 ();
 sg13g2_fill_1 FILLER_31_518 ();
 sg13g2_fill_2 FILLER_31_545 ();
 sg13g2_fill_1 FILLER_31_566 ();
 sg13g2_fill_2 FILLER_31_590 ();
 sg13g2_fill_1 FILLER_31_592 ();
 sg13g2_fill_1 FILLER_31_601 ();
 sg13g2_fill_2 FILLER_31_626 ();
 sg13g2_fill_1 FILLER_31_628 ();
 sg13g2_fill_2 FILLER_31_638 ();
 sg13g2_fill_1 FILLER_31_640 ();
 sg13g2_fill_1 FILLER_31_663 ();
 sg13g2_fill_1 FILLER_31_682 ();
 sg13g2_fill_2 FILLER_31_711 ();
 sg13g2_decap_4 FILLER_31_727 ();
 sg13g2_fill_1 FILLER_31_731 ();
 sg13g2_fill_1 FILLER_31_754 ();
 sg13g2_fill_2 FILLER_31_842 ();
 sg13g2_fill_1 FILLER_31_844 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_4 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_128 ();
 sg13g2_fill_1 FILLER_32_130 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_fill_1 FILLER_32_297 ();
 sg13g2_fill_2 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_315 ();
 sg13g2_fill_2 FILLER_32_326 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_fill_2 FILLER_32_344 ();
 sg13g2_decap_4 FILLER_32_350 ();
 sg13g2_fill_1 FILLER_32_354 ();
 sg13g2_decap_8 FILLER_32_359 ();
 sg13g2_decap_8 FILLER_32_366 ();
 sg13g2_fill_1 FILLER_32_382 ();
 sg13g2_fill_2 FILLER_32_396 ();
 sg13g2_fill_2 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_415 ();
 sg13g2_fill_1 FILLER_32_417 ();
 sg13g2_fill_2 FILLER_32_433 ();
 sg13g2_decap_8 FILLER_32_440 ();
 sg13g2_fill_1 FILLER_32_447 ();
 sg13g2_decap_4 FILLER_32_459 ();
 sg13g2_fill_1 FILLER_32_463 ();
 sg13g2_fill_1 FILLER_32_470 ();
 sg13g2_fill_2 FILLER_32_492 ();
 sg13g2_fill_1 FILLER_32_494 ();
 sg13g2_fill_2 FILLER_32_505 ();
 sg13g2_fill_2 FILLER_32_518 ();
 sg13g2_fill_1 FILLER_32_551 ();
 sg13g2_fill_2 FILLER_32_566 ();
 sg13g2_fill_2 FILLER_32_594 ();
 sg13g2_fill_1 FILLER_32_607 ();
 sg13g2_decap_8 FILLER_32_665 ();
 sg13g2_fill_2 FILLER_32_690 ();
 sg13g2_decap_8 FILLER_32_698 ();
 sg13g2_fill_2 FILLER_32_705 ();
 sg13g2_fill_1 FILLER_32_707 ();
 sg13g2_fill_2 FILLER_32_744 ();
 sg13g2_fill_2 FILLER_32_754 ();
 sg13g2_fill_1 FILLER_32_756 ();
 sg13g2_fill_1 FILLER_32_762 ();
 sg13g2_fill_2 FILLER_32_829 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_fill_2 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_44 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_71 ();
 sg13g2_decap_8 FILLER_33_78 ();
 sg13g2_decap_4 FILLER_33_85 ();
 sg13g2_fill_1 FILLER_33_99 ();
 sg13g2_fill_2 FILLER_33_110 ();
 sg13g2_fill_2 FILLER_33_132 ();
 sg13g2_fill_1 FILLER_33_134 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_fill_2 FILLER_33_165 ();
 sg13g2_fill_1 FILLER_33_167 ();
 sg13g2_fill_2 FILLER_33_200 ();
 sg13g2_decap_4 FILLER_33_215 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_257 ();
 sg13g2_decap_4 FILLER_33_280 ();
 sg13g2_decap_4 FILLER_33_294 ();
 sg13g2_fill_2 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_318 ();
 sg13g2_fill_1 FILLER_33_324 ();
 sg13g2_fill_2 FILLER_33_329 ();
 sg13g2_fill_1 FILLER_33_331 ();
 sg13g2_decap_4 FILLER_33_337 ();
 sg13g2_decap_4 FILLER_33_368 ();
 sg13g2_fill_1 FILLER_33_372 ();
 sg13g2_fill_2 FILLER_33_383 ();
 sg13g2_decap_8 FILLER_33_390 ();
 sg13g2_fill_1 FILLER_33_397 ();
 sg13g2_decap_4 FILLER_33_416 ();
 sg13g2_decap_4 FILLER_33_436 ();
 sg13g2_fill_1 FILLER_33_440 ();
 sg13g2_decap_8 FILLER_33_451 ();
 sg13g2_fill_1 FILLER_33_458 ();
 sg13g2_fill_2 FILLER_33_467 ();
 sg13g2_fill_1 FILLER_33_469 ();
 sg13g2_fill_2 FILLER_33_476 ();
 sg13g2_fill_1 FILLER_33_478 ();
 sg13g2_fill_2 FILLER_33_504 ();
 sg13g2_fill_2 FILLER_33_520 ();
 sg13g2_fill_1 FILLER_33_522 ();
 sg13g2_fill_2 FILLER_33_528 ();
 sg13g2_fill_1 FILLER_33_530 ();
 sg13g2_decap_4 FILLER_33_535 ();
 sg13g2_fill_2 FILLER_33_539 ();
 sg13g2_decap_8 FILLER_33_593 ();
 sg13g2_decap_8 FILLER_33_600 ();
 sg13g2_decap_8 FILLER_33_628 ();
 sg13g2_fill_2 FILLER_33_635 ();
 sg13g2_fill_1 FILLER_33_637 ();
 sg13g2_decap_4 FILLER_33_643 ();
 sg13g2_fill_1 FILLER_33_647 ();
 sg13g2_decap_4 FILLER_33_653 ();
 sg13g2_decap_4 FILLER_33_662 ();
 sg13g2_fill_1 FILLER_33_666 ();
 sg13g2_decap_8 FILLER_33_675 ();
 sg13g2_fill_2 FILLER_33_682 ();
 sg13g2_fill_2 FILLER_33_741 ();
 sg13g2_fill_1 FILLER_33_743 ();
 sg13g2_fill_2 FILLER_33_757 ();
 sg13g2_fill_1 FILLER_33_799 ();
 sg13g2_fill_2 FILLER_33_826 ();
 sg13g2_fill_1 FILLER_33_828 ();
 sg13g2_fill_2 FILLER_33_859 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_21 ();
 sg13g2_fill_1 FILLER_34_25 ();
 sg13g2_decap_4 FILLER_34_78 ();
 sg13g2_decap_8 FILLER_34_97 ();
 sg13g2_decap_4 FILLER_34_104 ();
 sg13g2_fill_2 FILLER_34_108 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_fill_1 FILLER_34_137 ();
 sg13g2_decap_4 FILLER_34_148 ();
 sg13g2_fill_1 FILLER_34_152 ();
 sg13g2_fill_2 FILLER_34_193 ();
 sg13g2_fill_1 FILLER_34_195 ();
 sg13g2_decap_8 FILLER_34_222 ();
 sg13g2_fill_2 FILLER_34_250 ();
 sg13g2_fill_2 FILLER_34_257 ();
 sg13g2_fill_2 FILLER_34_271 ();
 sg13g2_fill_1 FILLER_34_273 ();
 sg13g2_fill_2 FILLER_34_301 ();
 sg13g2_decap_4 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_337 ();
 sg13g2_decap_4 FILLER_34_348 ();
 sg13g2_fill_2 FILLER_34_366 ();
 sg13g2_fill_2 FILLER_34_380 ();
 sg13g2_fill_2 FILLER_34_411 ();
 sg13g2_fill_1 FILLER_34_413 ();
 sg13g2_fill_2 FILLER_34_424 ();
 sg13g2_fill_1 FILLER_34_430 ();
 sg13g2_decap_4 FILLER_34_451 ();
 sg13g2_fill_1 FILLER_34_455 ();
 sg13g2_fill_1 FILLER_34_464 ();
 sg13g2_decap_4 FILLER_34_471 ();
 sg13g2_decap_4 FILLER_34_492 ();
 sg13g2_fill_1 FILLER_34_496 ();
 sg13g2_fill_1 FILLER_34_523 ();
 sg13g2_decap_4 FILLER_34_628 ();
 sg13g2_fill_1 FILLER_34_645 ();
 sg13g2_fill_1 FILLER_34_661 ();
 sg13g2_decap_4 FILLER_34_677 ();
 sg13g2_fill_2 FILLER_34_684 ();
 sg13g2_decap_8 FILLER_34_692 ();
 sg13g2_decap_4 FILLER_34_699 ();
 sg13g2_decap_8 FILLER_34_714 ();
 sg13g2_fill_2 FILLER_34_774 ();
 sg13g2_fill_1 FILLER_34_776 ();
 sg13g2_fill_2 FILLER_34_834 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_4 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_25 ();
 sg13g2_fill_2 FILLER_35_45 ();
 sg13g2_fill_2 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_65 ();
 sg13g2_fill_2 FILLER_35_101 ();
 sg13g2_fill_1 FILLER_35_103 ();
 sg13g2_decap_8 FILLER_35_163 ();
 sg13g2_fill_2 FILLER_35_200 ();
 sg13g2_fill_1 FILLER_35_202 ();
 sg13g2_decap_8 FILLER_35_211 ();
 sg13g2_decap_8 FILLER_35_218 ();
 sg13g2_decap_8 FILLER_35_225 ();
 sg13g2_decap_8 FILLER_35_232 ();
 sg13g2_decap_8 FILLER_35_239 ();
 sg13g2_decap_8 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_253 ();
 sg13g2_decap_8 FILLER_35_265 ();
 sg13g2_decap_8 FILLER_35_296 ();
 sg13g2_fill_2 FILLER_35_303 ();
 sg13g2_fill_1 FILLER_35_329 ();
 sg13g2_fill_2 FILLER_35_349 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_fill_2 FILLER_35_371 ();
 sg13g2_fill_1 FILLER_35_373 ();
 sg13g2_fill_2 FILLER_35_379 ();
 sg13g2_fill_1 FILLER_35_381 ();
 sg13g2_decap_4 FILLER_35_395 ();
 sg13g2_fill_1 FILLER_35_410 ();
 sg13g2_decap_8 FILLER_35_421 ();
 sg13g2_fill_1 FILLER_35_432 ();
 sg13g2_decap_4 FILLER_35_442 ();
 sg13g2_fill_1 FILLER_35_446 ();
 sg13g2_fill_1 FILLER_35_456 ();
 sg13g2_fill_2 FILLER_35_466 ();
 sg13g2_fill_1 FILLER_35_468 ();
 sg13g2_decap_8 FILLER_35_495 ();
 sg13g2_fill_2 FILLER_35_502 ();
 sg13g2_fill_1 FILLER_35_504 ();
 sg13g2_decap_4 FILLER_35_519 ();
 sg13g2_fill_2 FILLER_35_535 ();
 sg13g2_fill_2 FILLER_35_546 ();
 sg13g2_fill_1 FILLER_35_548 ();
 sg13g2_fill_1 FILLER_35_553 ();
 sg13g2_fill_2 FILLER_35_559 ();
 sg13g2_fill_2 FILLER_35_571 ();
 sg13g2_fill_1 FILLER_35_608 ();
 sg13g2_decap_8 FILLER_35_628 ();
 sg13g2_decap_8 FILLER_35_635 ();
 sg13g2_decap_8 FILLER_35_642 ();
 sg13g2_decap_4 FILLER_35_661 ();
 sg13g2_fill_1 FILLER_35_665 ();
 sg13g2_fill_1 FILLER_35_674 ();
 sg13g2_fill_2 FILLER_35_679 ();
 sg13g2_fill_2 FILLER_35_685 ();
 sg13g2_decap_8 FILLER_35_697 ();
 sg13g2_fill_1 FILLER_35_704 ();
 sg13g2_decap_4 FILLER_35_721 ();
 sg13g2_fill_1 FILLER_35_798 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_11 ();
 sg13g2_decap_8 FILLER_36_16 ();
 sg13g2_fill_1 FILLER_36_23 ();
 sg13g2_fill_2 FILLER_36_54 ();
 sg13g2_fill_2 FILLER_36_77 ();
 sg13g2_fill_1 FILLER_36_79 ();
 sg13g2_decap_8 FILLER_36_123 ();
 sg13g2_fill_1 FILLER_36_130 ();
 sg13g2_fill_1 FILLER_36_141 ();
 sg13g2_fill_2 FILLER_36_152 ();
 sg13g2_fill_2 FILLER_36_264 ();
 sg13g2_fill_2 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_273 ();
 sg13g2_fill_2 FILLER_36_288 ();
 sg13g2_fill_1 FILLER_36_290 ();
 sg13g2_decap_4 FILLER_36_296 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_fill_1 FILLER_36_336 ();
 sg13g2_fill_2 FILLER_36_342 ();
 sg13g2_fill_1 FILLER_36_344 ();
 sg13g2_fill_1 FILLER_36_355 ();
 sg13g2_decap_4 FILLER_36_372 ();
 sg13g2_fill_2 FILLER_36_410 ();
 sg13g2_fill_1 FILLER_36_412 ();
 sg13g2_fill_1 FILLER_36_418 ();
 sg13g2_fill_2 FILLER_36_424 ();
 sg13g2_fill_1 FILLER_36_431 ();
 sg13g2_fill_2 FILLER_36_483 ();
 sg13g2_fill_1 FILLER_36_511 ();
 sg13g2_fill_2 FILLER_36_538 ();
 sg13g2_fill_2 FILLER_36_566 ();
 sg13g2_fill_1 FILLER_36_599 ();
 sg13g2_fill_1 FILLER_36_608 ();
 sg13g2_decap_4 FILLER_36_652 ();
 sg13g2_fill_2 FILLER_36_695 ();
 sg13g2_fill_1 FILLER_36_697 ();
 sg13g2_fill_2 FILLER_36_719 ();
 sg13g2_fill_1 FILLER_36_721 ();
 sg13g2_fill_1 FILLER_36_793 ();
 sg13g2_fill_2 FILLER_36_803 ();
 sg13g2_fill_1 FILLER_36_805 ();
 sg13g2_fill_1 FILLER_36_811 ();
 sg13g2_fill_1 FILLER_36_852 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_54 ();
 sg13g2_fill_1 FILLER_37_56 ();
 sg13g2_decap_4 FILLER_37_78 ();
 sg13g2_fill_2 FILLER_37_82 ();
 sg13g2_fill_2 FILLER_37_89 ();
 sg13g2_fill_1 FILLER_37_91 ();
 sg13g2_fill_2 FILLER_37_101 ();
 sg13g2_fill_1 FILLER_37_103 ();
 sg13g2_decap_4 FILLER_37_129 ();
 sg13g2_fill_2 FILLER_37_153 ();
 sg13g2_fill_1 FILLER_37_155 ();
 sg13g2_fill_1 FILLER_37_171 ();
 sg13g2_decap_4 FILLER_37_204 ();
 sg13g2_fill_2 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_220 ();
 sg13g2_fill_2 FILLER_37_244 ();
 sg13g2_fill_1 FILLER_37_246 ();
 sg13g2_fill_2 FILLER_37_265 ();
 sg13g2_fill_2 FILLER_37_322 ();
 sg13g2_fill_1 FILLER_37_352 ();
 sg13g2_fill_2 FILLER_37_363 ();
 sg13g2_fill_1 FILLER_37_369 ();
 sg13g2_fill_2 FILLER_37_375 ();
 sg13g2_fill_1 FILLER_37_377 ();
 sg13g2_fill_2 FILLER_37_382 ();
 sg13g2_decap_4 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_2 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_37_433 ();
 sg13g2_fill_2 FILLER_37_440 ();
 sg13g2_fill_1 FILLER_37_442 ();
 sg13g2_decap_8 FILLER_37_456 ();
 sg13g2_decap_8 FILLER_37_467 ();
 sg13g2_decap_8 FILLER_37_474 ();
 sg13g2_fill_1 FILLER_37_481 ();
 sg13g2_decap_4 FILLER_37_491 ();
 sg13g2_fill_1 FILLER_37_495 ();
 sg13g2_fill_1 FILLER_37_500 ();
 sg13g2_fill_2 FILLER_37_563 ();
 sg13g2_decap_4 FILLER_37_620 ();
 sg13g2_decap_8 FILLER_37_628 ();
 sg13g2_decap_4 FILLER_37_635 ();
 sg13g2_fill_2 FILLER_37_669 ();
 sg13g2_fill_1 FILLER_37_692 ();
 sg13g2_fill_1 FILLER_37_717 ();
 sg13g2_fill_2 FILLER_37_777 ();
 sg13g2_fill_1 FILLER_37_788 ();
 sg13g2_fill_2 FILLER_37_842 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_31 ();
 sg13g2_fill_2 FILLER_38_46 ();
 sg13g2_fill_2 FILLER_38_78 ();
 sg13g2_fill_1 FILLER_38_80 ();
 sg13g2_fill_2 FILLER_38_107 ();
 sg13g2_fill_1 FILLER_38_109 ();
 sg13g2_decap_8 FILLER_38_131 ();
 sg13g2_decap_4 FILLER_38_138 ();
 sg13g2_fill_2 FILLER_38_152 ();
 sg13g2_fill_1 FILLER_38_154 ();
 sg13g2_fill_2 FILLER_38_160 ();
 sg13g2_fill_1 FILLER_38_172 ();
 sg13g2_fill_2 FILLER_38_183 ();
 sg13g2_decap_4 FILLER_38_195 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_decap_4 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_328 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_4 FILLER_38_361 ();
 sg13g2_fill_2 FILLER_38_365 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_decap_8 FILLER_38_407 ();
 sg13g2_decap_4 FILLER_38_466 ();
 sg13g2_fill_1 FILLER_38_470 ();
 sg13g2_fill_1 FILLER_38_475 ();
 sg13g2_fill_2 FILLER_38_517 ();
 sg13g2_fill_2 FILLER_38_612 ();
 sg13g2_fill_2 FILLER_38_631 ();
 sg13g2_decap_4 FILLER_38_636 ();
 sg13g2_fill_2 FILLER_38_640 ();
 sg13g2_fill_1 FILLER_38_667 ();
 sg13g2_decap_4 FILLER_38_684 ();
 sg13g2_fill_2 FILLER_38_688 ();
 sg13g2_fill_1 FILLER_38_722 ();
 sg13g2_fill_2 FILLER_38_732 ();
 sg13g2_fill_1 FILLER_38_800 ();
 sg13g2_fill_1 FILLER_38_814 ();
 sg13g2_fill_2 FILLER_38_829 ();
 sg13g2_fill_1 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_78 ();
 sg13g2_fill_1 FILLER_39_96 ();
 sg13g2_fill_2 FILLER_39_106 ();
 sg13g2_decap_8 FILLER_39_129 ();
 sg13g2_decap_8 FILLER_39_136 ();
 sg13g2_fill_1 FILLER_39_147 ();
 sg13g2_fill_1 FILLER_39_174 ();
 sg13g2_decap_8 FILLER_39_193 ();
 sg13g2_decap_4 FILLER_39_200 ();
 sg13g2_fill_1 FILLER_39_218 ();
 sg13g2_fill_1 FILLER_39_236 ();
 sg13g2_decap_8 FILLER_39_330 ();
 sg13g2_fill_1 FILLER_39_337 ();
 sg13g2_fill_1 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_374 ();
 sg13g2_fill_1 FILLER_39_386 ();
 sg13g2_decap_4 FILLER_39_391 ();
 sg13g2_fill_2 FILLER_39_395 ();
 sg13g2_fill_2 FILLER_39_507 ();
 sg13g2_decap_8 FILLER_39_512 ();
 sg13g2_fill_1 FILLER_39_557 ();
 sg13g2_decap_8 FILLER_39_620 ();
 sg13g2_decap_4 FILLER_39_627 ();
 sg13g2_fill_2 FILLER_39_631 ();
 sg13g2_fill_1 FILLER_39_644 ();
 sg13g2_fill_2 FILLER_39_649 ();
 sg13g2_fill_2 FILLER_39_666 ();
 sg13g2_fill_1 FILLER_39_668 ();
 sg13g2_fill_1 FILLER_39_687 ();
 sg13g2_fill_2 FILLER_39_708 ();
 sg13g2_fill_1 FILLER_39_758 ();
 sg13g2_fill_2 FILLER_39_768 ();
 sg13g2_fill_1 FILLER_39_770 ();
 sg13g2_fill_2 FILLER_39_811 ();
 sg13g2_fill_1 FILLER_39_813 ();
 sg13g2_fill_1 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_36 ();
 sg13g2_fill_1 FILLER_40_47 ();
 sg13g2_decap_8 FILLER_40_78 ();
 sg13g2_fill_2 FILLER_40_85 ();
 sg13g2_decap_4 FILLER_40_122 ();
 sg13g2_fill_2 FILLER_40_126 ();
 sg13g2_fill_2 FILLER_40_146 ();
 sg13g2_fill_1 FILLER_40_148 ();
 sg13g2_decap_8 FILLER_40_155 ();
 sg13g2_decap_8 FILLER_40_162 ();
 sg13g2_decap_4 FILLER_40_169 ();
 sg13g2_decap_8 FILLER_40_194 ();
 sg13g2_fill_1 FILLER_40_201 ();
 sg13g2_fill_1 FILLER_40_212 ();
 sg13g2_fill_1 FILLER_40_221 ();
 sg13g2_fill_2 FILLER_40_246 ();
 sg13g2_fill_1 FILLER_40_248 ();
 sg13g2_decap_4 FILLER_40_260 ();
 sg13g2_fill_2 FILLER_40_264 ();
 sg13g2_decap_4 FILLER_40_276 ();
 sg13g2_fill_2 FILLER_40_309 ();
 sg13g2_fill_1 FILLER_40_311 ();
 sg13g2_decap_8 FILLER_40_325 ();
 sg13g2_fill_1 FILLER_40_332 ();
 sg13g2_fill_2 FILLER_40_402 ();
 sg13g2_fill_1 FILLER_40_422 ();
 sg13g2_fill_1 FILLER_40_428 ();
 sg13g2_fill_2 FILLER_40_450 ();
 sg13g2_fill_1 FILLER_40_452 ();
 sg13g2_fill_1 FILLER_40_467 ();
 sg13g2_fill_1 FILLER_40_478 ();
 sg13g2_fill_2 FILLER_40_484 ();
 sg13g2_fill_1 FILLER_40_486 ();
 sg13g2_fill_2 FILLER_40_517 ();
 sg13g2_decap_4 FILLER_40_549 ();
 sg13g2_fill_2 FILLER_40_594 ();
 sg13g2_fill_1 FILLER_40_614 ();
 sg13g2_decap_8 FILLER_40_619 ();
 sg13g2_decap_4 FILLER_40_626 ();
 sg13g2_decap_4 FILLER_40_633 ();
 sg13g2_fill_1 FILLER_40_637 ();
 sg13g2_fill_2 FILLER_40_661 ();
 sg13g2_fill_1 FILLER_40_663 ();
 sg13g2_fill_2 FILLER_40_668 ();
 sg13g2_fill_1 FILLER_40_670 ();
 sg13g2_fill_1 FILLER_40_737 ();
 sg13g2_fill_2 FILLER_40_765 ();
 sg13g2_fill_2 FILLER_40_798 ();
 sg13g2_fill_1 FILLER_40_800 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_4 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_11 ();
 sg13g2_fill_2 FILLER_41_25 ();
 sg13g2_decap_4 FILLER_41_53 ();
 sg13g2_decap_8 FILLER_41_78 ();
 sg13g2_fill_1 FILLER_41_85 ();
 sg13g2_decap_8 FILLER_41_138 ();
 sg13g2_decap_4 FILLER_41_145 ();
 sg13g2_decap_4 FILLER_41_170 ();
 sg13g2_fill_1 FILLER_41_174 ();
 sg13g2_fill_2 FILLER_41_181 ();
 sg13g2_fill_1 FILLER_41_183 ();
 sg13g2_decap_4 FILLER_41_194 ();
 sg13g2_decap_4 FILLER_41_214 ();
 sg13g2_fill_2 FILLER_41_218 ();
 sg13g2_fill_1 FILLER_41_230 ();
 sg13g2_decap_8 FILLER_41_242 ();
 sg13g2_decap_4 FILLER_41_249 ();
 sg13g2_fill_2 FILLER_41_253 ();
 sg13g2_fill_1 FILLER_41_277 ();
 sg13g2_decap_8 FILLER_41_288 ();
 sg13g2_decap_8 FILLER_41_331 ();
 sg13g2_fill_1 FILLER_41_338 ();
 sg13g2_fill_1 FILLER_41_366 ();
 sg13g2_fill_2 FILLER_41_397 ();
 sg13g2_fill_1 FILLER_41_404 ();
 sg13g2_fill_2 FILLER_41_413 ();
 sg13g2_fill_2 FILLER_41_440 ();
 sg13g2_fill_1 FILLER_41_442 ();
 sg13g2_fill_1 FILLER_41_461 ();
 sg13g2_fill_2 FILLER_41_479 ();
 sg13g2_fill_1 FILLER_41_481 ();
 sg13g2_fill_1 FILLER_41_580 ();
 sg13g2_fill_2 FILLER_41_597 ();
 sg13g2_fill_2 FILLER_41_631 ();
 sg13g2_fill_1 FILLER_41_633 ();
 sg13g2_fill_1 FILLER_41_835 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_28 ();
 sg13g2_fill_1 FILLER_42_30 ();
 sg13g2_fill_2 FILLER_42_40 ();
 sg13g2_decap_4 FILLER_42_51 ();
 sg13g2_fill_2 FILLER_42_55 ();
 sg13g2_decap_8 FILLER_42_78 ();
 sg13g2_fill_1 FILLER_42_85 ();
 sg13g2_fill_2 FILLER_42_95 ();
 sg13g2_fill_1 FILLER_42_101 ();
 sg13g2_fill_1 FILLER_42_111 ();
 sg13g2_fill_2 FILLER_42_121 ();
 sg13g2_fill_1 FILLER_42_127 ();
 sg13g2_fill_1 FILLER_42_137 ();
 sg13g2_decap_8 FILLER_42_159 ();
 sg13g2_decap_8 FILLER_42_166 ();
 sg13g2_fill_2 FILLER_42_173 ();
 sg13g2_fill_1 FILLER_42_175 ();
 sg13g2_fill_2 FILLER_42_181 ();
 sg13g2_decap_8 FILLER_42_187 ();
 sg13g2_decap_8 FILLER_42_194 ();
 sg13g2_fill_2 FILLER_42_201 ();
 sg13g2_fill_1 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_213 ();
 sg13g2_fill_2 FILLER_42_220 ();
 sg13g2_decap_4 FILLER_42_227 ();
 sg13g2_fill_1 FILLER_42_231 ();
 sg13g2_decap_4 FILLER_42_242 ();
 sg13g2_decap_4 FILLER_42_274 ();
 sg13g2_fill_1 FILLER_42_278 ();
 sg13g2_decap_8 FILLER_42_289 ();
 sg13g2_decap_4 FILLER_42_296 ();
 sg13g2_decap_8 FILLER_42_304 ();
 sg13g2_decap_8 FILLER_42_328 ();
 sg13g2_decap_4 FILLER_42_357 ();
 sg13g2_fill_1 FILLER_42_410 ();
 sg13g2_fill_2 FILLER_42_441 ();
 sg13g2_decap_4 FILLER_42_489 ();
 sg13g2_fill_1 FILLER_42_493 ();
 sg13g2_fill_2 FILLER_42_498 ();
 sg13g2_decap_8 FILLER_42_540 ();
 sg13g2_fill_2 FILLER_42_547 ();
 sg13g2_fill_1 FILLER_42_549 ();
 sg13g2_decap_4 FILLER_42_564 ();
 sg13g2_decap_8 FILLER_42_621 ();
 sg13g2_decap_8 FILLER_42_628 ();
 sg13g2_fill_2 FILLER_42_635 ();
 sg13g2_fill_1 FILLER_42_637 ();
 sg13g2_fill_1 FILLER_42_659 ();
 sg13g2_fill_1 FILLER_42_700 ();
 sg13g2_fill_2 FILLER_42_763 ();
 sg13g2_fill_2 FILLER_42_801 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_7 ();
 sg13g2_fill_2 FILLER_43_27 ();
 sg13g2_fill_2 FILLER_43_56 ();
 sg13g2_decap_4 FILLER_43_79 ();
 sg13g2_fill_2 FILLER_43_83 ();
 sg13g2_fill_1 FILLER_43_90 ();
 sg13g2_decap_4 FILLER_43_95 ();
 sg13g2_fill_2 FILLER_43_134 ();
 sg13g2_decap_4 FILLER_43_166 ();
 sg13g2_fill_1 FILLER_43_222 ();
 sg13g2_decap_4 FILLER_43_227 ();
 sg13g2_decap_8 FILLER_43_261 ();
 sg13g2_decap_8 FILLER_43_268 ();
 sg13g2_fill_2 FILLER_43_275 ();
 sg13g2_fill_1 FILLER_43_277 ();
 sg13g2_fill_1 FILLER_43_298 ();
 sg13g2_fill_2 FILLER_43_335 ();
 sg13g2_fill_1 FILLER_43_337 ();
 sg13g2_fill_2 FILLER_43_373 ();
 sg13g2_fill_1 FILLER_43_385 ();
 sg13g2_fill_2 FILLER_43_395 ();
 sg13g2_fill_1 FILLER_43_397 ();
 sg13g2_fill_1 FILLER_43_407 ();
 sg13g2_decap_4 FILLER_43_418 ();
 sg13g2_fill_2 FILLER_43_426 ();
 sg13g2_fill_1 FILLER_43_428 ();
 sg13g2_decap_8 FILLER_43_437 ();
 sg13g2_decap_4 FILLER_43_444 ();
 sg13g2_fill_1 FILLER_43_448 ();
 sg13g2_fill_1 FILLER_43_462 ();
 sg13g2_fill_1 FILLER_43_475 ();
 sg13g2_decap_4 FILLER_43_516 ();
 sg13g2_decap_4 FILLER_43_546 ();
 sg13g2_fill_2 FILLER_43_558 ();
 sg13g2_fill_1 FILLER_43_560 ();
 sg13g2_fill_2 FILLER_43_587 ();
 sg13g2_fill_1 FILLER_43_593 ();
 sg13g2_decap_4 FILLER_43_624 ();
 sg13g2_fill_2 FILLER_43_628 ();
 sg13g2_fill_1 FILLER_43_634 ();
 sg13g2_decap_8 FILLER_43_645 ();
 sg13g2_fill_2 FILLER_43_652 ();
 sg13g2_fill_1 FILLER_43_654 ();
 sg13g2_fill_1 FILLER_43_659 ();
 sg13g2_fill_2 FILLER_43_680 ();
 sg13g2_fill_1 FILLER_43_682 ();
 sg13g2_fill_2 FILLER_43_718 ();
 sg13g2_fill_2 FILLER_43_788 ();
 sg13g2_fill_2 FILLER_43_816 ();
 sg13g2_fill_1 FILLER_43_818 ();
 sg13g2_decap_4 FILLER_43_858 ();
 sg13g2_fill_1 FILLER_44_31 ();
 sg13g2_decap_4 FILLER_44_79 ();
 sg13g2_fill_1 FILLER_44_118 ();
 sg13g2_decap_8 FILLER_44_123 ();
 sg13g2_decap_8 FILLER_44_130 ();
 sg13g2_fill_2 FILLER_44_137 ();
 sg13g2_decap_8 FILLER_44_160 ();
 sg13g2_fill_2 FILLER_44_167 ();
 sg13g2_fill_1 FILLER_44_169 ();
 sg13g2_decap_4 FILLER_44_188 ();
 sg13g2_fill_2 FILLER_44_210 ();
 sg13g2_fill_1 FILLER_44_261 ();
 sg13g2_fill_1 FILLER_44_295 ();
 sg13g2_fill_2 FILLER_44_341 ();
 sg13g2_decap_4 FILLER_44_408 ();
 sg13g2_fill_2 FILLER_44_412 ();
 sg13g2_fill_2 FILLER_44_440 ();
 sg13g2_fill_2 FILLER_44_480 ();
 sg13g2_fill_2 FILLER_44_527 ();
 sg13g2_fill_1 FILLER_44_529 ();
 sg13g2_fill_2 FILLER_44_534 ();
 sg13g2_decap_8 FILLER_44_572 ();
 sg13g2_fill_2 FILLER_44_579 ();
 sg13g2_fill_1 FILLER_44_581 ();
 sg13g2_fill_2 FILLER_44_594 ();
 sg13g2_decap_4 FILLER_44_614 ();
 sg13g2_fill_1 FILLER_44_618 ();
 sg13g2_decap_8 FILLER_44_678 ();
 sg13g2_decap_8 FILLER_44_685 ();
 sg13g2_fill_1 FILLER_44_692 ();
 sg13g2_decap_8 FILLER_44_760 ();
 sg13g2_fill_2 FILLER_44_767 ();
 sg13g2_fill_2 FILLER_44_818 ();
 sg13g2_decap_4 FILLER_44_842 ();
 sg13g2_fill_1 FILLER_44_846 ();
 sg13g2_decap_8 FILLER_44_851 ();
 sg13g2_decap_4 FILLER_44_858 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_15 ();
 sg13g2_fill_2 FILLER_45_34 ();
 sg13g2_fill_1 FILLER_45_36 ();
 sg13g2_decap_8 FILLER_45_46 ();
 sg13g2_decap_4 FILLER_45_62 ();
 sg13g2_fill_1 FILLER_45_66 ();
 sg13g2_fill_2 FILLER_45_76 ();
 sg13g2_fill_2 FILLER_45_95 ();
 sg13g2_fill_1 FILLER_45_97 ();
 sg13g2_fill_2 FILLER_45_116 ();
 sg13g2_fill_1 FILLER_45_118 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_fill_1 FILLER_45_147 ();
 sg13g2_decap_4 FILLER_45_169 ();
 sg13g2_fill_2 FILLER_45_199 ();
 sg13g2_fill_1 FILLER_45_201 ();
 sg13g2_fill_1 FILLER_45_245 ();
 sg13g2_fill_2 FILLER_45_298 ();
 sg13g2_fill_1 FILLER_45_300 ();
 sg13g2_fill_1 FILLER_45_318 ();
 sg13g2_fill_1 FILLER_45_328 ();
 sg13g2_fill_2 FILLER_45_390 ();
 sg13g2_fill_1 FILLER_45_392 ();
 sg13g2_fill_1 FILLER_45_424 ();
 sg13g2_fill_2 FILLER_45_429 ();
 sg13g2_decap_8 FILLER_45_440 ();
 sg13g2_decap_4 FILLER_45_447 ();
 sg13g2_fill_1 FILLER_45_451 ();
 sg13g2_fill_2 FILLER_45_456 ();
 sg13g2_fill_1 FILLER_45_489 ();
 sg13g2_fill_2 FILLER_45_499 ();
 sg13g2_fill_1 FILLER_45_501 ();
 sg13g2_fill_2 FILLER_45_517 ();
 sg13g2_fill_2 FILLER_45_554 ();
 sg13g2_fill_2 FILLER_45_583 ();
 sg13g2_decap_8 FILLER_45_613 ();
 sg13g2_decap_8 FILLER_45_620 ();
 sg13g2_fill_1 FILLER_45_627 ();
 sg13g2_fill_2 FILLER_45_646 ();
 sg13g2_fill_1 FILLER_45_648 ();
 sg13g2_fill_2 FILLER_45_663 ();
 sg13g2_fill_1 FILLER_45_665 ();
 sg13g2_fill_1 FILLER_45_697 ();
 sg13g2_fill_2 FILLER_45_711 ();
 sg13g2_fill_2 FILLER_45_793 ();
 sg13g2_fill_1 FILLER_45_795 ();
 sg13g2_fill_2 FILLER_45_805 ();
 sg13g2_fill_1 FILLER_45_811 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_38 ();
 sg13g2_fill_1 FILLER_46_118 ();
 sg13g2_decap_4 FILLER_46_140 ();
 sg13g2_fill_2 FILLER_46_144 ();
 sg13g2_decap_8 FILLER_46_173 ();
 sg13g2_fill_1 FILLER_46_180 ();
 sg13g2_fill_1 FILLER_46_194 ();
 sg13g2_decap_4 FILLER_46_225 ();
 sg13g2_fill_1 FILLER_46_229 ();
 sg13g2_decap_8 FILLER_46_251 ();
 sg13g2_decap_8 FILLER_46_258 ();
 sg13g2_fill_2 FILLER_46_265 ();
 sg13g2_fill_2 FILLER_46_271 ();
 sg13g2_fill_1 FILLER_46_273 ();
 sg13g2_fill_2 FILLER_46_295 ();
 sg13g2_fill_1 FILLER_46_297 ();
 sg13g2_fill_1 FILLER_46_328 ();
 sg13g2_fill_2 FILLER_46_334 ();
 sg13g2_fill_2 FILLER_46_354 ();
 sg13g2_fill_1 FILLER_46_382 ();
 sg13g2_fill_2 FILLER_46_419 ();
 sg13g2_fill_1 FILLER_46_466 ();
 sg13g2_fill_2 FILLER_46_516 ();
 sg13g2_fill_2 FILLER_46_523 ();
 sg13g2_fill_2 FILLER_46_529 ();
 sg13g2_fill_1 FILLER_46_531 ();
 sg13g2_fill_2 FILLER_46_586 ();
 sg13g2_decap_4 FILLER_46_620 ();
 sg13g2_fill_1 FILLER_46_624 ();
 sg13g2_fill_1 FILLER_46_643 ();
 sg13g2_fill_1 FILLER_46_785 ();
 sg13g2_decap_8 FILLER_46_812 ();
 sg13g2_decap_8 FILLER_46_819 ();
 sg13g2_fill_1 FILLER_46_826 ();
 sg13g2_decap_4 FILLER_46_857 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_decap_4 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_4 ();
 sg13g2_fill_1 FILLER_47_44 ();
 sg13g2_fill_1 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_138 ();
 sg13g2_decap_4 FILLER_47_191 ();
 sg13g2_fill_2 FILLER_47_204 ();
 sg13g2_fill_1 FILLER_47_206 ();
 sg13g2_fill_1 FILLER_47_212 ();
 sg13g2_decap_8 FILLER_47_243 ();
 sg13g2_fill_2 FILLER_47_250 ();
 sg13g2_fill_1 FILLER_47_356 ();
 sg13g2_fill_2 FILLER_47_362 ();
 sg13g2_decap_8 FILLER_47_377 ();
 sg13g2_fill_2 FILLER_47_384 ();
 sg13g2_fill_2 FILLER_47_390 ();
 sg13g2_fill_1 FILLER_47_392 ();
 sg13g2_decap_4 FILLER_47_450 ();
 sg13g2_fill_1 FILLER_47_490 ();
 sg13g2_fill_2 FILLER_47_557 ();
 sg13g2_fill_1 FILLER_47_559 ();
 sg13g2_fill_2 FILLER_47_592 ();
 sg13g2_decap_4 FILLER_47_613 ();
 sg13g2_fill_1 FILLER_47_652 ();
 sg13g2_fill_2 FILLER_47_663 ();
 sg13g2_decap_4 FILLER_47_703 ();
 sg13g2_fill_1 FILLER_47_707 ();
 sg13g2_decap_4 FILLER_47_712 ();
 sg13g2_fill_1 FILLER_47_716 ();
 sg13g2_fill_2 FILLER_47_738 ();
 sg13g2_decap_8 FILLER_47_761 ();
 sg13g2_decap_4 FILLER_47_768 ();
 sg13g2_fill_1 FILLER_47_772 ();
 sg13g2_fill_2 FILLER_47_797 ();
 sg13g2_decap_8 FILLER_47_820 ();
 sg13g2_decap_8 FILLER_47_827 ();
 sg13g2_fill_2 FILLER_47_834 ();
 sg13g2_fill_1 FILLER_47_836 ();
 sg13g2_fill_2 FILLER_47_860 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_4 ();
 sg13g2_decap_4 FILLER_48_98 ();
 sg13g2_fill_2 FILLER_48_102 ();
 sg13g2_decap_8 FILLER_48_251 ();
 sg13g2_fill_2 FILLER_48_258 ();
 sg13g2_fill_1 FILLER_48_269 ();
 sg13g2_fill_1 FILLER_48_300 ();
 sg13g2_fill_1 FILLER_48_340 ();
 sg13g2_decap_8 FILLER_48_345 ();
 sg13g2_decap_8 FILLER_48_352 ();
 sg13g2_fill_1 FILLER_48_359 ();
 sg13g2_fill_2 FILLER_48_395 ();
 sg13g2_fill_1 FILLER_48_397 ();
 sg13g2_decap_4 FILLER_48_408 ();
 sg13g2_fill_2 FILLER_48_412 ();
 sg13g2_fill_1 FILLER_48_419 ();
 sg13g2_decap_8 FILLER_48_433 ();
 sg13g2_decap_4 FILLER_48_440 ();
 sg13g2_fill_1 FILLER_48_444 ();
 sg13g2_fill_1 FILLER_48_515 ();
 sg13g2_fill_2 FILLER_48_595 ();
 sg13g2_fill_1 FILLER_48_649 ();
 sg13g2_fill_2 FILLER_48_677 ();
 sg13g2_fill_1 FILLER_48_679 ();
 sg13g2_decap_8 FILLER_48_773 ();
 sg13g2_fill_2 FILLER_48_780 ();
 sg13g2_fill_1 FILLER_48_782 ();
 sg13g2_decap_4 FILLER_48_858 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_4 FILLER_49_7 ();
 sg13g2_fill_1 FILLER_49_11 ();
 sg13g2_fill_2 FILLER_49_29 ();
 sg13g2_fill_1 FILLER_49_31 ();
 sg13g2_decap_8 FILLER_49_50 ();
 sg13g2_fill_2 FILLER_49_57 ();
 sg13g2_decap_4 FILLER_49_68 ();
 sg13g2_fill_1 FILLER_49_76 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_fill_2 FILLER_49_105 ();
 sg13g2_fill_2 FILLER_49_128 ();
 sg13g2_fill_1 FILLER_49_130 ();
 sg13g2_decap_4 FILLER_49_139 ();
 sg13g2_fill_1 FILLER_49_143 ();
 sg13g2_fill_2 FILLER_49_171 ();
 sg13g2_fill_1 FILLER_49_178 ();
 sg13g2_fill_2 FILLER_49_224 ();
 sg13g2_fill_1 FILLER_49_226 ();
 sg13g2_fill_2 FILLER_49_252 ();
 sg13g2_decap_4 FILLER_49_280 ();
 sg13g2_fill_1 FILLER_49_284 ();
 sg13g2_fill_2 FILLER_49_311 ();
 sg13g2_decap_4 FILLER_49_317 ();
 sg13g2_decap_8 FILLER_49_356 ();
 sg13g2_fill_2 FILLER_49_363 ();
 sg13g2_fill_2 FILLER_49_384 ();
 sg13g2_fill_1 FILLER_49_386 ();
 sg13g2_decap_4 FILLER_49_392 ();
 sg13g2_fill_1 FILLER_49_396 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_fill_1 FILLER_49_409 ();
 sg13g2_fill_2 FILLER_49_428 ();
 sg13g2_fill_1 FILLER_49_430 ();
 sg13g2_fill_1 FILLER_49_467 ();
 sg13g2_fill_1 FILLER_49_477 ();
 sg13g2_fill_1 FILLER_49_514 ();
 sg13g2_fill_1 FILLER_49_532 ();
 sg13g2_fill_2 FILLER_49_595 ();
 sg13g2_fill_2 FILLER_49_638 ();
 sg13g2_fill_1 FILLER_49_640 ();
 sg13g2_fill_2 FILLER_49_676 ();
 sg13g2_fill_2 FILLER_49_686 ();
 sg13g2_fill_1 FILLER_49_688 ();
 sg13g2_decap_8 FILLER_49_710 ();
 sg13g2_decap_8 FILLER_49_717 ();
 sg13g2_decap_8 FILLER_49_724 ();
 sg13g2_fill_2 FILLER_49_731 ();
 sg13g2_fill_1 FILLER_49_733 ();
 sg13g2_fill_1 FILLER_49_755 ();
 sg13g2_fill_2 FILLER_49_777 ();
 sg13g2_fill_1 FILLER_49_779 ();
 sg13g2_decap_8 FILLER_49_800 ();
 sg13g2_decap_8 FILLER_49_807 ();
 sg13g2_decap_4 FILLER_49_814 ();
 sg13g2_fill_1 FILLER_49_818 ();
 sg13g2_fill_2 FILLER_49_840 ();
 sg13g2_fill_1 FILLER_49_842 ();
 sg13g2_decap_4 FILLER_49_858 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_fill_2 FILLER_50_14 ();
 sg13g2_fill_1 FILLER_50_85 ();
 sg13g2_decap_4 FILLER_50_100 ();
 sg13g2_fill_1 FILLER_50_104 ();
 sg13g2_fill_1 FILLER_50_113 ();
 sg13g2_fill_1 FILLER_50_118 ();
 sg13g2_fill_2 FILLER_50_140 ();
 sg13g2_fill_1 FILLER_50_208 ();
 sg13g2_fill_2 FILLER_50_217 ();
 sg13g2_fill_1 FILLER_50_219 ();
 sg13g2_fill_2 FILLER_50_225 ();
 sg13g2_decap_8 FILLER_50_248 ();
 sg13g2_fill_2 FILLER_50_255 ();
 sg13g2_fill_2 FILLER_50_300 ();
 sg13g2_decap_4 FILLER_50_337 ();
 sg13g2_decap_8 FILLER_50_345 ();
 sg13g2_fill_1 FILLER_50_368 ();
 sg13g2_decap_4 FILLER_50_381 ();
 sg13g2_fill_2 FILLER_50_405 ();
 sg13g2_fill_2 FILLER_50_425 ();
 sg13g2_fill_1 FILLER_50_427 ();
 sg13g2_fill_1 FILLER_50_449 ();
 sg13g2_fill_2 FILLER_50_458 ();
 sg13g2_fill_1 FILLER_50_460 ();
 sg13g2_decap_4 FILLER_50_505 ();
 sg13g2_fill_2 FILLER_50_509 ();
 sg13g2_fill_2 FILLER_50_554 ();
 sg13g2_fill_2 FILLER_50_691 ();
 sg13g2_fill_1 FILLER_50_693 ();
 sg13g2_decap_8 FILLER_50_748 ();
 sg13g2_fill_2 FILLER_50_755 ();
 sg13g2_fill_2 FILLER_50_773 ();
 sg13g2_fill_2 FILLER_50_790 ();
 sg13g2_fill_1 FILLER_50_792 ();
 sg13g2_decap_8 FILLER_50_797 ();
 sg13g2_fill_2 FILLER_50_804 ();
 sg13g2_fill_2 FILLER_50_818 ();
 sg13g2_fill_2 FILLER_50_830 ();
 sg13g2_fill_1 FILLER_50_832 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_7 ();
 sg13g2_fill_2 FILLER_51_15 ();
 sg13g2_decap_4 FILLER_51_48 ();
 sg13g2_fill_2 FILLER_51_65 ();
 sg13g2_fill_1 FILLER_51_67 ();
 sg13g2_fill_2 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_124 ();
 sg13g2_fill_2 FILLER_51_131 ();
 sg13g2_fill_1 FILLER_51_133 ();
 sg13g2_fill_1 FILLER_51_155 ();
 sg13g2_fill_2 FILLER_51_169 ();
 sg13g2_fill_2 FILLER_51_198 ();
 sg13g2_fill_1 FILLER_51_200 ();
 sg13g2_fill_2 FILLER_51_252 ();
 sg13g2_fill_2 FILLER_51_284 ();
 sg13g2_fill_1 FILLER_51_286 ();
 sg13g2_fill_1 FILLER_51_326 ();
 sg13g2_decap_4 FILLER_51_336 ();
 sg13g2_fill_2 FILLER_51_340 ();
 sg13g2_fill_1 FILLER_51_359 ();
 sg13g2_fill_2 FILLER_51_386 ();
 sg13g2_decap_8 FILLER_51_403 ();
 sg13g2_fill_2 FILLER_51_431 ();
 sg13g2_decap_8 FILLER_51_461 ();
 sg13g2_decap_4 FILLER_51_468 ();
 sg13g2_fill_1 FILLER_51_476 ();
 sg13g2_fill_1 FILLER_51_481 ();
 sg13g2_decap_4 FILLER_51_496 ();
 sg13g2_fill_2 FILLER_51_513 ();
 sg13g2_fill_1 FILLER_51_515 ();
 sg13g2_fill_2 FILLER_51_590 ();
 sg13g2_fill_1 FILLER_51_592 ();
 sg13g2_fill_1 FILLER_51_597 ();
 sg13g2_fill_1 FILLER_51_607 ();
 sg13g2_fill_2 FILLER_51_621 ();
 sg13g2_fill_1 FILLER_51_631 ();
 sg13g2_fill_2 FILLER_51_690 ();
 sg13g2_fill_1 FILLER_51_711 ();
 sg13g2_fill_2 FILLER_51_729 ();
 sg13g2_fill_1 FILLER_51_731 ();
 sg13g2_fill_2 FILLER_51_741 ();
 sg13g2_fill_2 FILLER_51_748 ();
 sg13g2_fill_1 FILLER_51_750 ();
 sg13g2_decap_8 FILLER_51_776 ();
 sg13g2_decap_4 FILLER_51_783 ();
 sg13g2_fill_1 FILLER_51_787 ();
 sg13g2_fill_1 FILLER_51_807 ();
 sg13g2_fill_2 FILLER_51_818 ();
 sg13g2_fill_1 FILLER_51_820 ();
 sg13g2_fill_2 FILLER_51_831 ();
 sg13g2_fill_1 FILLER_51_833 ();
 sg13g2_fill_2 FILLER_51_859 ();
 sg13g2_fill_1 FILLER_51_861 ();
 sg13g2_decap_8 FILLER_52_57 ();
 sg13g2_fill_1 FILLER_52_64 ();
 sg13g2_decap_4 FILLER_52_69 ();
 sg13g2_fill_1 FILLER_52_99 ();
 sg13g2_fill_1 FILLER_52_109 ();
 sg13g2_fill_2 FILLER_52_140 ();
 sg13g2_fill_1 FILLER_52_142 ();
 sg13g2_fill_1 FILLER_52_164 ();
 sg13g2_fill_2 FILLER_52_171 ();
 sg13g2_fill_2 FILLER_52_197 ();
 sg13g2_fill_2 FILLER_52_212 ();
 sg13g2_fill_2 FILLER_52_219 ();
 sg13g2_fill_1 FILLER_52_221 ();
 sg13g2_fill_2 FILLER_52_240 ();
 sg13g2_fill_1 FILLER_52_242 ();
 sg13g2_fill_1 FILLER_52_248 ();
 sg13g2_fill_2 FILLER_52_254 ();
 sg13g2_fill_1 FILLER_52_256 ();
 sg13g2_decap_8 FILLER_52_275 ();
 sg13g2_decap_4 FILLER_52_282 ();
 sg13g2_fill_2 FILLER_52_291 ();
 sg13g2_fill_1 FILLER_52_306 ();
 sg13g2_decap_8 FILLER_52_311 ();
 sg13g2_decap_8 FILLER_52_318 ();
 sg13g2_fill_2 FILLER_52_325 ();
 sg13g2_fill_1 FILLER_52_327 ();
 sg13g2_fill_2 FILLER_52_371 ();
 sg13g2_fill_1 FILLER_52_373 ();
 sg13g2_decap_4 FILLER_52_387 ();
 sg13g2_decap_8 FILLER_52_396 ();
 sg13g2_decap_4 FILLER_52_403 ();
 sg13g2_decap_4 FILLER_52_429 ();
 sg13g2_fill_2 FILLER_52_433 ();
 sg13g2_decap_4 FILLER_52_455 ();
 sg13g2_fill_1 FILLER_52_459 ();
 sg13g2_fill_1 FILLER_52_522 ();
 sg13g2_decap_4 FILLER_52_561 ();
 sg13g2_fill_1 FILLER_52_565 ();
 sg13g2_fill_2 FILLER_52_570 ();
 sg13g2_fill_1 FILLER_52_637 ();
 sg13g2_fill_1 FILLER_52_660 ();
 sg13g2_fill_1 FILLER_52_665 ();
 sg13g2_fill_2 FILLER_52_695 ();
 sg13g2_fill_1 FILLER_52_697 ();
 sg13g2_fill_2 FILLER_52_733 ();
 sg13g2_fill_1 FILLER_52_756 ();
 sg13g2_fill_2 FILLER_52_775 ();
 sg13g2_fill_1 FILLER_52_777 ();
 sg13g2_fill_1 FILLER_52_782 ();
 sg13g2_decap_4 FILLER_52_806 ();
 sg13g2_decap_8 FILLER_52_819 ();
 sg13g2_fill_1 FILLER_52_826 ();
 sg13g2_fill_2 FILLER_52_842 ();
 sg13g2_decap_4 FILLER_52_858 ();
 sg13g2_fill_2 FILLER_53_26 ();
 sg13g2_fill_2 FILLER_53_41 ();
 sg13g2_fill_1 FILLER_53_73 ();
 sg13g2_fill_2 FILLER_53_96 ();
 sg13g2_fill_1 FILLER_53_98 ();
 sg13g2_fill_1 FILLER_53_108 ();
 sg13g2_decap_4 FILLER_53_135 ();
 sg13g2_fill_2 FILLER_53_139 ();
 sg13g2_decap_4 FILLER_53_254 ();
 sg13g2_fill_1 FILLER_53_310 ();
 sg13g2_fill_2 FILLER_53_382 ();
 sg13g2_fill_2 FILLER_53_411 ();
 sg13g2_fill_1 FILLER_53_413 ();
 sg13g2_decap_8 FILLER_53_419 ();
 sg13g2_decap_4 FILLER_53_426 ();
 sg13g2_fill_2 FILLER_53_430 ();
 sg13g2_decap_8 FILLER_53_445 ();
 sg13g2_fill_2 FILLER_53_472 ();
 sg13g2_fill_2 FILLER_53_503 ();
 sg13g2_fill_1 FILLER_53_505 ();
 sg13g2_decap_4 FILLER_53_526 ();
 sg13g2_fill_1 FILLER_53_592 ();
 sg13g2_fill_1 FILLER_53_611 ();
 sg13g2_fill_2 FILLER_53_624 ();
 sg13g2_fill_1 FILLER_53_626 ();
 sg13g2_fill_2 FILLER_53_641 ();
 sg13g2_fill_1 FILLER_53_643 ();
 sg13g2_fill_2 FILLER_53_655 ();
 sg13g2_fill_1 FILLER_53_657 ();
 sg13g2_fill_1 FILLER_53_677 ();
 sg13g2_fill_2 FILLER_53_695 ();
 sg13g2_fill_2 FILLER_53_722 ();
 sg13g2_fill_1 FILLER_53_724 ();
 sg13g2_fill_1 FILLER_53_730 ();
 sg13g2_fill_2 FILLER_53_755 ();
 sg13g2_fill_1 FILLER_53_766 ();
 sg13g2_fill_1 FILLER_53_789 ();
 sg13g2_fill_2 FILLER_53_795 ();
 sg13g2_fill_1 FILLER_53_797 ();
 sg13g2_decap_8 FILLER_53_813 ();
 sg13g2_fill_1 FILLER_53_830 ();
 sg13g2_fill_2 FILLER_53_841 ();
 sg13g2_decap_8 FILLER_53_853 ();
 sg13g2_fill_2 FILLER_53_860 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_decap_4 FILLER_54_72 ();
 sg13g2_fill_1 FILLER_54_76 ();
 sg13g2_fill_2 FILLER_54_103 ();
 sg13g2_fill_2 FILLER_54_141 ();
 sg13g2_decap_8 FILLER_54_206 ();
 sg13g2_decap_4 FILLER_54_218 ();
 sg13g2_fill_2 FILLER_54_222 ();
 sg13g2_fill_1 FILLER_54_229 ();
 sg13g2_fill_1 FILLER_54_238 ();
 sg13g2_decap_4 FILLER_54_257 ();
 sg13g2_fill_1 FILLER_54_266 ();
 sg13g2_fill_1 FILLER_54_275 ();
 sg13g2_fill_1 FILLER_54_285 ();
 sg13g2_fill_1 FILLER_54_290 ();
 sg13g2_fill_1 FILLER_54_330 ();
 sg13g2_decap_4 FILLER_54_397 ();
 sg13g2_fill_1 FILLER_54_410 ();
 sg13g2_decap_8 FILLER_54_432 ();
 sg13g2_fill_2 FILLER_54_439 ();
 sg13g2_fill_1 FILLER_54_441 ();
 sg13g2_decap_4 FILLER_54_452 ();
 sg13g2_fill_1 FILLER_54_456 ();
 sg13g2_fill_2 FILLER_54_483 ();
 sg13g2_fill_1 FILLER_54_485 ();
 sg13g2_fill_2 FILLER_54_522 ();
 sg13g2_fill_2 FILLER_54_550 ();
 sg13g2_decap_4 FILLER_54_561 ();
 sg13g2_fill_1 FILLER_54_565 ();
 sg13g2_fill_2 FILLER_54_627 ();
 sg13g2_fill_1 FILLER_54_629 ();
 sg13g2_decap_8 FILLER_54_689 ();
 sg13g2_decap_8 FILLER_54_696 ();
 sg13g2_decap_4 FILLER_54_712 ();
 sg13g2_decap_4 FILLER_54_724 ();
 sg13g2_decap_8 FILLER_54_752 ();
 sg13g2_decap_8 FILLER_54_759 ();
 sg13g2_decap_8 FILLER_54_766 ();
 sg13g2_fill_1 FILLER_54_773 ();
 sg13g2_fill_1 FILLER_54_788 ();
 sg13g2_fill_2 FILLER_54_798 ();
 sg13g2_fill_1 FILLER_54_800 ();
 sg13g2_fill_2 FILLER_54_816 ();
 sg13g2_fill_2 FILLER_54_828 ();
 sg13g2_fill_2 FILLER_54_860 ();
 sg13g2_fill_1 FILLER_55_26 ();
 sg13g2_fill_2 FILLER_55_32 ();
 sg13g2_fill_1 FILLER_55_34 ();
 sg13g2_fill_2 FILLER_55_39 ();
 sg13g2_fill_1 FILLER_55_50 ();
 sg13g2_decap_8 FILLER_55_72 ();
 sg13g2_decap_4 FILLER_55_79 ();
 sg13g2_fill_1 FILLER_55_83 ();
 sg13g2_fill_2 FILLER_55_92 ();
 sg13g2_fill_1 FILLER_55_94 ();
 sg13g2_fill_1 FILLER_55_99 ();
 sg13g2_decap_8 FILLER_55_109 ();
 sg13g2_fill_2 FILLER_55_116 ();
 sg13g2_fill_2 FILLER_55_148 ();
 sg13g2_fill_1 FILLER_55_158 ();
 sg13g2_decap_8 FILLER_55_165 ();
 sg13g2_fill_1 FILLER_55_172 ();
 sg13g2_fill_2 FILLER_55_187 ();
 sg13g2_fill_1 FILLER_55_189 ();
 sg13g2_fill_2 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_296 ();
 sg13g2_decap_4 FILLER_55_303 ();
 sg13g2_fill_1 FILLER_55_363 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_fill_1 FILLER_55_409 ();
 sg13g2_fill_1 FILLER_55_422 ();
 sg13g2_fill_1 FILLER_55_435 ();
 sg13g2_fill_2 FILLER_55_446 ();
 sg13g2_fill_2 FILLER_55_477 ();
 sg13g2_decap_8 FILLER_55_502 ();
 sg13g2_fill_1 FILLER_55_509 ();
 sg13g2_fill_1 FILLER_55_519 ();
 sg13g2_decap_4 FILLER_55_529 ();
 sg13g2_fill_2 FILLER_55_533 ();
 sg13g2_decap_4 FILLER_55_614 ();
 sg13g2_fill_2 FILLER_55_618 ();
 sg13g2_fill_2 FILLER_55_659 ();
 sg13g2_fill_2 FILLER_55_671 ();
 sg13g2_fill_2 FILLER_55_707 ();
 sg13g2_fill_1 FILLER_55_709 ();
 sg13g2_fill_2 FILLER_55_730 ();
 sg13g2_decap_4 FILLER_55_757 ();
 sg13g2_fill_2 FILLER_55_801 ();
 sg13g2_decap_4 FILLER_55_813 ();
 sg13g2_fill_2 FILLER_55_835 ();
 sg13g2_fill_1 FILLER_55_841 ();
 sg13g2_decap_4 FILLER_55_857 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_4 FILLER_56_11 ();
 sg13g2_decap_4 FILLER_56_45 ();
 sg13g2_fill_2 FILLER_56_70 ();
 sg13g2_fill_1 FILLER_56_72 ();
 sg13g2_decap_8 FILLER_56_107 ();
 sg13g2_decap_8 FILLER_56_114 ();
 sg13g2_decap_8 FILLER_56_121 ();
 sg13g2_decap_4 FILLER_56_128 ();
 sg13g2_decap_8 FILLER_56_165 ();
 sg13g2_fill_2 FILLER_56_178 ();
 sg13g2_fill_1 FILLER_56_180 ();
 sg13g2_fill_1 FILLER_56_189 ();
 sg13g2_decap_8 FILLER_56_213 ();
 sg13g2_fill_2 FILLER_56_239 ();
 sg13g2_fill_1 FILLER_56_241 ();
 sg13g2_fill_1 FILLER_56_276 ();
 sg13g2_fill_2 FILLER_56_298 ();
 sg13g2_fill_1 FILLER_56_300 ();
 sg13g2_fill_1 FILLER_56_327 ();
 sg13g2_fill_2 FILLER_56_354 ();
 sg13g2_decap_4 FILLER_56_398 ();
 sg13g2_fill_1 FILLER_56_402 ();
 sg13g2_fill_1 FILLER_56_417 ();
 sg13g2_decap_4 FILLER_56_433 ();
 sg13g2_fill_2 FILLER_56_437 ();
 sg13g2_decap_8 FILLER_56_447 ();
 sg13g2_decap_4 FILLER_56_528 ();
 sg13g2_fill_1 FILLER_56_562 ();
 sg13g2_fill_2 FILLER_56_572 ();
 sg13g2_fill_2 FILLER_56_587 ();
 sg13g2_fill_1 FILLER_56_589 ();
 sg13g2_fill_1 FILLER_56_636 ();
 sg13g2_fill_1 FILLER_56_656 ();
 sg13g2_fill_2 FILLER_56_662 ();
 sg13g2_fill_2 FILLER_56_681 ();
 sg13g2_fill_1 FILLER_56_683 ();
 sg13g2_decap_8 FILLER_56_688 ();
 sg13g2_decap_8 FILLER_56_695 ();
 sg13g2_fill_1 FILLER_56_711 ();
 sg13g2_fill_2 FILLER_56_731 ();
 sg13g2_fill_1 FILLER_56_733 ();
 sg13g2_decap_8 FILLER_56_744 ();
 sg13g2_decap_8 FILLER_56_751 ();
 sg13g2_fill_1 FILLER_56_758 ();
 sg13g2_fill_2 FILLER_56_764 ();
 sg13g2_decap_4 FILLER_56_788 ();
 sg13g2_decap_4 FILLER_56_796 ();
 sg13g2_fill_2 FILLER_56_800 ();
 sg13g2_decap_4 FILLER_56_827 ();
 sg13g2_fill_1 FILLER_56_831 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_7 ();
 sg13g2_fill_1 FILLER_57_30 ();
 sg13g2_fill_2 FILLER_57_79 ();
 sg13g2_fill_1 FILLER_57_81 ();
 sg13g2_fill_2 FILLER_57_91 ();
 sg13g2_decap_4 FILLER_57_123 ();
 sg13g2_fill_1 FILLER_57_127 ();
 sg13g2_fill_1 FILLER_57_197 ();
 sg13g2_decap_8 FILLER_57_206 ();
 sg13g2_decap_8 FILLER_57_221 ();
 sg13g2_decap_8 FILLER_57_228 ();
 sg13g2_decap_4 FILLER_57_235 ();
 sg13g2_fill_1 FILLER_57_239 ();
 sg13g2_decap_4 FILLER_57_270 ();
 sg13g2_fill_1 FILLER_57_295 ();
 sg13g2_decap_4 FILLER_57_304 ();
 sg13g2_fill_2 FILLER_57_346 ();
 sg13g2_fill_2 FILLER_57_365 ();
 sg13g2_fill_1 FILLER_57_367 ();
 sg13g2_decap_8 FILLER_57_393 ();
 sg13g2_decap_8 FILLER_57_400 ();
 sg13g2_fill_1 FILLER_57_407 ();
 sg13g2_fill_1 FILLER_57_425 ();
 sg13g2_fill_2 FILLER_57_435 ();
 sg13g2_decap_4 FILLER_57_452 ();
 sg13g2_fill_2 FILLER_57_456 ();
 sg13g2_fill_2 FILLER_57_468 ();
 sg13g2_decap_4 FILLER_57_506 ();
 sg13g2_fill_2 FILLER_57_519 ();
 sg13g2_fill_2 FILLER_57_547 ();
 sg13g2_fill_1 FILLER_57_549 ();
 sg13g2_fill_1 FILLER_57_565 ();
 sg13g2_fill_2 FILLER_57_575 ();
 sg13g2_decap_4 FILLER_57_613 ();
 sg13g2_fill_1 FILLER_57_617 ();
 sg13g2_decap_8 FILLER_57_629 ();
 sg13g2_decap_4 FILLER_57_636 ();
 sg13g2_fill_1 FILLER_57_640 ();
 sg13g2_fill_1 FILLER_57_645 ();
 sg13g2_fill_2 FILLER_57_664 ();
 sg13g2_decap_4 FILLER_57_697 ();
 sg13g2_fill_1 FILLER_57_701 ();
 sg13g2_fill_1 FILLER_57_732 ();
 sg13g2_decap_8 FILLER_57_743 ();
 sg13g2_decap_4 FILLER_57_750 ();
 sg13g2_fill_1 FILLER_57_767 ();
 sg13g2_fill_2 FILLER_57_774 ();
 sg13g2_fill_1 FILLER_57_776 ();
 sg13g2_fill_2 FILLER_57_781 ();
 sg13g2_fill_1 FILLER_57_783 ();
 sg13g2_fill_1 FILLER_57_789 ();
 sg13g2_decap_4 FILLER_57_808 ();
 sg13g2_decap_4 FILLER_57_817 ();
 sg13g2_decap_8 FILLER_57_831 ();
 sg13g2_fill_2 FILLER_57_838 ();
 sg13g2_decap_8 FILLER_57_844 ();
 sg13g2_decap_8 FILLER_57_851 ();
 sg13g2_decap_4 FILLER_57_858 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_4 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_29 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_fill_1 FILLER_58_63 ();
 sg13g2_fill_2 FILLER_58_90 ();
 sg13g2_fill_1 FILLER_58_92 ();
 sg13g2_fill_2 FILLER_58_123 ();
 sg13g2_fill_1 FILLER_58_125 ();
 sg13g2_fill_2 FILLER_58_152 ();
 sg13g2_fill_1 FILLER_58_154 ();
 sg13g2_fill_1 FILLER_58_164 ();
 sg13g2_fill_1 FILLER_58_171 ();
 sg13g2_fill_1 FILLER_58_213 ();
 sg13g2_fill_2 FILLER_58_245 ();
 sg13g2_decap_4 FILLER_58_255 ();
 sg13g2_fill_1 FILLER_58_259 ();
 sg13g2_decap_8 FILLER_58_342 ();
 sg13g2_fill_2 FILLER_58_349 ();
 sg13g2_decap_8 FILLER_58_386 ();
 sg13g2_decap_8 FILLER_58_393 ();
 sg13g2_decap_8 FILLER_58_400 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_fill_1 FILLER_58_409 ();
 sg13g2_fill_2 FILLER_58_440 ();
 sg13g2_decap_8 FILLER_58_452 ();
 sg13g2_decap_4 FILLER_58_459 ();
 sg13g2_fill_1 FILLER_58_463 ();
 sg13g2_decap_8 FILLER_58_503 ();
 sg13g2_decap_4 FILLER_58_510 ();
 sg13g2_fill_1 FILLER_58_514 ();
 sg13g2_fill_1 FILLER_58_541 ();
 sg13g2_fill_2 FILLER_58_550 ();
 sg13g2_fill_2 FILLER_58_610 ();
 sg13g2_decap_4 FILLER_58_625 ();
 sg13g2_fill_2 FILLER_58_654 ();
 sg13g2_fill_1 FILLER_58_656 ();
 sg13g2_decap_8 FILLER_58_681 ();
 sg13g2_decap_4 FILLER_58_688 ();
 sg13g2_decap_8 FILLER_58_701 ();
 sg13g2_fill_2 FILLER_58_708 ();
 sg13g2_fill_2 FILLER_58_729 ();
 sg13g2_fill_1 FILLER_58_731 ();
 sg13g2_fill_2 FILLER_58_741 ();
 sg13g2_fill_2 FILLER_58_751 ();
 sg13g2_fill_1 FILLER_58_753 ();
 sg13g2_decap_4 FILLER_58_762 ();
 sg13g2_fill_2 FILLER_58_782 ();
 sg13g2_fill_1 FILLER_58_784 ();
 sg13g2_decap_8 FILLER_58_803 ();
 sg13g2_decap_4 FILLER_58_810 ();
 sg13g2_fill_1 FILLER_58_839 ();
 sg13g2_decap_8 FILLER_58_855 ();
 sg13g2_fill_2 FILLER_59_39 ();
 sg13g2_fill_2 FILLER_59_45 ();
 sg13g2_fill_1 FILLER_59_47 ();
 sg13g2_fill_2 FILLER_59_82 ();
 sg13g2_fill_1 FILLER_59_84 ();
 sg13g2_fill_2 FILLER_59_137 ();
 sg13g2_fill_1 FILLER_59_139 ();
 sg13g2_decap_4 FILLER_59_180 ();
 sg13g2_fill_1 FILLER_59_184 ();
 sg13g2_fill_2 FILLER_59_190 ();
 sg13g2_decap_8 FILLER_59_197 ();
 sg13g2_decap_8 FILLER_59_204 ();
 sg13g2_decap_4 FILLER_59_211 ();
 sg13g2_decap_4 FILLER_59_228 ();
 sg13g2_fill_2 FILLER_59_232 ();
 sg13g2_decap_8 FILLER_59_263 ();
 sg13g2_decap_4 FILLER_59_270 ();
 sg13g2_decap_4 FILLER_59_295 ();
 sg13g2_fill_2 FILLER_59_299 ();
 sg13g2_fill_1 FILLER_59_323 ();
 sg13g2_fill_2 FILLER_59_350 ();
 sg13g2_decap_8 FILLER_59_403 ();
 sg13g2_fill_2 FILLER_59_410 ();
 sg13g2_fill_1 FILLER_59_412 ();
 sg13g2_fill_1 FILLER_59_418 ();
 sg13g2_decap_4 FILLER_59_441 ();
 sg13g2_fill_1 FILLER_59_445 ();
 sg13g2_fill_2 FILLER_59_557 ();
 sg13g2_fill_2 FILLER_59_581 ();
 sg13g2_decap_8 FILLER_59_630 ();
 sg13g2_decap_4 FILLER_59_637 ();
 sg13g2_fill_1 FILLER_59_641 ();
 sg13g2_fill_2 FILLER_59_659 ();
 sg13g2_fill_1 FILLER_59_661 ();
 sg13g2_fill_2 FILLER_59_667 ();
 sg13g2_fill_2 FILLER_59_723 ();
 sg13g2_fill_1 FILLER_59_725 ();
 sg13g2_decap_8 FILLER_59_736 ();
 sg13g2_fill_2 FILLER_59_743 ();
 sg13g2_fill_1 FILLER_59_745 ();
 sg13g2_fill_1 FILLER_59_750 ();
 sg13g2_fill_1 FILLER_59_759 ();
 sg13g2_fill_1 FILLER_59_769 ();
 sg13g2_decap_4 FILLER_59_800 ();
 sg13g2_fill_1 FILLER_59_804 ();
 sg13g2_decap_4 FILLER_59_810 ();
 sg13g2_fill_1 FILLER_59_814 ();
 sg13g2_decap_4 FILLER_59_834 ();
 sg13g2_fill_1 FILLER_59_838 ();
 sg13g2_fill_2 FILLER_59_859 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_fill_2 FILLER_60_26 ();
 sg13g2_fill_1 FILLER_60_28 ();
 sg13g2_fill_2 FILLER_60_50 ();
 sg13g2_fill_1 FILLER_60_73 ();
 sg13g2_fill_2 FILLER_60_82 ();
 sg13g2_fill_1 FILLER_60_84 ();
 sg13g2_fill_1 FILLER_60_95 ();
 sg13g2_fill_1 FILLER_60_101 ();
 sg13g2_fill_2 FILLER_60_116 ();
 sg13g2_fill_1 FILLER_60_118 ();
 sg13g2_fill_1 FILLER_60_164 ();
 sg13g2_decap_8 FILLER_60_173 ();
 sg13g2_fill_2 FILLER_60_180 ();
 sg13g2_fill_2 FILLER_60_192 ();
 sg13g2_decap_8 FILLER_60_208 ();
 sg13g2_fill_1 FILLER_60_215 ();
 sg13g2_fill_2 FILLER_60_226 ();
 sg13g2_decap_8 FILLER_60_236 ();
 sg13g2_decap_4 FILLER_60_269 ();
 sg13g2_fill_1 FILLER_60_273 ();
 sg13g2_decap_4 FILLER_60_295 ();
 sg13g2_fill_1 FILLER_60_329 ();
 sg13g2_fill_1 FILLER_60_369 ();
 sg13g2_fill_1 FILLER_60_441 ();
 sg13g2_fill_2 FILLER_60_462 ();
 sg13g2_fill_1 FILLER_60_503 ();
 sg13g2_fill_1 FILLER_60_610 ();
 sg13g2_fill_1 FILLER_60_624 ();
 sg13g2_decap_8 FILLER_60_641 ();
 sg13g2_fill_1 FILLER_60_648 ();
 sg13g2_fill_1 FILLER_60_669 ();
 sg13g2_fill_2 FILLER_60_701 ();
 sg13g2_fill_2 FILLER_60_712 ();
 sg13g2_fill_2 FILLER_60_719 ();
 sg13g2_fill_1 FILLER_60_744 ();
 sg13g2_fill_1 FILLER_60_750 ();
 sg13g2_decap_4 FILLER_60_756 ();
 sg13g2_decap_4 FILLER_60_776 ();
 sg13g2_fill_2 FILLER_60_780 ();
 sg13g2_fill_2 FILLER_60_791 ();
 sg13g2_decap_8 FILLER_60_804 ();
 sg13g2_fill_2 FILLER_60_841 ();
 sg13g2_fill_1 FILLER_60_843 ();
 sg13g2_decap_4 FILLER_60_857 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_7 ();
 sg13g2_fill_1 FILLER_61_15 ();
 sg13g2_fill_2 FILLER_61_47 ();
 sg13g2_fill_1 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_71 ();
 sg13g2_fill_1 FILLER_61_78 ();
 sg13g2_fill_1 FILLER_61_113 ();
 sg13g2_fill_1 FILLER_61_124 ();
 sg13g2_fill_2 FILLER_61_130 ();
 sg13g2_fill_2 FILLER_61_161 ();
 sg13g2_fill_1 FILLER_61_163 ();
 sg13g2_fill_1 FILLER_61_174 ();
 sg13g2_decap_8 FILLER_61_179 ();
 sg13g2_fill_1 FILLER_61_186 ();
 sg13g2_decap_8 FILLER_61_231 ();
 sg13g2_fill_1 FILLER_61_238 ();
 sg13g2_fill_1 FILLER_61_253 ();
 sg13g2_decap_8 FILLER_61_271 ();
 sg13g2_decap_4 FILLER_61_278 ();
 sg13g2_fill_1 FILLER_61_282 ();
 sg13g2_decap_4 FILLER_61_304 ();
 sg13g2_fill_2 FILLER_61_308 ();
 sg13g2_fill_1 FILLER_61_314 ();
 sg13g2_decap_4 FILLER_61_346 ();
 sg13g2_fill_2 FILLER_61_350 ();
 sg13g2_fill_2 FILLER_61_408 ();
 sg13g2_fill_1 FILLER_61_410 ();
 sg13g2_decap_8 FILLER_61_433 ();
 sg13g2_decap_8 FILLER_61_440 ();
 sg13g2_fill_2 FILLER_61_447 ();
 sg13g2_fill_1 FILLER_61_449 ();
 sg13g2_fill_1 FILLER_61_465 ();
 sg13g2_fill_2 FILLER_61_475 ();
 sg13g2_fill_2 FILLER_61_518 ();
 sg13g2_fill_2 FILLER_61_533 ();
 sg13g2_fill_1 FILLER_61_535 ();
 sg13g2_fill_1 FILLER_61_546 ();
 sg13g2_fill_1 FILLER_61_580 ();
 sg13g2_fill_2 FILLER_61_654 ();
 sg13g2_decap_4 FILLER_61_699 ();
 sg13g2_fill_2 FILLER_61_703 ();
 sg13g2_fill_1 FILLER_61_728 ();
 sg13g2_decap_8 FILLER_61_740 ();
 sg13g2_fill_2 FILLER_61_771 ();
 sg13g2_fill_1 FILLER_61_773 ();
 sg13g2_fill_1 FILLER_61_820 ();
 sg13g2_decap_4 FILLER_61_832 ();
 sg13g2_decap_4 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_4 FILLER_62_77 ();
 sg13g2_fill_2 FILLER_62_81 ();
 sg13g2_fill_1 FILLER_62_113 ();
 sg13g2_decap_4 FILLER_62_131 ();
 sg13g2_fill_1 FILLER_62_160 ();
 sg13g2_fill_1 FILLER_62_171 ();
 sg13g2_fill_1 FILLER_62_178 ();
 sg13g2_decap_4 FILLER_62_187 ();
 sg13g2_decap_4 FILLER_62_201 ();
 sg13g2_fill_1 FILLER_62_205 ();
 sg13g2_fill_1 FILLER_62_228 ();
 sg13g2_fill_2 FILLER_62_234 ();
 sg13g2_fill_1 FILLER_62_236 ();
 sg13g2_fill_1 FILLER_62_273 ();
 sg13g2_decap_4 FILLER_62_278 ();
 sg13g2_fill_1 FILLER_62_282 ();
 sg13g2_fill_2 FILLER_62_308 ();
 sg13g2_fill_1 FILLER_62_310 ();
 sg13g2_fill_2 FILLER_62_341 ();
 sg13g2_fill_1 FILLER_62_343 ();
 sg13g2_fill_2 FILLER_62_349 ();
 sg13g2_fill_1 FILLER_62_403 ();
 sg13g2_fill_2 FILLER_62_408 ();
 sg13g2_fill_1 FILLER_62_410 ();
 sg13g2_fill_2 FILLER_62_419 ();
 sg13g2_fill_1 FILLER_62_473 ();
 sg13g2_fill_1 FILLER_62_492 ();
 sg13g2_fill_2 FILLER_62_595 ();
 sg13g2_fill_1 FILLER_62_597 ();
 sg13g2_fill_2 FILLER_62_624 ();
 sg13g2_fill_1 FILLER_62_626 ();
 sg13g2_fill_1 FILLER_62_632 ();
 sg13g2_decap_4 FILLER_62_689 ();
 sg13g2_decap_8 FILLER_62_717 ();
 sg13g2_fill_2 FILLER_62_724 ();
 sg13g2_fill_2 FILLER_62_741 ();
 sg13g2_decap_8 FILLER_62_753 ();
 sg13g2_fill_2 FILLER_62_764 ();
 sg13g2_decap_8 FILLER_62_776 ();
 sg13g2_decap_8 FILLER_62_783 ();
 sg13g2_decap_8 FILLER_62_790 ();
 sg13g2_decap_4 FILLER_62_797 ();
 sg13g2_decap_4 FILLER_62_825 ();
 sg13g2_decap_8 FILLER_62_855 ();
 sg13g2_decap_4 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_76 ();
 sg13g2_fill_1 FILLER_63_104 ();
 sg13g2_fill_2 FILLER_63_110 ();
 sg13g2_fill_1 FILLER_63_131 ();
 sg13g2_fill_1 FILLER_63_162 ();
 sg13g2_fill_2 FILLER_63_185 ();
 sg13g2_fill_1 FILLER_63_187 ();
 sg13g2_fill_2 FILLER_63_196 ();
 sg13g2_fill_1 FILLER_63_198 ();
 sg13g2_fill_2 FILLER_63_207 ();
 sg13g2_fill_1 FILLER_63_209 ();
 sg13g2_decap_8 FILLER_63_230 ();
 sg13g2_fill_2 FILLER_63_317 ();
 sg13g2_fill_1 FILLER_63_319 ();
 sg13g2_decap_8 FILLER_63_346 ();
 sg13g2_fill_2 FILLER_63_353 ();
 sg13g2_fill_1 FILLER_63_355 ();
 sg13g2_fill_2 FILLER_63_385 ();
 sg13g2_fill_2 FILLER_63_408 ();
 sg13g2_fill_1 FILLER_63_442 ();
 sg13g2_fill_2 FILLER_63_459 ();
 sg13g2_fill_1 FILLER_63_461 ();
 sg13g2_fill_1 FILLER_63_498 ();
 sg13g2_fill_2 FILLER_63_508 ();
 sg13g2_fill_1 FILLER_63_510 ();
 sg13g2_fill_2 FILLER_63_551 ();
 sg13g2_fill_2 FILLER_63_589 ();
 sg13g2_fill_1 FILLER_63_591 ();
 sg13g2_fill_2 FILLER_63_642 ();
 sg13g2_fill_1 FILLER_63_644 ();
 sg13g2_fill_1 FILLER_63_658 ();
 sg13g2_decap_4 FILLER_63_707 ();
 sg13g2_fill_2 FILLER_63_758 ();
 sg13g2_decap_4 FILLER_63_773 ();
 sg13g2_fill_1 FILLER_63_777 ();
 sg13g2_fill_1 FILLER_63_800 ();
 sg13g2_fill_2 FILLER_64_26 ();
 sg13g2_fill_1 FILLER_64_75 ();
 sg13g2_fill_1 FILLER_64_135 ();
 sg13g2_fill_2 FILLER_64_150 ();
 sg13g2_decap_8 FILLER_64_207 ();
 sg13g2_fill_1 FILLER_64_214 ();
 sg13g2_decap_4 FILLER_64_235 ();
 sg13g2_decap_4 FILLER_64_265 ();
 sg13g2_fill_1 FILLER_64_269 ();
 sg13g2_fill_1 FILLER_64_279 ();
 sg13g2_fill_1 FILLER_64_293 ();
 sg13g2_fill_1 FILLER_64_323 ();
 sg13g2_fill_1 FILLER_64_338 ();
 sg13g2_fill_2 FILLER_64_463 ();
 sg13g2_fill_1 FILLER_64_465 ();
 sg13g2_fill_1 FILLER_64_473 ();
 sg13g2_fill_1 FILLER_64_478 ();
 sg13g2_fill_1 FILLER_64_531 ();
 sg13g2_fill_1 FILLER_64_541 ();
 sg13g2_fill_1 FILLER_64_572 ();
 sg13g2_fill_1 FILLER_64_617 ();
 sg13g2_fill_2 FILLER_64_681 ();
 sg13g2_fill_1 FILLER_64_683 ();
 sg13g2_fill_2 FILLER_64_697 ();
 sg13g2_decap_4 FILLER_64_722 ();
 sg13g2_fill_2 FILLER_64_726 ();
 sg13g2_fill_2 FILLER_64_748 ();
 sg13g2_fill_1 FILLER_64_750 ();
 sg13g2_decap_4 FILLER_64_757 ();
 sg13g2_fill_2 FILLER_64_761 ();
 sg13g2_fill_1 FILLER_64_767 ();
 sg13g2_fill_1 FILLER_64_773 ();
 sg13g2_fill_1 FILLER_64_778 ();
 sg13g2_fill_2 FILLER_64_791 ();
 sg13g2_fill_2 FILLER_64_812 ();
 sg13g2_fill_1 FILLER_64_814 ();
 sg13g2_fill_2 FILLER_64_825 ();
 sg13g2_fill_2 FILLER_64_837 ();
 sg13g2_fill_1 FILLER_64_839 ();
 sg13g2_decap_4 FILLER_64_857 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_39 ();
 sg13g2_fill_1 FILLER_65_41 ();
 sg13g2_fill_2 FILLER_65_117 ();
 sg13g2_fill_1 FILLER_65_154 ();
 sg13g2_fill_2 FILLER_65_218 ();
 sg13g2_fill_2 FILLER_65_223 ();
 sg13g2_fill_1 FILLER_65_225 ();
 sg13g2_decap_8 FILLER_65_233 ();
 sg13g2_fill_2 FILLER_65_240 ();
 sg13g2_fill_2 FILLER_65_255 ();
 sg13g2_fill_2 FILLER_65_266 ();
 sg13g2_fill_1 FILLER_65_268 ();
 sg13g2_fill_2 FILLER_65_287 ();
 sg13g2_fill_2 FILLER_65_320 ();
 sg13g2_fill_1 FILLER_65_322 ();
 sg13g2_fill_2 FILLER_65_372 ();
 sg13g2_fill_1 FILLER_65_374 ();
 sg13g2_fill_1 FILLER_65_384 ();
 sg13g2_fill_2 FILLER_65_394 ();
 sg13g2_fill_1 FILLER_65_396 ();
 sg13g2_fill_1 FILLER_65_416 ();
 sg13g2_fill_2 FILLER_65_443 ();
 sg13g2_fill_1 FILLER_65_445 ();
 sg13g2_fill_1 FILLER_65_484 ();
 sg13g2_fill_2 FILLER_65_498 ();
 sg13g2_fill_1 FILLER_65_500 ();
 sg13g2_fill_1 FILLER_65_505 ();
 sg13g2_fill_2 FILLER_65_540 ();
 sg13g2_fill_1 FILLER_65_542 ();
 sg13g2_fill_2 FILLER_65_552 ();
 sg13g2_fill_2 FILLER_65_647 ();
 sg13g2_fill_1 FILLER_65_649 ();
 sg13g2_decap_4 FILLER_65_654 ();
 sg13g2_fill_1 FILLER_65_658 ();
 sg13g2_fill_2 FILLER_65_664 ();
 sg13g2_decap_8 FILLER_65_671 ();
 sg13g2_fill_1 FILLER_65_678 ();
 sg13g2_decap_8 FILLER_65_709 ();
 sg13g2_decap_4 FILLER_65_716 ();
 sg13g2_decap_4 FILLER_65_760 ();
 sg13g2_fill_1 FILLER_65_764 ();
 sg13g2_decap_8 FILLER_65_769 ();
 sg13g2_fill_1 FILLER_65_776 ();
 sg13g2_fill_2 FILLER_65_794 ();
 sg13g2_fill_2 FILLER_65_830 ();
 sg13g2_fill_1 FILLER_66_26 ();
 sg13g2_fill_1 FILLER_66_53 ();
 sg13g2_fill_2 FILLER_66_105 ();
 sg13g2_fill_1 FILLER_66_107 ();
 sg13g2_fill_2 FILLER_66_134 ();
 sg13g2_fill_1 FILLER_66_140 ();
 sg13g2_fill_2 FILLER_66_167 ();
 sg13g2_decap_4 FILLER_66_223 ();
 sg13g2_fill_1 FILLER_66_227 ();
 sg13g2_fill_1 FILLER_66_306 ();
 sg13g2_fill_1 FILLER_66_386 ();
 sg13g2_fill_2 FILLER_66_482 ();
 sg13g2_fill_1 FILLER_66_489 ();
 sg13g2_fill_2 FILLER_66_564 ();
 sg13g2_fill_2 FILLER_66_574 ();
 sg13g2_fill_1 FILLER_66_576 ();
 sg13g2_fill_2 FILLER_66_594 ();
 sg13g2_decap_4 FILLER_66_616 ();
 sg13g2_fill_2 FILLER_66_620 ();
 sg13g2_fill_1 FILLER_66_631 ();
 sg13g2_fill_2 FILLER_66_636 ();
 sg13g2_decap_8 FILLER_66_647 ();
 sg13g2_fill_1 FILLER_66_680 ();
 sg13g2_fill_1 FILLER_66_710 ();
 sg13g2_decap_4 FILLER_66_726 ();
 sg13g2_fill_1 FILLER_66_730 ();
 sg13g2_decap_4 FILLER_66_736 ();
 sg13g2_fill_1 FILLER_66_740 ();
 sg13g2_decap_4 FILLER_66_751 ();
 sg13g2_fill_2 FILLER_66_755 ();
 sg13g2_fill_2 FILLER_66_762 ();
 sg13g2_decap_8 FILLER_66_769 ();
 sg13g2_fill_1 FILLER_66_776 ();
 sg13g2_fill_2 FILLER_66_797 ();
 sg13g2_fill_2 FILLER_66_818 ();
 sg13g2_fill_1 FILLER_66_820 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_decap_4 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_30 ();
 sg13g2_fill_2 FILLER_67_36 ();
 sg13g2_fill_1 FILLER_67_61 ();
 sg13g2_fill_1 FILLER_67_71 ();
 sg13g2_fill_1 FILLER_67_108 ();
 sg13g2_fill_1 FILLER_67_118 ();
 sg13g2_decap_4 FILLER_67_216 ();
 sg13g2_fill_2 FILLER_67_220 ();
 sg13g2_fill_2 FILLER_67_277 ();
 sg13g2_fill_1 FILLER_67_279 ();
 sg13g2_fill_2 FILLER_67_321 ();
 sg13g2_fill_2 FILLER_67_367 ();
 sg13g2_fill_1 FILLER_67_369 ();
 sg13g2_fill_1 FILLER_67_374 ();
 sg13g2_decap_8 FILLER_67_379 ();
 sg13g2_fill_2 FILLER_67_422 ();
 sg13g2_fill_2 FILLER_67_468 ();
 sg13g2_fill_1 FILLER_67_470 ();
 sg13g2_fill_2 FILLER_67_497 ();
 sg13g2_fill_1 FILLER_67_499 ();
 sg13g2_fill_2 FILLER_67_514 ();
 sg13g2_fill_1 FILLER_67_516 ();
 sg13g2_fill_1 FILLER_67_574 ();
 sg13g2_decap_8 FILLER_67_643 ();
 sg13g2_fill_2 FILLER_67_650 ();
 sg13g2_fill_1 FILLER_67_652 ();
 sg13g2_fill_2 FILLER_67_663 ();
 sg13g2_fill_1 FILLER_67_669 ();
 sg13g2_fill_2 FILLER_67_719 ();
 sg13g2_fill_1 FILLER_67_721 ();
 sg13g2_decap_4 FILLER_67_752 ();
 sg13g2_decap_4 FILLER_67_776 ();
 sg13g2_fill_1 FILLER_67_797 ();
 sg13g2_fill_2 FILLER_67_808 ();
 sg13g2_fill_1 FILLER_67_810 ();
 sg13g2_fill_2 FILLER_67_824 ();
 sg13g2_fill_1 FILLER_67_826 ();
 sg13g2_decap_4 FILLER_67_857 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_4 FILLER_68_14 ();
 sg13g2_fill_1 FILLER_68_18 ();
 sg13g2_fill_2 FILLER_68_45 ();
 sg13g2_fill_1 FILLER_68_47 ();
 sg13g2_fill_2 FILLER_68_80 ();
 sg13g2_fill_2 FILLER_68_97 ();
 sg13g2_fill_2 FILLER_68_105 ();
 sg13g2_fill_2 FILLER_68_139 ();
 sg13g2_fill_1 FILLER_68_171 ();
 sg13g2_fill_2 FILLER_68_220 ();
 sg13g2_fill_1 FILLER_68_222 ();
 sg13g2_fill_2 FILLER_68_228 ();
 sg13g2_fill_2 FILLER_68_326 ();
 sg13g2_fill_2 FILLER_68_350 ();
 sg13g2_fill_2 FILLER_68_365 ();
 sg13g2_fill_1 FILLER_68_367 ();
 sg13g2_fill_2 FILLER_68_389 ();
 sg13g2_fill_1 FILLER_68_391 ();
 sg13g2_fill_2 FILLER_68_433 ();
 sg13g2_fill_1 FILLER_68_435 ();
 sg13g2_fill_1 FILLER_68_445 ();
 sg13g2_fill_1 FILLER_68_569 ();
 sg13g2_fill_1 FILLER_68_578 ();
 sg13g2_fill_2 FILLER_68_599 ();
 sg13g2_fill_2 FILLER_68_695 ();
 sg13g2_fill_1 FILLER_68_719 ();
 sg13g2_fill_1 FILLER_68_729 ();
 sg13g2_decap_4 FILLER_68_734 ();
 sg13g2_fill_2 FILLER_68_738 ();
 sg13g2_fill_1 FILLER_68_744 ();
 sg13g2_fill_1 FILLER_68_756 ();
 sg13g2_decap_4 FILLER_68_762 ();
 sg13g2_fill_1 FILLER_68_766 ();
 sg13g2_fill_1 FILLER_68_778 ();
 sg13g2_fill_2 FILLER_68_783 ();
 sg13g2_fill_2 FILLER_68_789 ();
 sg13g2_fill_1 FILLER_68_791 ();
 sg13g2_fill_2 FILLER_68_803 ();
 sg13g2_fill_1 FILLER_68_805 ();
 sg13g2_fill_2 FILLER_68_832 ();
 sg13g2_fill_1 FILLER_68_834 ();
 sg13g2_decap_8 FILLER_68_848 ();
 sg13g2_decap_8 FILLER_68_855 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_4 FILLER_69_21 ();
 sg13g2_fill_2 FILLER_69_49 ();
 sg13g2_fill_1 FILLER_69_51 ();
 sg13g2_fill_1 FILLER_69_58 ();
 sg13g2_fill_1 FILLER_69_84 ();
 sg13g2_fill_1 FILLER_69_108 ();
 sg13g2_fill_2 FILLER_69_141 ();
 sg13g2_decap_8 FILLER_69_206 ();
 sg13g2_fill_2 FILLER_69_213 ();
 sg13g2_fill_1 FILLER_69_237 ();
 sg13g2_fill_1 FILLER_69_264 ();
 sg13g2_fill_1 FILLER_69_314 ();
 sg13g2_fill_1 FILLER_69_324 ();
 sg13g2_fill_2 FILLER_69_347 ();
 sg13g2_fill_1 FILLER_69_349 ();
 sg13g2_fill_1 FILLER_69_358 ();
 sg13g2_decap_8 FILLER_69_377 ();
 sg13g2_decap_8 FILLER_69_384 ();
 sg13g2_fill_2 FILLER_69_391 ();
 sg13g2_fill_1 FILLER_69_393 ();
 sg13g2_fill_1 FILLER_69_402 ();
 sg13g2_decap_8 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_69_415 ();
 sg13g2_fill_2 FILLER_69_422 ();
 sg13g2_fill_1 FILLER_69_424 ();
 sg13g2_fill_1 FILLER_69_451 ();
 sg13g2_fill_1 FILLER_69_544 ();
 sg13g2_fill_1 FILLER_69_582 ();
 sg13g2_fill_1 FILLER_69_603 ();
 sg13g2_decap_8 FILLER_69_657 ();
 sg13g2_fill_2 FILLER_69_664 ();
 sg13g2_fill_2 FILLER_69_670 ();
 sg13g2_fill_1 FILLER_69_672 ();
 sg13g2_decap_8 FILLER_69_689 ();
 sg13g2_fill_1 FILLER_69_722 ();
 sg13g2_fill_1 FILLER_69_737 ();
 sg13g2_fill_1 FILLER_69_759 ();
 sg13g2_fill_1 FILLER_69_799 ();
 sg13g2_fill_2 FILLER_69_804 ();
 sg13g2_decap_8 FILLER_69_845 ();
 sg13g2_decap_8 FILLER_69_852 ();
 sg13g2_fill_2 FILLER_69_859 ();
 sg13g2_fill_1 FILLER_69_861 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_4 FILLER_70_28 ();
 sg13g2_fill_2 FILLER_70_32 ();
 sg13g2_fill_1 FILLER_70_103 ();
 sg13g2_fill_1 FILLER_70_116 ();
 sg13g2_fill_2 FILLER_70_187 ();
 sg13g2_fill_2 FILLER_70_204 ();
 sg13g2_fill_2 FILLER_70_216 ();
 sg13g2_fill_2 FILLER_70_284 ();
 sg13g2_fill_1 FILLER_70_286 ();
 sg13g2_fill_2 FILLER_70_295 ();
 sg13g2_fill_1 FILLER_70_297 ();
 sg13g2_fill_2 FILLER_70_341 ();
 sg13g2_fill_2 FILLER_70_363 ();
 sg13g2_fill_1 FILLER_70_365 ();
 sg13g2_decap_4 FILLER_70_371 ();
 sg13g2_fill_1 FILLER_70_380 ();
 sg13g2_fill_2 FILLER_70_412 ();
 sg13g2_fill_1 FILLER_70_414 ();
 sg13g2_fill_1 FILLER_70_450 ();
 sg13g2_fill_1 FILLER_70_475 ();
 sg13g2_fill_2 FILLER_70_485 ();
 sg13g2_fill_1 FILLER_70_575 ();
 sg13g2_fill_2 FILLER_70_584 ();
 sg13g2_fill_2 FILLER_70_602 ();
 sg13g2_fill_1 FILLER_70_617 ();
 sg13g2_fill_1 FILLER_70_674 ();
 sg13g2_fill_1 FILLER_70_710 ();
 sg13g2_fill_1 FILLER_70_763 ();
 sg13g2_fill_2 FILLER_70_829 ();
 sg13g2_fill_1 FILLER_70_831 ();
 sg13g2_decap_8 FILLER_70_841 ();
 sg13g2_decap_8 FILLER_70_848 ();
 sg13g2_decap_8 FILLER_70_855 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_fill_2 FILLER_71_58 ();
 sg13g2_fill_1 FILLER_71_68 ();
 sg13g2_fill_2 FILLER_71_86 ();
 sg13g2_fill_1 FILLER_71_121 ();
 sg13g2_fill_1 FILLER_71_208 ();
 sg13g2_decap_8 FILLER_71_267 ();
 sg13g2_decap_4 FILLER_71_274 ();
 sg13g2_fill_1 FILLER_71_278 ();
 sg13g2_decap_4 FILLER_71_284 ();
 sg13g2_fill_2 FILLER_71_288 ();
 sg13g2_fill_1 FILLER_71_312 ();
 sg13g2_fill_2 FILLER_71_340 ();
 sg13g2_fill_1 FILLER_71_342 ();
 sg13g2_fill_1 FILLER_71_353 ();
 sg13g2_fill_2 FILLER_71_373 ();
 sg13g2_fill_2 FILLER_71_405 ();
 sg13g2_fill_1 FILLER_71_457 ();
 sg13g2_fill_1 FILLER_71_489 ();
 sg13g2_fill_1 FILLER_71_540 ();
 sg13g2_fill_2 FILLER_71_555 ();
 sg13g2_fill_1 FILLER_71_576 ();
 sg13g2_fill_2 FILLER_71_582 ();
 sg13g2_fill_2 FILLER_71_592 ();
 sg13g2_fill_1 FILLER_71_594 ();
 sg13g2_fill_2 FILLER_71_608 ();
 sg13g2_fill_1 FILLER_71_610 ();
 sg13g2_fill_1 FILLER_71_617 ();
 sg13g2_decap_4 FILLER_71_623 ();
 sg13g2_fill_2 FILLER_71_627 ();
 sg13g2_fill_1 FILLER_71_643 ();
 sg13g2_fill_2 FILLER_71_648 ();
 sg13g2_fill_1 FILLER_71_650 ();
 sg13g2_fill_1 FILLER_71_677 ();
 sg13g2_fill_1 FILLER_71_696 ();
 sg13g2_fill_2 FILLER_71_708 ();
 sg13g2_fill_1 FILLER_71_710 ();
 sg13g2_decap_4 FILLER_71_736 ();
 sg13g2_decap_8 FILLER_71_762 ();
 sg13g2_decap_8 FILLER_71_809 ();
 sg13g2_decap_8 FILLER_71_816 ();
 sg13g2_decap_8 FILLER_71_823 ();
 sg13g2_decap_8 FILLER_71_830 ();
 sg13g2_decap_8 FILLER_71_837 ();
 sg13g2_decap_8 FILLER_71_844 ();
 sg13g2_decap_8 FILLER_71_851 ();
 sg13g2_decap_4 FILLER_71_858 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_4 FILLER_72_28 ();
 sg13g2_fill_1 FILLER_72_45 ();
 sg13g2_fill_1 FILLER_72_54 ();
 sg13g2_fill_1 FILLER_72_78 ();
 sg13g2_fill_2 FILLER_72_103 ();
 sg13g2_fill_1 FILLER_72_187 ();
 sg13g2_fill_2 FILLER_72_204 ();
 sg13g2_fill_1 FILLER_72_216 ();
 sg13g2_fill_1 FILLER_72_222 ();
 sg13g2_decap_8 FILLER_72_267 ();
 sg13g2_decap_4 FILLER_72_274 ();
 sg13g2_fill_2 FILLER_72_283 ();
 sg13g2_decap_8 FILLER_72_289 ();
 sg13g2_decap_4 FILLER_72_296 ();
 sg13g2_fill_1 FILLER_72_300 ();
 sg13g2_fill_2 FILLER_72_310 ();
 sg13g2_fill_2 FILLER_72_324 ();
 sg13g2_fill_2 FILLER_72_349 ();
 sg13g2_fill_2 FILLER_72_356 ();
 sg13g2_fill_1 FILLER_72_471 ();
 sg13g2_fill_1 FILLER_72_504 ();
 sg13g2_fill_2 FILLER_72_548 ();
 sg13g2_decap_4 FILLER_72_627 ();
 sg13g2_fill_2 FILLER_72_684 ();
 sg13g2_fill_1 FILLER_72_686 ();
 sg13g2_fill_2 FILLER_72_713 ();
 sg13g2_fill_2 FILLER_72_741 ();
 sg13g2_fill_1 FILLER_72_743 ();
 sg13g2_decap_8 FILLER_72_809 ();
 sg13g2_decap_8 FILLER_72_816 ();
 sg13g2_decap_8 FILLER_72_823 ();
 sg13g2_decap_8 FILLER_72_830 ();
 sg13g2_decap_8 FILLER_72_837 ();
 sg13g2_decap_8 FILLER_72_844 ();
 sg13g2_decap_8 FILLER_72_851 ();
 sg13g2_decap_4 FILLER_72_858 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_4 FILLER_73_14 ();
 sg13g2_fill_1 FILLER_73_109 ();
 sg13g2_fill_1 FILLER_73_147 ();
 sg13g2_fill_1 FILLER_73_158 ();
 sg13g2_fill_2 FILLER_73_187 ();
 sg13g2_fill_1 FILLER_73_189 ();
 sg13g2_fill_1 FILLER_73_214 ();
 sg13g2_fill_2 FILLER_73_220 ();
 sg13g2_fill_1 FILLER_73_227 ();
 sg13g2_fill_2 FILLER_73_237 ();
 sg13g2_fill_2 FILLER_73_249 ();
 sg13g2_fill_1 FILLER_73_296 ();
 sg13g2_fill_1 FILLER_73_312 ();
 sg13g2_fill_2 FILLER_73_326 ();
 sg13g2_fill_1 FILLER_73_328 ();
 sg13g2_fill_2 FILLER_73_357 ();
 sg13g2_fill_1 FILLER_73_377 ();
 sg13g2_fill_1 FILLER_73_409 ();
 sg13g2_fill_1 FILLER_73_549 ();
 sg13g2_fill_1 FILLER_73_597 ();
 sg13g2_decap_4 FILLER_73_611 ();
 sg13g2_fill_1 FILLER_73_615 ();
 sg13g2_decap_8 FILLER_73_633 ();
 sg13g2_fill_2 FILLER_73_640 ();
 sg13g2_decap_8 FILLER_73_646 ();
 sg13g2_fill_2 FILLER_73_653 ();
 sg13g2_fill_1 FILLER_73_678 ();
 sg13g2_fill_1 FILLER_73_684 ();
 sg13g2_fill_2 FILLER_73_698 ();
 sg13g2_fill_2 FILLER_73_751 ();
 sg13g2_fill_1 FILLER_73_775 ();
 sg13g2_fill_1 FILLER_73_780 ();
 sg13g2_decap_8 FILLER_73_795 ();
 sg13g2_decap_8 FILLER_73_802 ();
 sg13g2_decap_8 FILLER_73_809 ();
 sg13g2_decap_8 FILLER_73_816 ();
 sg13g2_decap_8 FILLER_73_823 ();
 sg13g2_decap_8 FILLER_73_830 ();
 sg13g2_decap_8 FILLER_73_837 ();
 sg13g2_decap_8 FILLER_73_844 ();
 sg13g2_decap_8 FILLER_73_851 ();
 sg13g2_decap_4 FILLER_73_858 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_4 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_51 ();
 sg13g2_fill_1 FILLER_74_75 ();
 sg13g2_fill_2 FILLER_74_81 ();
 sg13g2_fill_2 FILLER_74_168 ();
 sg13g2_fill_1 FILLER_74_170 ();
 sg13g2_fill_2 FILLER_74_286 ();
 sg13g2_fill_1 FILLER_74_288 ();
 sg13g2_fill_2 FILLER_74_297 ();
 sg13g2_fill_1 FILLER_74_330 ();
 sg13g2_fill_1 FILLER_74_348 ();
 sg13g2_fill_1 FILLER_74_368 ();
 sg13g2_fill_2 FILLER_74_382 ();
 sg13g2_fill_1 FILLER_74_394 ();
 sg13g2_fill_2 FILLER_74_421 ();
 sg13g2_fill_1 FILLER_74_463 ();
 sg13g2_fill_1 FILLER_74_494 ();
 sg13g2_decap_4 FILLER_74_600 ();
 sg13g2_fill_2 FILLER_74_604 ();
 sg13g2_fill_2 FILLER_74_623 ();
 sg13g2_fill_2 FILLER_74_652 ();
 sg13g2_fill_1 FILLER_74_654 ();
 sg13g2_fill_2 FILLER_74_681 ();
 sg13g2_fill_1 FILLER_74_683 ();
 sg13g2_fill_2 FILLER_74_739 ();
 sg13g2_fill_1 FILLER_74_741 ();
 sg13g2_fill_1 FILLER_74_752 ();
 sg13g2_decap_8 FILLER_74_779 ();
 sg13g2_decap_8 FILLER_74_786 ();
 sg13g2_decap_8 FILLER_74_793 ();
 sg13g2_decap_8 FILLER_74_800 ();
 sg13g2_decap_8 FILLER_74_807 ();
 sg13g2_decap_8 FILLER_74_814 ();
 sg13g2_decap_8 FILLER_74_821 ();
 sg13g2_decap_8 FILLER_74_828 ();
 sg13g2_decap_8 FILLER_74_835 ();
 sg13g2_decap_8 FILLER_74_842 ();
 sg13g2_decap_8 FILLER_74_849 ();
 sg13g2_decap_4 FILLER_74_856 ();
 sg13g2_fill_2 FILLER_74_860 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_4 FILLER_75_42 ();
 sg13g2_fill_1 FILLER_75_46 ();
 sg13g2_fill_2 FILLER_75_99 ();
 sg13g2_fill_2 FILLER_75_119 ();
 sg13g2_fill_1 FILLER_75_152 ();
 sg13g2_fill_2 FILLER_75_180 ();
 sg13g2_fill_1 FILLER_75_187 ();
 sg13g2_fill_1 FILLER_75_211 ();
 sg13g2_fill_2 FILLER_75_242 ();
 sg13g2_fill_1 FILLER_75_244 ();
 sg13g2_fill_2 FILLER_75_285 ();
 sg13g2_fill_1 FILLER_75_287 ();
 sg13g2_fill_2 FILLER_75_302 ();
 sg13g2_fill_2 FILLER_75_313 ();
 sg13g2_decap_8 FILLER_75_322 ();
 sg13g2_fill_2 FILLER_75_384 ();
 sg13g2_fill_1 FILLER_75_421 ();
 sg13g2_fill_2 FILLER_75_445 ();
 sg13g2_fill_2 FILLER_75_466 ();
 sg13g2_fill_1 FILLER_75_494 ();
 sg13g2_fill_1 FILLER_75_509 ();
 sg13g2_fill_1 FILLER_75_519 ();
 sg13g2_fill_2 FILLER_75_567 ();
 sg13g2_fill_2 FILLER_75_594 ();
 sg13g2_fill_2 FILLER_75_632 ();
 sg13g2_fill_2 FILLER_75_639 ();
 sg13g2_decap_8 FILLER_75_646 ();
 sg13g2_decap_4 FILLER_75_653 ();
 sg13g2_fill_2 FILLER_75_657 ();
 sg13g2_fill_1 FILLER_75_667 ();
 sg13g2_fill_2 FILLER_75_682 ();
 sg13g2_fill_1 FILLER_75_684 ();
 sg13g2_fill_2 FILLER_75_693 ();
 sg13g2_fill_1 FILLER_75_706 ();
 sg13g2_fill_1 FILLER_75_747 ();
 sg13g2_decap_8 FILLER_75_774 ();
 sg13g2_decap_8 FILLER_75_781 ();
 sg13g2_decap_8 FILLER_75_788 ();
 sg13g2_decap_8 FILLER_75_795 ();
 sg13g2_decap_8 FILLER_75_802 ();
 sg13g2_decap_8 FILLER_75_809 ();
 sg13g2_decap_8 FILLER_75_816 ();
 sg13g2_decap_8 FILLER_75_823 ();
 sg13g2_decap_8 FILLER_75_830 ();
 sg13g2_decap_8 FILLER_75_837 ();
 sg13g2_decap_8 FILLER_75_844 ();
 sg13g2_decap_8 FILLER_75_851 ();
 sg13g2_decap_4 FILLER_75_858 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_4 FILLER_76_56 ();
 sg13g2_fill_1 FILLER_76_60 ();
 sg13g2_decap_4 FILLER_76_65 ();
 sg13g2_fill_1 FILLER_76_69 ();
 sg13g2_fill_2 FILLER_76_84 ();
 sg13g2_fill_2 FILLER_76_164 ();
 sg13g2_fill_2 FILLER_76_200 ();
 sg13g2_fill_1 FILLER_76_210 ();
 sg13g2_fill_2 FILLER_76_279 ();
 sg13g2_fill_1 FILLER_76_311 ();
 sg13g2_decap_4 FILLER_76_338 ();
 sg13g2_fill_1 FILLER_76_342 ();
 sg13g2_fill_1 FILLER_76_356 ();
 sg13g2_fill_1 FILLER_76_484 ();
 sg13g2_fill_2 FILLER_76_587 ();
 sg13g2_fill_2 FILLER_76_607 ();
 sg13g2_fill_1 FILLER_76_609 ();
 sg13g2_fill_2 FILLER_76_634 ();
 sg13g2_fill_1 FILLER_76_636 ();
 sg13g2_fill_2 FILLER_76_644 ();
 sg13g2_fill_2 FILLER_76_684 ();
 sg13g2_decap_4 FILLER_76_699 ();
 sg13g2_fill_1 FILLER_76_703 ();
 sg13g2_decap_4 FILLER_76_709 ();
 sg13g2_fill_2 FILLER_76_731 ();
 sg13g2_fill_2 FILLER_76_746 ();
 sg13g2_fill_2 FILLER_76_757 ();
 sg13g2_decap_8 FILLER_76_763 ();
 sg13g2_decap_8 FILLER_76_770 ();
 sg13g2_decap_8 FILLER_76_777 ();
 sg13g2_decap_8 FILLER_76_784 ();
 sg13g2_decap_8 FILLER_76_791 ();
 sg13g2_decap_8 FILLER_76_798 ();
 sg13g2_decap_8 FILLER_76_805 ();
 sg13g2_decap_8 FILLER_76_812 ();
 sg13g2_decap_8 FILLER_76_819 ();
 sg13g2_decap_8 FILLER_76_826 ();
 sg13g2_decap_8 FILLER_76_833 ();
 sg13g2_decap_8 FILLER_76_840 ();
 sg13g2_decap_8 FILLER_76_847 ();
 sg13g2_decap_8 FILLER_76_854 ();
 sg13g2_fill_1 FILLER_76_861 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_4 FILLER_77_77 ();
 sg13g2_fill_2 FILLER_77_102 ();
 sg13g2_fill_1 FILLER_77_104 ();
 sg13g2_fill_1 FILLER_77_143 ();
 sg13g2_fill_2 FILLER_77_294 ();
 sg13g2_fill_1 FILLER_77_368 ();
 sg13g2_fill_2 FILLER_77_379 ();
 sg13g2_fill_1 FILLER_77_463 ();
 sg13g2_fill_1 FILLER_77_561 ();
 sg13g2_fill_2 FILLER_77_620 ();
 sg13g2_fill_1 FILLER_77_640 ();
 sg13g2_fill_2 FILLER_77_645 ();
 sg13g2_fill_1 FILLER_77_647 ();
 sg13g2_fill_2 FILLER_77_656 ();
 sg13g2_fill_1 FILLER_77_702 ();
 sg13g2_decap_8 FILLER_77_771 ();
 sg13g2_decap_8 FILLER_77_778 ();
 sg13g2_decap_8 FILLER_77_785 ();
 sg13g2_decap_8 FILLER_77_792 ();
 sg13g2_decap_8 FILLER_77_799 ();
 sg13g2_decap_8 FILLER_77_806 ();
 sg13g2_decap_8 FILLER_77_813 ();
 sg13g2_decap_8 FILLER_77_820 ();
 sg13g2_decap_8 FILLER_77_827 ();
 sg13g2_decap_8 FILLER_77_834 ();
 sg13g2_decap_8 FILLER_77_841 ();
 sg13g2_decap_8 FILLER_77_848 ();
 sg13g2_decap_8 FILLER_77_855 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_fill_2 FILLER_78_70 ();
 sg13g2_fill_1 FILLER_78_119 ();
 sg13g2_fill_2 FILLER_78_217 ();
 sg13g2_fill_1 FILLER_78_233 ();
 sg13g2_fill_2 FILLER_78_244 ();
 sg13g2_fill_1 FILLER_78_341 ();
 sg13g2_fill_2 FILLER_78_395 ();
 sg13g2_fill_2 FILLER_78_426 ();
 sg13g2_fill_1 FILLER_78_473 ();
 sg13g2_fill_2 FILLER_78_510 ();
 sg13g2_fill_1 FILLER_78_557 ();
 sg13g2_fill_1 FILLER_78_571 ();
 sg13g2_fill_1 FILLER_78_585 ();
 sg13g2_fill_2 FILLER_78_595 ();
 sg13g2_fill_1 FILLER_78_597 ();
 sg13g2_fill_1 FILLER_78_640 ();
 sg13g2_fill_1 FILLER_78_655 ();
 sg13g2_fill_1 FILLER_78_672 ();
 sg13g2_fill_2 FILLER_78_682 ();
 sg13g2_decap_4 FILLER_78_710 ();
 sg13g2_decap_8 FILLER_78_762 ();
 sg13g2_decap_8 FILLER_78_769 ();
 sg13g2_decap_8 FILLER_78_776 ();
 sg13g2_decap_8 FILLER_78_783 ();
 sg13g2_decap_8 FILLER_78_790 ();
 sg13g2_decap_8 FILLER_78_797 ();
 sg13g2_decap_8 FILLER_78_804 ();
 sg13g2_decap_8 FILLER_78_811 ();
 sg13g2_decap_8 FILLER_78_818 ();
 sg13g2_decap_8 FILLER_78_825 ();
 sg13g2_decap_8 FILLER_78_832 ();
 sg13g2_decap_8 FILLER_78_839 ();
 sg13g2_decap_8 FILLER_78_846 ();
 sg13g2_decap_8 FILLER_78_853 ();
 sg13g2_fill_2 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_fill_2 FILLER_79_56 ();
 sg13g2_fill_2 FILLER_79_124 ();
 sg13g2_fill_1 FILLER_79_135 ();
 sg13g2_fill_2 FILLER_79_150 ();
 sg13g2_fill_1 FILLER_79_189 ();
 sg13g2_fill_2 FILLER_79_216 ();
 sg13g2_fill_2 FILLER_79_305 ();
 sg13g2_fill_1 FILLER_79_307 ();
 sg13g2_fill_1 FILLER_79_349 ();
 sg13g2_fill_2 FILLER_79_414 ();
 sg13g2_fill_2 FILLER_79_500 ();
 sg13g2_fill_1 FILLER_79_502 ();
 sg13g2_decap_8 FILLER_79_584 ();
 sg13g2_decap_4 FILLER_79_591 ();
 sg13g2_fill_1 FILLER_79_595 ();
 sg13g2_fill_1 FILLER_79_600 ();
 sg13g2_fill_1 FILLER_79_609 ();
 sg13g2_fill_1 FILLER_79_615 ();
 sg13g2_fill_2 FILLER_79_632 ();
 sg13g2_fill_2 FILLER_79_647 ();
 sg13g2_fill_1 FILLER_79_649 ();
 sg13g2_fill_2 FILLER_79_656 ();
 sg13g2_fill_2 FILLER_79_691 ();
 sg13g2_fill_1 FILLER_79_693 ();
 sg13g2_decap_8 FILLER_79_698 ();
 sg13g2_decap_8 FILLER_79_705 ();
 sg13g2_decap_8 FILLER_79_712 ();
 sg13g2_decap_4 FILLER_79_719 ();
 sg13g2_fill_2 FILLER_79_723 ();
 sg13g2_decap_8 FILLER_79_733 ();
 sg13g2_decap_8 FILLER_79_740 ();
 sg13g2_decap_8 FILLER_79_747 ();
 sg13g2_decap_8 FILLER_79_754 ();
 sg13g2_decap_8 FILLER_79_761 ();
 sg13g2_decap_8 FILLER_79_768 ();
 sg13g2_decap_8 FILLER_79_775 ();
 sg13g2_decap_8 FILLER_79_782 ();
 sg13g2_decap_8 FILLER_79_789 ();
 sg13g2_decap_8 FILLER_79_796 ();
 sg13g2_decap_8 FILLER_79_803 ();
 sg13g2_decap_8 FILLER_79_810 ();
 sg13g2_decap_8 FILLER_79_817 ();
 sg13g2_decap_8 FILLER_79_824 ();
 sg13g2_decap_8 FILLER_79_831 ();
 sg13g2_decap_8 FILLER_79_838 ();
 sg13g2_decap_8 FILLER_79_845 ();
 sg13g2_decap_8 FILLER_79_852 ();
 sg13g2_fill_2 FILLER_79_859 ();
 sg13g2_fill_1 FILLER_79_861 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_fill_2 FILLER_80_98 ();
 sg13g2_fill_1 FILLER_80_126 ();
 sg13g2_fill_1 FILLER_80_153 ();
 sg13g2_fill_2 FILLER_80_210 ();
 sg13g2_fill_1 FILLER_80_232 ();
 sg13g2_fill_1 FILLER_80_276 ();
 sg13g2_fill_2 FILLER_80_313 ();
 sg13g2_fill_1 FILLER_80_315 ();
 sg13g2_fill_1 FILLER_80_410 ();
 sg13g2_fill_1 FILLER_80_420 ();
 sg13g2_fill_1 FILLER_80_506 ();
 sg13g2_fill_2 FILLER_80_541 ();
 sg13g2_fill_1 FILLER_80_543 ();
 sg13g2_fill_2 FILLER_80_583 ();
 sg13g2_fill_1 FILLER_80_611 ();
 sg13g2_fill_2 FILLER_80_651 ();
 sg13g2_fill_1 FILLER_80_653 ();
 sg13g2_decap_4 FILLER_80_658 ();
 sg13g2_fill_2 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_694 ();
 sg13g2_decap_8 FILLER_80_701 ();
 sg13g2_decap_8 FILLER_80_708 ();
 sg13g2_decap_8 FILLER_80_715 ();
 sg13g2_decap_8 FILLER_80_722 ();
 sg13g2_decap_8 FILLER_80_729 ();
 sg13g2_decap_8 FILLER_80_736 ();
 sg13g2_decap_8 FILLER_80_743 ();
 sg13g2_decap_8 FILLER_80_750 ();
 sg13g2_decap_8 FILLER_80_757 ();
 sg13g2_decap_8 FILLER_80_764 ();
 sg13g2_decap_8 FILLER_80_771 ();
 sg13g2_decap_8 FILLER_80_778 ();
 sg13g2_decap_8 FILLER_80_785 ();
 sg13g2_decap_8 FILLER_80_792 ();
 sg13g2_decap_8 FILLER_80_799 ();
 sg13g2_decap_8 FILLER_80_806 ();
 sg13g2_decap_8 FILLER_80_813 ();
 sg13g2_decap_8 FILLER_80_820 ();
 sg13g2_decap_8 FILLER_80_827 ();
 sg13g2_decap_8 FILLER_80_834 ();
 sg13g2_decap_8 FILLER_80_841 ();
 sg13g2_decap_8 FILLER_80_848 ();
 sg13g2_decap_8 FILLER_80_855 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
 assign uo_out[1] = net20;
 assign uo_out[2] = net21;
 assign uo_out[3] = net22;
 assign uo_out[4] = net23;
 assign uo_out[5] = net24;
 assign uo_out[6] = net25;
 assign uo_out[7] = net26;
endmodule

module tt_um_pid_controller (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire clknet_0_clk;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire \pid.Kd[0] ;
 wire \pid.Kd[1] ;
 wire \pid.Kd[2] ;
 wire \pid.Kd[3] ;
 wire \pid.Kd[4] ;
 wire \pid.Kd[5] ;
 wire \pid.Kd[6] ;
 wire \pid.Kd[7] ;
 wire \pid.Kd[8] ;
 wire \pid.Ki[0] ;
 wire \pid.Ki[1] ;
 wire \pid.Ki[2] ;
 wire \pid.Ki[3] ;
 wire \pid.Ki[4] ;
 wire \pid.Ki[5] ;
 wire \pid.Ki[6] ;
 wire \pid.Ki[7] ;
 wire \pid.Ki[8] ;
 wire \pid.Kp[0] ;
 wire \pid.Kp[1] ;
 wire \pid.Kp[2] ;
 wire \pid.Kp[3] ;
 wire \pid.Kp[4] ;
 wire \pid.Kp[5] ;
 wire \pid.Kp[6] ;
 wire \pid.Kp[7] ;
 wire \pid.Kp[8] ;
 wire \pid.integral[0] ;
 wire \pid.integral[10] ;
 wire \pid.integral[11] ;
 wire \pid.integral[12] ;
 wire \pid.integral[13] ;
 wire \pid.integral[14] ;
 wire \pid.integral[15] ;
 wire \pid.integral[1] ;
 wire \pid.integral[2] ;
 wire \pid.integral[3] ;
 wire \pid.integral[4] ;
 wire \pid.integral[5] ;
 wire \pid.integral[6] ;
 wire \pid.integral[7] ;
 wire \pid.integral[8] ;
 wire \pid.integral[9] ;
 wire \pid.prev_error[0] ;
 wire \pid.prev_error[1] ;
 wire \pid.prev_error[2] ;
 wire \pid.prev_error[3] ;
 wire \pid.prev_error[4] ;
 wire \pid.prev_error[5] ;
 wire \pid.prev_error[6] ;
 wire \pid.prev_error[7] ;
 wire \pid.prev_error[8] ;
 wire \pid.state[0] ;
 wire \pid.state[1] ;
 wire \pid.state[2] ;
 wire \pid.state[3] ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;

 sg13g2_inv_1 _2764_ (.Y(_0821_),
    .A(net4));
 sg13g2_inv_1 _2765_ (.Y(_0832_),
    .A(net461));
 sg13g2_inv_1 _2766_ (.Y(_0843_),
    .A(net135));
 sg13g2_inv_1 _2767_ (.Y(_0854_),
    .A(net434));
 sg13g2_inv_1 _2768_ (.Y(_0865_),
    .A(_0024_));
 sg13g2_inv_1 _2769_ (.Y(_0876_),
    .A(_0002_));
 sg13g2_inv_2 _2770_ (.Y(_0887_),
    .A(net444));
 sg13g2_inv_2 _2771_ (.Y(_0898_),
    .A(_0003_));
 sg13g2_inv_1 _2772_ (.Y(_0909_),
    .A(net446));
 sg13g2_inv_1 _2773_ (.Y(_0920_),
    .A(_0004_));
 sg13g2_inv_1 _2774_ (.Y(_0931_),
    .A(_0005_));
 sg13g2_inv_1 _2775_ (.Y(_0942_),
    .A(\pid.integral[14] ));
 sg13g2_inv_1 _2776_ (.Y(_0953_),
    .A(_0012_));
 sg13g2_or2_1 _2777_ (.X(_0000_),
    .B(net123),
    .A(net451));
 sg13g2_nor2_1 _2778_ (.A(net456),
    .B(net470),
    .Y(_0974_));
 sg13g2_and2_1 _2779_ (.A(net4),
    .B(net475),
    .X(_0985_));
 sg13g2_nand2_1 _2780_ (.Y(_0996_),
    .A(net4),
    .B(net474));
 sg13g2_nand3b_1 _2781_ (.B(_0996_),
    .C(net1),
    .Y(_1007_),
    .A_N(_0985_));
 sg13g2_a21oi_1 _2782_ (.A1(net456),
    .A2(_1007_),
    .Y(_0031_),
    .B1(_0974_));
 sg13g2_nor2b_1 _2783_ (.A(net1),
    .B_N(net475),
    .Y(_1028_));
 sg13g2_a21oi_1 _2784_ (.A1(net4),
    .A2(net474),
    .Y(_1039_),
    .B1(net475));
 sg13g2_a21o_2 _2785_ (.A2(_0985_),
    .A1(net1),
    .B1(_1039_),
    .X(_1050_));
 sg13g2_nor2_1 _2786_ (.A(net456),
    .B(net468),
    .Y(_1061_));
 sg13g2_a21oi_1 _2787_ (.A1(net456),
    .A2(_1050_),
    .Y(_0032_),
    .B1(_1061_));
 sg13g2_nor2_1 _2788_ (.A(net456),
    .B(net466),
    .Y(_1082_));
 sg13g2_or2_1 _2789_ (.X(_1093_),
    .B(net474),
    .A(net1));
 sg13g2_nand2_1 _2790_ (.Y(_1104_),
    .A(net1),
    .B(net474));
 sg13g2_o21ai_1 _2791_ (.B1(_1093_),
    .Y(_1115_),
    .A1(_0985_),
    .A2(_1104_));
 sg13g2_a21oi_1 _2792_ (.A1(net456),
    .A2(_1115_),
    .Y(_0033_),
    .B1(_1082_));
 sg13g2_nor2_1 _2793_ (.A(net456),
    .B(net138),
    .Y(_1136_));
 sg13g2_or2_1 _2794_ (.X(_1147_),
    .B(net474),
    .A(net4));
 sg13g2_o21ai_1 _2795_ (.B1(_1104_),
    .Y(_1158_),
    .A1(_0821_),
    .A2(net474));
 sg13g2_xnor2_1 _2796_ (.Y(_1169_),
    .A(net475),
    .B(_1158_));
 sg13g2_a21oi_1 _2797_ (.A1(net456),
    .A2(_1169_),
    .Y(_0034_),
    .B1(_1136_));
 sg13g2_nand2_1 _2798_ (.Y(_1190_),
    .A(_0821_),
    .B(net475));
 sg13g2_a22oi_1 _2799_ (.Y(_1201_),
    .B1(_1190_),
    .B2(net474),
    .A2(_1147_),
    .A1(_1028_));
 sg13g2_nor2_1 _2800_ (.A(net457),
    .B(net465),
    .Y(_1212_));
 sg13g2_a21oi_1 _2801_ (.A1(net457),
    .A2(_1201_),
    .Y(_0035_),
    .B1(_1212_));
 sg13g2_nor2_1 _2802_ (.A(net455),
    .B(net464),
    .Y(_1233_));
 sg13g2_o21ai_1 _2803_ (.B1(_1158_),
    .Y(_1244_),
    .A1(net4),
    .A2(net475));
 sg13g2_a21oi_1 _2804_ (.A1(net455),
    .A2(_1244_),
    .Y(_0036_),
    .B1(_1233_));
 sg13g2_nor2_1 _2805_ (.A(net455),
    .B(net463),
    .Y(_1265_));
 sg13g2_nand2b_1 _2806_ (.Y(_1276_),
    .B(_1104_),
    .A_N(net475));
 sg13g2_nand3_1 _2807_ (.B(_1093_),
    .C(_1276_),
    .A(net4),
    .Y(_1287_));
 sg13g2_a21oi_1 _2808_ (.A1(net455),
    .A2(_1287_),
    .Y(_0037_),
    .B1(_1265_));
 sg13g2_nor2_1 _2809_ (.A(net455),
    .B(net462),
    .Y(_1308_));
 sg13g2_or2_2 _2810_ (.X(_1319_),
    .B(_1028_),
    .A(_0996_));
 sg13g2_a21oi_1 _2811_ (.A1(net455),
    .A2(_1319_),
    .Y(_0038_),
    .B1(_1308_));
 sg13g2_nor2_1 _2812_ (.A(net455),
    .B(net461),
    .Y(_1340_));
 sg13g2_nand2_2 _2813_ (.Y(_1351_),
    .A(net474),
    .B(_0985_));
 sg13g2_a21oi_1 _2814_ (.A1(net455),
    .A2(_1351_),
    .Y(_0039_),
    .B1(_1340_));
 sg13g2_nor2_1 _2815_ (.A(net454),
    .B(net142),
    .Y(_1372_));
 sg13g2_a21oi_1 _2816_ (.A1(net453),
    .A2(_1007_),
    .Y(_0040_),
    .B1(_1372_));
 sg13g2_nor2_1 _2817_ (.A(net453),
    .B(net98),
    .Y(_1393_));
 sg13g2_a21oi_1 _2818_ (.A1(net453),
    .A2(_1050_),
    .Y(_0041_),
    .B1(_1393_));
 sg13g2_nor2_1 _2819_ (.A(net453),
    .B(net157),
    .Y(_1414_));
 sg13g2_a21oi_1 _2820_ (.A1(net453),
    .A2(_1115_),
    .Y(_0042_),
    .B1(_1414_));
 sg13g2_nor2_1 _2821_ (.A(net454),
    .B(net146),
    .Y(_1435_));
 sg13g2_a21oi_1 _2822_ (.A1(net453),
    .A2(_1169_),
    .Y(_0043_),
    .B1(_1435_));
 sg13g2_nor2_1 _2823_ (.A(net452),
    .B(net153),
    .Y(_1456_));
 sg13g2_a21oi_1 _2824_ (.A1(net452),
    .A2(_1201_),
    .Y(_0044_),
    .B1(_1456_));
 sg13g2_nor2_1 _2825_ (.A(net454),
    .B(\pid.Ki[5] ),
    .Y(_1477_));
 sg13g2_a21oi_1 _2826_ (.A1(net454),
    .A2(_1244_),
    .Y(_0045_),
    .B1(_1477_));
 sg13g2_nor2_1 _2827_ (.A(net452),
    .B(net155),
    .Y(_1498_));
 sg13g2_a21oi_1 _2828_ (.A1(net452),
    .A2(_1287_),
    .Y(_0046_),
    .B1(_1498_));
 sg13g2_nor2_1 _2829_ (.A(net452),
    .B(net158),
    .Y(_1519_));
 sg13g2_a21oi_1 _2830_ (.A1(net452),
    .A2(_1319_),
    .Y(_0047_),
    .B1(_1519_));
 sg13g2_nor2_1 _2831_ (.A(net452),
    .B(net149),
    .Y(_1540_));
 sg13g2_a21oi_1 _2832_ (.A1(net452),
    .A2(_1351_),
    .Y(_0048_),
    .B1(_1540_));
 sg13g2_nor3_1 _2833_ (.A(net457),
    .B(\pid.state[0] ),
    .C(net453),
    .Y(_1561_));
 sg13g2_nor2_1 _2834_ (.A(net134),
    .B(net426),
    .Y(_1572_));
 sg13g2_nand2b_1 _2835_ (.Y(_1583_),
    .B(net9),
    .A_N(net1));
 sg13g2_xnor2_1 _2836_ (.Y(_1594_),
    .A(net9),
    .B(net1));
 sg13g2_xor2_1 _2837_ (.B(net1),
    .A(net9),
    .X(_1605_));
 sg13g2_a21oi_1 _2838_ (.A1(net426),
    .A2(net471),
    .Y(_0049_),
    .B1(_1572_));
 sg13g2_nor2_1 _2839_ (.A(net110),
    .B(net426),
    .Y(_1626_));
 sg13g2_nor2b_1 _2840_ (.A(net10),
    .B_N(net2),
    .Y(_1637_));
 sg13g2_xnor2_1 _2841_ (.Y(_1648_),
    .A(net10),
    .B(net475));
 sg13g2_xor2_1 _2842_ (.B(net83),
    .A(_1583_),
    .X(_1659_));
 sg13g2_inv_1 _2843_ (.Y(_1670_),
    .A(net422));
 sg13g2_a21oi_1 _2844_ (.A1(net426),
    .A2(_1670_),
    .Y(_0050_),
    .B1(_1626_));
 sg13g2_nor2_1 _2845_ (.A(net119),
    .B(net426),
    .Y(_1691_));
 sg13g2_a21oi_2 _2846_ (.B1(_1637_),
    .Y(_1702_),
    .A2(_1583_),
    .A1(_1648_));
 sg13g2_nand2b_1 _2847_ (.Y(_1713_),
    .B(net3),
    .A_N(net11));
 sg13g2_xnor2_1 _2848_ (.Y(_1724_),
    .A(net11),
    .B(net3));
 sg13g2_inv_1 _2849_ (.Y(_1735_),
    .A(_1724_));
 sg13g2_xnor2_1 _2850_ (.Y(_1746_),
    .A(_1702_),
    .B(_1724_));
 sg13g2_xnor2_1 _2851_ (.Y(_1757_),
    .A(_1702_),
    .B(_1735_));
 sg13g2_a21oi_1 _2852_ (.A1(net430),
    .A2(net417),
    .Y(_0051_),
    .B1(_1691_));
 sg13g2_nand2b_1 _2853_ (.Y(_1778_),
    .B(net4),
    .A_N(net12));
 sg13g2_nand2_2 _2854_ (.Y(_1789_),
    .A(net12),
    .B(_0821_));
 sg13g2_nand2_1 _2855_ (.Y(_1800_),
    .A(_1778_),
    .B(_1789_));
 sg13g2_o21ai_1 _2856_ (.B1(_1713_),
    .Y(_1811_),
    .A1(_1702_),
    .A2(_1735_));
 sg13g2_xnor2_1 _2857_ (.Y(_1822_),
    .A(_1800_),
    .B(_1811_));
 sg13g2_mux2_1 _2858_ (.A0(net126),
    .A1(net414),
    .S(net426),
    .X(_0052_));
 sg13g2_nor2b_1 _2859_ (.A(net13),
    .B_N(net5),
    .Y(_1843_));
 sg13g2_xnor2_1 _2860_ (.Y(_1854_),
    .A(net13),
    .B(net5));
 sg13g2_and2_1 _2861_ (.A(_1713_),
    .B(_1778_),
    .X(_1865_));
 sg13g2_o21ai_1 _2862_ (.B1(_1865_),
    .Y(_1876_),
    .A1(_1735_),
    .A2(_1702_));
 sg13g2_and2_1 _2863_ (.A(_1789_),
    .B(net36),
    .X(_1887_));
 sg13g2_and3_2 _2864_ (.X(_1898_),
    .A(_1789_),
    .B(_1854_),
    .C(net37));
 sg13g2_nand3_1 _2865_ (.B(_1854_),
    .C(_1789_),
    .A(net67),
    .Y(_1909_));
 sg13g2_a21oi_2 _2866_ (.B1(_1854_),
    .Y(_1920_),
    .A2(net38),
    .A1(_1789_));
 sg13g2_nor2_1 _2867_ (.A(_1898_),
    .B(_1920_),
    .Y(_1931_));
 sg13g2_mux2_1 _2868_ (.A0(net111),
    .A1(net408),
    .S(net426),
    .X(_0053_));
 sg13g2_nor2b_1 _2869_ (.A(net14),
    .B_N(net6),
    .Y(_1952_));
 sg13g2_xnor2_1 _2870_ (.Y(_1963_),
    .A(net14),
    .B(net6));
 sg13g2_nor2_1 _2871_ (.A(_1843_),
    .B(_1963_),
    .Y(_1974_));
 sg13g2_and2_1 _2872_ (.A(_1843_),
    .B(_1963_),
    .X(_1985_));
 sg13g2_and2_1 _2873_ (.A(_1854_),
    .B(_1963_),
    .X(_1993_));
 sg13g2_and3_1 _2874_ (.X(_2001_),
    .A(net66),
    .B(_1789_),
    .C(_1993_));
 sg13g2_a21oi_1 _2875_ (.A1(net46),
    .A2(_1974_),
    .Y(_2007_),
    .B1(net50));
 sg13g2_nand2b_2 _2876_ (.Y(_2013_),
    .B(_2007_),
    .A_N(_1985_));
 sg13g2_a221oi_1 _2877_ (.B2(_1887_),
    .C1(_1985_),
    .B1(_1993_),
    .A1(_1974_),
    .Y(_2016_),
    .A2(_1909_));
 sg13g2_nand2_1 _2878_ (.Y(_2020_),
    .A(net425),
    .B(net404));
 sg13g2_o21ai_1 _2879_ (.B1(_2020_),
    .Y(_0054_),
    .A1(_0843_),
    .A2(net425));
 sg13g2_nand2b_1 _2880_ (.Y(_2021_),
    .B(net7),
    .A_N(net15));
 sg13g2_xnor2_1 _2881_ (.Y(_2022_),
    .A(net15),
    .B(net7));
 sg13g2_or2_1 _2882_ (.X(_2023_),
    .B(_1985_),
    .A(_1952_));
 sg13g2_or2_1 _2883_ (.X(_2024_),
    .B(_2023_),
    .A(net82));
 sg13g2_o21ai_1 _2884_ (.B1(_2022_),
    .Y(_2025_),
    .A1(_2023_),
    .A2(_2001_));
 sg13g2_xor2_1 _2885_ (.B(_2024_),
    .A(_2022_),
    .X(_2026_));
 sg13g2_xnor2_1 _2886_ (.Y(_2027_),
    .A(_2022_),
    .B(_2024_));
 sg13g2_nor2_1 _2887_ (.A(net122),
    .B(net425),
    .Y(_2028_));
 sg13g2_a21oi_1 _2888_ (.A1(net425),
    .A2(_2027_),
    .Y(_0055_),
    .B1(_2028_));
 sg13g2_nor2_1 _2889_ (.A(net95),
    .B(net425),
    .Y(_2029_));
 sg13g2_nor2b_2 _2890_ (.A(net16),
    .B_N(net8),
    .Y(_2030_));
 sg13g2_xor2_1 _2891_ (.B(net16),
    .A(net8),
    .X(_2031_));
 sg13g2_a21oi_2 _2892_ (.B1(_2031_),
    .Y(_2032_),
    .A2(_2025_),
    .A1(_2021_));
 sg13g2_a21o_2 _2893_ (.A2(_2021_),
    .A1(net80),
    .B1(_2031_),
    .X(_2033_));
 sg13g2_nand3_1 _2894_ (.B(_2021_),
    .C(_2031_),
    .A(net69),
    .Y(_2034_));
 sg13g2_and2_1 _2895_ (.A(_2033_),
    .B(_2034_),
    .X(_2035_));
 sg13g2_nand2_2 _2896_ (.Y(_2036_),
    .A(net62),
    .B(net54));
 sg13g2_a21oi_1 _2897_ (.A1(net425),
    .A2(_2036_),
    .Y(_0056_),
    .B1(_2029_));
 sg13g2_nor2_1 _2898_ (.A(_2030_),
    .B(_2032_),
    .Y(_2037_));
 sg13g2_nand2b_2 _2899_ (.Y(_2038_),
    .B(net60),
    .A_N(_2030_));
 sg13g2_nor2_1 _2900_ (.A(net100),
    .B(net425),
    .Y(_2039_));
 sg13g2_a21oi_1 _2901_ (.A1(net425),
    .A2(_2038_),
    .Y(_0057_),
    .B1(_2039_));
 sg13g2_nand2b_1 _2902_ (.Y(_2040_),
    .B(net101),
    .A_N(\pid.state[3] ));
 sg13g2_nand2b_1 _2903_ (.Y(_2041_),
    .B(net414),
    .A_N(\pid.prev_error[3] ));
 sg13g2_nor2_1 _2904_ (.A(\pid.prev_error[2] ),
    .B(net417),
    .Y(_2042_));
 sg13g2_nor2b_1 _2905_ (.A(\pid.prev_error[1] ),
    .B_N(net422),
    .Y(_2043_));
 sg13g2_nand2_1 _2906_ (.Y(_2044_),
    .A(\pid.prev_error[0] ),
    .B(net471));
 sg13g2_xnor2_1 _2907_ (.Y(_2045_),
    .A(\pid.prev_error[1] ),
    .B(net422));
 sg13g2_a21o_1 _2908_ (.A2(_2045_),
    .A1(_2044_),
    .B1(_2043_),
    .X(_2046_));
 sg13g2_xnor2_1 _2909_ (.Y(_2047_),
    .A(\pid.prev_error[2] ),
    .B(net419));
 sg13g2_a21oi_2 _2910_ (.B1(_2042_),
    .Y(_2048_),
    .A2(_2047_),
    .A1(_2046_));
 sg13g2_nor2b_1 _2911_ (.A(net414),
    .B_N(\pid.prev_error[3] ),
    .Y(_2049_));
 sg13g2_xnor2_1 _2912_ (.Y(_2050_),
    .A(\pid.prev_error[3] ),
    .B(net414));
 sg13g2_o21ai_1 _2913_ (.B1(_2041_),
    .Y(_2051_),
    .A1(_2048_),
    .A2(_2049_));
 sg13g2_nor3_1 _2914_ (.A(\pid.prev_error[4] ),
    .B(_1898_),
    .C(_1920_),
    .Y(_2052_));
 sg13g2_xnor2_1 _2915_ (.Y(_2053_),
    .A(\pid.prev_error[4] ),
    .B(net408));
 sg13g2_xor2_1 _2916_ (.B(_2053_),
    .A(_2051_),
    .X(_2054_));
 sg13g2_xnor2_1 _2917_ (.Y(_2055_),
    .A(_2048_),
    .B(_2050_));
 sg13g2_nand2_1 _2918_ (.Y(_2056_),
    .A(net461),
    .B(net397));
 sg13g2_nand3_1 _2919_ (.B(net388),
    .C(net397),
    .A(\pid.Kd[8] ),
    .Y(_2057_));
 sg13g2_o21ai_1 _2920_ (.B1(net461),
    .Y(_2058_),
    .A1(net388),
    .A2(net397));
 sg13g2_nand2b_2 _2921_ (.Y(_2059_),
    .B(_2057_),
    .A_N(_2058_));
 sg13g2_a21oi_1 _2922_ (.A1(_2051_),
    .A2(_2053_),
    .Y(_2060_),
    .B1(_2052_));
 sg13g2_nor2_1 _2923_ (.A(_0843_),
    .B(net404),
    .Y(_2061_));
 sg13g2_xnor2_1 _2924_ (.Y(_2062_),
    .A(\pid.prev_error[5] ),
    .B(net404));
 sg13g2_xnor2_1 _2925_ (.Y(_2063_),
    .A(_2060_),
    .B(_2062_));
 sg13g2_nand2_1 _2926_ (.Y(_2064_),
    .A(\pid.Kd[7] ),
    .B(net386));
 sg13g2_o21ai_1 _2927_ (.B1(_2057_),
    .Y(_2065_),
    .A1(_2059_),
    .A2(_2064_));
 sg13g2_nor2_1 _2928_ (.A(\pid.prev_error[7] ),
    .B(_2036_),
    .Y(_2066_));
 sg13g2_nor2_1 _2929_ (.A(\pid.prev_error[6] ),
    .B(_2027_),
    .Y(_2067_));
 sg13g2_xnor2_1 _2930_ (.Y(_2068_),
    .A(\pid.prev_error[6] ),
    .B(_2027_));
 sg13g2_a221oi_1 _2931_ (.B2(_2053_),
    .C1(_2052_),
    .B1(_2051_),
    .A1(_0843_),
    .Y(_2069_),
    .A2(net404));
 sg13g2_nor3_2 _2932_ (.A(_2061_),
    .B(_2068_),
    .C(_2069_),
    .Y(_2070_));
 sg13g2_nor2_1 _2933_ (.A(_2067_),
    .B(_2070_),
    .Y(_2071_));
 sg13g2_nand2_1 _2934_ (.Y(_2072_),
    .A(\pid.prev_error[7] ),
    .B(_2036_));
 sg13g2_or3_1 _2935_ (.A(_2066_),
    .B(_2067_),
    .C(_2070_),
    .X(_2073_));
 sg13g2_xnor2_1 _2936_ (.Y(_2074_),
    .A(\pid.prev_error[8] ),
    .B(net390));
 sg13g2_nand3_1 _2937_ (.B(_2073_),
    .C(_2074_),
    .A(_2072_),
    .Y(_2075_));
 sg13g2_a21o_1 _2938_ (.A2(_2073_),
    .A1(_2072_),
    .B1(_2074_),
    .X(_2076_));
 sg13g2_and2_2 _2939_ (.A(_2075_),
    .B(_2076_),
    .X(_2077_));
 sg13g2_inv_1 _2940_ (.Y(_2078_),
    .A(net379));
 sg13g2_nand2_1 _2941_ (.Y(_2079_),
    .A(_0015_),
    .B(net379));
 sg13g2_o21ai_1 _2942_ (.B1(_2068_),
    .Y(_2080_),
    .A1(_2061_),
    .A2(_2069_));
 sg13g2_nor2b_1 _2943_ (.A(_2070_),
    .B_N(_2080_),
    .Y(_2081_));
 sg13g2_nor2b_1 _2944_ (.A(_0013_),
    .B_N(net382),
    .Y(_2082_));
 sg13g2_nand2b_1 _2945_ (.Y(_2083_),
    .B(_2072_),
    .A_N(_2066_));
 sg13g2_xor2_1 _2946_ (.B(_2083_),
    .A(_2071_),
    .X(_2084_));
 sg13g2_nand3_1 _2947_ (.B(_2082_),
    .C(net380),
    .A(net463),
    .Y(_2085_));
 sg13g2_a21o_1 _2948_ (.A2(net380),
    .A1(net463),
    .B1(_2082_),
    .X(_2086_));
 sg13g2_and2_1 _2949_ (.A(_2085_),
    .B(_2086_),
    .X(_2087_));
 sg13g2_nand2b_1 _2950_ (.Y(_2088_),
    .B(_2087_),
    .A_N(_2079_));
 sg13g2_xnor2_1 _2951_ (.Y(_2089_),
    .A(_2079_),
    .B(_2087_));
 sg13g2_nor2b_1 _2952_ (.A(_0014_),
    .B_N(net382),
    .Y(_2090_));
 sg13g2_nand3_1 _2953_ (.B(net380),
    .C(_2090_),
    .A(net464),
    .Y(_2091_));
 sg13g2_nand2_1 _2954_ (.Y(_2092_),
    .A(_0016_),
    .B(net379));
 sg13g2_a21o_1 _2955_ (.A2(net380),
    .A1(net464),
    .B1(_2090_),
    .X(_2093_));
 sg13g2_and2_1 _2956_ (.A(_2091_),
    .B(_2093_),
    .X(_2094_));
 sg13g2_nand2b_1 _2957_ (.Y(_2095_),
    .B(_2094_),
    .A_N(_2092_));
 sg13g2_nand2_1 _2958_ (.Y(_2096_),
    .A(_2091_),
    .B(_2095_));
 sg13g2_xnor2_1 _2959_ (.Y(_2097_),
    .A(_2065_),
    .B(_2089_));
 sg13g2_nor2b_1 _2960_ (.A(_2097_),
    .B_N(_2096_),
    .Y(_2098_));
 sg13g2_a21o_1 _2961_ (.A2(_2089_),
    .A1(_2065_),
    .B1(_2098_),
    .X(_2099_));
 sg13g2_xor2_1 _2962_ (.B(_2047_),
    .A(_2046_),
    .X(_2100_));
 sg13g2_xor2_1 _2963_ (.B(_2045_),
    .A(_2044_),
    .X(_2101_));
 sg13g2_xnor2_1 _2964_ (.Y(_2102_),
    .A(\pid.prev_error[0] ),
    .B(_1605_));
 sg13g2_xnor2_1 _2965_ (.Y(_2103_),
    .A(\pid.prev_error[0] ),
    .B(net471));
 sg13g2_nor2_1 _2966_ (.A(_0832_),
    .B(_2102_),
    .Y(_2104_));
 sg13g2_and2_1 _2967_ (.A(net410),
    .B(_2104_),
    .X(_2105_));
 sg13g2_inv_1 _2968_ (.Y(_2106_),
    .A(_2105_));
 sg13g2_nand2_2 _2969_ (.Y(_2107_),
    .A(net401),
    .B(_2105_));
 sg13g2_a21oi_1 _2970_ (.A1(_2045_),
    .A2(_2102_),
    .Y(_2108_),
    .B1(_0832_));
 sg13g2_nand2_2 _2971_ (.Y(_2109_),
    .A(_2106_),
    .B(_2108_));
 sg13g2_nand2_1 _2972_ (.Y(_2110_),
    .A(\pid.Kd[8] ),
    .B(net401));
 sg13g2_nand3_1 _2973_ (.B(_2109_),
    .C(_2110_),
    .A(_2106_),
    .Y(_2111_));
 sg13g2_and2_2 _2974_ (.A(_2107_),
    .B(_2111_),
    .X(_2112_));
 sg13g2_xor2_1 _2975_ (.B(_2064_),
    .A(_2059_),
    .X(_2113_));
 sg13g2_nand2_1 _2976_ (.Y(_2114_),
    .A(_2112_),
    .B(_2113_));
 sg13g2_nand2_1 _2977_ (.Y(_2115_),
    .A(\pid.Kd[8] ),
    .B(net386));
 sg13g2_xor2_1 _2978_ (.B(_2115_),
    .A(_2059_),
    .X(_2116_));
 sg13g2_xnor2_1 _2979_ (.Y(_2117_),
    .A(_2112_),
    .B(_2116_));
 sg13g2_a21oi_1 _2980_ (.A1(_2107_),
    .A2(_2114_),
    .Y(_2118_),
    .B1(_2117_));
 sg13g2_nand3_1 _2981_ (.B(_2114_),
    .C(_2117_),
    .A(_2107_),
    .Y(_2119_));
 sg13g2_nor2b_1 _2982_ (.A(_2118_),
    .B_N(_2119_),
    .Y(_2120_));
 sg13g2_inv_1 _2983_ (.Y(_2121_),
    .A(_2120_));
 sg13g2_xor2_1 _2984_ (.B(_2097_),
    .A(_2096_),
    .X(_2122_));
 sg13g2_nor2_1 _2985_ (.A(_2121_),
    .B(_2122_),
    .Y(_2123_));
 sg13g2_or2_1 _2986_ (.X(_2124_),
    .B(_2123_),
    .A(_2118_));
 sg13g2_nor2b_2 _2987_ (.A(_2107_),
    .B_N(_2116_),
    .Y(_2125_));
 sg13g2_nor2_1 _2988_ (.A(_2111_),
    .B(_2116_),
    .Y(_2126_));
 sg13g2_nor2_2 _2989_ (.A(_2125_),
    .B(_2126_),
    .Y(_2127_));
 sg13g2_nand2_1 _2990_ (.Y(_2128_),
    .A(_2085_),
    .B(_2088_));
 sg13g2_o21ai_1 _2991_ (.B1(_2057_),
    .Y(_2129_),
    .A1(_2059_),
    .A2(_2115_));
 sg13g2_a22oi_1 _2992_ (.Y(_2130_),
    .B1(net380),
    .B2(net462),
    .A2(net382),
    .A1(net461));
 sg13g2_and3_1 _2993_ (.X(_2131_),
    .A(net461),
    .B(net382),
    .C(net380));
 sg13g2_inv_1 _2994_ (.Y(_2132_),
    .A(_2131_));
 sg13g2_nand2_1 _2995_ (.Y(_2133_),
    .A(net462),
    .B(_2131_));
 sg13g2_a21oi_1 _2996_ (.A1(net462),
    .A2(_2131_),
    .Y(_2134_),
    .B1(_2130_));
 sg13g2_nand2_1 _2997_ (.Y(_2135_),
    .A(_0014_),
    .B(net379));
 sg13g2_xor2_1 _2998_ (.B(_2135_),
    .A(_2134_),
    .X(_2136_));
 sg13g2_nand2b_1 _2999_ (.Y(_2137_),
    .B(_2129_),
    .A_N(_2136_));
 sg13g2_xor2_1 _3000_ (.B(_2136_),
    .A(_2129_),
    .X(_2138_));
 sg13g2_nand2b_1 _3001_ (.Y(_2139_),
    .B(_2128_),
    .A_N(_2138_));
 sg13g2_xor2_1 _3002_ (.B(_2138_),
    .A(_2128_),
    .X(_2140_));
 sg13g2_inv_1 _3003_ (.Y(_2141_),
    .A(_2140_));
 sg13g2_xor2_1 _3004_ (.B(_2140_),
    .A(_2127_),
    .X(_2142_));
 sg13g2_nor2b_1 _3005_ (.A(_2142_),
    .B_N(_2124_),
    .Y(_2143_));
 sg13g2_xor2_1 _3006_ (.B(_2142_),
    .A(_2124_),
    .X(_2144_));
 sg13g2_nor2b_1 _3007_ (.A(_2144_),
    .B_N(_2099_),
    .Y(_2145_));
 sg13g2_xnor2_1 _3008_ (.Y(_2146_),
    .A(_2099_),
    .B(_2144_));
 sg13g2_nand2_2 _3009_ (.Y(_2147_),
    .A(net462),
    .B(net388));
 sg13g2_xor2_1 _3010_ (.B(_2147_),
    .A(_2056_),
    .X(_2148_));
 sg13g2_nand3_1 _3011_ (.B(net386),
    .C(_2148_),
    .A(net463),
    .Y(_2149_));
 sg13g2_a21o_1 _3012_ (.A2(net386),
    .A1(net463),
    .B1(_2148_),
    .X(_2150_));
 sg13g2_and2_1 _3013_ (.A(_2149_),
    .B(_2150_),
    .X(_2151_));
 sg13g2_nand2_1 _3014_ (.Y(_2152_),
    .A(_2112_),
    .B(_2151_));
 sg13g2_xnor2_1 _3015_ (.Y(_2153_),
    .A(_2112_),
    .B(_2113_));
 sg13g2_a21oi_1 _3016_ (.A1(_2107_),
    .A2(_2152_),
    .Y(_2154_),
    .B1(_2153_));
 sg13g2_nand3_1 _3017_ (.B(_2152_),
    .C(_2153_),
    .A(_2107_),
    .Y(_2155_));
 sg13g2_nor2b_1 _3018_ (.A(_2154_),
    .B_N(_2155_),
    .Y(_2156_));
 sg13g2_inv_1 _3019_ (.Y(_2157_),
    .A(_2156_));
 sg13g2_nor2b_1 _3020_ (.A(_0015_),
    .B_N(net382),
    .Y(_2158_));
 sg13g2_nand3_1 _3021_ (.B(net381),
    .C(_2158_),
    .A(net465),
    .Y(_2159_));
 sg13g2_nand2_1 _3022_ (.Y(_2160_),
    .A(_0017_),
    .B(_2077_));
 sg13g2_a21o_1 _3023_ (.A2(net380),
    .A1(net465),
    .B1(_2158_),
    .X(_2161_));
 sg13g2_and2_1 _3024_ (.A(_2159_),
    .B(_2161_),
    .X(_2162_));
 sg13g2_nand2b_1 _3025_ (.Y(_2163_),
    .B(_2162_),
    .A_N(_2160_));
 sg13g2_nand2_1 _3026_ (.Y(_2164_),
    .A(_2159_),
    .B(_2163_));
 sg13g2_o21ai_1 _3027_ (.B1(_2149_),
    .Y(_2165_),
    .A1(_2056_),
    .A2(_2147_));
 sg13g2_xnor2_1 _3028_ (.Y(_2166_),
    .A(_2092_),
    .B(_2094_));
 sg13g2_xnor2_1 _3029_ (.Y(_2167_),
    .A(_2165_),
    .B(_2166_));
 sg13g2_nor2b_1 _3030_ (.A(_2167_),
    .B_N(_2164_),
    .Y(_2168_));
 sg13g2_xor2_1 _3031_ (.B(_2167_),
    .A(_2164_),
    .X(_2169_));
 sg13g2_nor2_1 _3032_ (.A(_2157_),
    .B(_2169_),
    .Y(_2170_));
 sg13g2_or2_1 _3033_ (.X(_2171_),
    .B(_2170_),
    .A(_2154_));
 sg13g2_xnor2_1 _3034_ (.Y(_2172_),
    .A(_2121_),
    .B(_2122_));
 sg13g2_nor2b_1 _3035_ (.A(_2172_),
    .B_N(_2171_),
    .Y(_2173_));
 sg13g2_a21o_1 _3036_ (.A2(_2166_),
    .A1(_2165_),
    .B1(_2168_),
    .X(_2174_));
 sg13g2_xor2_1 _3037_ (.B(_2172_),
    .A(_2171_),
    .X(_2175_));
 sg13g2_nor2b_1 _3038_ (.A(_2175_),
    .B_N(_2174_),
    .Y(_2176_));
 sg13g2_o21ai_1 _3039_ (.B1(_2146_),
    .Y(_2177_),
    .A1(_2173_),
    .A2(_2176_));
 sg13g2_nor2_1 _3040_ (.A(_2143_),
    .B(_2145_),
    .Y(_2178_));
 sg13g2_nand2_1 _3041_ (.Y(_2179_),
    .A(_2137_),
    .B(_2139_));
 sg13g2_a21oi_1 _3042_ (.A1(_2127_),
    .A2(_2141_),
    .Y(_2180_),
    .B1(_2125_));
 sg13g2_o21ai_1 _3043_ (.B1(_2133_),
    .Y(_2181_),
    .A1(_2130_),
    .A2(_2135_));
 sg13g2_nand2_1 _3044_ (.Y(_2182_),
    .A(_0013_),
    .B(net379));
 sg13g2_o21ai_1 _3045_ (.B1(net461),
    .Y(_2183_),
    .A1(net382),
    .A2(net380));
 sg13g2_or2_1 _3046_ (.X(_2184_),
    .B(_2183_),
    .A(_2131_));
 sg13g2_xor2_1 _3047_ (.B(_2184_),
    .A(_2182_),
    .X(_2185_));
 sg13g2_nand2_1 _3048_ (.Y(_2186_),
    .A(_2129_),
    .B(_2185_));
 sg13g2_xnor2_1 _3049_ (.Y(_2187_),
    .A(_2129_),
    .B(_2185_));
 sg13g2_nand2b_1 _3050_ (.Y(_2188_),
    .B(_2181_),
    .A_N(_2187_));
 sg13g2_xor2_1 _3051_ (.B(_2187_),
    .A(_2181_),
    .X(_2189_));
 sg13g2_inv_1 _3052_ (.Y(_2190_),
    .A(_2189_));
 sg13g2_xor2_1 _3053_ (.B(_2189_),
    .A(_2127_),
    .X(_2191_));
 sg13g2_nor2_1 _3054_ (.A(_2180_),
    .B(_2191_),
    .Y(_2192_));
 sg13g2_xnor2_1 _3055_ (.Y(_2193_),
    .A(_2180_),
    .B(_2191_));
 sg13g2_nor2b_1 _3056_ (.A(_2193_),
    .B_N(_2179_),
    .Y(_2194_));
 sg13g2_xnor2_1 _3057_ (.Y(_2195_),
    .A(_2179_),
    .B(_2193_));
 sg13g2_o21ai_1 _3058_ (.B1(_2195_),
    .Y(_2196_),
    .A1(_2143_),
    .A2(_2145_));
 sg13g2_xor2_1 _3059_ (.B(_2195_),
    .A(_2178_),
    .X(_2197_));
 sg13g2_or2_1 _3060_ (.X(_2198_),
    .B(_2197_),
    .A(_2177_));
 sg13g2_nand2_1 _3061_ (.Y(_2199_),
    .A(net463),
    .B(net397));
 sg13g2_nand2_1 _3062_ (.Y(_2200_),
    .A(net463),
    .B(net388));
 sg13g2_nand2_1 _3063_ (.Y(_2201_),
    .A(net462),
    .B(net397));
 sg13g2_xor2_1 _3064_ (.B(_2201_),
    .A(_2200_),
    .X(_2202_));
 sg13g2_nand3_1 _3065_ (.B(net386),
    .C(_2202_),
    .A(net464),
    .Y(_2203_));
 sg13g2_a21o_1 _3066_ (.A2(net386),
    .A1(net464),
    .B1(_2202_),
    .X(_2204_));
 sg13g2_and2_1 _3067_ (.A(_2203_),
    .B(_2204_),
    .X(_2205_));
 sg13g2_inv_1 _3068_ (.Y(_2206_),
    .A(_2205_));
 sg13g2_xor2_1 _3069_ (.B(_2110_),
    .A(_2109_),
    .X(_2207_));
 sg13g2_nand2_1 _3070_ (.Y(_2208_),
    .A(net462),
    .B(net401));
 sg13g2_o21ai_1 _3071_ (.B1(_2106_),
    .Y(_2209_),
    .A1(_2109_),
    .A2(_2208_));
 sg13g2_o21ai_1 _3072_ (.B1(_2107_),
    .Y(_2210_),
    .A1(_2207_),
    .A2(_2209_));
 sg13g2_o21ai_1 _3073_ (.B1(_2107_),
    .Y(_2211_),
    .A1(_2206_),
    .A2(_2210_));
 sg13g2_xor2_1 _3074_ (.B(_2151_),
    .A(_2112_),
    .X(_2212_));
 sg13g2_nand2_1 _3075_ (.Y(_2213_),
    .A(_2211_),
    .B(_2212_));
 sg13g2_xor2_1 _3076_ (.B(_2212_),
    .A(_2211_),
    .X(_2214_));
 sg13g2_inv_1 _3077_ (.Y(_2215_),
    .A(_2214_));
 sg13g2_nor2b_1 _3078_ (.A(_0016_),
    .B_N(net383),
    .Y(_2216_));
 sg13g2_nand3_1 _3079_ (.B(net381),
    .C(_2216_),
    .A(\pid.Kd[3] ),
    .Y(_2217_));
 sg13g2_nand2_1 _3080_ (.Y(_2218_),
    .A(_0018_),
    .B(net379));
 sg13g2_a21o_1 _3081_ (.A2(net381),
    .A1(\pid.Kd[3] ),
    .B1(_2216_),
    .X(_2219_));
 sg13g2_and2_1 _3082_ (.A(_2217_),
    .B(_2219_),
    .X(_2220_));
 sg13g2_nand2b_1 _3083_ (.Y(_2221_),
    .B(_2220_),
    .A_N(_2218_));
 sg13g2_nand2_1 _3084_ (.Y(_2222_),
    .A(_2217_),
    .B(_2221_));
 sg13g2_o21ai_1 _3085_ (.B1(_2203_),
    .Y(_2223_),
    .A1(_2147_),
    .A2(_2199_));
 sg13g2_xnor2_1 _3086_ (.Y(_2224_),
    .A(_2160_),
    .B(_2162_));
 sg13g2_nand2_1 _3087_ (.Y(_2225_),
    .A(_2223_),
    .B(_2224_));
 sg13g2_xnor2_1 _3088_ (.Y(_2226_),
    .A(_2223_),
    .B(_2224_));
 sg13g2_nand2b_1 _3089_ (.Y(_2227_),
    .B(_2222_),
    .A_N(_2226_));
 sg13g2_xor2_1 _3090_ (.B(_2226_),
    .A(_2222_),
    .X(_2228_));
 sg13g2_o21ai_1 _3091_ (.B1(_2213_),
    .Y(_2229_),
    .A1(_2215_),
    .A2(_2228_));
 sg13g2_xnor2_1 _3092_ (.Y(_2230_),
    .A(_2157_),
    .B(_2169_));
 sg13g2_nand2b_1 _3093_ (.Y(_2231_),
    .B(_2229_),
    .A_N(_2230_));
 sg13g2_nand2_1 _3094_ (.Y(_2232_),
    .A(_2225_),
    .B(_2227_));
 sg13g2_xor2_1 _3095_ (.B(_2230_),
    .A(_2229_),
    .X(_2233_));
 sg13g2_nand2b_1 _3096_ (.Y(_2234_),
    .B(_2232_),
    .A_N(_2233_));
 sg13g2_nand2_1 _3097_ (.Y(_2235_),
    .A(_2231_),
    .B(_2234_));
 sg13g2_xor2_1 _3098_ (.B(_2175_),
    .A(_2174_),
    .X(_2236_));
 sg13g2_nand2b_1 _3099_ (.Y(_2237_),
    .B(_2235_),
    .A_N(_2236_));
 sg13g2_or3_1 _3100_ (.A(_2146_),
    .B(_2173_),
    .C(_2176_),
    .X(_2238_));
 sg13g2_nand2_1 _3101_ (.Y(_2239_),
    .A(_2177_),
    .B(_2238_));
 sg13g2_nor2_1 _3102_ (.A(_2237_),
    .B(_2239_),
    .Y(_2240_));
 sg13g2_nand3_1 _3103_ (.B(_2076_),
    .C(_2104_),
    .A(_2075_),
    .Y(_2241_));
 sg13g2_a21o_1 _3104_ (.A2(_2076_),
    .A1(_2075_),
    .B1(_2104_),
    .X(_2242_));
 sg13g2_and4_1 _3105_ (.A(\pid.Kd[7] ),
    .B(net410),
    .C(_2241_),
    .D(_2242_),
    .X(_2243_));
 sg13g2_a21o_1 _3106_ (.A2(_2104_),
    .A1(net379),
    .B1(_2243_),
    .X(_2244_));
 sg13g2_xor2_1 _3107_ (.B(_2208_),
    .A(_2109_),
    .X(_2245_));
 sg13g2_and2_1 _3108_ (.A(_2244_),
    .B(_2245_),
    .X(_2246_));
 sg13g2_xor2_1 _3109_ (.B(_2245_),
    .A(_2244_),
    .X(_2247_));
 sg13g2_nand2_1 _3110_ (.Y(_2248_),
    .A(net464),
    .B(net397));
 sg13g2_nand2_1 _3111_ (.Y(_2249_),
    .A(net464),
    .B(net388));
 sg13g2_xor2_1 _3112_ (.B(_2249_),
    .A(_2199_),
    .X(_2250_));
 sg13g2_nand3_1 _3113_ (.B(net386),
    .C(_2250_),
    .A(net465),
    .Y(_2251_));
 sg13g2_a21o_1 _3114_ (.A2(net386),
    .A1(net465),
    .B1(_2250_),
    .X(_2252_));
 sg13g2_and2_1 _3115_ (.A(_2251_),
    .B(_2252_),
    .X(_2253_));
 sg13g2_a21oi_1 _3116_ (.A1(_2247_),
    .A2(_2253_),
    .Y(_2254_),
    .B1(_2246_));
 sg13g2_xor2_1 _3117_ (.B(_2210_),
    .A(_2205_),
    .X(_2255_));
 sg13g2_nor2_1 _3118_ (.A(_2254_),
    .B(_2255_),
    .Y(_2256_));
 sg13g2_xor2_1 _3119_ (.B(_2255_),
    .A(_2254_),
    .X(_2257_));
 sg13g2_nor2b_1 _3120_ (.A(_0017_),
    .B_N(net383),
    .Y(_2258_));
 sg13g2_nand3_1 _3121_ (.B(net381),
    .C(_2258_),
    .A(net466),
    .Y(_2259_));
 sg13g2_a21o_1 _3122_ (.A2(net381),
    .A1(net466),
    .B1(_2258_),
    .X(_2260_));
 sg13g2_and2_1 _3123_ (.A(_2259_),
    .B(_2260_),
    .X(_2261_));
 sg13g2_nand3_1 _3124_ (.B(_2077_),
    .C(_2261_),
    .A(_0019_),
    .Y(_2262_));
 sg13g2_nand2_1 _3125_ (.Y(_2263_),
    .A(_2259_),
    .B(_2262_));
 sg13g2_o21ai_1 _3126_ (.B1(_2251_),
    .Y(_2264_),
    .A1(_2200_),
    .A2(_2248_));
 sg13g2_xnor2_1 _3127_ (.Y(_2265_),
    .A(_2218_),
    .B(_2220_));
 sg13g2_xnor2_1 _3128_ (.Y(_2266_),
    .A(_2264_),
    .B(_2265_));
 sg13g2_nor2b_1 _3129_ (.A(_2266_),
    .B_N(_2263_),
    .Y(_2267_));
 sg13g2_xor2_1 _3130_ (.B(_2266_),
    .A(_2263_),
    .X(_2268_));
 sg13g2_inv_1 _3131_ (.Y(_2269_),
    .A(_2268_));
 sg13g2_a21oi_1 _3132_ (.A1(_2257_),
    .A2(_2269_),
    .Y(_2270_),
    .B1(_2256_));
 sg13g2_xnor2_1 _3133_ (.Y(_2271_),
    .A(_2215_),
    .B(_2228_));
 sg13g2_or2_1 _3134_ (.X(_2272_),
    .B(_2271_),
    .A(_2270_));
 sg13g2_a21o_1 _3135_ (.A2(_2265_),
    .A1(_2264_),
    .B1(_2267_),
    .X(_2273_));
 sg13g2_xor2_1 _3136_ (.B(_2271_),
    .A(_2270_),
    .X(_2274_));
 sg13g2_nand2_1 _3137_ (.Y(_2275_),
    .A(_2273_),
    .B(_2274_));
 sg13g2_xor2_1 _3138_ (.B(_2233_),
    .A(_2232_),
    .X(_2276_));
 sg13g2_a21oi_2 _3139_ (.B1(_2276_),
    .Y(_2277_),
    .A2(_2275_),
    .A1(_2272_));
 sg13g2_xnor2_1 _3140_ (.Y(_2278_),
    .A(_2235_),
    .B(_2236_));
 sg13g2_nand2_1 _3141_ (.Y(_2279_),
    .A(_2277_),
    .B(_2278_));
 sg13g2_nor2_1 _3142_ (.A(_0013_),
    .B(_2102_),
    .Y(_2280_));
 sg13g2_nand3_1 _3143_ (.B(net410),
    .C(_2280_),
    .A(\pid.Kd[6] ),
    .Y(_2281_));
 sg13g2_nand2_2 _3144_ (.Y(_2282_),
    .A(net464),
    .B(net401));
 sg13g2_a21o_1 _3145_ (.A2(net410),
    .A1(\pid.Kd[6] ),
    .B1(_2280_),
    .X(_2283_));
 sg13g2_nand2_1 _3146_ (.Y(_2284_),
    .A(_2281_),
    .B(_2283_));
 sg13g2_o21ai_1 _3147_ (.B1(_2281_),
    .Y(_2285_),
    .A1(_2282_),
    .A2(_2284_));
 sg13g2_inv_1 _3148_ (.Y(_2286_),
    .A(_2285_));
 sg13g2_a22oi_1 _3149_ (.Y(_2287_),
    .B1(_2241_),
    .B2(_2242_),
    .A2(net410),
    .A1(net462));
 sg13g2_or3_1 _3150_ (.A(_2243_),
    .B(_2286_),
    .C(_2287_),
    .X(_2288_));
 sg13g2_o21ai_1 _3151_ (.B1(_2286_),
    .Y(_2289_),
    .A1(_2243_),
    .A2(_2287_));
 sg13g2_nand2_1 _3152_ (.Y(_2290_),
    .A(net465),
    .B(net388));
 sg13g2_nand2_1 _3153_ (.Y(_2291_),
    .A(net463),
    .B(net401));
 sg13g2_xor2_1 _3154_ (.B(_2291_),
    .A(_2248_),
    .X(_2292_));
 sg13g2_nand2b_1 _3155_ (.Y(_2293_),
    .B(_2292_),
    .A_N(_2290_));
 sg13g2_xnor2_1 _3156_ (.Y(_2294_),
    .A(_2290_),
    .B(_2292_));
 sg13g2_nand3_1 _3157_ (.B(_2289_),
    .C(_2294_),
    .A(_2288_),
    .Y(_2295_));
 sg13g2_nand2_2 _3158_ (.Y(_2296_),
    .A(_2288_),
    .B(_2295_));
 sg13g2_xnor2_1 _3159_ (.Y(_2297_),
    .A(_2247_),
    .B(_2253_));
 sg13g2_nand2b_1 _3160_ (.Y(_2298_),
    .B(_2296_),
    .A_N(_2297_));
 sg13g2_xor2_1 _3161_ (.B(_2297_),
    .A(_2296_),
    .X(_2299_));
 sg13g2_nor2b_1 _3162_ (.A(_0017_),
    .B_N(net387),
    .Y(_2300_));
 sg13g2_nand3_1 _3163_ (.B(net383),
    .C(_2300_),
    .A(net466),
    .Y(_2301_));
 sg13g2_nand2_1 _3164_ (.Y(_2302_),
    .A(net468),
    .B(net381));
 sg13g2_a21o_1 _3165_ (.A2(net383),
    .A1(net466),
    .B1(_2300_),
    .X(_2303_));
 sg13g2_and2_1 _3166_ (.A(_2301_),
    .B(_2303_),
    .X(_2304_));
 sg13g2_nand2b_1 _3167_ (.Y(_2305_),
    .B(_2304_),
    .A_N(_2302_));
 sg13g2_nand2_1 _3168_ (.Y(_2306_),
    .A(_2301_),
    .B(_2305_));
 sg13g2_inv_1 _3169_ (.Y(_2307_),
    .A(_2306_));
 sg13g2_o21ai_1 _3170_ (.B1(_2293_),
    .Y(_2308_),
    .A1(_2199_),
    .A2(_2282_));
 sg13g2_a21o_1 _3171_ (.A2(net379),
    .A1(_0019_),
    .B1(_2261_),
    .X(_2309_));
 sg13g2_and2_1 _3172_ (.A(_2262_),
    .B(_2309_),
    .X(_2310_));
 sg13g2_nand2_1 _3173_ (.Y(_2311_),
    .A(_2308_),
    .B(_2310_));
 sg13g2_xnor2_1 _3174_ (.Y(_2312_),
    .A(_2308_),
    .B(_2310_));
 sg13g2_xnor2_1 _3175_ (.Y(_2313_),
    .A(_2307_),
    .B(_2312_));
 sg13g2_o21ai_1 _3176_ (.B1(_2298_),
    .Y(_2314_),
    .A1(_2299_),
    .A2(_2313_));
 sg13g2_xnor2_1 _3177_ (.Y(_2315_),
    .A(_2257_),
    .B(_2269_));
 sg13g2_inv_1 _3178_ (.Y(_2316_),
    .A(_2315_));
 sg13g2_o21ai_1 _3179_ (.B1(_2311_),
    .Y(_2317_),
    .A1(_2307_),
    .A2(_2312_));
 sg13g2_xor2_1 _3180_ (.B(_2315_),
    .A(_2314_),
    .X(_2318_));
 sg13g2_nor2b_1 _3181_ (.A(_2318_),
    .B_N(_2317_),
    .Y(_2319_));
 sg13g2_a21oi_1 _3182_ (.A1(_2314_),
    .A2(_2316_),
    .Y(_2320_),
    .B1(_2319_));
 sg13g2_xnor2_1 _3183_ (.Y(_2321_),
    .A(_2273_),
    .B(_2274_));
 sg13g2_nor2_1 _3184_ (.A(_2320_),
    .B(_2321_),
    .Y(_2322_));
 sg13g2_nand3_1 _3185_ (.B(_2275_),
    .C(_2276_),
    .A(_2272_),
    .Y(_2323_));
 sg13g2_nor2b_1 _3186_ (.A(_2277_),
    .B_N(_2323_),
    .Y(_2324_));
 sg13g2_and2_1 _3187_ (.A(_2322_),
    .B(_2324_),
    .X(_2325_));
 sg13g2_or2_1 _3188_ (.X(_2326_),
    .B(_2324_),
    .A(_2322_));
 sg13g2_nand2b_1 _3189_ (.Y(_2327_),
    .B(_2326_),
    .A_N(_2325_));
 sg13g2_nor2_1 _3190_ (.A(_0014_),
    .B(_2102_),
    .Y(_2328_));
 sg13g2_nand3_1 _3191_ (.B(net410),
    .C(_2328_),
    .A(\pid.Kd[5] ),
    .Y(_2329_));
 sg13g2_nand2_1 _3192_ (.Y(_2330_),
    .A(net465),
    .B(net401));
 sg13g2_a21o_1 _3193_ (.A2(net410),
    .A1(\pid.Kd[5] ),
    .B1(_2328_),
    .X(_2331_));
 sg13g2_nand2_1 _3194_ (.Y(_2332_),
    .A(_2329_),
    .B(_2331_));
 sg13g2_o21ai_1 _3195_ (.B1(_2329_),
    .Y(_2333_),
    .A1(_2330_),
    .A2(_2332_));
 sg13g2_xor2_1 _3196_ (.B(_2284_),
    .A(_2282_),
    .X(_2334_));
 sg13g2_xnor2_1 _3197_ (.Y(_2335_),
    .A(_2333_),
    .B(_2334_));
 sg13g2_nand2_1 _3198_ (.Y(_2336_),
    .A(\pid.Kd[3] ),
    .B(_2055_));
 sg13g2_nand2_1 _3199_ (.Y(_2337_),
    .A(\pid.Kd[3] ),
    .B(_2054_));
 sg13g2_nand2_1 _3200_ (.Y(_2338_),
    .A(\pid.Kd[4] ),
    .B(net397));
 sg13g2_xor2_1 _3201_ (.B(_2338_),
    .A(_2337_),
    .X(_2339_));
 sg13g2_nand3_1 _3202_ (.B(net387),
    .C(_2339_),
    .A(net466),
    .Y(_2340_));
 sg13g2_a21o_1 _3203_ (.A2(net387),
    .A1(net466),
    .B1(_2339_),
    .X(_2341_));
 sg13g2_and2_1 _3204_ (.A(_2340_),
    .B(_2341_),
    .X(_2342_));
 sg13g2_nor2b_1 _3205_ (.A(_2335_),
    .B_N(_2342_),
    .Y(_2343_));
 sg13g2_a21o_1 _3206_ (.A2(_2334_),
    .A1(_2333_),
    .B1(_2343_),
    .X(_2344_));
 sg13g2_a21o_1 _3207_ (.A2(_2289_),
    .A1(_2288_),
    .B1(_2294_),
    .X(_2345_));
 sg13g2_nand3_1 _3208_ (.B(_2344_),
    .C(_2345_),
    .A(_2295_),
    .Y(_2346_));
 sg13g2_a21o_1 _3209_ (.A2(_2345_),
    .A1(_2295_),
    .B1(_2344_),
    .X(_2347_));
 sg13g2_nand2_1 _3210_ (.Y(_2348_),
    .A(net469),
    .B(net381));
 sg13g2_nand2b_1 _3211_ (.Y(_2349_),
    .B(net382),
    .A_N(_0019_));
 sg13g2_or2_1 _3212_ (.X(_2350_),
    .B(_2349_),
    .A(_2348_));
 sg13g2_o21ai_1 _3213_ (.B1(_2340_),
    .Y(_2351_),
    .A1(_2337_),
    .A2(_2338_));
 sg13g2_xnor2_1 _3214_ (.Y(_2352_),
    .A(_2302_),
    .B(_2304_));
 sg13g2_nand2_1 _3215_ (.Y(_2353_),
    .A(_2351_),
    .B(_2352_));
 sg13g2_xnor2_1 _3216_ (.Y(_2354_),
    .A(_2351_),
    .B(_2352_));
 sg13g2_xor2_1 _3217_ (.B(_2354_),
    .A(_2350_),
    .X(_2355_));
 sg13g2_nand3_1 _3218_ (.B(_2347_),
    .C(_2355_),
    .A(_2346_),
    .Y(_2356_));
 sg13g2_nand2_1 _3219_ (.Y(_2357_),
    .A(_2346_),
    .B(_2356_));
 sg13g2_xor2_1 _3220_ (.B(_2313_),
    .A(_2299_),
    .X(_2358_));
 sg13g2_o21ai_1 _3221_ (.B1(_2353_),
    .Y(_2359_),
    .A1(_2350_),
    .A2(_2354_));
 sg13g2_xnor2_1 _3222_ (.Y(_2360_),
    .A(_2357_),
    .B(_2358_));
 sg13g2_nor2b_1 _3223_ (.A(_2360_),
    .B_N(_2359_),
    .Y(_2361_));
 sg13g2_a21oi_1 _3224_ (.A1(_2357_),
    .A2(_2358_),
    .Y(_2362_),
    .B1(_2361_));
 sg13g2_xor2_1 _3225_ (.B(_2318_),
    .A(_2317_),
    .X(_2363_));
 sg13g2_nor2_1 _3226_ (.A(_2362_),
    .B(_2363_),
    .Y(_2364_));
 sg13g2_xor2_1 _3227_ (.B(_2321_),
    .A(_2320_),
    .X(_2365_));
 sg13g2_and2_1 _3228_ (.A(_2364_),
    .B(_2365_),
    .X(_2366_));
 sg13g2_nor2_1 _3229_ (.A(_0015_),
    .B(_2102_),
    .Y(_2367_));
 sg13g2_nand3_1 _3230_ (.B(net411),
    .C(_2367_),
    .A(\pid.Kd[4] ),
    .Y(_2368_));
 sg13g2_nand2_1 _3231_ (.Y(_2369_),
    .A(\pid.Kd[3] ),
    .B(_2100_));
 sg13g2_a21o_1 _3232_ (.A2(net410),
    .A1(net465),
    .B1(_2367_),
    .X(_2370_));
 sg13g2_nand2_1 _3233_ (.Y(_2371_),
    .A(_2368_),
    .B(_2370_));
 sg13g2_o21ai_1 _3234_ (.B1(_2368_),
    .Y(_2372_),
    .A1(_2369_),
    .A2(_2371_));
 sg13g2_xor2_1 _3235_ (.B(_2332_),
    .A(_2330_),
    .X(_2373_));
 sg13g2_xnor2_1 _3236_ (.Y(_2374_),
    .A(_2372_),
    .B(_2373_));
 sg13g2_nand2_1 _3237_ (.Y(_2375_),
    .A(net467),
    .B(_2055_));
 sg13g2_nand2_1 _3238_ (.Y(_2376_),
    .A(net467),
    .B(_2054_));
 sg13g2_xor2_1 _3239_ (.B(_2376_),
    .A(_2336_),
    .X(_2377_));
 sg13g2_nand3_1 _3240_ (.B(net387),
    .C(_2377_),
    .A(net468),
    .Y(_2378_));
 sg13g2_a21o_1 _3241_ (.A2(net387),
    .A1(net468),
    .B1(_2377_),
    .X(_2379_));
 sg13g2_and2_1 _3242_ (.A(_2378_),
    .B(_2379_),
    .X(_2380_));
 sg13g2_nor2b_1 _3243_ (.A(_2374_),
    .B_N(_2380_),
    .Y(_2381_));
 sg13g2_a21o_1 _3244_ (.A2(_2373_),
    .A1(_2372_),
    .B1(_2381_),
    .X(_2382_));
 sg13g2_xnor2_1 _3245_ (.Y(_2383_),
    .A(_2335_),
    .B(_2342_));
 sg13g2_and2_1 _3246_ (.A(_2382_),
    .B(_2383_),
    .X(_2384_));
 sg13g2_xor2_1 _3247_ (.B(_2349_),
    .A(_2348_),
    .X(_2385_));
 sg13g2_o21ai_1 _3248_ (.B1(_2378_),
    .Y(_2386_),
    .A1(_2336_),
    .A2(_2376_));
 sg13g2_nand2_1 _3249_ (.Y(_2387_),
    .A(_2385_),
    .B(_2386_));
 sg13g2_inv_1 _3250_ (.Y(_2388_),
    .A(_2387_));
 sg13g2_xor2_1 _3251_ (.B(_2386_),
    .A(_2385_),
    .X(_2389_));
 sg13g2_xor2_1 _3252_ (.B(_2383_),
    .A(_2382_),
    .X(_2390_));
 sg13g2_a21o_1 _3253_ (.A2(_2390_),
    .A1(_2389_),
    .B1(_2384_),
    .X(_2391_));
 sg13g2_a21o_1 _3254_ (.A2(_2347_),
    .A1(_2346_),
    .B1(_2355_),
    .X(_2392_));
 sg13g2_nand3_1 _3255_ (.B(_2391_),
    .C(_2392_),
    .A(_2356_),
    .Y(_2393_));
 sg13g2_a21o_1 _3256_ (.A2(_2392_),
    .A1(_2356_),
    .B1(_2391_),
    .X(_2394_));
 sg13g2_nand3_1 _3257_ (.B(_2393_),
    .C(_2394_),
    .A(_2388_),
    .Y(_2395_));
 sg13g2_nand2_1 _3258_ (.Y(_2396_),
    .A(_2393_),
    .B(_2395_));
 sg13g2_xor2_1 _3259_ (.B(_2360_),
    .A(_2359_),
    .X(_2397_));
 sg13g2_nand2b_1 _3260_ (.Y(_2398_),
    .B(_2396_),
    .A_N(_2397_));
 sg13g2_xor2_1 _3261_ (.B(_2363_),
    .A(_2362_),
    .X(_2399_));
 sg13g2_nor2b_1 _3262_ (.A(_2398_),
    .B_N(_2399_),
    .Y(_2400_));
 sg13g2_nor2_1 _3263_ (.A(_0016_),
    .B(_2102_),
    .Y(_2401_));
 sg13g2_nand3_1 _3264_ (.B(net411),
    .C(_2401_),
    .A(\pid.Kd[3] ),
    .Y(_2402_));
 sg13g2_nand2_1 _3265_ (.Y(_2403_),
    .A(net467),
    .B(_2100_));
 sg13g2_a21o_1 _3266_ (.A2(_2101_),
    .A1(\pid.Kd[3] ),
    .B1(_2401_),
    .X(_2404_));
 sg13g2_and2_1 _3267_ (.A(_2402_),
    .B(_2404_),
    .X(_2405_));
 sg13g2_nand2b_1 _3268_ (.Y(_2406_),
    .B(_2405_),
    .A_N(_2403_));
 sg13g2_nand2_1 _3269_ (.Y(_2407_),
    .A(_2402_),
    .B(_2406_));
 sg13g2_xor2_1 _3270_ (.B(_2371_),
    .A(_2369_),
    .X(_2408_));
 sg13g2_nand2_1 _3271_ (.Y(_2409_),
    .A(_2407_),
    .B(_2408_));
 sg13g2_xnor2_1 _3272_ (.Y(_2410_),
    .A(_2407_),
    .B(_2408_));
 sg13g2_nand2_2 _3273_ (.Y(_2411_),
    .A(\pid.Kd[1] ),
    .B(net388));
 sg13g2_xor2_1 _3274_ (.B(_2411_),
    .A(_2375_),
    .X(_2412_));
 sg13g2_nand3_1 _3275_ (.B(net387),
    .C(_2412_),
    .A(net469),
    .Y(_2413_));
 sg13g2_a21o_1 _3276_ (.A2(net387),
    .A1(net469),
    .B1(_2412_),
    .X(_2414_));
 sg13g2_nand2_1 _3277_ (.Y(_2415_),
    .A(_2413_),
    .B(_2414_));
 sg13g2_o21ai_1 _3278_ (.B1(_2409_),
    .Y(_2416_),
    .A1(_2410_),
    .A2(_2415_));
 sg13g2_xnor2_1 _3279_ (.Y(_2417_),
    .A(_2374_),
    .B(_2380_));
 sg13g2_nand2_1 _3280_ (.Y(_2418_),
    .A(net469),
    .B(net382));
 sg13g2_o21ai_1 _3281_ (.B1(_2413_),
    .Y(_2419_),
    .A1(_2375_),
    .A2(_2411_));
 sg13g2_nor2b_1 _3282_ (.A(_2418_),
    .B_N(_2419_),
    .Y(_2420_));
 sg13g2_xor2_1 _3283_ (.B(_2419_),
    .A(_2418_),
    .X(_2421_));
 sg13g2_xnor2_1 _3284_ (.Y(_2422_),
    .A(_2416_),
    .B(_2417_));
 sg13g2_nor2_1 _3285_ (.A(_2421_),
    .B(_2422_),
    .Y(_2423_));
 sg13g2_a21oi_1 _3286_ (.A1(_2416_),
    .A2(_2417_),
    .Y(_2424_),
    .B1(_2423_));
 sg13g2_xnor2_1 _3287_ (.Y(_2425_),
    .A(_2389_),
    .B(_2390_));
 sg13g2_xor2_1 _3288_ (.B(_2425_),
    .A(_2424_),
    .X(_2426_));
 sg13g2_nand2_1 _3289_ (.Y(_2427_),
    .A(_2420_),
    .B(_2426_));
 sg13g2_o21ai_1 _3290_ (.B1(_2427_),
    .Y(_2428_),
    .A1(_2424_),
    .A2(_2425_));
 sg13g2_a21o_1 _3291_ (.A2(_2394_),
    .A1(_2393_),
    .B1(_2388_),
    .X(_2429_));
 sg13g2_nand3_1 _3292_ (.B(_2428_),
    .C(_2429_),
    .A(_2395_),
    .Y(_2430_));
 sg13g2_nand2b_1 _3293_ (.Y(_2431_),
    .B(_2077_),
    .A_N(net469));
 sg13g2_inv_1 _3294_ (.Y(_2432_),
    .A(_2431_));
 sg13g2_a21o_1 _3295_ (.A2(_2429_),
    .A1(_2395_),
    .B1(_2428_),
    .X(_2433_));
 sg13g2_nand3_1 _3296_ (.B(_2432_),
    .C(_2433_),
    .A(_2430_),
    .Y(_2434_));
 sg13g2_nand2_1 _3297_ (.Y(_2435_),
    .A(_2430_),
    .B(_2434_));
 sg13g2_xor2_1 _3298_ (.B(_2397_),
    .A(_2396_),
    .X(_2436_));
 sg13g2_a21oi_1 _3299_ (.A1(_2430_),
    .A2(_2434_),
    .Y(_2437_),
    .B1(_2436_));
 sg13g2_xnor2_1 _3300_ (.Y(_2438_),
    .A(_2420_),
    .B(_2426_));
 sg13g2_nor2_1 _3301_ (.A(_0017_),
    .B(_2102_),
    .Y(_2439_));
 sg13g2_nand3_1 _3302_ (.B(net411),
    .C(_2439_),
    .A(net467),
    .Y(_2440_));
 sg13g2_nand2_1 _3303_ (.Y(_2441_),
    .A(\pid.Kd[1] ),
    .B(net401));
 sg13g2_a21o_1 _3304_ (.A2(net411),
    .A1(net466),
    .B1(_2439_),
    .X(_2442_));
 sg13g2_and2_1 _3305_ (.A(_2440_),
    .B(_2442_),
    .X(_2443_));
 sg13g2_nand2b_1 _3306_ (.Y(_2444_),
    .B(_2443_),
    .A_N(_2441_));
 sg13g2_nand2_1 _3307_ (.Y(_2445_),
    .A(_2440_),
    .B(_2444_));
 sg13g2_xnor2_1 _3308_ (.Y(_2446_),
    .A(_2403_),
    .B(_2405_));
 sg13g2_a22oi_1 _3309_ (.Y(_2447_),
    .B1(_2055_),
    .B2(net468),
    .A2(net388),
    .A1(net469));
 sg13g2_nand2_2 _3310_ (.Y(_2448_),
    .A(net470),
    .B(net397));
 sg13g2_nor2_2 _3311_ (.A(_2411_),
    .B(_2448_),
    .Y(_2449_));
 sg13g2_xnor2_1 _3312_ (.Y(_2450_),
    .A(_2445_),
    .B(_2446_));
 sg13g2_nor3_1 _3313_ (.A(_2447_),
    .B(_2449_),
    .C(_2450_),
    .Y(_2451_));
 sg13g2_a21oi_1 _3314_ (.A1(_2445_),
    .A2(_2446_),
    .Y(_2452_),
    .B1(_2451_));
 sg13g2_xor2_1 _3315_ (.B(_2415_),
    .A(_2410_),
    .X(_2453_));
 sg13g2_nor2b_1 _3316_ (.A(_2452_),
    .B_N(_2453_),
    .Y(_2454_));
 sg13g2_xnor2_1 _3317_ (.Y(_2455_),
    .A(_2452_),
    .B(_2453_));
 sg13g2_a21o_1 _3318_ (.A2(_2455_),
    .A1(_2449_),
    .B1(_2454_),
    .X(_2456_));
 sg13g2_xor2_1 _3319_ (.B(_2422_),
    .A(_2421_),
    .X(_2457_));
 sg13g2_nand2_1 _3320_ (.Y(_2458_),
    .A(_2456_),
    .B(_2457_));
 sg13g2_nor2_1 _3321_ (.A(_2438_),
    .B(_2458_),
    .Y(_2459_));
 sg13g2_a21o_1 _3322_ (.A2(_2433_),
    .A1(_2430_),
    .B1(_2432_),
    .X(_2460_));
 sg13g2_nand3_1 _3323_ (.B(_2459_),
    .C(_2460_),
    .A(_2434_),
    .Y(_2461_));
 sg13g2_xor2_1 _3324_ (.B(_2458_),
    .A(_2438_),
    .X(_2462_));
 sg13g2_nor2_1 _3325_ (.A(_0018_),
    .B(_2102_),
    .Y(_2463_));
 sg13g2_nand3_1 _3326_ (.B(net411),
    .C(_2463_),
    .A(net468),
    .Y(_2464_));
 sg13g2_nand2_1 _3327_ (.Y(_2465_),
    .A(net470),
    .B(net401));
 sg13g2_a21o_1 _3328_ (.A2(net411),
    .A1(net468),
    .B1(_2463_),
    .X(_2466_));
 sg13g2_and2_1 _3329_ (.A(_2464_),
    .B(_2466_),
    .X(_2467_));
 sg13g2_nand2b_1 _3330_ (.Y(_2468_),
    .B(_2467_),
    .A_N(_2465_));
 sg13g2_nand2_1 _3331_ (.Y(_2469_),
    .A(_2464_),
    .B(_2468_));
 sg13g2_xnor2_1 _3332_ (.Y(_2470_),
    .A(_2441_),
    .B(_2443_));
 sg13g2_nand2_1 _3333_ (.Y(_2471_),
    .A(_2469_),
    .B(_2470_));
 sg13g2_xnor2_1 _3334_ (.Y(_2472_),
    .A(_2469_),
    .B(_2470_));
 sg13g2_o21ai_1 _3335_ (.B1(_2471_),
    .Y(_2473_),
    .A1(_2448_),
    .A2(_2472_));
 sg13g2_o21ai_1 _3336_ (.B1(_2450_),
    .Y(_2474_),
    .A1(_2447_),
    .A2(_2449_));
 sg13g2_nand2b_1 _3337_ (.Y(_2475_),
    .B(_2474_),
    .A_N(_2451_));
 sg13g2_nand2b_1 _3338_ (.Y(_2476_),
    .B(_2473_),
    .A_N(_2475_));
 sg13g2_xnor2_1 _3339_ (.Y(_2477_),
    .A(_2449_),
    .B(_2455_));
 sg13g2_or2_1 _3340_ (.X(_2478_),
    .B(_2477_),
    .A(_2476_));
 sg13g2_xnor2_1 _3341_ (.Y(_2479_),
    .A(_2456_),
    .B(_2457_));
 sg13g2_nor2_1 _3342_ (.A(_2478_),
    .B(_2479_),
    .Y(_2480_));
 sg13g2_and2_1 _3343_ (.A(_2462_),
    .B(_2480_),
    .X(_2481_));
 sg13g2_nand2_1 _3344_ (.Y(_2482_),
    .A(net469),
    .B(_2103_));
 sg13g2_nand2_2 _3345_ (.Y(_2483_),
    .A(net469),
    .B(net411));
 sg13g2_nand2_2 _3346_ (.Y(_2484_),
    .A(net468),
    .B(_2103_));
 sg13g2_or2_1 _3347_ (.X(_2485_),
    .B(_2484_),
    .A(_2483_));
 sg13g2_xnor2_1 _3348_ (.Y(_2486_),
    .A(_2465_),
    .B(_2467_));
 sg13g2_nor2b_1 _3349_ (.A(_2485_),
    .B_N(_2486_),
    .Y(_2487_));
 sg13g2_xor2_1 _3350_ (.B(_2472_),
    .A(_2448_),
    .X(_2488_));
 sg13g2_nand2_1 _3351_ (.Y(_2489_),
    .A(_2487_),
    .B(_2488_));
 sg13g2_xor2_1 _3352_ (.B(_2475_),
    .A(_2473_),
    .X(_2490_));
 sg13g2_nor2_1 _3353_ (.A(_2489_),
    .B(_2490_),
    .Y(_2491_));
 sg13g2_xor2_1 _3354_ (.B(_2477_),
    .A(_2476_),
    .X(_2492_));
 sg13g2_nand2_1 _3355_ (.Y(_2493_),
    .A(_2491_),
    .B(_2492_));
 sg13g2_nor2_1 _3356_ (.A(_2479_),
    .B(_2493_),
    .Y(_2494_));
 sg13g2_xor2_1 _3357_ (.B(_2480_),
    .A(_2462_),
    .X(_2495_));
 sg13g2_a21oi_1 _3358_ (.A1(_2494_),
    .A2(_2495_),
    .Y(_2496_),
    .B1(_2481_));
 sg13g2_inv_1 _3359_ (.Y(_2497_),
    .A(_2496_));
 sg13g2_a21oi_1 _3360_ (.A1(_2434_),
    .A2(_2460_),
    .Y(_2498_),
    .B1(_2459_));
 sg13g2_a21o_1 _3361_ (.A2(_2460_),
    .A1(_2434_),
    .B1(_2459_),
    .X(_2499_));
 sg13g2_nand3_1 _3362_ (.B(_2497_),
    .C(_2499_),
    .A(_2461_),
    .Y(_2500_));
 sg13g2_o21ai_1 _3363_ (.B1(_2461_),
    .Y(_2501_),
    .A1(_2496_),
    .A2(_2498_));
 sg13g2_xnor2_1 _3364_ (.Y(_2502_),
    .A(_2435_),
    .B(_2436_));
 sg13g2_a21o_1 _3365_ (.A2(_2502_),
    .A1(_2501_),
    .B1(_2437_),
    .X(_2503_));
 sg13g2_xnor2_1 _3366_ (.Y(_2504_),
    .A(_2398_),
    .B(_2399_));
 sg13g2_a21o_1 _3367_ (.A2(_2504_),
    .A1(_2503_),
    .B1(_2400_),
    .X(_2505_));
 sg13g2_xnor2_1 _3368_ (.Y(_2506_),
    .A(_2364_),
    .B(_2365_));
 sg13g2_inv_1 _3369_ (.Y(_2507_),
    .A(_2506_));
 sg13g2_a21o_1 _3370_ (.A2(_2507_),
    .A1(_2505_),
    .B1(_2366_),
    .X(_2508_));
 sg13g2_a21oi_1 _3371_ (.A1(_2326_),
    .A2(_2508_),
    .Y(_2509_),
    .B1(_2325_));
 sg13g2_xnor2_1 _3372_ (.Y(_2510_),
    .A(_2277_),
    .B(_2278_));
 sg13g2_o21ai_1 _3373_ (.B1(_2279_),
    .Y(_2511_),
    .A1(_2509_),
    .A2(_2510_));
 sg13g2_xor2_1 _3374_ (.B(_2239_),
    .A(_2237_),
    .X(_2512_));
 sg13g2_a21oi_1 _3375_ (.A1(_2511_),
    .A2(_2512_),
    .Y(_2513_),
    .B1(_2240_));
 sg13g2_xor2_1 _3376_ (.B(_2197_),
    .A(_2177_),
    .X(_2514_));
 sg13g2_inv_1 _3377_ (.Y(_2515_),
    .A(_2514_));
 sg13g2_o21ai_1 _3378_ (.B1(_2198_),
    .Y(_2516_),
    .A1(_2515_),
    .A2(_2513_));
 sg13g2_nand2_1 _3379_ (.Y(_2517_),
    .A(_2186_),
    .B(_2188_));
 sg13g2_a21oi_1 _3380_ (.A1(_2127_),
    .A2(_2190_),
    .Y(_2518_),
    .B1(_2125_));
 sg13g2_o21ai_1 _3381_ (.B1(_2132_),
    .Y(_2519_),
    .A1(_2182_),
    .A2(_2184_));
 sg13g2_o21ai_1 _3382_ (.B1(_2184_),
    .Y(_2520_),
    .A1(net461),
    .A2(_2078_));
 sg13g2_and2_1 _3383_ (.A(_2129_),
    .B(_2520_),
    .X(_2521_));
 sg13g2_xor2_1 _3384_ (.B(_2520_),
    .A(_2129_),
    .X(_2522_));
 sg13g2_xor2_1 _3385_ (.B(_2522_),
    .A(_2519_),
    .X(_2523_));
 sg13g2_xnor2_1 _3386_ (.Y(_2524_),
    .A(_2127_),
    .B(_2523_));
 sg13g2_xnor2_1 _3387_ (.Y(_2525_),
    .A(_2518_),
    .B(_2524_));
 sg13g2_nand2b_1 _3388_ (.Y(_2526_),
    .B(_2517_),
    .A_N(_2525_));
 sg13g2_xnor2_1 _3389_ (.Y(_2527_),
    .A(_2517_),
    .B(_2525_));
 sg13g2_o21ai_1 _3390_ (.B1(_2527_),
    .Y(_2528_),
    .A1(_2192_),
    .A2(_2194_));
 sg13g2_or3_1 _3391_ (.A(_2192_),
    .B(_2194_),
    .C(_2527_),
    .X(_2529_));
 sg13g2_nand2_1 _3392_ (.Y(_2530_),
    .A(_2528_),
    .B(_2529_));
 sg13g2_xor2_1 _3393_ (.B(_2530_),
    .A(_2196_),
    .X(_2531_));
 sg13g2_nand2_1 _3394_ (.Y(_2532_),
    .A(net87),
    .B(_2531_));
 sg13g2_o21ai_1 _3395_ (.B1(_2526_),
    .Y(_2533_),
    .A1(_2518_),
    .A2(_2524_));
 sg13g2_a21oi_1 _3396_ (.A1(_2127_),
    .A2(_2523_),
    .Y(_2534_),
    .B1(_2125_));
 sg13g2_a21oi_1 _3397_ (.A1(_2519_),
    .A2(_2522_),
    .Y(_2535_),
    .B1(_2521_));
 sg13g2_xnor2_1 _3398_ (.Y(_2536_),
    .A(_2127_),
    .B(_2132_));
 sg13g2_xnor2_1 _3399_ (.Y(_2537_),
    .A(_2522_),
    .B(_2536_));
 sg13g2_xnor2_1 _3400_ (.Y(_2538_),
    .A(_2535_),
    .B(_2537_));
 sg13g2_xnor2_1 _3401_ (.Y(_2539_),
    .A(_2534_),
    .B(_2538_));
 sg13g2_xnor2_1 _3402_ (.Y(_2540_),
    .A(_2533_),
    .B(_2539_));
 sg13g2_xnor2_1 _3403_ (.Y(_2541_),
    .A(_2528_),
    .B(_2540_));
 sg13g2_o21ai_1 _3404_ (.B1(_2541_),
    .Y(_2542_),
    .A1(_2196_),
    .A2(_2530_));
 sg13g2_nand2b_1 _3405_ (.Y(_2543_),
    .B(_2532_),
    .A_N(_2542_));
 sg13g2_inv_1 _3406_ (.Y(_2544_),
    .A(net372));
 sg13g2_or2_1 _3407_ (.X(_2545_),
    .B(_2531_),
    .A(net87));
 sg13g2_xnor2_1 _3408_ (.Y(_2546_),
    .A(_2509_),
    .B(_2510_));
 sg13g2_xor2_1 _3409_ (.B(_2508_),
    .A(_2327_),
    .X(_2547_));
 sg13g2_xnor2_1 _3410_ (.Y(_2548_),
    .A(_2505_),
    .B(_2507_));
 sg13g2_xnor2_1 _3411_ (.Y(_2549_),
    .A(_2503_),
    .B(_2504_));
 sg13g2_xnor2_1 _3412_ (.Y(_2550_),
    .A(_2501_),
    .B(_2502_));
 sg13g2_nand3_1 _3413_ (.B(_2483_),
    .C(_2484_),
    .A(_2482_),
    .Y(_2551_));
 sg13g2_xnor2_1 _3414_ (.Y(_2552_),
    .A(_2485_),
    .B(_2486_));
 sg13g2_or2_1 _3415_ (.X(_2553_),
    .B(_2552_),
    .A(_2551_));
 sg13g2_xnor2_1 _3416_ (.Y(_2554_),
    .A(_2487_),
    .B(_2488_));
 sg13g2_nand2b_1 _3417_ (.Y(_2555_),
    .B(_2554_),
    .A_N(_2553_));
 sg13g2_xor2_1 _3418_ (.B(_2490_),
    .A(_2489_),
    .X(_2556_));
 sg13g2_nor2_1 _3419_ (.A(_2555_),
    .B(_2556_),
    .Y(_2557_));
 sg13g2_xnor2_1 _3420_ (.Y(_2558_),
    .A(_2491_),
    .B(_2492_));
 sg13g2_or2_1 _3421_ (.X(_2559_),
    .B(_2557_),
    .A(net372));
 sg13g2_or2_1 _3422_ (.X(_2560_),
    .B(_2559_),
    .A(_2558_));
 sg13g2_nand2_1 _3423_ (.Y(_2561_),
    .A(_2558_),
    .B(_2559_));
 sg13g2_and2_1 _3424_ (.A(_2560_),
    .B(_2561_),
    .X(_2562_));
 sg13g2_nand2_1 _3425_ (.Y(_2563_),
    .A(_2557_),
    .B(_2558_));
 sg13g2_nand2_1 _3426_ (.Y(_2564_),
    .A(_2478_),
    .B(_2493_));
 sg13g2_xor2_1 _3427_ (.B(_2564_),
    .A(_2479_),
    .X(_2565_));
 sg13g2_nand2b_1 _3428_ (.Y(_2566_),
    .B(_2565_),
    .A_N(_2563_));
 sg13g2_xnor2_1 _3429_ (.Y(_2567_),
    .A(_2494_),
    .B(_2495_));
 sg13g2_nand2_1 _3430_ (.Y(_2568_),
    .A(net371),
    .B(_2566_));
 sg13g2_or2_1 _3431_ (.X(_2569_),
    .B(_2568_),
    .A(_2567_));
 sg13g2_nand2_1 _3432_ (.Y(_2570_),
    .A(_2567_),
    .B(_2568_));
 sg13g2_and2_1 _3433_ (.A(_2569_),
    .B(_2570_),
    .X(_2571_));
 sg13g2_nand2b_1 _3434_ (.Y(_2572_),
    .B(_2567_),
    .A_N(_2566_));
 sg13g2_a21o_1 _3435_ (.A2(_2499_),
    .A1(_2461_),
    .B1(_2497_),
    .X(_2573_));
 sg13g2_nand2_1 _3436_ (.Y(_2574_),
    .A(_2500_),
    .B(_2573_));
 sg13g2_nand2_1 _3437_ (.Y(_2575_),
    .A(net371),
    .B(_2572_));
 sg13g2_or2_1 _3438_ (.X(_2576_),
    .B(_2575_),
    .A(_2574_));
 sg13g2_nand2_1 _3439_ (.Y(_2577_),
    .A(_2574_),
    .B(_2575_));
 sg13g2_nand2_1 _3440_ (.Y(_2578_),
    .A(_2576_),
    .B(_2577_));
 sg13g2_a21oi_1 _3441_ (.A1(_2500_),
    .A2(_2573_),
    .Y(_2579_),
    .B1(_2572_));
 sg13g2_and2_1 _3442_ (.A(_2550_),
    .B(_2579_),
    .X(_2580_));
 sg13g2_and2_1 _3443_ (.A(_2549_),
    .B(_2580_),
    .X(_2581_));
 sg13g2_and2_1 _3444_ (.A(_2548_),
    .B(_2581_),
    .X(_2582_));
 sg13g2_and2_1 _3445_ (.A(_2547_),
    .B(_2582_),
    .X(_2583_));
 sg13g2_a221oi_1 _3446_ (.B2(_2582_),
    .C1(_2542_),
    .B1(_2547_),
    .A1(net87),
    .Y(_2584_),
    .A2(_2531_));
 sg13g2_xnor2_1 _3447_ (.Y(_2585_),
    .A(_2546_),
    .B(_2584_));
 sg13g2_a221oi_1 _3448_ (.B2(_2581_),
    .C1(_2542_),
    .B1(_2548_),
    .A1(net87),
    .Y(_2586_),
    .A2(_2531_));
 sg13g2_xnor2_1 _3449_ (.Y(_2587_),
    .A(_2547_),
    .B(_2586_));
 sg13g2_a221oi_1 _3450_ (.B2(_2580_),
    .C1(_2542_),
    .B1(_2549_),
    .A1(net87),
    .Y(_2588_),
    .A2(_2531_));
 sg13g2_xnor2_1 _3451_ (.Y(_2589_),
    .A(_2588_),
    .B(_2548_));
 sg13g2_xnor2_1 _3452_ (.Y(_2590_),
    .A(_2513_),
    .B(_2514_));
 sg13g2_xnor2_1 _3453_ (.Y(_2591_),
    .A(_2511_),
    .B(_2512_));
 sg13g2_and2_1 _3454_ (.A(_2546_),
    .B(_2583_),
    .X(_2592_));
 sg13g2_a221oi_1 _3455_ (.B2(_2583_),
    .C1(_2542_),
    .B1(_2546_),
    .A1(net87),
    .Y(_2593_),
    .A2(_2531_));
 sg13g2_a221oi_1 _3456_ (.B2(_2592_),
    .C1(_2542_),
    .B1(_2591_),
    .A1(net87),
    .Y(_2594_),
    .A2(_2531_));
 sg13g2_xor2_1 _3457_ (.B(_2594_),
    .A(_2590_),
    .X(_2595_));
 sg13g2_or2_1 _3458_ (.X(_2596_),
    .B(_2589_),
    .A(_2587_));
 sg13g2_nor3_1 _3459_ (.A(_2585_),
    .B(_2587_),
    .C(_2589_),
    .Y(_2597_));
 sg13g2_or3_1 _3460_ (.A(_2585_),
    .B(_2587_),
    .C(_2589_),
    .X(_2598_));
 sg13g2_xor2_1 _3461_ (.B(_2593_),
    .A(_2591_),
    .X(_2599_));
 sg13g2_nor2b_1 _3462_ (.A(_2599_),
    .B_N(_2595_),
    .Y(_2600_));
 sg13g2_nand2b_1 _3463_ (.Y(_2601_),
    .B(_2595_),
    .A_N(_2599_));
 sg13g2_nand2_1 _3464_ (.Y(_2602_),
    .A(_2598_),
    .B(_2600_));
 sg13g2_nand3_1 _3465_ (.B(_2542_),
    .C(_2545_),
    .A(_2532_),
    .Y(_2603_));
 sg13g2_a22oi_1 _3466_ (.Y(_2604_),
    .B1(_2598_),
    .B2(_2600_),
    .A2(_2545_),
    .A1(_2542_));
 sg13g2_o21ai_1 _3467_ (.B1(_2603_),
    .Y(_2605_),
    .A1(_2597_),
    .A2(_2601_));
 sg13g2_nand2b_1 _3468_ (.Y(_2606_),
    .B(_2605_),
    .A_N(_2589_));
 sg13g2_o21ai_1 _3469_ (.B1(_2585_),
    .Y(_2607_),
    .A1(_2596_),
    .A2(_2604_));
 sg13g2_nand2_1 _3470_ (.Y(_2608_),
    .A(_2603_),
    .B(_2607_));
 sg13g2_xnor2_1 _3471_ (.Y(_2609_),
    .A(_2589_),
    .B(_2605_));
 sg13g2_xnor2_1 _3472_ (.Y(_2610_),
    .A(_2589_),
    .B(_2604_));
 sg13g2_nor2_1 _3473_ (.A(net372),
    .B(_2580_),
    .Y(_2611_));
 sg13g2_xor2_1 _3474_ (.B(_2611_),
    .A(_2549_),
    .X(_2612_));
 sg13g2_nor2b_1 _3475_ (.A(_2587_),
    .B_N(_2612_),
    .Y(_2613_));
 sg13g2_and2_1 _3476_ (.A(_2609_),
    .B(_2612_),
    .X(_2614_));
 sg13g2_nand2_1 _3477_ (.Y(_2615_),
    .A(_2609_),
    .B(_2613_));
 sg13g2_and2_1 _3478_ (.A(_2595_),
    .B(_2602_),
    .X(_2616_));
 sg13g2_nand2b_1 _3479_ (.Y(_2617_),
    .B(_2602_),
    .A_N(_2599_));
 sg13g2_a221oi_1 _3480_ (.B2(_2609_),
    .C1(_2617_),
    .B1(_2613_),
    .A1(_2603_),
    .Y(_2618_),
    .A2(_2607_));
 sg13g2_nor2_1 _3481_ (.A(_2616_),
    .B(_2618_),
    .Y(_2619_));
 sg13g2_o21ai_1 _3482_ (.B1(_2615_),
    .Y(_2620_),
    .A1(_2616_),
    .A2(_2618_));
 sg13g2_nand2b_1 _3483_ (.Y(_2621_),
    .B(_2608_),
    .A_N(_2620_));
 sg13g2_xor2_1 _3484_ (.B(_2620_),
    .A(_2608_),
    .X(_2622_));
 sg13g2_o21ai_1 _3485_ (.B1(_2612_),
    .Y(_2623_),
    .A1(_2616_),
    .A2(_2618_));
 sg13g2_o21ai_1 _3486_ (.B1(_2614_),
    .Y(_2624_),
    .A1(_2616_),
    .A2(_2618_));
 sg13g2_xor2_1 _3487_ (.B(_2606_),
    .A(_2587_),
    .X(_2625_));
 sg13g2_xnor2_1 _3488_ (.Y(_2626_),
    .A(_2624_),
    .B(_2625_));
 sg13g2_or3_1 _3489_ (.A(_2612_),
    .B(_2616_),
    .C(_2618_),
    .X(_2627_));
 sg13g2_and2_1 _3490_ (.A(_2623_),
    .B(_2627_),
    .X(_2628_));
 sg13g2_inv_1 _3491_ (.Y(_2629_),
    .A(_2628_));
 sg13g2_or3_1 _3492_ (.A(net372),
    .B(_2550_),
    .C(_2579_),
    .X(_2630_));
 sg13g2_o21ai_1 _3493_ (.B1(_2550_),
    .Y(_2631_),
    .A1(net372),
    .A2(_2579_));
 sg13g2_and2_1 _3494_ (.A(_2630_),
    .B(_2631_),
    .X(_2632_));
 sg13g2_nor2_1 _3495_ (.A(_2610_),
    .B(_2632_),
    .Y(_2633_));
 sg13g2_and3_1 _3496_ (.X(_2634_),
    .A(_2623_),
    .B(_2627_),
    .C(_2633_));
 sg13g2_or2_1 _3497_ (.X(_2635_),
    .B(_2634_),
    .A(_2626_));
 sg13g2_nor2_1 _3498_ (.A(_2622_),
    .B(_2635_),
    .Y(_2636_));
 sg13g2_or3_1 _3499_ (.A(_2622_),
    .B(_2626_),
    .C(_2634_),
    .X(_2637_));
 sg13g2_xnor2_1 _3500_ (.Y(_2638_),
    .A(_2617_),
    .B(_2621_));
 sg13g2_and2_1 _3501_ (.A(_2637_),
    .B(_2638_),
    .X(_2639_));
 sg13g2_a21oi_2 _3502_ (.B1(_2632_),
    .Y(_2640_),
    .A2(_2638_),
    .A1(_2637_));
 sg13g2_a221oi_1 _3503_ (.B2(_2638_),
    .C1(_2629_),
    .B1(_2637_),
    .A1(_2630_),
    .Y(_2641_),
    .A2(_2631_));
 sg13g2_xnor2_1 _3504_ (.Y(_2642_),
    .A(_2609_),
    .B(_2623_));
 sg13g2_xor2_1 _3505_ (.B(_2642_),
    .A(_2641_),
    .X(_2643_));
 sg13g2_o21ai_1 _3506_ (.B1(_2626_),
    .Y(_2644_),
    .A1(_2634_),
    .A2(_2638_));
 sg13g2_or2_1 _3507_ (.X(_2645_),
    .B(_2639_),
    .A(_2635_));
 sg13g2_o21ai_1 _3508_ (.B1(_2644_),
    .Y(_2646_),
    .A1(_2635_),
    .A2(_2639_));
 sg13g2_and3_1 _3509_ (.X(_2647_),
    .A(_2632_),
    .B(_2637_),
    .C(_2638_));
 sg13g2_or2_1 _3510_ (.X(_2648_),
    .B(_2647_),
    .A(_2640_));
 sg13g2_nand2_1 _3511_ (.Y(_2649_),
    .A(_2578_),
    .B(_2628_));
 sg13g2_nor3_1 _3512_ (.A(_2640_),
    .B(_2647_),
    .C(_2649_),
    .Y(_2650_));
 sg13g2_nor3_1 _3513_ (.A(_2643_),
    .B(_2646_),
    .C(_2650_),
    .Y(_2651_));
 sg13g2_or3_1 _3514_ (.A(_2643_),
    .B(_2646_),
    .C(_2650_),
    .X(_2652_));
 sg13g2_a21oi_1 _3515_ (.A1(_2622_),
    .A2(_2645_),
    .Y(_2653_),
    .B1(_2636_));
 sg13g2_a21o_1 _3516_ (.A2(_2645_),
    .A1(_2622_),
    .B1(_2636_),
    .X(_2654_));
 sg13g2_nor2_1 _3517_ (.A(_2651_),
    .B(_2653_),
    .Y(_2655_));
 sg13g2_inv_1 _3518_ (.Y(_2656_),
    .A(_2655_));
 sg13g2_o21ai_1 _3519_ (.B1(_2578_),
    .Y(_2657_),
    .A1(_2651_),
    .A2(_2653_));
 sg13g2_nand4_1 _3520_ (.B(_2577_),
    .C(_2652_),
    .A(_2576_),
    .Y(_2658_),
    .D(_2654_));
 sg13g2_nand2_2 _3521_ (.Y(_2659_),
    .A(_2657_),
    .B(_2658_));
 sg13g2_inv_1 _3522_ (.Y(_2660_),
    .A(_2659_));
 sg13g2_a21oi_1 _3523_ (.A1(_2652_),
    .A2(_2654_),
    .Y(_2661_),
    .B1(_2650_));
 sg13g2_nand2b_1 _3524_ (.Y(_2662_),
    .B(_2661_),
    .A_N(_2643_));
 sg13g2_xnor2_1 _3525_ (.Y(_2663_),
    .A(_2643_),
    .B(_2661_));
 sg13g2_nor2_1 _3526_ (.A(_2571_),
    .B(_2648_),
    .Y(_2664_));
 sg13g2_nor2b_1 _3527_ (.A(_2659_),
    .B_N(_2664_),
    .Y(_2665_));
 sg13g2_nand3_1 _3528_ (.B(_2658_),
    .C(_2664_),
    .A(_2657_),
    .Y(_2666_));
 sg13g2_a221oi_1 _3529_ (.B2(_2654_),
    .C1(_2648_),
    .B1(_2652_),
    .A1(_2576_),
    .Y(_2667_),
    .A2(_2577_));
 sg13g2_o21ai_1 _3530_ (.B1(_2629_),
    .Y(_2668_),
    .A1(_2640_),
    .A2(_2667_));
 sg13g2_or3_1 _3531_ (.A(_2629_),
    .B(_2640_),
    .C(_2667_),
    .X(_2669_));
 sg13g2_nand2_1 _3532_ (.Y(_2670_),
    .A(_2668_),
    .B(_2669_));
 sg13g2_nor2_1 _3533_ (.A(_2665_),
    .B(_2670_),
    .Y(_2671_));
 sg13g2_and2_1 _3534_ (.A(_2663_),
    .B(_2671_),
    .X(_2672_));
 sg13g2_nand4_1 _3535_ (.B(_2669_),
    .C(_2668_),
    .A(_2663_),
    .Y(_2673_),
    .D(_2666_));
 sg13g2_xnor2_1 _3536_ (.Y(_2674_),
    .A(_2646_),
    .B(_2662_));
 sg13g2_nand2_2 _3537_ (.Y(_2675_),
    .A(_2673_),
    .B(_2674_));
 sg13g2_nand3_1 _3538_ (.B(_2673_),
    .C(_2674_),
    .A(_2571_),
    .Y(_2676_));
 sg13g2_a21o_1 _3539_ (.A2(_2674_),
    .A1(_2673_),
    .B1(_2571_),
    .X(_2677_));
 sg13g2_nand2_1 _3540_ (.Y(_2678_),
    .A(net371),
    .B(_2563_));
 sg13g2_or2_1 _3541_ (.X(_2679_),
    .B(_2678_),
    .A(_2565_));
 sg13g2_nand2_1 _3542_ (.Y(_2680_),
    .A(_2565_),
    .B(_2678_));
 sg13g2_and2_1 _3543_ (.A(_2679_),
    .B(_2680_),
    .X(_2681_));
 sg13g2_a21oi_1 _3544_ (.A1(_2673_),
    .A2(_2674_),
    .Y(_2682_),
    .B1(_2665_));
 sg13g2_a21oi_1 _3545_ (.A1(_2671_),
    .A2(_2675_),
    .Y(_2683_),
    .B1(_2663_));
 sg13g2_nor2_1 _3546_ (.A(_2672_),
    .B(_2683_),
    .Y(_2684_));
 sg13g2_or2_1 _3547_ (.X(_2685_),
    .B(_2683_),
    .A(_2672_));
 sg13g2_a221oi_1 _3548_ (.B2(_2674_),
    .C1(_2659_),
    .B1(_2673_),
    .A1(_2569_),
    .Y(_2686_),
    .A2(_2570_));
 sg13g2_xor2_1 _3549_ (.B(_2657_),
    .A(_2648_),
    .X(_2687_));
 sg13g2_or2_1 _3550_ (.X(_2688_),
    .B(_2674_),
    .A(_2666_));
 sg13g2_o21ai_1 _3551_ (.B1(_2688_),
    .Y(_2689_),
    .A1(_2686_),
    .A2(_2687_));
 sg13g2_nand2_1 _3552_ (.Y(_2690_),
    .A(_2676_),
    .B(_2677_));
 sg13g2_nor2_1 _3553_ (.A(_2659_),
    .B(_2681_),
    .Y(_2691_));
 sg13g2_nand3_1 _3554_ (.B(_2677_),
    .C(_2691_),
    .A(_2676_),
    .Y(_2692_));
 sg13g2_xnor2_1 _3555_ (.Y(_2693_),
    .A(_2670_),
    .B(_2682_));
 sg13g2_and3_1 _3556_ (.X(_2694_),
    .A(_2689_),
    .B(_2692_),
    .C(_2693_));
 sg13g2_nand3_1 _3557_ (.B(_2692_),
    .C(_2693_),
    .A(_2689_),
    .Y(_2695_));
 sg13g2_nor2_2 _3558_ (.A(_2684_),
    .B(_2694_),
    .Y(_2696_));
 sg13g2_a21oi_2 _3559_ (.B1(_2681_),
    .Y(_2697_),
    .A2(_2695_),
    .A1(_2685_));
 sg13g2_a221oi_1 _3560_ (.B2(_2695_),
    .C1(_2690_),
    .B1(_2685_),
    .A1(_2679_),
    .Y(_2698_),
    .A2(_2680_));
 sg13g2_xnor2_1 _3561_ (.Y(_2699_),
    .A(_2659_),
    .B(_2677_));
 sg13g2_mux2_1 _3562_ (.A0(_2699_),
    .A1(_2660_),
    .S(_2698_),
    .X(_2700_));
 sg13g2_and3_1 _3563_ (.X(_2701_),
    .A(_2681_),
    .B(_2685_),
    .C(_2695_));
 sg13g2_or2_1 _3564_ (.X(_2702_),
    .B(_2701_),
    .A(_2697_));
 sg13g2_nor4_1 _3565_ (.A(_2562_),
    .B(_2690_),
    .C(_2697_),
    .D(_2701_),
    .Y(_2703_));
 sg13g2_o21ai_1 _3566_ (.B1(_2692_),
    .Y(_2704_),
    .A1(_2684_),
    .A2(_2694_));
 sg13g2_nand3b_1 _3567_ (.B(_2689_),
    .C(_2692_),
    .Y(_2705_),
    .A_N(_2696_));
 sg13g2_xnor2_1 _3568_ (.Y(_2706_),
    .A(_2689_),
    .B(_2704_));
 sg13g2_nand3b_1 _3569_ (.B(_2706_),
    .C(_2700_),
    .Y(_2707_),
    .A_N(_2703_));
 sg13g2_xor2_1 _3570_ (.B(_2705_),
    .A(_2693_),
    .X(_2708_));
 sg13g2_and2_1 _3571_ (.A(_2707_),
    .B(_2708_),
    .X(_2709_));
 sg13g2_a21oi_1 _3572_ (.A1(_2707_),
    .A2(_2708_),
    .Y(_2710_),
    .B1(_2703_));
 sg13g2_and2_1 _3573_ (.A(_2700_),
    .B(_2710_),
    .X(_2711_));
 sg13g2_o21ai_1 _3574_ (.B1(_2707_),
    .Y(_2712_),
    .A1(_2706_),
    .A2(_2711_));
 sg13g2_nor2_1 _3575_ (.A(_2562_),
    .B(_2709_),
    .Y(_2713_));
 sg13g2_a21o_1 _3576_ (.A2(_2708_),
    .A1(_2707_),
    .B1(_2562_),
    .X(_2714_));
 sg13g2_a221oi_1 _3577_ (.B2(_2708_),
    .C1(_2702_),
    .B1(_2707_),
    .A1(_2560_),
    .Y(_2715_),
    .A2(_2561_));
 sg13g2_o21ai_1 _3578_ (.B1(_2690_),
    .Y(_2716_),
    .A1(_2697_),
    .A2(_2715_));
 sg13g2_or3_1 _3579_ (.A(_2690_),
    .B(_2697_),
    .C(_2715_),
    .X(_2717_));
 sg13g2_and2_1 _3580_ (.A(_2716_),
    .B(_2717_),
    .X(_2718_));
 sg13g2_xor2_1 _3581_ (.B(_2710_),
    .A(_2700_),
    .X(_2719_));
 sg13g2_nand3_1 _3582_ (.B(_2707_),
    .C(_2708_),
    .A(_2562_),
    .Y(_2720_));
 sg13g2_nand2_1 _3583_ (.Y(_2721_),
    .A(_2714_),
    .B(_2720_));
 sg13g2_inv_1 _3584_ (.Y(_2722_),
    .A(_2721_));
 sg13g2_nand2_1 _3585_ (.Y(_2723_),
    .A(net371),
    .B(_2555_));
 sg13g2_xor2_1 _3586_ (.B(_2723_),
    .A(_2556_),
    .X(_2724_));
 sg13g2_inv_1 _3587_ (.Y(_2725_),
    .A(_2724_));
 sg13g2_nor2_1 _3588_ (.A(_2702_),
    .B(_2725_),
    .Y(_2726_));
 sg13g2_nand3_1 _3589_ (.B(_2720_),
    .C(_2726_),
    .A(_2714_),
    .Y(_2727_));
 sg13g2_nand4_1 _3590_ (.B(_2719_),
    .C(_2717_),
    .A(_2716_),
    .Y(_2728_),
    .D(_2727_));
 sg13g2_nand2_1 _3591_ (.Y(_0091_),
    .A(_2712_),
    .B(_2728_));
 sg13g2_a21o_1 _3592_ (.A2(_2728_),
    .A1(_2712_),
    .B1(_2725_),
    .X(_0092_));
 sg13g2_a221oi_1 _3593_ (.B2(_2728_),
    .C1(_2725_),
    .B1(_2712_),
    .A1(_2562_),
    .Y(_0093_),
    .A2(_2709_));
 sg13g2_or3_1 _3594_ (.A(_2702_),
    .B(_2713_),
    .C(_0093_),
    .X(_0094_));
 sg13g2_o21ai_1 _3595_ (.B1(_2702_),
    .Y(_0095_),
    .A1(_2713_),
    .A2(_0093_));
 sg13g2_and2_1 _3596_ (.A(_0094_),
    .B(_0095_),
    .X(_0096_));
 sg13g2_nand3_1 _3597_ (.B(_2725_),
    .C(_2728_),
    .A(_2712_),
    .Y(_0097_));
 sg13g2_nand2_1 _3598_ (.Y(_0098_),
    .A(_0092_),
    .B(_0097_));
 sg13g2_nand2_1 _3599_ (.Y(_0099_),
    .A(net371),
    .B(_2553_));
 sg13g2_xor2_1 _3600_ (.B(_0099_),
    .A(_2554_),
    .X(_0100_));
 sg13g2_nor2_1 _3601_ (.A(_2721_),
    .B(_0100_),
    .Y(_0101_));
 sg13g2_nor2_1 _3602_ (.A(_0098_),
    .B(_0100_),
    .Y(_0102_));
 sg13g2_nand3_1 _3603_ (.B(_0097_),
    .C(_0101_),
    .A(_0092_),
    .Y(_0103_));
 sg13g2_a22oi_1 _3604_ (.Y(_0104_),
    .B1(_2712_),
    .B2(_2728_),
    .A2(_2726_),
    .A1(_2722_));
 sg13g2_nand2_1 _3605_ (.Y(_0105_),
    .A(_2718_),
    .B(_0104_));
 sg13g2_xor2_1 _3606_ (.B(_0104_),
    .A(_2718_),
    .X(_0106_));
 sg13g2_xnor2_1 _3607_ (.Y(_0107_),
    .A(_2718_),
    .B(_0104_));
 sg13g2_and4_1 _3608_ (.A(_0094_),
    .B(_0095_),
    .C(_0103_),
    .D(_0106_),
    .X(_0108_));
 sg13g2_nand4_1 _3609_ (.B(_0095_),
    .C(_0103_),
    .A(_0094_),
    .Y(_0109_),
    .D(_0106_));
 sg13g2_xnor2_1 _3610_ (.Y(_0110_),
    .A(_2719_),
    .B(_0105_));
 sg13g2_xor2_1 _3611_ (.B(_0105_),
    .A(_2719_),
    .X(_0111_));
 sg13g2_nand2_2 _3612_ (.Y(_0112_),
    .A(_0109_),
    .B(_0111_));
 sg13g2_nand3_1 _3613_ (.B(_0103_),
    .C(_0112_),
    .A(_0096_),
    .Y(_0113_));
 sg13g2_a21oi_2 _3614_ (.B1(_0108_),
    .Y(_0114_),
    .A2(_0113_),
    .A1(_0107_));
 sg13g2_a21o_1 _3615_ (.A2(_0112_),
    .A1(_0103_),
    .B1(_0096_),
    .X(_0115_));
 sg13g2_and2_1 _3616_ (.A(_0113_),
    .B(_0115_),
    .X(_0116_));
 sg13g2_a21oi_1 _3617_ (.A1(_0109_),
    .A2(_0111_),
    .Y(_0117_),
    .B1(_0100_));
 sg13g2_and3_1 _3618_ (.X(_0118_),
    .A(_0100_),
    .B(_0109_),
    .C(_0111_));
 sg13g2_nor2_1 _3619_ (.A(_0117_),
    .B(_0118_),
    .Y(_0119_));
 sg13g2_nand2_1 _3620_ (.Y(_0120_),
    .A(net371),
    .B(_2551_));
 sg13g2_xor2_1 _3621_ (.B(_0120_),
    .A(_2552_),
    .X(_0121_));
 sg13g2_xnor2_1 _3622_ (.Y(_0122_),
    .A(_2552_),
    .B(_0120_));
 sg13g2_nand2_1 _3623_ (.Y(_0123_),
    .A(_0119_),
    .B(_0121_));
 sg13g2_o21ai_1 _3624_ (.B1(_0102_),
    .Y(_0124_),
    .A1(_0108_),
    .A2(_0110_));
 sg13g2_xor2_1 _3625_ (.B(_0117_),
    .A(_0098_),
    .X(_0125_));
 sg13g2_or4_1 _3626_ (.A(_0098_),
    .B(_0117_),
    .C(_0118_),
    .D(_0122_),
    .X(_0126_));
 sg13g2_nand3_1 _3627_ (.B(_0092_),
    .C(_0124_),
    .A(_2722_),
    .Y(_0127_));
 sg13g2_a21o_1 _3628_ (.A2(_0124_),
    .A1(_0092_),
    .B1(_2722_),
    .X(_0128_));
 sg13g2_and2_1 _3629_ (.A(_0127_),
    .B(_0128_),
    .X(_0129_));
 sg13g2_nand2_1 _3630_ (.Y(_0130_),
    .A(_0126_),
    .B(_0129_));
 sg13g2_and4_1 _3631_ (.A(_0107_),
    .B(_0126_),
    .C(_0127_),
    .D(_0128_),
    .X(_0131_));
 sg13g2_a21oi_2 _3632_ (.B1(_0114_),
    .Y(_0132_),
    .A2(_0131_),
    .A1(_0116_));
 sg13g2_nand3_1 _3633_ (.B(_0126_),
    .C(_0129_),
    .A(_0114_),
    .Y(_0133_));
 sg13g2_nand2b_1 _3634_ (.Y(_0134_),
    .B(_0116_),
    .A_N(_0131_));
 sg13g2_nor2_1 _3635_ (.A(_2482_),
    .B(net372),
    .Y(_0135_));
 sg13g2_xor2_1 _3636_ (.B(_2484_),
    .A(_2483_),
    .X(_0136_));
 sg13g2_xnor2_1 _3637_ (.Y(_0137_),
    .A(_0135_),
    .B(_0136_));
 sg13g2_nand3_1 _3638_ (.B(_0121_),
    .C(_0137_),
    .A(_0119_),
    .Y(_0138_));
 sg13g2_nand4_1 _3639_ (.B(_0129_),
    .C(_0132_),
    .A(_0125_),
    .Y(_0139_),
    .D(_0138_));
 sg13g2_a21o_1 _3640_ (.A2(_0125_),
    .A1(_0123_),
    .B1(_0129_),
    .X(_0140_));
 sg13g2_nand3_1 _3641_ (.B(_0122_),
    .C(_0137_),
    .A(_0119_),
    .Y(_0141_));
 sg13g2_nand4_1 _3642_ (.B(_0130_),
    .C(_0140_),
    .A(_0114_),
    .Y(_0142_),
    .D(_0141_));
 sg13g2_and4_2 _3643_ (.A(_0133_),
    .B(_0134_),
    .C(_0139_),
    .D(_0142_),
    .X(_0143_));
 sg13g2_a21oi_1 _3644_ (.A1(_0132_),
    .A2(_0143_),
    .Y(_0144_),
    .B1(net373));
 sg13g2_a21o_1 _3645_ (.A2(_0112_),
    .A1(_2544_),
    .B1(_0144_),
    .X(_0145_));
 sg13g2_a21oi_1 _3646_ (.A1(_2544_),
    .A2(_0091_),
    .Y(_0146_),
    .B1(_0145_));
 sg13g2_o21ai_1 _3647_ (.B1(_0146_),
    .Y(_0147_),
    .A1(net373),
    .A2(_2709_));
 sg13g2_nor2_1 _3648_ (.A(net373),
    .B(_2696_),
    .Y(_0148_));
 sg13g2_or2_1 _3649_ (.X(_0149_),
    .B(_0148_),
    .A(_0147_));
 sg13g2_a21o_1 _3650_ (.A2(_2675_),
    .A1(net371),
    .B1(_0149_),
    .X(_0150_));
 sg13g2_nor2_1 _3651_ (.A(_2656_),
    .B(_0150_),
    .Y(_0151_));
 sg13g2_nor2_1 _3652_ (.A(net373),
    .B(_0151_),
    .Y(_0152_));
 sg13g2_a21o_1 _3653_ (.A2(_0151_),
    .A1(_2639_),
    .B1(net372),
    .X(_0153_));
 sg13g2_o21ai_1 _3654_ (.B1(_0153_),
    .Y(_0154_),
    .A1(net372),
    .A2(_2619_));
 sg13g2_a21o_2 _3655_ (.A2(_2605_),
    .A1(net371),
    .B1(_0154_),
    .X(_0155_));
 sg13g2_nor2_2 _3656_ (.A(_0020_),
    .B(net473),
    .Y(_0156_));
 sg13g2_inv_2 _3657_ (.Y(_0157_),
    .A(_0156_));
 sg13g2_and3_1 _3658_ (.X(_0158_),
    .A(net431),
    .B(net420),
    .C(net418));
 sg13g2_o21ai_1 _3659_ (.B1(net431),
    .Y(_0159_),
    .A1(net420),
    .A2(net418));
 sg13g2_nor2_1 _3660_ (.A(_0158_),
    .B(_0159_),
    .Y(_0160_));
 sg13g2_xnor2_1 _3661_ (.Y(_0161_),
    .A(_0157_),
    .B(_0160_));
 sg13g2_nand3_1 _3662_ (.B(net407),
    .C(net402),
    .A(net432),
    .Y(_0162_));
 sg13g2_nand2_2 _3663_ (.Y(_0163_),
    .A(net432),
    .B(net412));
 sg13g2_o21ai_1 _3664_ (.B1(net432),
    .Y(_0164_),
    .A1(net406),
    .A2(net402));
 sg13g2_nand2b_1 _3665_ (.Y(_0165_),
    .B(_0162_),
    .A_N(_0164_));
 sg13g2_o21ai_1 _3666_ (.B1(_0162_),
    .Y(_0166_),
    .A1(_0163_),
    .A2(_0164_));
 sg13g2_a21o_2 _3667_ (.A2(_0160_),
    .A1(_0156_),
    .B1(_0158_),
    .X(_0167_));
 sg13g2_xor2_1 _3668_ (.B(_0166_),
    .A(_0161_),
    .X(_0168_));
 sg13g2_and2_1 _3669_ (.A(_0167_),
    .B(_0168_),
    .X(_0169_));
 sg13g2_a21o_2 _3670_ (.A2(_0166_),
    .A1(_0161_),
    .B1(_0169_),
    .X(_0170_));
 sg13g2_inv_1 _3671_ (.Y(_0171_),
    .A(_0170_));
 sg13g2_nor2_1 _3672_ (.A(net436),
    .B(net389),
    .Y(_0172_));
 sg13g2_nand3_1 _3673_ (.B(net393),
    .C(_0172_),
    .A(\pid.Kp[5] ),
    .Y(_0173_));
 sg13g2_nand2_1 _3674_ (.Y(_0174_),
    .A(net435),
    .B(net399));
 sg13g2_a21o_1 _3675_ (.A2(net393),
    .A1(\pid.Kp[5] ),
    .B1(_0172_),
    .X(_0175_));
 sg13g2_and2_1 _3676_ (.A(_0173_),
    .B(_0175_),
    .X(_0176_));
 sg13g2_nand2b_1 _3677_ (.Y(_0177_),
    .B(_0176_),
    .A_N(_0174_));
 sg13g2_nand2_1 _3678_ (.Y(_0178_),
    .A(_0173_),
    .B(_0177_));
 sg13g2_nand2_1 _3679_ (.Y(_0179_),
    .A(net433),
    .B(net399));
 sg13g2_nand2_1 _3680_ (.Y(_0180_),
    .A(net435),
    .B(net393));
 sg13g2_nor2_1 _3681_ (.A(\pid.Kp[5] ),
    .B(net389),
    .Y(_0181_));
 sg13g2_nand2b_1 _3682_ (.Y(_0182_),
    .B(_0181_),
    .A_N(_0180_));
 sg13g2_xnor2_1 _3683_ (.Y(_0183_),
    .A(_0180_),
    .B(_0181_));
 sg13g2_nand2b_1 _3684_ (.Y(_0184_),
    .B(_0183_),
    .A_N(_0179_));
 sg13g2_xnor2_1 _3685_ (.Y(_0185_),
    .A(_0179_),
    .B(_0183_));
 sg13g2_nand2_1 _3686_ (.Y(_0186_),
    .A(_0178_),
    .B(_0185_));
 sg13g2_xnor2_1 _3687_ (.Y(_0187_),
    .A(_0178_),
    .B(_0185_));
 sg13g2_xor2_1 _3688_ (.B(_0165_),
    .A(_0163_),
    .X(_0188_));
 sg13g2_inv_1 _3689_ (.Y(_0189_),
    .A(_0188_));
 sg13g2_o21ai_1 _3690_ (.B1(_0186_),
    .Y(_0190_),
    .A1(_0187_),
    .A2(_0189_));
 sg13g2_nand2_1 _3691_ (.Y(_0191_),
    .A(_0182_),
    .B(_0184_));
 sg13g2_and2_1 _3692_ (.A(net431),
    .B(net398),
    .X(_0192_));
 sg13g2_nand2_1 _3693_ (.Y(_0193_),
    .A(net431),
    .B(net399));
 sg13g2_nand2_1 _3694_ (.Y(_0194_),
    .A(net433),
    .B(net393));
 sg13g2_nor2_1 _3695_ (.A(net435),
    .B(net389),
    .Y(_0195_));
 sg13g2_nor2b_1 _3696_ (.A(_0194_),
    .B_N(_0195_),
    .Y(_0196_));
 sg13g2_xnor2_1 _3697_ (.Y(_0197_),
    .A(_0194_),
    .B(_0195_));
 sg13g2_xnor2_1 _3698_ (.Y(_0198_),
    .A(_0193_),
    .B(_0197_));
 sg13g2_nand2_1 _3699_ (.Y(_0199_),
    .A(_0191_),
    .B(_0198_));
 sg13g2_xnor2_1 _3700_ (.Y(_0200_),
    .A(_0191_),
    .B(_0198_));
 sg13g2_xnor2_1 _3701_ (.Y(_0201_),
    .A(_0189_),
    .B(_0200_));
 sg13g2_nand2b_1 _3702_ (.Y(_0202_),
    .B(_0190_),
    .A_N(_0201_));
 sg13g2_xnor2_1 _3703_ (.Y(_0203_),
    .A(_0167_),
    .B(_0168_));
 sg13g2_xor2_1 _3704_ (.B(_0201_),
    .A(_0190_),
    .X(_0204_));
 sg13g2_o21ai_1 _3705_ (.B1(_0202_),
    .Y(_0205_),
    .A1(_0203_),
    .A2(_0204_));
 sg13g2_o21ai_1 _3706_ (.B1(_0199_),
    .Y(_0206_),
    .A1(_0189_),
    .A2(_0200_));
 sg13g2_a21oi_1 _3707_ (.A1(_0192_),
    .A2(_0197_),
    .Y(_0207_),
    .B1(_0196_));
 sg13g2_nor2_2 _3708_ (.A(_0020_),
    .B(_2036_),
    .Y(_0208_));
 sg13g2_and3_1 _3709_ (.X(_0209_),
    .A(_0021_),
    .B(net391),
    .C(_0208_));
 sg13g2_a21oi_1 _3710_ (.A1(_0021_),
    .A2(net391),
    .Y(_0210_),
    .B1(_0208_));
 sg13g2_nor2_1 _3711_ (.A(_0209_),
    .B(_0210_),
    .Y(_0211_));
 sg13g2_xnor2_1 _3712_ (.Y(_0212_),
    .A(_0193_),
    .B(_0211_));
 sg13g2_nor2b_1 _3713_ (.A(_0207_),
    .B_N(_0212_),
    .Y(_0213_));
 sg13g2_xnor2_1 _3714_ (.Y(_0214_),
    .A(_0207_),
    .B(_0212_));
 sg13g2_xnor2_1 _3715_ (.Y(_0215_),
    .A(_0188_),
    .B(_0214_));
 sg13g2_nand2b_1 _3716_ (.Y(_0216_),
    .B(_0206_),
    .A_N(_0215_));
 sg13g2_xnor2_1 _3717_ (.Y(_0217_),
    .A(_0206_),
    .B(_0215_));
 sg13g2_inv_1 _3718_ (.Y(_0218_),
    .A(_0217_));
 sg13g2_xnor2_1 _3719_ (.Y(_0219_),
    .A(_0203_),
    .B(_0217_));
 sg13g2_nand2_1 _3720_ (.Y(_0220_),
    .A(_0205_),
    .B(_0219_));
 sg13g2_xnor2_1 _3721_ (.Y(_0221_),
    .A(_0205_),
    .B(_0219_));
 sg13g2_xnor2_1 _3722_ (.Y(_0222_),
    .A(_0171_),
    .B(_0221_));
 sg13g2_nor2_1 _3723_ (.A(net438),
    .B(net389),
    .Y(_0223_));
 sg13g2_nand3_1 _3724_ (.B(net392),
    .C(_0223_),
    .A(net436),
    .Y(_0224_));
 sg13g2_nand2_1 _3725_ (.Y(_0225_),
    .A(\pid.Kp[5] ),
    .B(net398));
 sg13g2_a21o_1 _3726_ (.A2(net392),
    .A1(net436),
    .B1(_0223_),
    .X(_0226_));
 sg13g2_and2_1 _3727_ (.A(_0224_),
    .B(_0226_),
    .X(_0227_));
 sg13g2_nand2b_1 _3728_ (.Y(_0228_),
    .B(_0227_),
    .A_N(_0225_));
 sg13g2_nand2_1 _3729_ (.Y(_0229_),
    .A(_0224_),
    .B(_0228_));
 sg13g2_xnor2_1 _3730_ (.Y(_0230_),
    .A(_0174_),
    .B(_0176_));
 sg13g2_nand2_1 _3731_ (.Y(_0231_),
    .A(_0229_),
    .B(_0230_));
 sg13g2_nor2_1 _3732_ (.A(_0854_),
    .B(_0162_),
    .Y(_0232_));
 sg13g2_or2_1 _3733_ (.X(_0233_),
    .B(_0162_),
    .A(_0854_));
 sg13g2_a22oi_1 _3734_ (.Y(_0234_),
    .B1(net402),
    .B2(net434),
    .A2(net407),
    .A1(net431));
 sg13g2_nor2_1 _3735_ (.A(_0232_),
    .B(_0234_),
    .Y(_0235_));
 sg13g2_xnor2_1 _3736_ (.Y(_0236_),
    .A(_0163_),
    .B(_0235_));
 sg13g2_inv_1 _3737_ (.Y(_0237_),
    .A(_0236_));
 sg13g2_xnor2_1 _3738_ (.Y(_0238_),
    .A(_0229_),
    .B(_0230_));
 sg13g2_o21ai_1 _3739_ (.B1(_0231_),
    .Y(_0239_),
    .A1(_0237_),
    .A2(_0238_));
 sg13g2_xnor2_1 _3740_ (.Y(_0240_),
    .A(_0187_),
    .B(_0188_));
 sg13g2_nand2_1 _3741_ (.Y(_0241_),
    .A(_0239_),
    .B(_0240_));
 sg13g2_o21ai_1 _3742_ (.B1(_0233_),
    .Y(_0242_),
    .A1(_0163_),
    .A2(_0234_));
 sg13g2_nand2_1 _3743_ (.Y(_0243_),
    .A(net396),
    .B(_0242_));
 sg13g2_xnor2_1 _3744_ (.Y(_0244_),
    .A(net396),
    .B(_0242_));
 sg13g2_nand2b_1 _3745_ (.Y(_0245_),
    .B(_0167_),
    .A_N(_0244_));
 sg13g2_xor2_1 _3746_ (.B(_0244_),
    .A(_0167_),
    .X(_0246_));
 sg13g2_xnor2_1 _3747_ (.Y(_0247_),
    .A(_0239_),
    .B(_0240_));
 sg13g2_o21ai_1 _3748_ (.B1(_0241_),
    .Y(_0248_),
    .A1(_0246_),
    .A2(_0247_));
 sg13g2_xor2_1 _3749_ (.B(_0204_),
    .A(_0203_),
    .X(_0249_));
 sg13g2_nand2_1 _3750_ (.Y(_0250_),
    .A(_0243_),
    .B(_0245_));
 sg13g2_xnor2_1 _3751_ (.Y(_0251_),
    .A(_0248_),
    .B(_0249_));
 sg13g2_nor2b_1 _3752_ (.A(_0251_),
    .B_N(_0250_),
    .Y(_0252_));
 sg13g2_a21oi_2 _3753_ (.B1(_0252_),
    .Y(_0253_),
    .A2(_0249_),
    .A1(_0248_));
 sg13g2_nor2_1 _3754_ (.A(_0222_),
    .B(_0253_),
    .Y(_0254_));
 sg13g2_o21ai_1 _3755_ (.B1(_0220_),
    .Y(_0255_),
    .A1(_0171_),
    .A2(_0221_));
 sg13g2_o21ai_1 _3756_ (.B1(_0216_),
    .Y(_0256_),
    .A1(_0203_),
    .A2(_0218_));
 sg13g2_a21oi_2 _3757_ (.B1(_0213_),
    .Y(_0257_),
    .A2(_0214_),
    .A1(_0188_));
 sg13g2_a21oi_1 _3758_ (.A1(_0192_),
    .A2(_0211_),
    .Y(_0258_),
    .B1(_0209_));
 sg13g2_nand2_1 _3759_ (.Y(_0259_),
    .A(net393),
    .B(_0192_));
 sg13g2_nor2_1 _3760_ (.A(net431),
    .B(net389),
    .Y(_0260_));
 sg13g2_o21ai_1 _3761_ (.B1(net431),
    .Y(_0261_),
    .A1(net399),
    .A2(net393));
 sg13g2_nand2b_1 _3762_ (.Y(_0262_),
    .B(_0261_),
    .A_N(_0260_));
 sg13g2_nand3_1 _3763_ (.B(_0259_),
    .C(_0262_),
    .A(_0188_),
    .Y(_0263_));
 sg13g2_inv_1 _3764_ (.Y(_0264_),
    .A(_0263_));
 sg13g2_a21oi_1 _3765_ (.A1(_0259_),
    .A2(_0262_),
    .Y(_0265_),
    .B1(_0188_));
 sg13g2_inv_1 _3766_ (.Y(_0266_),
    .A(_0265_));
 sg13g2_nand2_1 _3767_ (.Y(_0267_),
    .A(_0263_),
    .B(_0266_));
 sg13g2_xnor2_1 _3768_ (.Y(_0268_),
    .A(_0258_),
    .B(_0267_));
 sg13g2_xnor2_1 _3769_ (.Y(_0269_),
    .A(_0257_),
    .B(_0268_));
 sg13g2_xor2_1 _3770_ (.B(_0269_),
    .A(_0203_),
    .X(_0270_));
 sg13g2_and2_1 _3771_ (.A(_0256_),
    .B(_0270_),
    .X(_0271_));
 sg13g2_xor2_1 _3772_ (.B(_0270_),
    .A(_0256_),
    .X(_0272_));
 sg13g2_xnor2_1 _3773_ (.Y(_0273_),
    .A(_0170_),
    .B(_0272_));
 sg13g2_nand2b_1 _3774_ (.Y(_0274_),
    .B(_0255_),
    .A_N(_0273_));
 sg13g2_xor2_1 _3775_ (.B(_0273_),
    .A(_0255_),
    .X(_0275_));
 sg13g2_nor3_2 _3776_ (.A(_0222_),
    .B(_0253_),
    .C(_0275_),
    .Y(_0276_));
 sg13g2_inv_1 _3777_ (.Y(_0277_),
    .A(_0276_));
 sg13g2_xor2_1 _3778_ (.B(_0275_),
    .A(_0254_),
    .X(_0278_));
 sg13g2_inv_1 _3779_ (.Y(_0279_),
    .A(_0278_));
 sg13g2_xor2_1 _3780_ (.B(_0251_),
    .A(_0250_),
    .X(_0280_));
 sg13g2_nor2_1 _3781_ (.A(net439),
    .B(net389),
    .Y(_0281_));
 sg13g2_nand3_1 _3782_ (.B(net392),
    .C(_0281_),
    .A(net438),
    .Y(_0282_));
 sg13g2_nand2_1 _3783_ (.Y(_0283_),
    .A(net436),
    .B(net398));
 sg13g2_a21o_1 _3784_ (.A2(net392),
    .A1(net438),
    .B1(_0281_),
    .X(_0284_));
 sg13g2_and2_1 _3785_ (.A(_0282_),
    .B(_0284_),
    .X(_0285_));
 sg13g2_nand2b_1 _3786_ (.Y(_0286_),
    .B(_0285_),
    .A_N(_0283_));
 sg13g2_nand2_1 _3787_ (.Y(_0287_),
    .A(_0282_),
    .B(_0286_));
 sg13g2_xnor2_1 _3788_ (.Y(_0288_),
    .A(_0225_),
    .B(_0227_));
 sg13g2_nand2_1 _3789_ (.Y(_0289_),
    .A(_0287_),
    .B(_0288_));
 sg13g2_nand2_1 _3790_ (.Y(_0290_),
    .A(net433),
    .B(net407));
 sg13g2_nand2b_2 _3791_ (.Y(_0291_),
    .B(net403),
    .A_N(_0022_));
 sg13g2_xor2_1 _3792_ (.B(_0291_),
    .A(_0290_),
    .X(_0292_));
 sg13g2_nand2b_1 _3793_ (.Y(_0293_),
    .B(_0292_),
    .A_N(_0163_));
 sg13g2_xnor2_1 _3794_ (.Y(_0294_),
    .A(_0163_),
    .B(_0292_));
 sg13g2_inv_1 _3795_ (.Y(_0295_),
    .A(_0294_));
 sg13g2_xnor2_1 _3796_ (.Y(_0296_),
    .A(_0287_),
    .B(_0288_));
 sg13g2_o21ai_1 _3797_ (.B1(_0289_),
    .Y(_0297_),
    .A1(_0295_),
    .A2(_0296_));
 sg13g2_xnor2_1 _3798_ (.Y(_0298_),
    .A(_0237_),
    .B(_0238_));
 sg13g2_nand2b_1 _3799_ (.Y(_0299_),
    .B(_0297_),
    .A_N(_0298_));
 sg13g2_o21ai_1 _3800_ (.B1(_0293_),
    .Y(_0300_),
    .A1(_0290_),
    .A2(_0291_));
 sg13g2_nand2_1 _3801_ (.Y(_0301_),
    .A(net396),
    .B(_0300_));
 sg13g2_xnor2_1 _3802_ (.Y(_0302_),
    .A(net396),
    .B(_0300_));
 sg13g2_nand2b_1 _3803_ (.Y(_0303_),
    .B(_0167_),
    .A_N(_0302_));
 sg13g2_xor2_1 _3804_ (.B(_0302_),
    .A(_0167_),
    .X(_0304_));
 sg13g2_xor2_1 _3805_ (.B(_0298_),
    .A(_0297_),
    .X(_0305_));
 sg13g2_o21ai_1 _3806_ (.B1(_0299_),
    .Y(_0306_),
    .A1(_0304_),
    .A2(_0305_));
 sg13g2_xor2_1 _3807_ (.B(_0247_),
    .A(_0246_),
    .X(_0307_));
 sg13g2_nand2_1 _3808_ (.Y(_0308_),
    .A(_0301_),
    .B(_0303_));
 sg13g2_xnor2_1 _3809_ (.Y(_0309_),
    .A(_0306_),
    .B(_0307_));
 sg13g2_nor2b_1 _3810_ (.A(_0309_),
    .B_N(_0308_),
    .Y(_0310_));
 sg13g2_a21oi_2 _3811_ (.B1(_0310_),
    .Y(_0311_),
    .A2(_0307_),
    .A1(_0306_));
 sg13g2_nor2_1 _3812_ (.A(_0280_),
    .B(_0311_),
    .Y(_0312_));
 sg13g2_xnor2_1 _3813_ (.Y(_0313_),
    .A(_0222_),
    .B(_0253_));
 sg13g2_or3_1 _3814_ (.A(_0280_),
    .B(_0311_),
    .C(_0313_),
    .X(_0314_));
 sg13g2_inv_1 _3815_ (.Y(_0315_),
    .A(_0314_));
 sg13g2_xnor2_1 _3816_ (.Y(_0316_),
    .A(_0280_),
    .B(_0311_));
 sg13g2_xor2_1 _3817_ (.B(_0309_),
    .A(_0308_),
    .X(_0317_));
 sg13g2_nor2_1 _3818_ (.A(net440),
    .B(net389),
    .Y(_0318_));
 sg13g2_nand2_1 _3819_ (.Y(_0319_),
    .A(net439),
    .B(net392));
 sg13g2_nand3_1 _3820_ (.B(net392),
    .C(_0318_),
    .A(net439),
    .Y(_0320_));
 sg13g2_nand2_1 _3821_ (.Y(_0321_),
    .A(net438),
    .B(net398));
 sg13g2_xnor2_1 _3822_ (.Y(_0322_),
    .A(_0318_),
    .B(_0319_));
 sg13g2_nand2b_1 _3823_ (.Y(_0323_),
    .B(_0322_),
    .A_N(_0321_));
 sg13g2_nand2_1 _3824_ (.Y(_0324_),
    .A(_0320_),
    .B(_0323_));
 sg13g2_xnor2_1 _3825_ (.Y(_0325_),
    .A(_0283_),
    .B(_0285_));
 sg13g2_nand2_1 _3826_ (.Y(_0326_),
    .A(_0324_),
    .B(_0325_));
 sg13g2_nand2_1 _3827_ (.Y(_0327_),
    .A(net433),
    .B(net412));
 sg13g2_and2_1 _3828_ (.A(\pid.Kp[5] ),
    .B(net402),
    .X(_0328_));
 sg13g2_nand3_1 _3829_ (.B(net406),
    .C(_0328_),
    .A(net435),
    .Y(_0329_));
 sg13g2_a21o_1 _3830_ (.A2(net406),
    .A1(net435),
    .B1(_0328_),
    .X(_0330_));
 sg13g2_nand2_1 _3831_ (.Y(_0331_),
    .A(_0329_),
    .B(_0330_));
 sg13g2_xor2_1 _3832_ (.B(_0331_),
    .A(_0327_),
    .X(_0332_));
 sg13g2_inv_1 _3833_ (.Y(_0333_),
    .A(_0332_));
 sg13g2_xnor2_1 _3834_ (.Y(_0334_),
    .A(_0324_),
    .B(_0325_));
 sg13g2_o21ai_1 _3835_ (.B1(_0326_),
    .Y(_0335_),
    .A1(_0333_),
    .A2(_0334_));
 sg13g2_xnor2_1 _3836_ (.Y(_0336_),
    .A(_0295_),
    .B(_0296_));
 sg13g2_nand2b_1 _3837_ (.Y(_0337_),
    .B(_0335_),
    .A_N(_0336_));
 sg13g2_o21ai_1 _3838_ (.B1(_0329_),
    .Y(_0338_),
    .A1(_0327_),
    .A2(_0331_));
 sg13g2_nand2_1 _3839_ (.Y(_0339_),
    .A(net396),
    .B(_0338_));
 sg13g2_xnor2_1 _3840_ (.Y(_0340_),
    .A(net396),
    .B(_0338_));
 sg13g2_nand2b_1 _3841_ (.Y(_0341_),
    .B(_0167_),
    .A_N(_0340_));
 sg13g2_xor2_1 _3842_ (.B(_0340_),
    .A(_0167_),
    .X(_0342_));
 sg13g2_xor2_1 _3843_ (.B(_0336_),
    .A(_0335_),
    .X(_0343_));
 sg13g2_o21ai_1 _3844_ (.B1(_0337_),
    .Y(_0344_),
    .A1(_0342_),
    .A2(_0343_));
 sg13g2_xor2_1 _3845_ (.B(_0305_),
    .A(_0304_),
    .X(_0345_));
 sg13g2_nand2_1 _3846_ (.Y(_0346_),
    .A(_0339_),
    .B(_0341_));
 sg13g2_xnor2_1 _3847_ (.Y(_0347_),
    .A(_0344_),
    .B(_0345_));
 sg13g2_nor2b_1 _3848_ (.A(_0347_),
    .B_N(_0346_),
    .Y(_0348_));
 sg13g2_a21oi_1 _3849_ (.A1(_0344_),
    .A2(_0345_),
    .Y(_0349_),
    .B1(_0348_));
 sg13g2_nor2_1 _3850_ (.A(_0317_),
    .B(_0349_),
    .Y(_0350_));
 sg13g2_nor2b_1 _3851_ (.A(_0316_),
    .B_N(_0350_),
    .Y(_0351_));
 sg13g2_inv_1 _3852_ (.Y(_0352_),
    .A(_0351_));
 sg13g2_xnor2_1 _3853_ (.Y(_0353_),
    .A(_0316_),
    .B(_0350_));
 sg13g2_inv_1 _3854_ (.Y(_0354_),
    .A(_0353_));
 sg13g2_xor2_1 _3855_ (.B(_0347_),
    .A(_0346_),
    .X(_0355_));
 sg13g2_nand3_1 _3856_ (.B(net60),
    .C(net53),
    .A(net440),
    .Y(_0356_));
 sg13g2_nor3_2 _3857_ (.A(\pid.Kp[0] ),
    .B(_2030_),
    .C(_2032_),
    .Y(_0357_));
 sg13g2_nand2b_1 _3858_ (.Y(_0358_),
    .B(_0357_),
    .A_N(_0356_));
 sg13g2_nand2_1 _3859_ (.Y(_0359_),
    .A(net439),
    .B(net400));
 sg13g2_a21oi_1 _3860_ (.A1(\pid.Kp[1] ),
    .A2(net394),
    .Y(_0360_),
    .B1(_0357_));
 sg13g2_xnor2_1 _3861_ (.Y(_0361_),
    .A(_0356_),
    .B(_0357_));
 sg13g2_o21ai_1 _3862_ (.B1(_0358_),
    .Y(_0362_),
    .A1(_0360_),
    .A2(_0359_));
 sg13g2_xnor2_1 _3863_ (.Y(_0363_),
    .A(_0321_),
    .B(_0322_));
 sg13g2_nand2_1 _3864_ (.Y(_0364_),
    .A(net78),
    .B(_0363_));
 sg13g2_nand2_2 _3865_ (.Y(_0365_),
    .A(net435),
    .B(net412));
 sg13g2_and2_1 _3866_ (.A(net436),
    .B(net406),
    .X(_0366_));
 sg13g2_nand2_1 _3867_ (.Y(_0367_),
    .A(net436),
    .B(net406));
 sg13g2_nand2_1 _3868_ (.Y(_0368_),
    .A(_0328_),
    .B(_0366_));
 sg13g2_a22oi_1 _3869_ (.Y(_0369_),
    .B1(net402),
    .B2(net436),
    .A2(net406),
    .A1(\pid.Kp[5] ));
 sg13g2_a21oi_1 _3870_ (.A1(_0328_),
    .A2(_0366_),
    .Y(_0370_),
    .B1(_0369_));
 sg13g2_xnor2_1 _3871_ (.Y(_0371_),
    .A(_0365_),
    .B(_0370_));
 sg13g2_inv_1 _3872_ (.Y(_0372_),
    .A(_0371_));
 sg13g2_xnor2_1 _3873_ (.Y(_0373_),
    .A(net78),
    .B(_0363_));
 sg13g2_o21ai_1 _3874_ (.B1(_0364_),
    .Y(_0374_),
    .A1(_0372_),
    .A2(_0373_));
 sg13g2_xnor2_1 _3875_ (.Y(_0375_),
    .A(_0333_),
    .B(_0334_));
 sg13g2_nand2b_1 _3876_ (.Y(_0376_),
    .B(_0374_),
    .A_N(_0375_));
 sg13g2_nand2_1 _3877_ (.Y(_0377_),
    .A(net433),
    .B(_0158_));
 sg13g2_a22oi_1 _3878_ (.Y(_0378_),
    .B1(net418),
    .B2(net433),
    .A2(net420),
    .A1(net431));
 sg13g2_a21oi_1 _3879_ (.A1(net433),
    .A2(_0158_),
    .Y(_0379_),
    .B1(_0378_));
 sg13g2_o21ai_1 _3880_ (.B1(_0377_),
    .Y(_0380_),
    .A1(_0157_),
    .A2(_0378_));
 sg13g2_inv_1 _3881_ (.Y(_0381_),
    .A(_0380_));
 sg13g2_o21ai_1 _3882_ (.B1(_0368_),
    .Y(_0382_),
    .A1(_0365_),
    .A2(_0369_));
 sg13g2_nand2_1 _3883_ (.Y(_0383_),
    .A(net396),
    .B(_0382_));
 sg13g2_xnor2_1 _3884_ (.Y(_0384_),
    .A(net396),
    .B(_0382_));
 sg13g2_xnor2_1 _3885_ (.Y(_0385_),
    .A(_0381_),
    .B(_0384_));
 sg13g2_xor2_1 _3886_ (.B(_0375_),
    .A(_0374_),
    .X(_0386_));
 sg13g2_o21ai_1 _3887_ (.B1(_0376_),
    .Y(_0387_),
    .A1(_0385_),
    .A2(_0386_));
 sg13g2_xor2_1 _3888_ (.B(_0343_),
    .A(_0342_),
    .X(_0388_));
 sg13g2_o21ai_1 _3889_ (.B1(_0383_),
    .Y(_0389_),
    .A1(_0381_),
    .A2(_0384_));
 sg13g2_xnor2_1 _3890_ (.Y(_0390_),
    .A(_0387_),
    .B(_0388_));
 sg13g2_nor2b_1 _3891_ (.A(_0390_),
    .B_N(_0389_),
    .Y(_0391_));
 sg13g2_a21oi_1 _3892_ (.A1(_0387_),
    .A2(_0388_),
    .Y(_0392_),
    .B1(_0391_));
 sg13g2_nor2_1 _3893_ (.A(_0355_),
    .B(_0392_),
    .Y(_0393_));
 sg13g2_xor2_1 _3894_ (.B(_0349_),
    .A(_0317_),
    .X(_0394_));
 sg13g2_or2_1 _3895_ (.X(_0395_),
    .B(_0394_),
    .A(_0393_));
 sg13g2_inv_1 _3896_ (.Y(_0396_),
    .A(_0395_));
 sg13g2_nand2_1 _3897_ (.Y(_0397_),
    .A(net441),
    .B(net398));
 sg13g2_and3_1 _3898_ (.X(_0398_),
    .A(net440),
    .B(net441),
    .C(net392));
 sg13g2_nand2_1 _3899_ (.Y(_0399_),
    .A(net398),
    .B(_0398_));
 sg13g2_xnor2_1 _3900_ (.Y(_0400_),
    .A(_0359_),
    .B(_0361_));
 sg13g2_nor2b_1 _3901_ (.A(_0399_),
    .B_N(_0400_),
    .Y(_0401_));
 sg13g2_nand2b_1 _3902_ (.Y(_0402_),
    .B(net402),
    .A_N(_0023_));
 sg13g2_xnor2_1 _3903_ (.Y(_0403_),
    .A(net391),
    .B(_0402_));
 sg13g2_nand2_1 _3904_ (.Y(_0404_),
    .A(_0366_),
    .B(_0403_));
 sg13g2_xnor2_1 _3905_ (.Y(_0405_),
    .A(_0367_),
    .B(_0403_));
 sg13g2_xnor2_1 _3906_ (.Y(_0406_),
    .A(_0399_),
    .B(_0400_));
 sg13g2_a21oi_1 _3907_ (.A1(_0405_),
    .A2(net71),
    .Y(_0407_),
    .B1(_0401_));
 sg13g2_xnor2_1 _3908_ (.Y(_0408_),
    .A(_0372_),
    .B(_0373_));
 sg13g2_nor2_1 _3909_ (.A(_0407_),
    .B(_0408_),
    .Y(_0409_));
 sg13g2_nor3_1 _3910_ (.A(_0024_),
    .B(net416),
    .C(_0365_),
    .Y(_0410_));
 sg13g2_nand2_1 _3911_ (.Y(_0411_),
    .A(net433),
    .B(net420));
 sg13g2_a22oi_1 _3912_ (.Y(_0412_),
    .B1(net412),
    .B2(_0865_),
    .A2(net418),
    .A1(net435));
 sg13g2_or2_1 _3913_ (.X(_0413_),
    .B(_0412_),
    .A(_0410_));
 sg13g2_nor2_1 _3914_ (.A(_0411_),
    .B(_0413_),
    .Y(_0414_));
 sg13g2_nor2_1 _3915_ (.A(_0410_),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_o21ai_1 _3916_ (.B1(_0404_),
    .Y(_0416_),
    .A1(net389),
    .A2(_0402_));
 sg13g2_xnor2_1 _3917_ (.Y(_0417_),
    .A(_0156_),
    .B(_0379_));
 sg13g2_nand2b_1 _3918_ (.Y(_0418_),
    .B(_0416_),
    .A_N(_0417_));
 sg13g2_xor2_1 _3919_ (.B(_0417_),
    .A(_0416_),
    .X(_0419_));
 sg13g2_xor2_1 _3920_ (.B(_0419_),
    .A(_0415_),
    .X(_0420_));
 sg13g2_xor2_1 _3921_ (.B(_0407_),
    .A(_0408_),
    .X(_0421_));
 sg13g2_a21oi_1 _3922_ (.A1(_0420_),
    .A2(_0421_),
    .Y(_0422_),
    .B1(_0409_));
 sg13g2_xor2_1 _3923_ (.B(_0386_),
    .A(_0385_),
    .X(_0423_));
 sg13g2_nor2b_1 _3924_ (.A(_0422_),
    .B_N(_0423_),
    .Y(_0424_));
 sg13g2_o21ai_1 _3925_ (.B1(_0418_),
    .Y(_0425_),
    .A1(_0415_),
    .A2(_0419_));
 sg13g2_xnor2_1 _3926_ (.Y(_0426_),
    .A(_0422_),
    .B(_0423_));
 sg13g2_a21oi_1 _3927_ (.A1(_0425_),
    .A2(_0426_),
    .Y(_0427_),
    .B1(_0424_));
 sg13g2_xor2_1 _3928_ (.B(_0390_),
    .A(_0389_),
    .X(_0428_));
 sg13g2_nor2_1 _3929_ (.A(_0427_),
    .B(_0428_),
    .Y(_0429_));
 sg13g2_inv_1 _3930_ (.Y(_0430_),
    .A(_0429_));
 sg13g2_xnor2_1 _3931_ (.Y(_0431_),
    .A(_0355_),
    .B(_0392_));
 sg13g2_nor2_1 _3932_ (.A(_0430_),
    .B(_0431_),
    .Y(_0432_));
 sg13g2_xor2_1 _3933_ (.B(_0428_),
    .A(_0427_),
    .X(_0433_));
 sg13g2_nand2_2 _3934_ (.Y(_0434_),
    .A(net439),
    .B(net402));
 sg13g2_nand2_1 _3935_ (.Y(_0435_),
    .A(net438),
    .B(net406));
 sg13g2_xor2_1 _3936_ (.B(_0435_),
    .A(_0434_),
    .X(_0436_));
 sg13g2_nand3_1 _3937_ (.B(net412),
    .C(net437),
    .A(_0436_),
    .Y(_0437_));
 sg13g2_a21o_1 _3938_ (.A2(net412),
    .A1(net436),
    .B1(_0436_),
    .X(_0438_));
 sg13g2_and2_1 _3939_ (.A(_0438_),
    .B(_0437_),
    .X(_0439_));
 sg13g2_a22oi_1 _3940_ (.Y(_0440_),
    .B1(net392),
    .B2(net441),
    .A2(net398),
    .A1(net440));
 sg13g2_a21oi_1 _3941_ (.A1(net398),
    .A2(_0398_),
    .Y(_0441_),
    .B1(_0440_));
 sg13g2_nand2_1 _3942_ (.Y(_0442_),
    .A(_0439_),
    .B(_0441_));
 sg13g2_xnor2_1 _3943_ (.Y(_0443_),
    .A(_0405_),
    .B(_0406_));
 sg13g2_nor2_1 _3944_ (.A(_0442_),
    .B(net70),
    .Y(_0444_));
 sg13g2_nand2_1 _3945_ (.Y(_0445_),
    .A(\pid.Kp[6] ),
    .B(net420));
 sg13g2_nor3_1 _3946_ (.A(_0024_),
    .B(net416),
    .C(_0445_),
    .Y(_0446_));
 sg13g2_nor2_1 _3947_ (.A(_0021_),
    .B(net473),
    .Y(_0447_));
 sg13g2_o21ai_1 _3948_ (.B1(_0445_),
    .Y(_0448_),
    .A1(_0024_),
    .A2(net416));
 sg13g2_nor2b_1 _3949_ (.A(_0446_),
    .B_N(_0448_),
    .Y(_0449_));
 sg13g2_a21oi_2 _3950_ (.B1(_0446_),
    .Y(_0450_),
    .A2(_0448_),
    .A1(_0447_));
 sg13g2_o21ai_1 _3951_ (.B1(_0437_),
    .Y(_0451_),
    .A1(_0434_),
    .A2(_0435_));
 sg13g2_xor2_1 _3952_ (.B(_0413_),
    .A(_0411_),
    .X(_0452_));
 sg13g2_xnor2_1 _3953_ (.Y(_0453_),
    .A(_0452_),
    .B(_0451_));
 sg13g2_nor2_1 _3954_ (.A(_0450_),
    .B(_0453_),
    .Y(_0454_));
 sg13g2_xor2_1 _3955_ (.B(_0450_),
    .A(_0453_),
    .X(_0455_));
 sg13g2_xor2_1 _3956_ (.B(_0442_),
    .A(_0443_),
    .X(_0456_));
 sg13g2_a21oi_1 _3957_ (.A1(net42),
    .A2(net68),
    .Y(_0457_),
    .B1(_0444_));
 sg13g2_xnor2_1 _3958_ (.Y(_0458_),
    .A(_0420_),
    .B(_0421_));
 sg13g2_a21oi_2 _3959_ (.B1(_0454_),
    .Y(_0459_),
    .A2(_0452_),
    .A1(_0451_));
 sg13g2_xor2_1 _3960_ (.B(_0458_),
    .A(_0457_),
    .X(_0460_));
 sg13g2_nand2b_1 _3961_ (.Y(_0461_),
    .B(_0460_),
    .A_N(_0459_));
 sg13g2_o21ai_1 _3962_ (.B1(_0461_),
    .Y(_0462_),
    .A1(_0457_),
    .A2(_0458_));
 sg13g2_xnor2_1 _3963_ (.Y(_0463_),
    .A(_0425_),
    .B(_0426_));
 sg13g2_nor2b_1 _3964_ (.A(_0463_),
    .B_N(_0462_),
    .Y(_0464_));
 sg13g2_nand2_1 _3965_ (.Y(_0465_),
    .A(_0433_),
    .B(_0464_));
 sg13g2_nand2_2 _3966_ (.Y(_0466_),
    .A(net440),
    .B(net407));
 sg13g2_nand2_1 _3967_ (.Y(_0467_),
    .A(net440),
    .B(net402));
 sg13g2_nand2_1 _3968_ (.Y(_0468_),
    .A(net439),
    .B(net406));
 sg13g2_xor2_1 _3969_ (.B(_0468_),
    .A(_0467_),
    .X(_0469_));
 sg13g2_nand3_1 _3970_ (.B(net412),
    .C(net438),
    .A(_0469_),
    .Y(_0470_));
 sg13g2_a21o_1 _3971_ (.A2(net412),
    .A1(net438),
    .B1(_0469_),
    .X(_0471_));
 sg13g2_and2_1 _3972_ (.A(_0470_),
    .B(_0471_),
    .X(_0472_));
 sg13g2_nand2b_1 _3973_ (.Y(_0473_),
    .B(_0472_),
    .A_N(_0397_));
 sg13g2_xnor2_1 _3974_ (.Y(_0474_),
    .A(_0439_),
    .B(_0441_));
 sg13g2_nor2_1 _3975_ (.A(_0473_),
    .B(_0474_),
    .Y(_0475_));
 sg13g2_xor2_1 _3976_ (.B(_0473_),
    .A(_0474_),
    .X(_0476_));
 sg13g2_nand2_1 _3977_ (.Y(_0477_),
    .A(\pid.Kp[5] ),
    .B(net420));
 sg13g2_nor3_1 _3978_ (.A(_0025_),
    .B(net416),
    .C(_0477_),
    .Y(_0478_));
 sg13g2_o21ai_1 _3979_ (.B1(_0477_),
    .Y(_0479_),
    .A1(_0025_),
    .A2(net416));
 sg13g2_nand2b_1 _3980_ (.Y(_0480_),
    .B(_0479_),
    .A_N(_0478_));
 sg13g2_nor3_1 _3981_ (.A(_0022_),
    .B(net473),
    .C(_0480_),
    .Y(_0481_));
 sg13g2_nor2_1 _3982_ (.A(_0478_),
    .B(_0481_),
    .Y(_0482_));
 sg13g2_o21ai_1 _3983_ (.B1(_0470_),
    .Y(_0483_),
    .A1(_0434_),
    .A2(_0466_));
 sg13g2_xnor2_1 _3984_ (.Y(_0484_),
    .A(_0447_),
    .B(_0449_));
 sg13g2_nand2b_1 _3985_ (.Y(_0485_),
    .B(_0483_),
    .A_N(_0484_));
 sg13g2_xor2_1 _3986_ (.B(_0483_),
    .A(_0484_),
    .X(_0486_));
 sg13g2_xor2_1 _3987_ (.B(_0486_),
    .A(_0482_),
    .X(_0487_));
 sg13g2_a21oi_1 _3988_ (.A1(_0476_),
    .A2(_0487_),
    .Y(_0488_),
    .B1(_0475_));
 sg13g2_xnor2_1 _3989_ (.Y(_0489_),
    .A(_0455_),
    .B(_0456_));
 sg13g2_o21ai_1 _3990_ (.B1(_0485_),
    .Y(_0490_),
    .A1(_0482_),
    .A2(net59));
 sg13g2_xor2_1 _3991_ (.B(_0489_),
    .A(_0488_),
    .X(_0491_));
 sg13g2_nand2_1 _3992_ (.Y(_0492_),
    .A(_0490_),
    .B(net49));
 sg13g2_o21ai_1 _3993_ (.B1(_0492_),
    .Y(_0493_),
    .A1(_0488_),
    .A2(_0489_));
 sg13g2_xor2_1 _3994_ (.B(_0460_),
    .A(_0459_),
    .X(_0494_));
 sg13g2_nor2b_1 _3995_ (.A(_0494_),
    .B_N(_0493_),
    .Y(_0495_));
 sg13g2_xnor2_1 _3996_ (.Y(_0496_),
    .A(_0462_),
    .B(_0463_));
 sg13g2_and2_1 _3997_ (.A(_0495_),
    .B(_0496_),
    .X(_0497_));
 sg13g2_xnor2_1 _3998_ (.Y(_0498_),
    .A(_0397_),
    .B(_0472_));
 sg13g2_nand2_1 _3999_ (.Y(_0499_),
    .A(net437),
    .B(net420));
 sg13g2_nor3_1 _4000_ (.A(_0023_),
    .B(net416),
    .C(_0499_),
    .Y(_0500_));
 sg13g2_nor2_1 _4001_ (.A(_0024_),
    .B(net473),
    .Y(_0501_));
 sg13g2_o21ai_1 _4002_ (.B1(_0499_),
    .Y(_0502_),
    .A1(_0023_),
    .A2(net416));
 sg13g2_nor2b_1 _4003_ (.A(_0500_),
    .B_N(_0502_),
    .Y(_0503_));
 sg13g2_a21o_1 _4004_ (.A2(_0502_),
    .A1(_0501_),
    .B1(_0500_),
    .X(_0504_));
 sg13g2_nand2_1 _4005_ (.Y(_0505_),
    .A(net441),
    .B(net403));
 sg13g2_nand2_1 _4006_ (.Y(_0506_),
    .A(net439),
    .B(net413));
 sg13g2_xor2_1 _4007_ (.B(_0505_),
    .A(_0466_),
    .X(_0507_));
 sg13g2_nand2b_1 _4008_ (.Y(_0508_),
    .B(_0507_),
    .A_N(_0506_));
 sg13g2_o21ai_1 _4009_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_0466_),
    .A2(_0505_));
 sg13g2_o21ai_1 _4010_ (.B1(_0480_),
    .Y(_0510_),
    .A1(_0022_),
    .A2(net473));
 sg13g2_nand2b_1 _4011_ (.Y(_0511_),
    .B(_0510_),
    .A_N(_0481_));
 sg13g2_nor2b_1 _4012_ (.A(_0511_),
    .B_N(_0509_),
    .Y(_0512_));
 sg13g2_xor2_1 _4013_ (.B(_0511_),
    .A(_0509_),
    .X(_0513_));
 sg13g2_nor2b_1 _4014_ (.A(_0513_),
    .B_N(_0504_),
    .Y(_0514_));
 sg13g2_xnor2_1 _4015_ (.Y(_0515_),
    .A(_0504_),
    .B(_0513_));
 sg13g2_nand2_1 _4016_ (.Y(_0516_),
    .A(_0498_),
    .B(_0515_));
 sg13g2_xnor2_1 _4017_ (.Y(_0517_),
    .A(_0487_),
    .B(_0476_));
 sg13g2_nor2_1 _4018_ (.A(_0512_),
    .B(_0514_),
    .Y(_0518_));
 sg13g2_xor2_1 _4019_ (.B(_0516_),
    .A(_0517_),
    .X(_0519_));
 sg13g2_nand2b_1 _4020_ (.Y(_0520_),
    .B(_0519_),
    .A_N(_0518_));
 sg13g2_o21ai_1 _4021_ (.B1(_0520_),
    .Y(_0521_),
    .A1(_0516_),
    .A2(_0517_));
 sg13g2_xnor2_1 _4022_ (.Y(_0522_),
    .A(_0490_),
    .B(_0491_));
 sg13g2_nand2b_1 _4023_ (.Y(_0523_),
    .B(_0521_),
    .A_N(_0522_));
 sg13g2_xor2_1 _4024_ (.B(_0521_),
    .A(_0522_),
    .X(_0524_));
 sg13g2_o21ai_1 _4025_ (.B1(_0523_),
    .Y(_0525_),
    .A1(net41),
    .A2(_0157_));
 sg13g2_xnor2_1 _4026_ (.Y(_0526_),
    .A(_0493_),
    .B(_0494_));
 sg13g2_nand2_1 _4027_ (.Y(_0527_),
    .A(_0525_),
    .B(_0526_));
 sg13g2_xnor2_1 _4028_ (.Y(_0528_),
    .A(_0518_),
    .B(net47));
 sg13g2_xnor2_1 _4029_ (.Y(_0529_),
    .A(_0498_),
    .B(_0515_));
 sg13g2_nand2_1 _4030_ (.Y(_0530_),
    .A(\pid.Kp[3] ),
    .B(net421));
 sg13g2_nor3_1 _4031_ (.A(_0026_),
    .B(net417),
    .C(_0530_),
    .Y(_0531_));
 sg13g2_nor2_1 _4032_ (.A(_0025_),
    .B(net473),
    .Y(_0532_));
 sg13g2_o21ai_1 _4033_ (.B1(_0530_),
    .Y(_0533_),
    .A1(_0026_),
    .A2(net417));
 sg13g2_nor2b_1 _4034_ (.A(_0531_),
    .B_N(_0533_),
    .Y(_0534_));
 sg13g2_a21o_1 _4035_ (.A2(_0533_),
    .A1(_0532_),
    .B1(_0531_),
    .X(_0535_));
 sg13g2_nand2_2 _4036_ (.Y(_0536_),
    .A(\pid.Kp[0] ),
    .B(net413));
 sg13g2_nor2_1 _4037_ (.A(_0466_),
    .B(_0536_),
    .Y(_0537_));
 sg13g2_xor2_1 _4038_ (.B(_0503_),
    .A(_0501_),
    .X(_0538_));
 sg13g2_xnor2_1 _4039_ (.Y(_0539_),
    .A(_0537_),
    .B(_0538_));
 sg13g2_nor2b_1 _4040_ (.A(_0539_),
    .B_N(_0535_),
    .Y(_0540_));
 sg13g2_xnor2_1 _4041_ (.Y(_0541_),
    .A(_0535_),
    .B(_0539_));
 sg13g2_xnor2_1 _4042_ (.Y(_0542_),
    .A(_0506_),
    .B(_0507_));
 sg13g2_nand2_1 _4043_ (.Y(_0543_),
    .A(_0541_),
    .B(_0542_));
 sg13g2_nor2_1 _4044_ (.A(_0529_),
    .B(_0543_),
    .Y(_0544_));
 sg13g2_a21oi_1 _4045_ (.A1(_0537_),
    .A2(_0538_),
    .Y(_0545_),
    .B1(_0540_));
 sg13g2_xor2_1 _4046_ (.B(_0543_),
    .A(_0529_),
    .X(_0546_));
 sg13g2_nor2b_1 _4047_ (.A(_0545_),
    .B_N(_0546_),
    .Y(_0547_));
 sg13g2_nor2_1 _4048_ (.A(_0544_),
    .B(_0547_),
    .Y(_0548_));
 sg13g2_nand2b_1 _4049_ (.Y(_0549_),
    .B(_0528_),
    .A_N(_0548_));
 sg13g2_xnor2_1 _4050_ (.Y(_0550_),
    .A(_0157_),
    .B(_0524_));
 sg13g2_nor2_1 _4051_ (.A(_0549_),
    .B(_0550_),
    .Y(_0551_));
 sg13g2_xnor2_1 _4052_ (.Y(_0552_),
    .A(_0528_),
    .B(_0548_));
 sg13g2_a22oi_1 _4053_ (.Y(_0553_),
    .B1(net407),
    .B2(net441),
    .A2(net413),
    .A1(net440));
 sg13g2_nor2_1 _4054_ (.A(_0537_),
    .B(_0553_),
    .Y(_0554_));
 sg13g2_nand2_1 _4055_ (.Y(_0555_),
    .A(\pid.Kp[2] ),
    .B(net421));
 sg13g2_nor2_1 _4056_ (.A(_0027_),
    .B(net417),
    .Y(_0556_));
 sg13g2_nand2b_1 _4057_ (.Y(_0557_),
    .B(_0556_),
    .A_N(_0555_));
 sg13g2_nor2_1 _4058_ (.A(_0023_),
    .B(net473),
    .Y(_0558_));
 sg13g2_xnor2_1 _4059_ (.Y(_0559_),
    .A(_0555_),
    .B(_0556_));
 sg13g2_nand2_1 _4060_ (.Y(_0560_),
    .A(_0558_),
    .B(_0559_));
 sg13g2_xnor2_1 _4061_ (.Y(_0561_),
    .A(_0532_),
    .B(_0534_));
 sg13g2_a21oi_2 _4062_ (.B1(_0561_),
    .Y(_0562_),
    .A2(_0560_),
    .A1(_0557_));
 sg13g2_nand3_1 _4063_ (.B(_0560_),
    .C(_0561_),
    .A(_0557_),
    .Y(_0563_));
 sg13g2_nor2b_1 _4064_ (.A(_0562_),
    .B_N(_0563_),
    .Y(_0564_));
 sg13g2_nand2_1 _4065_ (.Y(_0565_),
    .A(_0554_),
    .B(_0564_));
 sg13g2_xor2_1 _4066_ (.B(_0542_),
    .A(_0541_),
    .X(_0566_));
 sg13g2_nor2b_1 _4067_ (.A(_0565_),
    .B_N(_0566_),
    .Y(_0567_));
 sg13g2_xnor2_1 _4068_ (.Y(_0568_),
    .A(_0565_),
    .B(_0566_));
 sg13g2_a21oi_1 _4069_ (.A1(_0562_),
    .A2(_0568_),
    .Y(_0569_),
    .B1(_0567_));
 sg13g2_xnor2_1 _4070_ (.Y(_0570_),
    .A(_0545_),
    .B(_0546_));
 sg13g2_nor2b_1 _4071_ (.A(_0569_),
    .B_N(_0570_),
    .Y(_0571_));
 sg13g2_xnor2_1 _4072_ (.Y(_0572_),
    .A(_0569_),
    .B(_0570_));
 sg13g2_nand2_1 _4073_ (.Y(_0573_),
    .A(\pid.Kp[1] ),
    .B(net421));
 sg13g2_nor2_1 _4074_ (.A(_0028_),
    .B(net417),
    .Y(_0574_));
 sg13g2_nand2b_1 _4075_ (.Y(_0575_),
    .B(_0574_),
    .A_N(_0573_));
 sg13g2_nor2_1 _4076_ (.A(_0026_),
    .B(net473),
    .Y(_0576_));
 sg13g2_xnor2_1 _4077_ (.Y(_0577_),
    .A(_0573_),
    .B(_0574_));
 sg13g2_nand2_1 _4078_ (.Y(_0578_),
    .A(_0576_),
    .B(_0577_));
 sg13g2_xnor2_1 _4079_ (.Y(_0579_),
    .A(_0558_),
    .B(_0559_));
 sg13g2_a21oi_2 _4080_ (.B1(_0579_),
    .Y(_0580_),
    .A2(_0578_),
    .A1(_0575_));
 sg13g2_nand3_1 _4081_ (.B(_0578_),
    .C(_0579_),
    .A(_0575_),
    .Y(_0581_));
 sg13g2_nor2b_1 _4082_ (.A(_0580_),
    .B_N(_0581_),
    .Y(_0582_));
 sg13g2_nor2b_1 _4083_ (.A(_0536_),
    .B_N(_0582_),
    .Y(_0583_));
 sg13g2_xor2_1 _4084_ (.B(_0564_),
    .A(_0554_),
    .X(_0584_));
 sg13g2_xnor2_1 _4085_ (.Y(_0585_),
    .A(_0583_),
    .B(_0584_));
 sg13g2_o21ai_1 _4086_ (.B1(_0584_),
    .Y(_0586_),
    .A1(_0580_),
    .A2(_0583_));
 sg13g2_xnor2_1 _4087_ (.Y(_0587_),
    .A(_0562_),
    .B(_0568_));
 sg13g2_nor2_1 _4088_ (.A(_0586_),
    .B(_0587_),
    .Y(_0588_));
 sg13g2_nor2_1 _4089_ (.A(_0027_),
    .B(net471),
    .Y(_0589_));
 sg13g2_nand3_1 _4090_ (.B(net422),
    .C(_0589_),
    .A(net441),
    .Y(_0590_));
 sg13g2_xnor2_1 _4091_ (.Y(_0591_),
    .A(_0576_),
    .B(_0577_));
 sg13g2_nor2_1 _4092_ (.A(_0590_),
    .B(_0591_),
    .Y(_0592_));
 sg13g2_xnor2_1 _4093_ (.Y(_0593_),
    .A(_0536_),
    .B(_0582_));
 sg13g2_nand2_1 _4094_ (.Y(_0594_),
    .A(_0592_),
    .B(_0593_));
 sg13g2_xor2_1 _4095_ (.B(_0585_),
    .A(_0580_),
    .X(_0595_));
 sg13g2_nor2_1 _4096_ (.A(_0594_),
    .B(_0595_),
    .Y(_0596_));
 sg13g2_nand2_1 _4097_ (.Y(_0597_),
    .A(_0586_),
    .B(_0587_));
 sg13g2_nand2b_1 _4098_ (.Y(_0598_),
    .B(_0597_),
    .A_N(_0588_));
 sg13g2_a21oi_1 _4099_ (.A1(_0596_),
    .A2(_0597_),
    .Y(_0599_),
    .B1(_0588_));
 sg13g2_nor2b_1 _4100_ (.A(_0599_),
    .B_N(_0572_),
    .Y(_0600_));
 sg13g2_xnor2_1 _4101_ (.Y(_0601_),
    .A(_0552_),
    .B(_0571_));
 sg13g2_o21ai_1 _4102_ (.B1(_0552_),
    .Y(_0602_),
    .A1(_0571_),
    .A2(_0600_));
 sg13g2_inv_1 _4103_ (.Y(_0603_),
    .A(_0602_));
 sg13g2_xor2_1 _4104_ (.B(_0549_),
    .A(_0550_),
    .X(_0604_));
 sg13g2_a21oi_2 _4105_ (.B1(_0551_),
    .Y(_0605_),
    .A2(_0604_),
    .A1(_0603_));
 sg13g2_xnor2_1 _4106_ (.Y(_0606_),
    .A(_0526_),
    .B(_0525_));
 sg13g2_o21ai_1 _4107_ (.B1(_0527_),
    .Y(_0607_),
    .A1(_0606_),
    .A2(_0605_));
 sg13g2_xnor2_1 _4108_ (.Y(_0608_),
    .A(_0495_),
    .B(_0496_));
 sg13g2_inv_1 _4109_ (.Y(_0609_),
    .A(_0608_));
 sg13g2_a21oi_2 _4110_ (.B1(_0497_),
    .Y(_0610_),
    .A2(_0607_),
    .A1(_0609_));
 sg13g2_xnor2_1 _4111_ (.Y(_0611_),
    .A(_0433_),
    .B(_0464_));
 sg13g2_o21ai_1 _4112_ (.B1(_0465_),
    .Y(_0612_),
    .A1(_0611_),
    .A2(_0610_));
 sg13g2_xnor2_1 _4113_ (.Y(_0613_),
    .A(_0430_),
    .B(_0431_));
 sg13g2_inv_1 _4114_ (.Y(_0614_),
    .A(_0613_));
 sg13g2_a21o_1 _4115_ (.A2(_0614_),
    .A1(_0612_),
    .B1(_0432_),
    .X(_0615_));
 sg13g2_xor2_1 _4116_ (.B(_0394_),
    .A(_0393_),
    .X(_0616_));
 sg13g2_a221oi_1 _4117_ (.B2(_0612_),
    .C1(_0432_),
    .B1(_0614_),
    .A1(_0393_),
    .Y(_0617_),
    .A2(_0394_));
 sg13g2_nor3_2 _4118_ (.A(_0354_),
    .B(_0396_),
    .C(net45),
    .Y(_0618_));
 sg13g2_nand3b_1 _4119_ (.B(_0353_),
    .C(_0395_),
    .Y(_0619_),
    .A_N(_0617_));
 sg13g2_xor2_1 _4120_ (.B(_0313_),
    .A(_0312_),
    .X(_0620_));
 sg13g2_inv_1 _4121_ (.Y(_0621_),
    .A(_0620_));
 sg13g2_a21oi_2 _4122_ (.B1(_0620_),
    .Y(_0622_),
    .A2(_0619_),
    .A1(_0352_));
 sg13g2_o21ai_1 _4123_ (.B1(_0621_),
    .Y(_0623_),
    .A1(_0351_),
    .A2(_0618_));
 sg13g2_a21oi_2 _4124_ (.B1(_0278_),
    .Y(_0624_),
    .A2(_0623_),
    .A1(_0314_));
 sg13g2_o21ai_1 _4125_ (.B1(_0279_),
    .Y(_0625_),
    .A1(_0622_),
    .A2(_0315_));
 sg13g2_a21oi_1 _4126_ (.A1(_0170_),
    .A2(_0272_),
    .Y(_0626_),
    .B1(_0271_));
 sg13g2_a21oi_1 _4127_ (.A1(_0257_),
    .A2(_0268_),
    .Y(_0627_),
    .B1(_0203_));
 sg13g2_o21ai_1 _4128_ (.B1(_0203_),
    .Y(_0628_),
    .A1(_0257_),
    .A2(_0268_));
 sg13g2_nand2b_1 _4129_ (.Y(_0629_),
    .B(_0628_),
    .A_N(_0627_));
 sg13g2_a21oi_1 _4130_ (.A1(_0258_),
    .A2(_0266_),
    .Y(_0630_),
    .B1(_0264_));
 sg13g2_a22oi_1 _4131_ (.Y(_0631_),
    .B1(_0208_),
    .B2(_0260_),
    .A2(_0192_),
    .A1(net393));
 sg13g2_xnor2_1 _4132_ (.Y(_0632_),
    .A(_0170_),
    .B(_0631_));
 sg13g2_xnor2_1 _4133_ (.Y(_0633_),
    .A(_0630_),
    .B(_0632_));
 sg13g2_xnor2_1 _4134_ (.Y(_0634_),
    .A(_0629_),
    .B(_0633_));
 sg13g2_xnor2_1 _4135_ (.Y(_0635_),
    .A(_0626_),
    .B(_0634_));
 sg13g2_xnor2_1 _4136_ (.Y(_0636_),
    .A(_0274_),
    .B(_0635_));
 sg13g2_inv_1 _4137_ (.Y(_0637_),
    .A(_0636_));
 sg13g2_a21oi_2 _4138_ (.B1(_0636_),
    .Y(_0638_),
    .A2(_0277_),
    .A1(_0625_));
 sg13g2_o21ai_1 _4139_ (.B1(_0637_),
    .Y(_0639_),
    .A1(_0276_),
    .A2(_0624_));
 sg13g2_nor3_2 _4140_ (.A(_0276_),
    .B(_0637_),
    .C(_0624_),
    .Y(_0640_));
 sg13g2_nand3_1 _4141_ (.B(_0625_),
    .C(_0636_),
    .A(_0277_),
    .Y(_0641_));
 sg13g2_nor2_1 _4142_ (.A(_0638_),
    .B(_0640_),
    .Y(_0642_));
 sg13g2_inv_4 _4143_ (.A(net375),
    .Y(_0643_));
 sg13g2_nor3_1 _4144_ (.A(_0351_),
    .B(_0618_),
    .C(_0621_),
    .Y(_0644_));
 sg13g2_nor2_1 _4145_ (.A(_0622_),
    .B(_0644_),
    .Y(_0645_));
 sg13g2_o21ai_1 _4146_ (.B1(_0354_),
    .Y(_0646_),
    .A1(_0396_),
    .A2(net39));
 sg13g2_and2_1 _4147_ (.A(_0619_),
    .B(_0646_),
    .X(_0647_));
 sg13g2_xnor2_1 _4148_ (.Y(_0648_),
    .A(net40),
    .B(_0613_));
 sg13g2_xnor2_1 _4149_ (.Y(_0649_),
    .A(_0610_),
    .B(_0611_));
 sg13g2_xnor2_1 _4150_ (.Y(_0650_),
    .A(_0596_),
    .B(_0598_));
 sg13g2_a21o_1 _4151_ (.A2(net422),
    .A1(net441),
    .B1(_0589_),
    .X(_0651_));
 sg13g2_and2_1 _4152_ (.A(_0590_),
    .B(_0651_),
    .X(_0652_));
 sg13g2_nor2_1 _4153_ (.A(_0028_),
    .B(net471),
    .Y(_0653_));
 sg13g2_or2_1 _4154_ (.X(_0654_),
    .B(_0653_),
    .A(_0652_));
 sg13g2_xor2_1 _4155_ (.B(_0591_),
    .A(_0590_),
    .X(_0655_));
 sg13g2_nor2_1 _4156_ (.A(_0654_),
    .B(_0655_),
    .Y(_0656_));
 sg13g2_xor2_1 _4157_ (.B(_0593_),
    .A(_0592_),
    .X(_0657_));
 sg13g2_nor2b_1 _4158_ (.A(_0657_),
    .B_N(_0656_),
    .Y(_0658_));
 sg13g2_xnor2_1 _4159_ (.Y(_0659_),
    .A(_0594_),
    .B(_0595_));
 sg13g2_nand2_1 _4160_ (.Y(_0660_),
    .A(_0658_),
    .B(_0659_));
 sg13g2_or2_1 _4161_ (.X(_0661_),
    .B(_0660_),
    .A(_0650_));
 sg13g2_xnor2_1 _4162_ (.Y(_0662_),
    .A(_0572_),
    .B(_0599_));
 sg13g2_nand2_1 _4163_ (.Y(_0663_),
    .A(_0643_),
    .B(_0661_));
 sg13g2_xor2_1 _4164_ (.B(_0663_),
    .A(_0662_),
    .X(_0664_));
 sg13g2_inv_1 _4165_ (.Y(_0665_),
    .A(_0664_));
 sg13g2_nor2_1 _4166_ (.A(_0661_),
    .B(_0662_),
    .Y(_0666_));
 sg13g2_xnor2_1 _4167_ (.Y(_0667_),
    .A(_0600_),
    .B(_0601_));
 sg13g2_nor2_1 _4168_ (.A(net376),
    .B(_0666_),
    .Y(_0668_));
 sg13g2_xnor2_1 _4169_ (.Y(_0669_),
    .A(_0667_),
    .B(_0668_));
 sg13g2_inv_1 _4170_ (.Y(_0670_),
    .A(_0669_));
 sg13g2_nand2b_1 _4171_ (.Y(_0671_),
    .B(_0666_),
    .A_N(_0667_));
 sg13g2_xnor2_1 _4172_ (.Y(_0672_),
    .A(_0602_),
    .B(net57));
 sg13g2_or2_1 _4173_ (.X(_0673_),
    .B(_0672_),
    .A(_0671_));
 sg13g2_xor2_1 _4174_ (.B(_0606_),
    .A(_0605_),
    .X(_0674_));
 sg13g2_nand2_1 _4175_ (.Y(_0675_),
    .A(_0643_),
    .B(_0671_));
 sg13g2_nor2b_1 _4176_ (.A(net376),
    .B_N(_0673_),
    .Y(_0676_));
 sg13g2_nand2_1 _4177_ (.Y(_0677_),
    .A(_0674_),
    .B(_0676_));
 sg13g2_or2_1 _4178_ (.X(_0678_),
    .B(_0676_),
    .A(_0674_));
 sg13g2_nand2_1 _4179_ (.Y(_0679_),
    .A(_0677_),
    .B(_0678_));
 sg13g2_inv_1 _4180_ (.Y(_0680_),
    .A(_0679_));
 sg13g2_xor2_1 _4181_ (.B(_0675_),
    .A(_0672_),
    .X(_0681_));
 sg13g2_nor2_1 _4182_ (.A(_0673_),
    .B(_0674_),
    .Y(_0682_));
 sg13g2_xnor2_1 _4183_ (.Y(_0683_),
    .A(net43),
    .B(_0608_));
 sg13g2_nor2b_1 _4184_ (.A(_0683_),
    .B_N(_0682_),
    .Y(_0684_));
 sg13g2_nand2_1 _4185_ (.Y(_0685_),
    .A(_0649_),
    .B(_0684_));
 sg13g2_nor2_1 _4186_ (.A(_0648_),
    .B(_0685_),
    .Y(_0686_));
 sg13g2_xnor2_1 _4187_ (.Y(_0687_),
    .A(_0615_),
    .B(_0616_));
 sg13g2_nand2_1 _4188_ (.Y(_0688_),
    .A(_0686_),
    .B(_0687_));
 sg13g2_nor2_1 _4189_ (.A(_0647_),
    .B(_0688_),
    .Y(_0689_));
 sg13g2_a21oi_1 _4190_ (.A1(_0639_),
    .A2(_0641_),
    .Y(_0690_),
    .B1(_0689_));
 sg13g2_xor2_1 _4191_ (.B(_0690_),
    .A(_0645_),
    .X(_0691_));
 sg13g2_o21ai_1 _4192_ (.B1(_0688_),
    .Y(_0692_),
    .A1(_0638_),
    .A2(_0640_));
 sg13g2_xor2_1 _4193_ (.B(_0692_),
    .A(_0647_),
    .X(_0693_));
 sg13g2_o21ai_1 _4194_ (.B1(_0685_),
    .Y(_0694_),
    .A1(_0640_),
    .A2(_0638_));
 sg13g2_xor2_1 _4195_ (.B(_0694_),
    .A(_0648_),
    .X(_0695_));
 sg13g2_a21oi_2 _4196_ (.B1(_0686_),
    .Y(_0696_),
    .A2(_0641_),
    .A1(_0639_));
 sg13g2_xnor2_1 _4197_ (.Y(_0697_),
    .A(_0687_),
    .B(_0696_));
 sg13g2_xor2_1 _4198_ (.B(_0696_),
    .A(_0687_),
    .X(_0698_));
 sg13g2_nand3_1 _4199_ (.B(_0693_),
    .C(_0698_),
    .A(_0695_),
    .Y(_0699_));
 sg13g2_nor3_1 _4200_ (.A(_0279_),
    .B(_0315_),
    .C(_0622_),
    .Y(_0700_));
 sg13g2_nor2_1 _4201_ (.A(_0624_),
    .B(_0700_),
    .Y(_0701_));
 sg13g2_nand2b_1 _4202_ (.Y(_0702_),
    .B(_0689_),
    .A_N(_0645_));
 sg13g2_o21ai_1 _4203_ (.B1(_0702_),
    .Y(_0703_),
    .A1(_0638_),
    .A2(_0640_));
 sg13g2_xnor2_1 _4204_ (.Y(_0704_),
    .A(_0701_),
    .B(_0703_));
 sg13g2_and2_1 _4205_ (.A(_0691_),
    .B(_0704_),
    .X(_0705_));
 sg13g2_nand2_1 _4206_ (.Y(_0706_),
    .A(_0699_),
    .B(_0705_));
 sg13g2_nor3_1 _4207_ (.A(net376),
    .B(_0701_),
    .C(_0702_),
    .Y(_0707_));
 sg13g2_or3_1 _4208_ (.A(net376),
    .B(_0701_),
    .C(_0702_),
    .X(_0708_));
 sg13g2_a21o_2 _4209_ (.A2(_0699_),
    .A1(_0705_),
    .B1(_0707_),
    .X(_0709_));
 sg13g2_and2_1 _4210_ (.A(_0695_),
    .B(_0709_),
    .X(_0710_));
 sg13g2_xor2_1 _4211_ (.B(_0709_),
    .A(_0695_),
    .X(_0711_));
 sg13g2_xnor2_1 _4212_ (.Y(_0712_),
    .A(_0695_),
    .B(_0709_));
 sg13g2_nor2_1 _4213_ (.A(net376),
    .B(_0684_),
    .Y(_0713_));
 sg13g2_xnor2_1 _4214_ (.Y(_0714_),
    .A(_0649_),
    .B(_0713_));
 sg13g2_and3_1 _4215_ (.X(_0715_),
    .A(_0695_),
    .B(_0698_),
    .C(_0709_));
 sg13g2_nor2_1 _4216_ (.A(_0693_),
    .B(_0715_),
    .Y(_0716_));
 sg13g2_nor2_1 _4217_ (.A(_0707_),
    .B(_0716_),
    .Y(_0717_));
 sg13g2_o21ai_1 _4218_ (.B1(_0708_),
    .Y(_0718_),
    .A1(_0715_),
    .A2(_0693_));
 sg13g2_nor2_1 _4219_ (.A(_0697_),
    .B(_0714_),
    .Y(_0719_));
 sg13g2_nand2_1 _4220_ (.Y(_0720_),
    .A(_0691_),
    .B(_0706_));
 sg13g2_a21oi_1 _4221_ (.A1(_0711_),
    .A2(_0719_),
    .Y(_0721_),
    .B1(_0720_));
 sg13g2_a22oi_1 _4222_ (.Y(_0722_),
    .B1(_0721_),
    .B2(_0718_),
    .A2(_0706_),
    .A1(_0704_));
 sg13g2_nor2_1 _4223_ (.A(_0714_),
    .B(_0722_),
    .Y(_0723_));
 sg13g2_xnor2_1 _4224_ (.Y(_0724_),
    .A(_0722_),
    .B(_0714_));
 sg13g2_nor2_1 _4225_ (.A(net376),
    .B(_0682_),
    .Y(_0725_));
 sg13g2_nand2_1 _4226_ (.Y(_0726_),
    .A(_0683_),
    .B(_0725_));
 sg13g2_or2_1 _4227_ (.X(_0727_),
    .B(_0725_),
    .A(_0683_));
 sg13g2_nand2_1 _4228_ (.Y(_0728_),
    .A(_0726_),
    .B(_0727_));
 sg13g2_inv_1 _4229_ (.Y(_0729_),
    .A(_0728_));
 sg13g2_a21oi_2 _4230_ (.B1(_0722_),
    .Y(_0730_),
    .A2(_0719_),
    .A1(_0711_));
 sg13g2_a22oi_1 _4231_ (.Y(_0731_),
    .B1(_0718_),
    .B2(_0730_),
    .A2(_0706_),
    .A1(_0691_));
 sg13g2_a21o_2 _4232_ (.A2(_0721_),
    .A1(_0718_),
    .B1(_0731_),
    .X(_0732_));
 sg13g2_nor3_1 _4233_ (.A(_0712_),
    .B(_0714_),
    .C(_0722_),
    .Y(_0733_));
 sg13g2_or3_1 _4234_ (.A(_0697_),
    .B(_0710_),
    .C(_0733_),
    .X(_0734_));
 sg13g2_o21ai_1 _4235_ (.B1(_0697_),
    .Y(_0735_),
    .A1(_0710_),
    .A2(_0733_));
 sg13g2_and2_1 _4236_ (.A(_0734_),
    .B(_0735_),
    .X(_0736_));
 sg13g2_xnor2_1 _4237_ (.Y(_0737_),
    .A(_0717_),
    .B(_0730_));
 sg13g2_nand2_1 _4238_ (.Y(_0738_),
    .A(_0711_),
    .B(_0728_));
 sg13g2_nor2_1 _4239_ (.A(_0724_),
    .B(_0738_),
    .Y(_0739_));
 sg13g2_or2_1 _4240_ (.X(_0740_),
    .B(_0724_),
    .A(_0738_));
 sg13g2_nand4_1 _4241_ (.B(_0735_),
    .C(_0737_),
    .A(_0740_),
    .Y(_0741_),
    .D(_0734_));
 sg13g2_and2_2 _4242_ (.A(_0732_),
    .B(_0741_),
    .X(_0742_));
 sg13g2_a21o_1 _4243_ (.A2(_0741_),
    .A1(_0732_),
    .B1(_0729_),
    .X(_0743_));
 sg13g2_a221oi_1 _4244_ (.B2(_0732_),
    .C1(_0724_),
    .B1(_0741_),
    .A1(_0726_),
    .Y(_0744_),
    .A2(_0727_));
 sg13g2_o21ai_1 _4245_ (.B1(_0712_),
    .Y(_0745_),
    .A1(_0723_),
    .A2(_0744_));
 sg13g2_or3_1 _4246_ (.A(_0712_),
    .B(_0744_),
    .C(_0723_),
    .X(_0746_));
 sg13g2_nand2_1 _4247_ (.Y(_0747_),
    .A(_0745_),
    .B(_0746_));
 sg13g2_nand3_1 _4248_ (.B(_0732_),
    .C(net44),
    .A(_0729_),
    .Y(_0748_));
 sg13g2_and2_1 _4249_ (.A(_0743_),
    .B(_0748_),
    .X(_0749_));
 sg13g2_inv_1 _4250_ (.Y(_0750_),
    .A(_0749_));
 sg13g2_nor2_1 _4251_ (.A(_0680_),
    .B(_0724_),
    .Y(_0751_));
 sg13g2_nand3_1 _4252_ (.B(_0748_),
    .C(_0751_),
    .A(_0743_),
    .Y(_0752_));
 sg13g2_inv_1 _4253_ (.Y(_0753_),
    .A(_0752_));
 sg13g2_a21oi_2 _4254_ (.B1(_0739_),
    .Y(_0754_),
    .A2(_0741_),
    .A1(_0732_));
 sg13g2_nand2_1 _4255_ (.Y(_0755_),
    .A(_0736_),
    .B(_0754_));
 sg13g2_xor2_1 _4256_ (.B(_0754_),
    .A(_0736_),
    .X(_0756_));
 sg13g2_nand4_1 _4257_ (.B(_0756_),
    .C(_0752_),
    .A(_0745_),
    .Y(_0757_),
    .D(_0746_));
 sg13g2_xor2_1 _4258_ (.B(_0755_),
    .A(_0737_),
    .X(_0758_));
 sg13g2_and2_2 _4259_ (.A(_0757_),
    .B(_0758_),
    .X(_0759_));
 sg13g2_nor2_1 _4260_ (.A(_0753_),
    .B(_0759_),
    .Y(_0760_));
 sg13g2_nor3_1 _4261_ (.A(_0747_),
    .B(_0753_),
    .C(_0759_),
    .Y(_0761_));
 sg13g2_xor2_1 _4262_ (.B(_0760_),
    .A(_0747_),
    .X(_0762_));
 sg13g2_a21o_1 _4263_ (.A2(_0758_),
    .A1(_0757_),
    .B1(_0680_),
    .X(_0763_));
 sg13g2_nand3_1 _4264_ (.B(_0757_),
    .C(_0758_),
    .A(_0680_),
    .Y(_0764_));
 sg13g2_and2_1 _4265_ (.A(_0763_),
    .B(_0764_),
    .X(_0765_));
 sg13g2_inv_1 _4266_ (.Y(_0766_),
    .A(_0765_));
 sg13g2_nand3_1 _4267_ (.B(_0763_),
    .C(_0764_),
    .A(_0749_),
    .Y(_0767_));
 sg13g2_xnor2_1 _4268_ (.Y(_0768_),
    .A(_0724_),
    .B(_0743_));
 sg13g2_a221oi_1 _4269_ (.B2(_0757_),
    .C1(_0750_),
    .B1(_0758_),
    .A1(_0677_),
    .Y(_0769_),
    .A2(_0678_));
 sg13g2_xnor2_1 _4270_ (.Y(_0770_),
    .A(_0769_),
    .B(_0768_));
 sg13g2_nand2b_1 _4271_ (.Y(_0771_),
    .B(_0768_),
    .A_N(_0681_));
 sg13g2_mux2_1 _4272_ (.A0(_0771_),
    .A1(_0770_),
    .S(_0767_),
    .X(_0772_));
 sg13g2_or2_1 _4273_ (.X(_0773_),
    .B(_0772_),
    .A(_0762_));
 sg13g2_o21ai_1 _4274_ (.B1(_0757_),
    .Y(_0774_),
    .A1(_0756_),
    .A2(_0761_));
 sg13g2_o21ai_1 _4275_ (.B1(_0774_),
    .Y(_0775_),
    .A1(_0772_),
    .A2(_0762_));
 sg13g2_nand2_1 _4276_ (.Y(_0776_),
    .A(_0681_),
    .B(_0775_));
 sg13g2_xor2_1 _4277_ (.B(_0681_),
    .A(_0775_),
    .X(_0777_));
 sg13g2_nand2_1 _4278_ (.Y(_0778_),
    .A(_0669_),
    .B(_0777_));
 sg13g2_nor2_1 _4279_ (.A(_0670_),
    .B(_0766_),
    .Y(_0779_));
 sg13g2_nor2_1 _4280_ (.A(_0766_),
    .B(_0778_),
    .Y(_0780_));
 sg13g2_nand3_1 _4281_ (.B(_0765_),
    .C(_0775_),
    .A(_0681_),
    .Y(_0781_));
 sg13g2_xnor2_1 _4282_ (.Y(_0782_),
    .A(_0750_),
    .B(_0763_));
 sg13g2_xor2_1 _4283_ (.B(_0782_),
    .A(_0781_),
    .X(_0783_));
 sg13g2_xnor2_1 _4284_ (.Y(_0784_),
    .A(_0781_),
    .B(_0782_));
 sg13g2_nand2b_1 _4285_ (.Y(_0785_),
    .B(_0681_),
    .A_N(_0767_));
 sg13g2_nand3_1 _4286_ (.B(_0775_),
    .C(_0785_),
    .A(_0770_),
    .Y(_0786_));
 sg13g2_a21o_1 _4287_ (.A2(_0785_),
    .A1(_0775_),
    .B1(_0770_),
    .X(_0787_));
 sg13g2_a22oi_1 _4288_ (.Y(_0788_),
    .B1(_0786_),
    .B2(_0787_),
    .A2(_0777_),
    .A1(_0779_));
 sg13g2_o21ai_1 _4289_ (.B1(_0762_),
    .Y(_0789_),
    .A1(_0772_),
    .A2(_0774_));
 sg13g2_a22oi_1 _4290_ (.Y(_0790_),
    .B1(_0789_),
    .B2(_0773_),
    .A2(_0788_),
    .A1(_0784_));
 sg13g2_nor2_1 _4291_ (.A(_0670_),
    .B(net370),
    .Y(_0791_));
 sg13g2_o21ai_1 _4292_ (.B1(_0776_),
    .Y(_0792_),
    .A1(_0778_),
    .A2(net370));
 sg13g2_xnor2_1 _4293_ (.Y(_0793_),
    .A(_0792_),
    .B(_0766_));
 sg13g2_nand2b_1 _4294_ (.Y(_0794_),
    .B(_0670_),
    .A_N(net370));
 sg13g2_nand2_1 _4295_ (.Y(_0795_),
    .A(_0669_),
    .B(net370));
 sg13g2_xnor2_1 _4296_ (.Y(_0796_),
    .A(_0669_),
    .B(net370));
 sg13g2_inv_1 _4297_ (.Y(_0797_),
    .A(_0796_));
 sg13g2_and3_1 _4298_ (.X(_0798_),
    .A(_0664_),
    .B(_0777_),
    .C(_0796_));
 sg13g2_or3_1 _4299_ (.A(_0780_),
    .B(_0783_),
    .C(net370),
    .X(_0799_));
 sg13g2_o21ai_1 _4300_ (.B1(_0783_),
    .Y(_0800_),
    .A1(_0780_),
    .A2(net370));
 sg13g2_nand2_1 _4301_ (.Y(_0801_),
    .A(_0799_),
    .B(_0800_));
 sg13g2_nor3_1 _4302_ (.A(_0793_),
    .B(_0798_),
    .C(_0801_),
    .Y(_0802_));
 sg13g2_or3_2 _4303_ (.A(_0798_),
    .B(_0793_),
    .C(_0801_),
    .X(_0803_));
 sg13g2_and3_1 _4304_ (.X(_0804_),
    .A(_0786_),
    .B(_0787_),
    .C(_0799_));
 sg13g2_a21o_2 _4305_ (.A2(_0788_),
    .A1(_0784_),
    .B1(_0804_),
    .X(_0805_));
 sg13g2_nand2_2 _4306_ (.Y(_0806_),
    .A(_0803_),
    .B(_0805_));
 sg13g2_xnor2_1 _4307_ (.Y(_0807_),
    .A(_0777_),
    .B(_0791_));
 sg13g2_a21oi_2 _4308_ (.B1(_0665_),
    .Y(_0808_),
    .A2(_0805_),
    .A1(_0803_));
 sg13g2_a221oi_1 _4309_ (.B2(_0803_),
    .C1(_0665_),
    .B1(_0805_),
    .A1(_0794_),
    .Y(_0809_),
    .A2(_0795_));
 sg13g2_xnor2_1 _4310_ (.Y(_0810_),
    .A(_0809_),
    .B(_0807_));
 sg13g2_and3_1 _4311_ (.X(_0811_),
    .A(_0665_),
    .B(_0803_),
    .C(_0805_));
 sg13g2_nor2_1 _4312_ (.A(_0808_),
    .B(_0811_),
    .Y(_0812_));
 sg13g2_inv_1 _4313_ (.Y(_0813_),
    .A(_0812_));
 sg13g2_nor2b_1 _4314_ (.A(net375),
    .B_N(_0660_),
    .Y(_0814_));
 sg13g2_nand2_1 _4315_ (.Y(_0815_),
    .A(_0650_),
    .B(_0814_));
 sg13g2_or2_1 _4316_ (.X(_0816_),
    .B(_0814_),
    .A(_0650_));
 sg13g2_nand2_1 _4317_ (.Y(_0817_),
    .A(_0815_),
    .B(_0816_));
 sg13g2_and2_1 _4318_ (.A(_0796_),
    .B(_0817_),
    .X(_0818_));
 sg13g2_inv_1 _4319_ (.Y(_0819_),
    .A(_0818_));
 sg13g2_nor3_1 _4320_ (.A(_0808_),
    .B(_0811_),
    .C(_0819_),
    .Y(_0820_));
 sg13g2_a21o_1 _4321_ (.A2(_0805_),
    .A1(_0803_),
    .B1(_0798_),
    .X(_0822_));
 sg13g2_or2_1 _4322_ (.X(_0823_),
    .B(_0822_),
    .A(_0793_));
 sg13g2_xnor2_1 _4323_ (.Y(_0824_),
    .A(_0793_),
    .B(_0822_));
 sg13g2_inv_1 _4324_ (.Y(_0825_),
    .A(_0824_));
 sg13g2_nor3_1 _4325_ (.A(_0810_),
    .B(_0820_),
    .C(_0824_),
    .Y(_0826_));
 sg13g2_or3_2 _4326_ (.A(_0824_),
    .B(_0820_),
    .C(_0810_),
    .X(_0827_));
 sg13g2_a21oi_1 _4327_ (.A1(_0801_),
    .A2(_0823_),
    .Y(_0828_),
    .B1(_0802_));
 sg13g2_a21o_1 _4328_ (.A2(_0823_),
    .A1(_0801_),
    .B1(_0802_),
    .X(_0829_));
 sg13g2_nand2_2 _4329_ (.Y(_0830_),
    .A(_0827_),
    .B(_0829_));
 sg13g2_o21ai_1 _4330_ (.B1(_0817_),
    .Y(_0831_),
    .A1(_0826_),
    .A2(_0828_));
 sg13g2_a221oi_1 _4331_ (.B2(_0827_),
    .C1(_0813_),
    .B1(_0829_),
    .A1(_0815_),
    .Y(_0833_),
    .A2(_0816_));
 sg13g2_or3_1 _4332_ (.A(_0833_),
    .B(_0808_),
    .C(_0797_),
    .X(_0834_));
 sg13g2_o21ai_1 _4333_ (.B1(_0797_),
    .Y(_0835_),
    .A1(_0808_),
    .A2(_0833_));
 sg13g2_nand2_1 _4334_ (.Y(_0836_),
    .A(_0834_),
    .B(_0835_));
 sg13g2_a21oi_1 _4335_ (.A1(_0827_),
    .A2(_0829_),
    .Y(_0837_),
    .B1(_0820_));
 sg13g2_nor2b_1 _4336_ (.A(_0810_),
    .B_N(_0837_),
    .Y(_0838_));
 sg13g2_xnor2_1 _4337_ (.Y(_0839_),
    .A(_0810_),
    .B(_0837_));
 sg13g2_nand4_1 _4338_ (.B(_0816_),
    .C(_0827_),
    .A(_0815_),
    .Y(_0840_),
    .D(_0829_));
 sg13g2_nand2_2 _4339_ (.Y(_0841_),
    .A(_0831_),
    .B(_0840_));
 sg13g2_or2_1 _4340_ (.X(_0842_),
    .B(_0658_),
    .A(net375));
 sg13g2_or2_1 _4341_ (.X(_0844_),
    .B(_0842_),
    .A(_0659_));
 sg13g2_nand2_1 _4342_ (.Y(_0845_),
    .A(_0659_),
    .B(_0842_));
 sg13g2_and2_1 _4343_ (.A(_0844_),
    .B(_0845_),
    .X(_0846_));
 sg13g2_nor2_1 _4344_ (.A(_0813_),
    .B(_0846_),
    .Y(_0847_));
 sg13g2_nor2b_1 _4345_ (.A(_0841_),
    .B_N(_0847_),
    .Y(_0848_));
 sg13g2_nand3_1 _4346_ (.B(_0840_),
    .C(_0847_),
    .A(_0831_),
    .Y(_0849_));
 sg13g2_nor2_1 _4347_ (.A(_0836_),
    .B(_0848_),
    .Y(_0850_));
 sg13g2_nand4_1 _4348_ (.B(_0835_),
    .C(_0839_),
    .A(_0834_),
    .Y(_0851_),
    .D(_0849_));
 sg13g2_o21ai_1 _4349_ (.B1(_0827_),
    .Y(_0852_),
    .A1(_0825_),
    .A2(_0838_));
 sg13g2_nand2_2 _4350_ (.Y(_0853_),
    .A(_0851_),
    .B(_0852_));
 sg13g2_a21oi_1 _4351_ (.A1(_0851_),
    .A2(_0852_),
    .Y(_0855_),
    .B1(_0846_));
 sg13g2_a21o_1 _4352_ (.A2(_0852_),
    .A1(_0851_),
    .B1(_0846_),
    .X(_0856_));
 sg13g2_nand3_1 _4353_ (.B(_0851_),
    .C(_0852_),
    .A(_0846_),
    .Y(_0857_));
 sg13g2_and2_1 _4354_ (.A(_0856_),
    .B(_0857_),
    .X(_0858_));
 sg13g2_nor2_1 _4355_ (.A(net375),
    .B(_0656_),
    .Y(_0859_));
 sg13g2_xor2_1 _4356_ (.B(_0859_),
    .A(_0657_),
    .X(_0860_));
 sg13g2_a221oi_1 _4357_ (.B2(_0851_),
    .C1(_0841_),
    .B1(_0852_),
    .A1(_0844_),
    .Y(_0861_),
    .A2(_0845_));
 sg13g2_xnor2_1 _4358_ (.Y(_0862_),
    .A(_0813_),
    .B(_0831_));
 sg13g2_nand2_1 _4359_ (.Y(_0863_),
    .A(_0813_),
    .B(_0861_));
 sg13g2_o21ai_1 _4360_ (.B1(_0863_),
    .Y(_0864_),
    .A1(_0861_),
    .A2(_0862_));
 sg13g2_mux2_1 _4361_ (.A0(_0862_),
    .A1(_0812_),
    .S(_0861_),
    .X(_0866_));
 sg13g2_nor2_1 _4362_ (.A(_0841_),
    .B(_0860_),
    .Y(_0867_));
 sg13g2_nand3_1 _4363_ (.B(_0857_),
    .C(_0867_),
    .A(_0856_),
    .Y(_0868_));
 sg13g2_a21oi_1 _4364_ (.A1(_0851_),
    .A2(_0852_),
    .Y(_0869_),
    .B1(_0848_));
 sg13g2_xnor2_1 _4365_ (.Y(_0870_),
    .A(_0836_),
    .B(_0869_));
 sg13g2_nand3_1 _4366_ (.B(_0866_),
    .C(_0870_),
    .A(_0868_),
    .Y(_0871_));
 sg13g2_a21oi_1 _4367_ (.A1(_0850_),
    .A2(_0853_),
    .Y(_0872_),
    .B1(_0839_));
 sg13g2_a21o_2 _4368_ (.A2(_0850_),
    .A1(_0839_),
    .B1(_0872_),
    .X(_0873_));
 sg13g2_nand2_1 _4369_ (.Y(_0874_),
    .A(_0871_),
    .B(_0873_));
 sg13g2_a21oi_2 _4370_ (.B1(_0860_),
    .Y(_0875_),
    .A2(_0871_),
    .A1(_0873_));
 sg13g2_a21o_1 _4371_ (.A2(_0873_),
    .A1(_0871_),
    .B1(_0860_),
    .X(_0877_));
 sg13g2_a21oi_2 _4372_ (.B1(_0855_),
    .Y(_0878_),
    .A2(_0875_),
    .A1(_0858_));
 sg13g2_xnor2_1 _4373_ (.Y(_0879_),
    .A(_0878_),
    .B(_0841_));
 sg13g2_nand3_1 _4374_ (.B(_0871_),
    .C(_0873_),
    .A(_0860_),
    .Y(_0880_));
 sg13g2_nand2_1 _4375_ (.Y(_0881_),
    .A(_0877_),
    .B(_0880_));
 sg13g2_nand2_1 _4376_ (.Y(_0882_),
    .A(_0643_),
    .B(_0654_));
 sg13g2_xor2_1 _4377_ (.B(_0882_),
    .A(_0655_),
    .X(_0883_));
 sg13g2_nand2_1 _4378_ (.Y(_0884_),
    .A(_0643_),
    .B(_0653_));
 sg13g2_xor2_1 _4379_ (.B(_0884_),
    .A(_0652_),
    .X(_0885_));
 sg13g2_nand4_1 _4380_ (.B(_0880_),
    .C(_0883_),
    .A(_0877_),
    .Y(_0886_),
    .D(_0885_));
 sg13g2_xnor2_1 _4381_ (.Y(_0888_),
    .A(_0858_),
    .B(_0875_));
 sg13g2_and2_1 _4382_ (.A(_0886_),
    .B(_0888_),
    .X(_0889_));
 sg13g2_a22oi_1 _4383_ (.Y(_0890_),
    .B1(_0871_),
    .B2(_0873_),
    .A2(_0867_),
    .A1(_0858_));
 sg13g2_a221oi_1 _4384_ (.B2(_0873_),
    .C1(_0864_),
    .B1(_0871_),
    .A1(_0858_),
    .Y(_0891_),
    .A2(_0867_));
 sg13g2_xnor2_1 _4385_ (.Y(_0892_),
    .A(_0866_),
    .B(_0890_));
 sg13g2_o21ai_1 _4386_ (.B1(_0871_),
    .Y(_0893_),
    .A1(_0870_),
    .A2(_0891_));
 sg13g2_nand2_1 _4387_ (.Y(_0894_),
    .A(_0892_),
    .B(_0893_));
 sg13g2_a21oi_2 _4388_ (.B1(_0894_),
    .Y(_0895_),
    .A2(_0889_),
    .A1(_0879_));
 sg13g2_nor2_1 _4389_ (.A(net374),
    .B(_0895_),
    .Y(_0896_));
 sg13g2_a21oi_1 _4390_ (.A1(_0643_),
    .A2(_0874_),
    .Y(_0897_),
    .B1(_0896_));
 sg13g2_nand2b_1 _4391_ (.Y(_0899_),
    .B(_0897_),
    .A_N(_0853_));
 sg13g2_nor3_2 _4392_ (.A(_0806_),
    .B(_0830_),
    .C(_0899_),
    .Y(_0900_));
 sg13g2_and2_1 _4393_ (.A(_0643_),
    .B(_0899_),
    .X(_0901_));
 sg13g2_o21ai_1 _4394_ (.B1(_0643_),
    .Y(_0902_),
    .A1(_0830_),
    .A2(_0899_));
 sg13g2_o21ai_1 _4395_ (.B1(_0790_),
    .Y(_0903_),
    .A1(net374),
    .A2(_0900_));
 sg13g2_inv_1 _4396_ (.Y(_0904_),
    .A(_0903_));
 sg13g2_nor2_1 _4397_ (.A(net34),
    .B(_0903_),
    .Y(_0905_));
 sg13g2_nand2_1 _4398_ (.Y(_0906_),
    .A(_0643_),
    .B(_0903_));
 sg13g2_nor2_1 _4399_ (.A(net375),
    .B(_0905_),
    .Y(_0907_));
 sg13g2_a21o_1 _4400_ (.A2(_0905_),
    .A1(_0759_),
    .B1(net374),
    .X(_0908_));
 sg13g2_o21ai_1 _4401_ (.B1(_0908_),
    .Y(_0910_),
    .A1(net374),
    .A2(_0742_));
 sg13g2_nor2_1 _4402_ (.A(net374),
    .B(net35),
    .Y(_0911_));
 sg13g2_nor3_2 _4403_ (.A(net48),
    .B(_0910_),
    .C(_0911_),
    .Y(_0912_));
 sg13g2_nor2_2 _4404_ (.A(net374),
    .B(_0912_),
    .Y(_0913_));
 sg13g2_and2_1 _4405_ (.A(_0155_),
    .B(_0913_),
    .X(_0914_));
 sg13g2_nand2_1 _4406_ (.Y(_0915_),
    .A(_0155_),
    .B(_0913_));
 sg13g2_nor2_2 _4407_ (.A(_0155_),
    .B(_0913_),
    .Y(_0916_));
 sg13g2_nor2_2 _4408_ (.A(_0914_),
    .B(_0916_),
    .Y(_0917_));
 sg13g2_nand2_1 _4409_ (.Y(_0918_),
    .A(net442),
    .B(net416));
 sg13g2_nand2_1 _4410_ (.Y(_0919_),
    .A(\pid.Ki[7] ),
    .B(net413));
 sg13g2_nand2_1 _4411_ (.Y(_0921_),
    .A(net444),
    .B(net409));
 sg13g2_xor2_1 _4412_ (.B(_0919_),
    .A(_0918_),
    .X(_0922_));
 sg13g2_nand2b_1 _4413_ (.Y(_0923_),
    .B(_0922_),
    .A_N(_0921_));
 sg13g2_o21ai_1 _4414_ (.B1(_0923_),
    .Y(_0924_),
    .A1(_0918_),
    .A2(_0919_));
 sg13g2_nor2_1 _4415_ (.A(_0887_),
    .B(_2013_),
    .Y(_0925_));
 sg13g2_nand2b_1 _4416_ (.Y(_0926_),
    .B(net442),
    .A_N(net413));
 sg13g2_nand2_1 _4417_ (.Y(_0927_),
    .A(net443),
    .B(net409));
 sg13g2_nor2_1 _4418_ (.A(_0926_),
    .B(_0927_),
    .Y(_0928_));
 sg13g2_xor2_1 _4419_ (.B(_0927_),
    .A(_0926_),
    .X(_0929_));
 sg13g2_xor2_1 _4420_ (.B(_0929_),
    .A(_0925_),
    .X(_0930_));
 sg13g2_xnor2_1 _4421_ (.Y(_0932_),
    .A(_0924_),
    .B(_0930_));
 sg13g2_nand2_1 _4422_ (.Y(_0933_),
    .A(net449),
    .B(net390));
 sg13g2_nor2_1 _4423_ (.A(_0004_),
    .B(_2036_),
    .Y(_0934_));
 sg13g2_nor2_2 _4424_ (.A(_0004_),
    .B(_2027_),
    .Y(_0935_));
 sg13g2_nor2_1 _4425_ (.A(_0005_),
    .B(_2036_),
    .Y(_0936_));
 sg13g2_xnor2_1 _4426_ (.Y(_0937_),
    .A(_0935_),
    .B(_0936_));
 sg13g2_nor2_1 _4427_ (.A(net384),
    .B(_0937_),
    .Y(_0938_));
 sg13g2_xor2_1 _4428_ (.B(_0937_),
    .A(net384),
    .X(_0939_));
 sg13g2_nor2b_1 _4429_ (.A(_0932_),
    .B_N(_0939_),
    .Y(_0940_));
 sg13g2_a21o_1 _4430_ (.A2(_0930_),
    .A1(_0924_),
    .B1(_0940_),
    .X(_0941_));
 sg13g2_inv_1 _4431_ (.Y(_0943_),
    .A(_0941_));
 sg13g2_a21oi_1 _4432_ (.A1(_0925_),
    .A2(_0929_),
    .Y(_0944_),
    .B1(_0928_));
 sg13g2_nand2_1 _4433_ (.Y(_0945_),
    .A(net444),
    .B(_2026_));
 sg13g2_o21ai_1 _4434_ (.B1(\pid.Ki[8] ),
    .Y(_0946_),
    .A1(_1898_),
    .A2(_1920_));
 sg13g2_nand2_1 _4435_ (.Y(_0947_),
    .A(net443),
    .B(net403));
 sg13g2_xor2_1 _4436_ (.B(_0947_),
    .A(_0946_),
    .X(_0948_));
 sg13g2_nand2b_1 _4437_ (.Y(_0949_),
    .B(_0948_),
    .A_N(_0945_));
 sg13g2_xnor2_1 _4438_ (.Y(_0950_),
    .A(_0945_),
    .B(_0948_));
 sg13g2_nor2b_1 _4439_ (.A(_0944_),
    .B_N(_0950_),
    .Y(_0951_));
 sg13g2_xnor2_1 _4440_ (.Y(_0952_),
    .A(_0944_),
    .B(_0950_));
 sg13g2_nand3_1 _4441_ (.B(net390),
    .C(_0934_),
    .A(net445),
    .Y(_0954_));
 sg13g2_a21o_1 _4442_ (.A2(net391),
    .A1(net445),
    .B1(_0934_),
    .X(_0955_));
 sg13g2_nand2_1 _4443_ (.Y(_0956_),
    .A(_0954_),
    .B(_0955_));
 sg13g2_xor2_1 _4444_ (.B(_0956_),
    .A(net384),
    .X(_0957_));
 sg13g2_xnor2_1 _4445_ (.Y(_0958_),
    .A(_0952_),
    .B(_0957_));
 sg13g2_xor2_1 _4446_ (.B(_0958_),
    .A(_0941_),
    .X(_0959_));
 sg13g2_nor3_2 _4447_ (.A(_0003_),
    .B(_2030_),
    .C(_2032_),
    .Y(_0960_));
 sg13g2_nand2_1 _4448_ (.Y(_0961_),
    .A(net448),
    .B(_0960_));
 sg13g2_nand2b_1 _4449_ (.Y(_0962_),
    .B(_0003_),
    .A_N(net448));
 sg13g2_nand3_1 _4450_ (.B(_0961_),
    .C(_0962_),
    .A(net390),
    .Y(_0963_));
 sg13g2_nor2_1 _4451_ (.A(_0909_),
    .B(_0963_),
    .Y(_0964_));
 sg13g2_a21oi_2 _4452_ (.B1(_0964_),
    .Y(_0965_),
    .A2(_0960_),
    .A1(net448));
 sg13g2_nor2_1 _4453_ (.A(_0909_),
    .B(_2038_),
    .Y(_0966_));
 sg13g2_mux2_2 _4454_ (.A0(_0909_),
    .A1(_0966_),
    .S(_0963_),
    .X(_0967_));
 sg13g2_a21oi_1 _4455_ (.A1(_0935_),
    .A2(_0936_),
    .Y(_0968_),
    .B1(_0938_));
 sg13g2_nand2b_1 _4456_ (.Y(_0969_),
    .B(_0967_),
    .A_N(_0968_));
 sg13g2_xnor2_1 _4457_ (.Y(_0970_),
    .A(_0967_),
    .B(_0968_));
 sg13g2_nand2b_1 _4458_ (.Y(_0971_),
    .B(_0970_),
    .A_N(_0965_));
 sg13g2_xnor2_1 _4459_ (.Y(_0972_),
    .A(_0965_),
    .B(_0970_));
 sg13g2_nand2b_1 _4460_ (.Y(_0973_),
    .B(_0972_),
    .A_N(_0959_));
 sg13g2_o21ai_1 _4461_ (.B1(_0973_),
    .Y(_0975_),
    .A1(_0943_),
    .A2(_0958_));
 sg13g2_a21oi_1 _4462_ (.A1(_0952_),
    .A2(_0957_),
    .Y(_0976_),
    .B1(_0951_));
 sg13g2_o21ai_1 _4463_ (.B1(_0949_),
    .Y(_0977_),
    .A1(_0946_),
    .A2(_0947_));
 sg13g2_nand2_1 _4464_ (.Y(_0978_),
    .A(net443),
    .B(net400));
 sg13g2_nand2_1 _4465_ (.Y(_0979_),
    .A(net442),
    .B(_2013_));
 sg13g2_xor2_1 _4466_ (.B(_0979_),
    .A(_0978_),
    .X(_0980_));
 sg13g2_nand3_1 _4467_ (.B(net394),
    .C(_0980_),
    .A(net444),
    .Y(_0981_));
 sg13g2_a21o_1 _4468_ (.A2(net394),
    .A1(net444),
    .B1(_0980_),
    .X(_0982_));
 sg13g2_and2_1 _4469_ (.A(_0981_),
    .B(_0982_),
    .X(_0983_));
 sg13g2_nand2_1 _4470_ (.Y(_0984_),
    .A(_0977_),
    .B(_0983_));
 sg13g2_xnor2_1 _4471_ (.Y(_0986_),
    .A(_0977_),
    .B(_0983_));
 sg13g2_nand3_1 _4472_ (.B(net445),
    .C(net390),
    .A(\pid.Ki[5] ),
    .Y(_0987_));
 sg13g2_o21ai_1 _4473_ (.B1(net390),
    .Y(_0988_),
    .A1(\pid.Ki[5] ),
    .A2(net445));
 sg13g2_nand2b_1 _4474_ (.Y(_0989_),
    .B(_0987_),
    .A_N(_0988_));
 sg13g2_xor2_1 _4475_ (.B(_0989_),
    .A(net384),
    .X(_0990_));
 sg13g2_inv_2 _4476_ (.Y(_0991_),
    .A(_0990_));
 sg13g2_xnor2_1 _4477_ (.Y(_0992_),
    .A(_0986_),
    .B(_0990_));
 sg13g2_nor2b_1 _4478_ (.A(_0976_),
    .B_N(_0992_),
    .Y(_0993_));
 sg13g2_xnor2_1 _4479_ (.Y(_0994_),
    .A(_0976_),
    .B(_0992_));
 sg13g2_o21ai_1 _4480_ (.B1(_0954_),
    .Y(_0995_),
    .A1(net384),
    .A2(_0956_));
 sg13g2_xor2_1 _4481_ (.B(_0995_),
    .A(_0967_),
    .X(_0997_));
 sg13g2_nor2b_1 _4482_ (.A(_0965_),
    .B_N(_0997_),
    .Y(_0998_));
 sg13g2_xnor2_1 _4483_ (.Y(_0999_),
    .A(_0965_),
    .B(_0997_));
 sg13g2_xnor2_1 _4484_ (.Y(_1000_),
    .A(_0994_),
    .B(_0999_));
 sg13g2_nand2b_1 _4485_ (.Y(_1001_),
    .B(_0975_),
    .A_N(_1000_));
 sg13g2_nand2_1 _4486_ (.Y(_1002_),
    .A(_0969_),
    .B(_0971_));
 sg13g2_xor2_1 _4487_ (.B(_1000_),
    .A(_0975_),
    .X(_1003_));
 sg13g2_nand2b_1 _4488_ (.Y(_1004_),
    .B(_1002_),
    .A_N(_1003_));
 sg13g2_nand2_1 _4489_ (.Y(_1005_),
    .A(_1001_),
    .B(_1004_));
 sg13g2_a21o_1 _4490_ (.A2(_0995_),
    .A1(_0967_),
    .B1(_0998_),
    .X(_1006_));
 sg13g2_a21oi_1 _4491_ (.A1(_0994_),
    .A2(_0999_),
    .Y(_1008_),
    .B1(_0993_));
 sg13g2_o21ai_1 _4492_ (.B1(_0987_),
    .Y(_1009_),
    .A1(net384),
    .A2(_0988_));
 sg13g2_xor2_1 _4493_ (.B(_1009_),
    .A(_0967_),
    .X(_1010_));
 sg13g2_nor2b_1 _4494_ (.A(_0965_),
    .B_N(_1010_),
    .Y(_1011_));
 sg13g2_xnor2_1 _4495_ (.Y(_1012_),
    .A(_0965_),
    .B(_1010_));
 sg13g2_inv_1 _4496_ (.Y(_1013_),
    .A(_1012_));
 sg13g2_o21ai_1 _4497_ (.B1(_0984_),
    .Y(_1014_),
    .A1(_0986_),
    .A2(_0991_));
 sg13g2_o21ai_1 _4498_ (.B1(_0981_),
    .Y(_1015_),
    .A1(_0978_),
    .A2(_0979_));
 sg13g2_nand2_2 _4499_ (.Y(_1016_),
    .A(net444),
    .B(net391));
 sg13g2_nand2_1 _4500_ (.Y(_1017_),
    .A(net443),
    .B(net394));
 sg13g2_nand2_2 _4501_ (.Y(_1018_),
    .A(net442),
    .B(_2027_));
 sg13g2_xor2_1 _4502_ (.B(_1018_),
    .A(_1017_),
    .X(_1019_));
 sg13g2_nand2b_1 _4503_ (.Y(_1020_),
    .B(_1019_),
    .A_N(_1016_));
 sg13g2_xnor2_1 _4504_ (.Y(_1021_),
    .A(_1016_),
    .B(_1019_));
 sg13g2_nand2_1 _4505_ (.Y(_1022_),
    .A(_1015_),
    .B(_1021_));
 sg13g2_xnor2_1 _4506_ (.Y(_1023_),
    .A(_1015_),
    .B(_1021_));
 sg13g2_xnor2_1 _4507_ (.Y(_1024_),
    .A(_0991_),
    .B(_1023_));
 sg13g2_nand2b_1 _4508_ (.Y(_1025_),
    .B(_1014_),
    .A_N(_1024_));
 sg13g2_xor2_1 _4509_ (.B(_1024_),
    .A(_1014_),
    .X(_1026_));
 sg13g2_xnor2_1 _4510_ (.Y(_1027_),
    .A(_1013_),
    .B(_1026_));
 sg13g2_nor2_1 _4511_ (.A(_1008_),
    .B(_1027_),
    .Y(_1029_));
 sg13g2_xor2_1 _4512_ (.B(_1027_),
    .A(_1008_),
    .X(_1030_));
 sg13g2_xnor2_1 _4513_ (.Y(_1031_),
    .A(_1006_),
    .B(_1030_));
 sg13g2_a21oi_1 _4514_ (.A1(_1001_),
    .A2(_1004_),
    .Y(_1032_),
    .B1(_1031_));
 sg13g2_a21oi_1 _4515_ (.A1(_1006_),
    .A2(_1030_),
    .Y(_1033_),
    .B1(_1029_));
 sg13g2_a21oi_2 _4516_ (.B1(_1011_),
    .Y(_1034_),
    .A2(_1009_),
    .A1(_0967_));
 sg13g2_o21ai_1 _4517_ (.B1(_1025_),
    .Y(_1035_),
    .A1(_1013_),
    .A2(_1026_));
 sg13g2_o21ai_1 _4518_ (.B1(_1022_),
    .Y(_1036_),
    .A1(_0991_),
    .A2(_1023_));
 sg13g2_o21ai_1 _4519_ (.B1(_1020_),
    .Y(_1037_),
    .A1(_1017_),
    .A2(_1018_));
 sg13g2_nor2_1 _4520_ (.A(_0001_),
    .B(net394),
    .Y(_1038_));
 sg13g2_nor2_1 _4521_ (.A(_0002_),
    .B(_2038_),
    .Y(_1040_));
 sg13g2_nand2_1 _4522_ (.Y(_1041_),
    .A(_1038_),
    .B(_1040_));
 sg13g2_xnor2_1 _4523_ (.Y(_1042_),
    .A(_1038_),
    .B(_1040_));
 sg13g2_xor2_1 _4524_ (.B(_1042_),
    .A(_1016_),
    .X(_1043_));
 sg13g2_nand2_1 _4525_ (.Y(_1044_),
    .A(_1037_),
    .B(_1043_));
 sg13g2_xnor2_1 _4526_ (.Y(_1045_),
    .A(_1037_),
    .B(_1043_));
 sg13g2_or2_1 _4527_ (.X(_1046_),
    .B(_1045_),
    .A(_0991_));
 sg13g2_xnor2_1 _4528_ (.Y(_1047_),
    .A(_0991_),
    .B(_1045_));
 sg13g2_nand2b_1 _4529_ (.Y(_1048_),
    .B(_1036_),
    .A_N(_1047_));
 sg13g2_xor2_1 _4530_ (.B(_1047_),
    .A(_1036_),
    .X(_1049_));
 sg13g2_xnor2_1 _4531_ (.Y(_1051_),
    .A(_1012_),
    .B(_1049_));
 sg13g2_nand2_1 _4532_ (.Y(_1052_),
    .A(_1035_),
    .B(_1051_));
 sg13g2_xnor2_1 _4533_ (.Y(_1053_),
    .A(_1035_),
    .B(_1051_));
 sg13g2_xor2_1 _4534_ (.B(_1053_),
    .A(_1034_),
    .X(_1054_));
 sg13g2_nand2b_1 _4535_ (.Y(_1055_),
    .B(_1054_),
    .A_N(_1033_));
 sg13g2_xnor2_1 _4536_ (.Y(_1056_),
    .A(_1033_),
    .B(_1054_));
 sg13g2_and2_1 _4537_ (.A(_1032_),
    .B(_1056_),
    .X(_1057_));
 sg13g2_inv_1 _4538_ (.Y(_1058_),
    .A(_1057_));
 sg13g2_nand2_1 _4539_ (.Y(_1059_),
    .A(net442),
    .B(_1670_));
 sg13g2_nand2_1 _4540_ (.Y(_1060_),
    .A(net443),
    .B(net418));
 sg13g2_nand2_1 _4541_ (.Y(_1062_),
    .A(\pid.Ki[6] ),
    .B(net415));
 sg13g2_xor2_1 _4542_ (.B(_1060_),
    .A(_1059_),
    .X(_1063_));
 sg13g2_nand2b_1 _4543_ (.Y(_1064_),
    .B(_1063_),
    .A_N(_1062_));
 sg13g2_o21ai_1 _4544_ (.B1(_1064_),
    .Y(_1065_),
    .A1(_1059_),
    .A2(_1060_));
 sg13g2_xnor2_1 _4545_ (.Y(_1066_),
    .A(_0921_),
    .B(_0922_));
 sg13g2_xnor2_1 _4546_ (.Y(_1067_),
    .A(_1065_),
    .B(_1066_));
 sg13g2_nor2_2 _4547_ (.A(_0005_),
    .B(_2013_),
    .Y(_1068_));
 sg13g2_nand2_1 _4548_ (.Y(_1069_),
    .A(_0935_),
    .B(_1068_));
 sg13g2_a22oi_1 _4549_ (.Y(_1070_),
    .B1(net400),
    .B2(_0931_),
    .A2(net52),
    .A1(_0920_));
 sg13g2_a21oi_1 _4550_ (.A1(_0935_),
    .A2(_1068_),
    .Y(_1071_),
    .B1(_1070_));
 sg13g2_xnor2_1 _4551_ (.Y(_1072_),
    .A(net385),
    .B(_1071_));
 sg13g2_nor2b_1 _4552_ (.A(_1067_),
    .B_N(_1072_),
    .Y(_1073_));
 sg13g2_a21o_1 _4553_ (.A2(_1066_),
    .A1(_1065_),
    .B1(_1073_),
    .X(_1074_));
 sg13g2_xnor2_1 _4554_ (.Y(_1075_),
    .A(_0932_),
    .B(_0939_));
 sg13g2_xnor2_1 _4555_ (.Y(_1076_),
    .A(_1074_),
    .B(_1075_));
 sg13g2_nand2_1 _4556_ (.Y(_1077_),
    .A(net446),
    .B(net394));
 sg13g2_a22oi_1 _4557_ (.Y(_1078_),
    .B1(_0964_),
    .B2(net394),
    .A2(_0960_),
    .A1(net448));
 sg13g2_o21ai_1 _4558_ (.B1(_1069_),
    .Y(_1079_),
    .A1(net385),
    .A2(_1070_));
 sg13g2_nand2_1 _4559_ (.Y(_1080_),
    .A(_0967_),
    .B(_1079_));
 sg13g2_xor2_1 _4560_ (.B(_1079_),
    .A(_0967_),
    .X(_1081_));
 sg13g2_inv_1 _4561_ (.Y(_1083_),
    .A(_1081_));
 sg13g2_xnor2_1 _4562_ (.Y(_1084_),
    .A(_1078_),
    .B(_1081_));
 sg13g2_nor2b_1 _4563_ (.A(_1076_),
    .B_N(_1084_),
    .Y(_1085_));
 sg13g2_a21o_1 _4564_ (.A2(_1075_),
    .A1(_1074_),
    .B1(_1085_),
    .X(_1086_));
 sg13g2_xnor2_1 _4565_ (.Y(_1087_),
    .A(_0959_),
    .B(_0972_));
 sg13g2_o21ai_1 _4566_ (.B1(_1080_),
    .Y(_1088_),
    .A1(_1078_),
    .A2(_1083_));
 sg13g2_xnor2_1 _4567_ (.Y(_1089_),
    .A(_1086_),
    .B(_1087_));
 sg13g2_nor2b_1 _4568_ (.A(_1089_),
    .B_N(_1088_),
    .Y(_1090_));
 sg13g2_a21o_1 _4569_ (.A2(_1087_),
    .A1(_1086_),
    .B1(_1090_),
    .X(_1091_));
 sg13g2_xor2_1 _4570_ (.B(_1003_),
    .A(_1002_),
    .X(_1092_));
 sg13g2_nor2b_1 _4571_ (.A(_1092_),
    .B_N(_1091_),
    .Y(_1094_));
 sg13g2_xnor2_1 _4572_ (.Y(_1095_),
    .A(_1005_),
    .B(_1031_));
 sg13g2_nand2_1 _4573_ (.Y(_1096_),
    .A(_1094_),
    .B(_1095_));
 sg13g2_xor2_1 _4574_ (.B(_1095_),
    .A(_1094_),
    .X(_1097_));
 sg13g2_nor2_1 _4575_ (.A(_0001_),
    .B(_1605_),
    .Y(_1098_));
 sg13g2_nand3_1 _4576_ (.B(net421),
    .C(_1098_),
    .A(net443),
    .Y(_1099_));
 sg13g2_nand2_1 _4577_ (.Y(_1100_),
    .A(\pid.Ki[6] ),
    .B(net419));
 sg13g2_a21o_1 _4578_ (.A2(net420),
    .A1(net443),
    .B1(_1098_),
    .X(_1101_));
 sg13g2_nand2_1 _4579_ (.Y(_1102_),
    .A(_1099_),
    .B(_1101_));
 sg13g2_o21ai_1 _4580_ (.B1(_1099_),
    .Y(_1103_),
    .A1(_1100_),
    .A2(_1102_));
 sg13g2_xnor2_1 _4581_ (.Y(_1105_),
    .A(_1062_),
    .B(_1063_));
 sg13g2_xnor2_1 _4582_ (.Y(_1106_),
    .A(_1103_),
    .B(_1105_));
 sg13g2_nand2_1 _4583_ (.Y(_1107_),
    .A(\pid.Ki[5] ),
    .B(net409));
 sg13g2_nand3_1 _4584_ (.B(net409),
    .C(_1068_),
    .A(\pid.Ki[5] ),
    .Y(_1108_));
 sg13g2_xnor2_1 _4585_ (.Y(_1109_),
    .A(_1068_),
    .B(_1107_));
 sg13g2_nand2b_1 _4586_ (.Y(_1110_),
    .B(_1109_),
    .A_N(net385));
 sg13g2_xnor2_1 _4587_ (.Y(_1111_),
    .A(net385),
    .B(_1109_));
 sg13g2_nor2b_1 _4588_ (.A(_1106_),
    .B_N(_1111_),
    .Y(_1112_));
 sg13g2_a21oi_1 _4589_ (.A1(_1103_),
    .A2(_1105_),
    .Y(_1113_),
    .B1(_1112_));
 sg13g2_xnor2_1 _4590_ (.Y(_1114_),
    .A(_1067_),
    .B(_1072_));
 sg13g2_nor2b_1 _4591_ (.A(_1113_),
    .B_N(_1114_),
    .Y(_1116_));
 sg13g2_xnor2_1 _4592_ (.Y(_1117_),
    .A(_1113_),
    .B(_1114_));
 sg13g2_nand2_1 _4593_ (.Y(_1118_),
    .A(net448),
    .B(net395));
 sg13g2_nand2_1 _4594_ (.Y(_1119_),
    .A(net446),
    .B(net400));
 sg13g2_xnor2_1 _4595_ (.Y(_1120_),
    .A(_0960_),
    .B(_1118_));
 sg13g2_nand2b_1 _4596_ (.Y(_1121_),
    .B(_1120_),
    .A_N(_1119_));
 sg13g2_o21ai_1 _4597_ (.B1(_1121_),
    .Y(_1122_),
    .A1(_2036_),
    .A2(_0961_));
 sg13g2_nand2_1 _4598_ (.Y(_1123_),
    .A(_1108_),
    .B(_1110_));
 sg13g2_xor2_1 _4599_ (.B(_1077_),
    .A(_0963_),
    .X(_1124_));
 sg13g2_xnor2_1 _4600_ (.Y(_1125_),
    .A(_1123_),
    .B(_1124_));
 sg13g2_nor2b_1 _4601_ (.A(_1125_),
    .B_N(_1122_),
    .Y(_1126_));
 sg13g2_xor2_1 _4602_ (.B(_1125_),
    .A(_1122_),
    .X(_1127_));
 sg13g2_inv_1 _4603_ (.Y(_1128_),
    .A(_1127_));
 sg13g2_a21oi_1 _4604_ (.A1(_1117_),
    .A2(_1128_),
    .Y(_1129_),
    .B1(_1116_));
 sg13g2_xnor2_1 _4605_ (.Y(_1130_),
    .A(_1076_),
    .B(_1084_));
 sg13g2_nand2b_1 _4606_ (.Y(_1131_),
    .B(_1130_),
    .A_N(_1129_));
 sg13g2_a21oi_1 _4607_ (.A1(_1123_),
    .A2(_1124_),
    .Y(_1132_),
    .B1(_1126_));
 sg13g2_xnor2_1 _4608_ (.Y(_1133_),
    .A(_1129_),
    .B(_1130_));
 sg13g2_nand2b_1 _4609_ (.Y(_1134_),
    .B(_1133_),
    .A_N(_1132_));
 sg13g2_nand2_1 _4610_ (.Y(_1135_),
    .A(_1131_),
    .B(_1134_));
 sg13g2_xor2_1 _4611_ (.B(_1089_),
    .A(_1088_),
    .X(_1137_));
 sg13g2_nand2b_1 _4612_ (.Y(_1138_),
    .B(_1135_),
    .A_N(_1137_));
 sg13g2_xor2_1 _4613_ (.B(_1092_),
    .A(_1091_),
    .X(_1139_));
 sg13g2_nand2_1 _4614_ (.Y(_1140_),
    .A(_1138_),
    .B(_1139_));
 sg13g2_nor2_1 _4615_ (.A(_1138_),
    .B(_1139_),
    .Y(_1141_));
 sg13g2_nor4_2 _4616_ (.A(_0002_),
    .B(_0887_),
    .C(net472),
    .Y(_1142_),
    .D(_1670_));
 sg13g2_xor2_1 _4617_ (.B(_1102_),
    .A(_1100_),
    .X(_1143_));
 sg13g2_and2_1 _4618_ (.A(_0920_),
    .B(net415),
    .X(_1144_));
 sg13g2_nand3_1 _4619_ (.B(net409),
    .C(_1144_),
    .A(\pid.Ki[4] ),
    .Y(_1145_));
 sg13g2_a21o_1 _4620_ (.A2(net408),
    .A1(\pid.Ki[4] ),
    .B1(_1144_),
    .X(_1146_));
 sg13g2_and2_1 _4621_ (.A(_1145_),
    .B(_1146_),
    .X(_1148_));
 sg13g2_inv_1 _4622_ (.Y(_1149_),
    .A(_1148_));
 sg13g2_xnor2_1 _4623_ (.Y(_1150_),
    .A(net384),
    .B(_1149_));
 sg13g2_xnor2_1 _4624_ (.Y(_1151_),
    .A(_1142_),
    .B(_1143_));
 sg13g2_nor2_1 _4625_ (.A(_1150_),
    .B(_1151_),
    .Y(_1152_));
 sg13g2_a21oi_1 _4626_ (.A1(_1142_),
    .A2(_1143_),
    .Y(_1153_),
    .B1(_1152_));
 sg13g2_xnor2_1 _4627_ (.Y(_1154_),
    .A(_1106_),
    .B(_1111_));
 sg13g2_nor2b_1 _4628_ (.A(_1153_),
    .B_N(_1154_),
    .Y(_1155_));
 sg13g2_xnor2_1 _4629_ (.Y(_1156_),
    .A(_1153_),
    .B(_1154_));
 sg13g2_nand2_1 _4630_ (.Y(_1157_),
    .A(_0898_),
    .B(net400));
 sg13g2_nand2_1 _4631_ (.Y(_1159_),
    .A(net448),
    .B(net400));
 sg13g2_nand3_1 _4632_ (.B(net55),
    .C(net61),
    .A(_0898_),
    .Y(_1160_));
 sg13g2_nor2_1 _4633_ (.A(_1159_),
    .B(net75),
    .Y(_1161_));
 sg13g2_xor2_1 _4634_ (.B(_1159_),
    .A(_1160_),
    .X(_1162_));
 sg13g2_a21oi_1 _4635_ (.A1(net442),
    .A2(net79),
    .Y(_1163_),
    .B1(_1161_));
 sg13g2_o21ai_1 _4636_ (.B1(_1145_),
    .Y(_1164_),
    .A1(net384),
    .A2(_1149_));
 sg13g2_xnor2_1 _4637_ (.Y(_1165_),
    .A(_1119_),
    .B(_1120_));
 sg13g2_xnor2_1 _4638_ (.Y(_1166_),
    .A(_1164_),
    .B(_1165_));
 sg13g2_nor2_1 _4639_ (.A(_1163_),
    .B(_1166_),
    .Y(_1167_));
 sg13g2_xor2_1 _4640_ (.B(_1166_),
    .A(_1163_),
    .X(_1168_));
 sg13g2_a21oi_1 _4641_ (.A1(_1156_),
    .A2(_1168_),
    .Y(_1170_),
    .B1(_1155_));
 sg13g2_xor2_1 _4642_ (.B(_1127_),
    .A(_1117_),
    .X(_1171_));
 sg13g2_nor2_1 _4643_ (.A(_1170_),
    .B(_1171_),
    .Y(_1172_));
 sg13g2_a21oi_1 _4644_ (.A1(_1164_),
    .A2(_1165_),
    .Y(_1173_),
    .B1(_1167_));
 sg13g2_xor2_1 _4645_ (.B(_1171_),
    .A(_1170_),
    .X(_1174_));
 sg13g2_nor2b_1 _4646_ (.A(_1173_),
    .B_N(_1174_),
    .Y(_1175_));
 sg13g2_nor2_1 _4647_ (.A(_1172_),
    .B(_1175_),
    .Y(_1176_));
 sg13g2_xor2_1 _4648_ (.B(_1133_),
    .A(_1132_),
    .X(_1177_));
 sg13g2_nor2_1 _4649_ (.A(_1176_),
    .B(_1177_),
    .Y(_1178_));
 sg13g2_xnor2_1 _4650_ (.Y(_1179_),
    .A(_1135_),
    .B(_1137_));
 sg13g2_and2_1 _4651_ (.A(_1178_),
    .B(_1179_),
    .X(_1180_));
 sg13g2_a22oi_1 _4652_ (.Y(_1181_),
    .B1(net422),
    .B2(\pid.Ki[6] ),
    .A2(_1605_),
    .A1(_0876_));
 sg13g2_nor2_1 _4653_ (.A(_1142_),
    .B(_1181_),
    .Y(_1182_));
 sg13g2_nand2_1 _4654_ (.Y(_1183_),
    .A(\pid.Ki[5] ),
    .B(net419));
 sg13g2_nand2_1 _4655_ (.Y(_1184_),
    .A(net445),
    .B(net415));
 sg13g2_xor2_1 _4656_ (.B(_1184_),
    .A(_1183_),
    .X(_1185_));
 sg13g2_nand3_1 _4657_ (.B(net395),
    .C(_1185_),
    .A(net449),
    .Y(_1186_));
 sg13g2_a21o_1 _4658_ (.A2(net394),
    .A1(net449),
    .B1(_1185_),
    .X(_1187_));
 sg13g2_nand2_1 _4659_ (.Y(_1188_),
    .A(_1186_),
    .B(_1187_));
 sg13g2_or3_1 _4660_ (.A(_1142_),
    .B(_1181_),
    .C(_1188_),
    .X(_1189_));
 sg13g2_xnor2_1 _4661_ (.Y(_1191_),
    .A(_1150_),
    .B(_1151_));
 sg13g2_nor2_1 _4662_ (.A(_1189_),
    .B(_1191_),
    .Y(_1192_));
 sg13g2_xor2_1 _4663_ (.B(_1189_),
    .A(_1191_),
    .X(_1193_));
 sg13g2_nand2_1 _4664_ (.Y(_1194_),
    .A(_0898_),
    .B(net51));
 sg13g2_nand2_2 _4665_ (.Y(_1195_),
    .A(\pid.Ki[2] ),
    .B(net404));
 sg13g2_nand2_1 _4666_ (.Y(_1196_),
    .A(net446),
    .B(net408));
 sg13g2_xnor2_1 _4667_ (.Y(_1197_),
    .A(_1195_),
    .B(_1157_));
 sg13g2_or2_1 _4668_ (.X(_1198_),
    .B(_1197_),
    .A(_1196_));
 sg13g2_o21ai_1 _4669_ (.B1(_1198_),
    .Y(_1199_),
    .A1(_1157_),
    .A2(_1195_));
 sg13g2_inv_1 _4670_ (.Y(_1200_),
    .A(_1199_));
 sg13g2_o21ai_1 _4671_ (.B1(_1186_),
    .Y(_1202_),
    .A1(_1183_),
    .A2(_1184_));
 sg13g2_xnor2_1 _4672_ (.Y(_1203_),
    .A(_1162_),
    .B(net442));
 sg13g2_nand2b_1 _4673_ (.Y(_1204_),
    .B(_1202_),
    .A_N(_1203_));
 sg13g2_xor2_1 _4674_ (.B(_1203_),
    .A(_1202_),
    .X(_1205_));
 sg13g2_xnor2_1 _4675_ (.Y(_1206_),
    .A(_1199_),
    .B(_1205_));
 sg13g2_a21oi_1 _4676_ (.A1(net74),
    .A2(_1206_),
    .Y(_1207_),
    .B1(_1192_));
 sg13g2_xnor2_1 _4677_ (.Y(_1208_),
    .A(_1156_),
    .B(_1168_));
 sg13g2_nor2_1 _4678_ (.A(_1207_),
    .B(_1208_),
    .Y(_1209_));
 sg13g2_o21ai_1 _4679_ (.B1(_1204_),
    .Y(_1210_),
    .A1(_1200_),
    .A2(net77));
 sg13g2_xor2_1 _4680_ (.B(_1208_),
    .A(_1207_),
    .X(_1211_));
 sg13g2_a21oi_1 _4681_ (.A1(_1210_),
    .A2(_1211_),
    .Y(_1213_),
    .B1(_1209_));
 sg13g2_xor2_1 _4682_ (.B(_1174_),
    .A(_1173_),
    .X(_1214_));
 sg13g2_nor2_1 _4683_ (.A(_1213_),
    .B(_1214_),
    .Y(_1215_));
 sg13g2_xor2_1 _4684_ (.B(_1177_),
    .A(_1176_),
    .X(_1216_));
 sg13g2_nand2_1 _4685_ (.Y(_1217_),
    .A(_1215_),
    .B(_1216_));
 sg13g2_nor2_1 _4686_ (.A(_0006_),
    .B(_2027_),
    .Y(_1218_));
 sg13g2_nand2_1 _4687_ (.Y(_1219_),
    .A(net445),
    .B(net419));
 sg13g2_nand2_1 _4688_ (.Y(_1220_),
    .A(\pid.Ki[5] ),
    .B(net423));
 sg13g2_xor2_1 _4689_ (.B(_1220_),
    .A(_1219_),
    .X(_1221_));
 sg13g2_nand2_1 _4690_ (.Y(_1222_),
    .A(_1218_),
    .B(_1221_));
 sg13g2_xnor2_1 _4691_ (.Y(_1223_),
    .A(_1218_),
    .B(_1221_));
 sg13g2_nor3_2 _4692_ (.A(_0887_),
    .B(net472),
    .C(_1223_),
    .Y(_1224_));
 sg13g2_xnor2_1 _4693_ (.Y(_1225_),
    .A(_1188_),
    .B(_1182_));
 sg13g2_nand2_1 _4694_ (.Y(_1226_),
    .A(_1224_),
    .B(_1225_));
 sg13g2_xnor2_1 _4695_ (.Y(_1227_),
    .A(_1224_),
    .B(_1225_));
 sg13g2_nor3_1 _4696_ (.A(_0003_),
    .B(_1898_),
    .C(_1920_),
    .Y(_1228_));
 sg13g2_nand2_1 _4697_ (.Y(_1229_),
    .A(net447),
    .B(net408));
 sg13g2_nand2_1 _4698_ (.Y(_1230_),
    .A(\pid.Ki[3] ),
    .B(net415));
 sg13g2_xor2_1 _4699_ (.B(_1229_),
    .A(_1194_),
    .X(_1231_));
 sg13g2_nand2b_1 _4700_ (.Y(_1232_),
    .B(_1231_),
    .A_N(_1230_));
 sg13g2_o21ai_1 _4701_ (.B1(_1232_),
    .Y(_1234_),
    .A1(_1194_),
    .A2(_1229_));
 sg13g2_o21ai_1 _4702_ (.B1(_1222_),
    .Y(_1235_),
    .A1(_1219_),
    .A2(_1220_));
 sg13g2_xor2_1 _4703_ (.B(_1196_),
    .A(_1197_),
    .X(_1236_));
 sg13g2_and2_1 _4704_ (.A(_1235_),
    .B(net86),
    .X(_1237_));
 sg13g2_xor2_1 _4705_ (.B(_1236_),
    .A(_1235_),
    .X(_1238_));
 sg13g2_xnor2_1 _4706_ (.Y(_1239_),
    .A(_1234_),
    .B(_1238_));
 sg13g2_o21ai_1 _4707_ (.B1(_1226_),
    .Y(_1240_),
    .A1(_1239_),
    .A2(_1227_));
 sg13g2_xnor2_1 _4708_ (.Y(_1241_),
    .A(_1206_),
    .B(_1193_));
 sg13g2_nand2b_1 _4709_ (.Y(_1242_),
    .B(net65),
    .A_N(_1241_));
 sg13g2_a21oi_1 _4710_ (.A1(_1234_),
    .A2(net73),
    .Y(_1243_),
    .B1(_1237_));
 sg13g2_xor2_1 _4711_ (.B(_1240_),
    .A(_1241_),
    .X(_1245_));
 sg13g2_o21ai_1 _4712_ (.B1(_1242_),
    .Y(_1246_),
    .A1(_1243_),
    .A2(net63));
 sg13g2_xnor2_1 _4713_ (.Y(_1247_),
    .A(_1210_),
    .B(_1211_));
 sg13g2_nand2b_1 _4714_ (.Y(_1248_),
    .B(_1246_),
    .A_N(_1247_));
 sg13g2_xor2_1 _4715_ (.B(_1214_),
    .A(_1213_),
    .X(_1249_));
 sg13g2_nor2b_1 _4716_ (.A(_1248_),
    .B_N(_1249_),
    .Y(_1250_));
 sg13g2_xnor2_1 _4717_ (.Y(_1251_),
    .A(_1248_),
    .B(_1249_));
 sg13g2_o21ai_1 _4718_ (.B1(_1223_),
    .Y(_1252_),
    .A1(_0887_),
    .A2(net472));
 sg13g2_nor2b_1 _4719_ (.A(_1224_),
    .B_N(_1252_),
    .Y(_1253_));
 sg13g2_inv_1 _4720_ (.Y(_1254_),
    .A(_1253_));
 sg13g2_and2_1 _4721_ (.A(_0898_),
    .B(net414),
    .X(_1255_));
 sg13g2_nand2_1 _4722_ (.Y(_1256_),
    .A(net447),
    .B(net414));
 sg13g2_nand3_1 _4723_ (.B(net408),
    .C(_1255_),
    .A(\pid.Ki[2] ),
    .Y(_1257_));
 sg13g2_nand2_1 _4724_ (.Y(_1258_),
    .A(\pid.Ki[3] ),
    .B(net418));
 sg13g2_xor2_1 _4725_ (.B(_1256_),
    .A(_1228_),
    .X(_1259_));
 sg13g2_o21ai_1 _4726_ (.B1(_1257_),
    .Y(_1260_),
    .A1(_1258_),
    .A2(_1259_));
 sg13g2_nor2_1 _4727_ (.A(_0004_),
    .B(net471),
    .Y(_1261_));
 sg13g2_nand3_1 _4728_ (.B(net422),
    .C(_1261_),
    .A(\pid.Ki[4] ),
    .Y(_1262_));
 sg13g2_a21o_1 _4729_ (.A2(net422),
    .A1(net445),
    .B1(_1261_),
    .X(_1263_));
 sg13g2_and2_1 _4730_ (.A(_1262_),
    .B(_1263_),
    .X(_1264_));
 sg13g2_nand3_1 _4731_ (.B(net404),
    .C(_1264_),
    .A(net450),
    .Y(_1266_));
 sg13g2_nand2_1 _4732_ (.Y(_1267_),
    .A(_1262_),
    .B(_1266_));
 sg13g2_xnor2_1 _4733_ (.Y(_1268_),
    .A(_1230_),
    .B(_1231_));
 sg13g2_xnor2_1 _4734_ (.Y(_1269_),
    .A(_1267_),
    .B(_1268_));
 sg13g2_nor2b_1 _4735_ (.A(_1269_),
    .B_N(_1260_),
    .Y(_1270_));
 sg13g2_xor2_1 _4736_ (.B(_1269_),
    .A(_1260_),
    .X(_1271_));
 sg13g2_or2_1 _4737_ (.X(_1272_),
    .B(_1271_),
    .A(_1254_));
 sg13g2_xnor2_1 _4738_ (.Y(_1273_),
    .A(_1227_),
    .B(_1239_));
 sg13g2_nor2_1 _4739_ (.A(_1272_),
    .B(_1273_),
    .Y(_1274_));
 sg13g2_a21o_1 _4740_ (.A2(_1268_),
    .A1(_1267_),
    .B1(_1270_),
    .X(_1275_));
 sg13g2_xor2_1 _4741_ (.B(_1273_),
    .A(_1272_),
    .X(_1277_));
 sg13g2_a21oi_1 _4742_ (.A1(_1275_),
    .A2(_1277_),
    .Y(_1278_),
    .B1(_1274_));
 sg13g2_xor2_1 _4743_ (.B(_1245_),
    .A(_1243_),
    .X(_1279_));
 sg13g2_nand2b_1 _4744_ (.Y(_1280_),
    .B(_1279_),
    .A_N(_1278_));
 sg13g2_nand2_1 _4745_ (.Y(_1281_),
    .A(net446),
    .B(net404));
 sg13g2_nor2b_1 _4746_ (.A(_1279_),
    .B_N(_1278_),
    .Y(_1282_));
 sg13g2_xnor2_1 _4747_ (.Y(_1283_),
    .A(_1278_),
    .B(_1279_));
 sg13g2_o21ai_1 _4748_ (.B1(_1280_),
    .Y(_1284_),
    .A1(_1281_),
    .A2(_1282_));
 sg13g2_xnor2_1 _4749_ (.Y(_1285_),
    .A(_1246_),
    .B(_1247_));
 sg13g2_and2_1 _4750_ (.A(_1284_),
    .B(_1285_),
    .X(_1286_));
 sg13g2_or2_1 _4751_ (.X(_1288_),
    .B(_1285_),
    .A(_1284_));
 sg13g2_a21o_1 _4752_ (.A2(net404),
    .A1(net450),
    .B1(_1264_),
    .X(_1289_));
 sg13g2_and2_1 _4753_ (.A(_1266_),
    .B(_1289_),
    .X(_1290_));
 sg13g2_inv_1 _4754_ (.Y(_1291_),
    .A(_1290_));
 sg13g2_nor2_1 _4755_ (.A(_0003_),
    .B(net417),
    .Y(_1292_));
 sg13g2_nand3_1 _4756_ (.B(net414),
    .C(_1292_),
    .A(net447),
    .Y(_1293_));
 sg13g2_nand2_1 _4757_ (.Y(_1294_),
    .A(net446),
    .B(net424));
 sg13g2_a21o_1 _4758_ (.A2(net418),
    .A1(net447),
    .B1(_1255_),
    .X(_1295_));
 sg13g2_nand2_1 _4759_ (.Y(_1296_),
    .A(_1293_),
    .B(_1295_));
 sg13g2_o21ai_1 _4760_ (.B1(_1293_),
    .Y(_1297_),
    .A1(_1294_),
    .A2(_1296_));
 sg13g2_nor2_1 _4761_ (.A(_0005_),
    .B(net472),
    .Y(_1298_));
 sg13g2_nand3_1 _4762_ (.B(net408),
    .C(_1298_),
    .A(net450),
    .Y(_1299_));
 sg13g2_xor2_1 _4763_ (.B(_1259_),
    .A(_1258_),
    .X(_1300_));
 sg13g2_nor2b_1 _4764_ (.A(_1299_),
    .B_N(_1300_),
    .Y(_1301_));
 sg13g2_xnor2_1 _4765_ (.Y(_1302_),
    .A(_1299_),
    .B(_1300_));
 sg13g2_xnor2_1 _4766_ (.Y(_1303_),
    .A(_1297_),
    .B(_1302_));
 sg13g2_nor2_1 _4767_ (.A(_1291_),
    .B(_1303_),
    .Y(_1304_));
 sg13g2_xnor2_1 _4768_ (.Y(_1305_),
    .A(_1253_),
    .B(_1271_));
 sg13g2_and2_1 _4769_ (.A(_1304_),
    .B(_1305_),
    .X(_1306_));
 sg13g2_a21o_1 _4770_ (.A2(_1302_),
    .A1(_1297_),
    .B1(_1301_),
    .X(_1307_));
 sg13g2_xor2_1 _4771_ (.B(_1304_),
    .A(_1305_),
    .X(_1309_));
 sg13g2_a21oi_2 _4772_ (.B1(_1306_),
    .Y(_1310_),
    .A2(net58),
    .A1(_1307_));
 sg13g2_xnor2_1 _4773_ (.Y(_1311_),
    .A(_1275_),
    .B(_1277_));
 sg13g2_nor2_2 _4774_ (.A(_1310_),
    .B(_1311_),
    .Y(_1312_));
 sg13g2_xnor2_1 _4775_ (.Y(_1313_),
    .A(_1283_),
    .B(_1281_));
 sg13g2_nand2_1 _4776_ (.Y(_1314_),
    .A(_1312_),
    .B(_1313_));
 sg13g2_xnor2_1 _4777_ (.Y(_1315_),
    .A(_1291_),
    .B(_1303_));
 sg13g2_a21o_1 _4778_ (.A2(net408),
    .A1(net450),
    .B1(_1298_),
    .X(_1316_));
 sg13g2_nand2_1 _4779_ (.Y(_1317_),
    .A(_1299_),
    .B(_1316_));
 sg13g2_nand3_1 _4780_ (.B(net423),
    .C(_1292_),
    .A(net447),
    .Y(_1318_));
 sg13g2_nand2_1 _4781_ (.Y(_1320_),
    .A(net446),
    .B(_1605_));
 sg13g2_a21o_1 _4782_ (.A2(net423),
    .A1(net447),
    .B1(_1292_),
    .X(_1321_));
 sg13g2_and2_1 _4783_ (.A(_1318_),
    .B(_1321_),
    .X(_1322_));
 sg13g2_nand2b_1 _4784_ (.Y(_1323_),
    .B(_1322_),
    .A_N(_1320_));
 sg13g2_nand2_1 _4785_ (.Y(_1324_),
    .A(_1318_),
    .B(_1323_));
 sg13g2_xnor2_1 _4786_ (.Y(_1325_),
    .A(_1294_),
    .B(_1296_));
 sg13g2_nor2b_1 _4787_ (.A(_1325_),
    .B_N(_1324_),
    .Y(_1326_));
 sg13g2_xnor2_1 _4788_ (.Y(_1327_),
    .A(_1324_),
    .B(_1325_));
 sg13g2_nand2b_1 _4789_ (.Y(_1328_),
    .B(_1327_),
    .A_N(_1317_));
 sg13g2_xor2_1 _4790_ (.B(_1328_),
    .A(_1315_),
    .X(_1329_));
 sg13g2_nand2_1 _4791_ (.Y(_1330_),
    .A(_1326_),
    .B(_1329_));
 sg13g2_o21ai_1 _4792_ (.B1(_1330_),
    .Y(_1331_),
    .A1(_1315_),
    .A2(_1328_));
 sg13g2_xnor2_1 _4793_ (.Y(_1332_),
    .A(_1307_),
    .B(_1309_));
 sg13g2_nor2b_1 _4794_ (.A(_1332_),
    .B_N(_1331_),
    .Y(_1333_));
 sg13g2_xor2_1 _4795_ (.B(_1311_),
    .A(_1310_),
    .X(_1334_));
 sg13g2_and2_1 _4796_ (.A(_1333_),
    .B(_1334_),
    .X(_1335_));
 sg13g2_xor2_1 _4797_ (.B(_1332_),
    .A(_1331_),
    .X(_1336_));
 sg13g2_xnor2_1 _4798_ (.Y(_1337_),
    .A(_1326_),
    .B(_1329_));
 sg13g2_xnor2_1 _4799_ (.Y(_1338_),
    .A(_1317_),
    .B(_1327_));
 sg13g2_and4_1 _4800_ (.A(\pid.Ki[1] ),
    .B(net447),
    .C(_1605_),
    .D(net423),
    .X(_1339_));
 sg13g2_xnor2_1 _4801_ (.Y(_1341_),
    .A(_1320_),
    .B(_1322_));
 sg13g2_nand2_1 _4802_ (.Y(_1342_),
    .A(_1339_),
    .B(_1341_));
 sg13g2_nand2_1 _4803_ (.Y(_1343_),
    .A(net449),
    .B(net414));
 sg13g2_xnor2_1 _4804_ (.Y(_1344_),
    .A(_1339_),
    .B(_1341_));
 sg13g2_o21ai_1 _4805_ (.B1(_1342_),
    .Y(_1345_),
    .A1(_1343_),
    .A2(_1344_));
 sg13g2_nand2_1 _4806_ (.Y(_1346_),
    .A(_1338_),
    .B(_1345_));
 sg13g2_nor2_1 _4807_ (.A(_1337_),
    .B(_1346_),
    .Y(_1347_));
 sg13g2_nand2b_1 _4808_ (.Y(_1348_),
    .B(_1347_),
    .A_N(_1336_));
 sg13g2_xor2_1 _4809_ (.B(_1346_),
    .A(_1337_),
    .X(_1349_));
 sg13g2_nand2_1 _4810_ (.Y(_1350_),
    .A(net449),
    .B(net418));
 sg13g2_a22oi_1 _4811_ (.Y(_1352_),
    .B1(net423),
    .B2(\pid.Ki[1] ),
    .A2(_1605_),
    .A1(net447));
 sg13g2_nor2_1 _4812_ (.A(_1339_),
    .B(_1352_),
    .Y(_1353_));
 sg13g2_nor2b_1 _4813_ (.A(_1350_),
    .B_N(_1353_),
    .Y(_1354_));
 sg13g2_xor2_1 _4814_ (.B(_1344_),
    .A(_1343_),
    .X(_1355_));
 sg13g2_nand2_1 _4815_ (.Y(_1356_),
    .A(_1354_),
    .B(_1355_));
 sg13g2_xnor2_1 _4816_ (.Y(_1357_),
    .A(_1338_),
    .B(_1345_));
 sg13g2_nor2_1 _4817_ (.A(_1356_),
    .B(_1357_),
    .Y(_1358_));
 sg13g2_and2_1 _4818_ (.A(_1349_),
    .B(_1358_),
    .X(_1359_));
 sg13g2_nor2_1 _4819_ (.A(_0003_),
    .B(net471),
    .Y(_1360_));
 sg13g2_nand3_1 _4820_ (.B(net423),
    .C(_1360_),
    .A(net449),
    .Y(_1361_));
 sg13g2_xnor2_1 _4821_ (.Y(_1362_),
    .A(_1350_),
    .B(_1353_));
 sg13g2_nor2b_1 _4822_ (.A(_1361_),
    .B_N(_1362_),
    .Y(_1363_));
 sg13g2_xnor2_1 _4823_ (.Y(_1364_),
    .A(_1354_),
    .B(_1355_));
 sg13g2_inv_1 _4824_ (.Y(_1365_),
    .A(_1364_));
 sg13g2_nand2_1 _4825_ (.Y(_1366_),
    .A(_1363_),
    .B(_1365_));
 sg13g2_nor2_1 _4826_ (.A(_1357_),
    .B(_1366_),
    .Y(_1367_));
 sg13g2_or2_1 _4827_ (.X(_1368_),
    .B(_1358_),
    .A(_1349_));
 sg13g2_nand2b_1 _4828_ (.Y(_1369_),
    .B(_1368_),
    .A_N(_1359_));
 sg13g2_a21oi_1 _4829_ (.A1(_1367_),
    .A2(_1368_),
    .Y(_1370_),
    .B1(_1359_));
 sg13g2_xor2_1 _4830_ (.B(_1336_),
    .A(_1347_),
    .X(_1371_));
 sg13g2_o21ai_1 _4831_ (.B1(_1348_),
    .Y(_1373_),
    .A1(_1370_),
    .A2(_1371_));
 sg13g2_or2_1 _4832_ (.X(_1374_),
    .B(_1334_),
    .A(_1333_));
 sg13g2_nand2b_1 _4833_ (.Y(_1375_),
    .B(_1374_),
    .A_N(_1335_));
 sg13g2_a21oi_2 _4834_ (.B1(_1335_),
    .Y(_1376_),
    .A2(_1374_),
    .A1(_1373_));
 sg13g2_xnor2_1 _4835_ (.Y(_1377_),
    .A(_1313_),
    .B(_1312_));
 sg13g2_o21ai_1 _4836_ (.B1(_1314_),
    .Y(_1378_),
    .A1(_1376_),
    .A2(_1377_));
 sg13g2_a22oi_1 _4837_ (.Y(_1379_),
    .B1(_1312_),
    .B2(_1313_),
    .A2(_1285_),
    .A1(_1284_));
 sg13g2_o21ai_1 _4838_ (.B1(_1379_),
    .Y(_1380_),
    .A1(_1377_),
    .A2(_1376_));
 sg13g2_nand2_1 _4839_ (.Y(_1381_),
    .A(_1288_),
    .B(_1380_));
 sg13g2_and3_1 _4840_ (.X(_1382_),
    .A(_1251_),
    .B(_1380_),
    .C(_1288_));
 sg13g2_xor2_1 _4841_ (.B(_1216_),
    .A(_1215_),
    .X(_1383_));
 sg13g2_o21ai_1 _4842_ (.B1(_1383_),
    .Y(_1384_),
    .A1(_1382_),
    .A2(_1250_));
 sg13g2_nand2_1 _4843_ (.Y(_1385_),
    .A(_1217_),
    .B(_1384_));
 sg13g2_xnor2_1 _4844_ (.Y(_1386_),
    .A(_1178_),
    .B(_1179_));
 sg13g2_inv_1 _4845_ (.Y(_1387_),
    .A(_1386_));
 sg13g2_a21oi_1 _4846_ (.A1(_1385_),
    .A2(_1387_),
    .Y(_1388_),
    .B1(_1180_));
 sg13g2_a21o_1 _4847_ (.A2(_1180_),
    .A1(_1140_),
    .B1(_1141_),
    .X(_1389_));
 sg13g2_xor2_1 _4848_ (.B(_1139_),
    .A(_1138_),
    .X(_1390_));
 sg13g2_nand2b_1 _4849_ (.Y(_1391_),
    .B(_1390_),
    .A_N(_1386_));
 sg13g2_a21oi_2 _4850_ (.B1(_1391_),
    .Y(_1392_),
    .A2(_1217_),
    .A1(_1384_));
 sg13g2_nor2_1 _4851_ (.A(_1389_),
    .B(_1392_),
    .Y(_1394_));
 sg13g2_o21ai_1 _4852_ (.B1(_1097_),
    .Y(_1395_),
    .A1(_1392_),
    .A2(_1389_));
 sg13g2_xnor2_1 _4853_ (.Y(_1396_),
    .A(_1032_),
    .B(_1056_));
 sg13g2_a21o_1 _4854_ (.A2(_1096_),
    .A1(_1395_),
    .B1(_1396_),
    .X(_1397_));
 sg13g2_o21ai_1 _4855_ (.B1(_1052_),
    .Y(_1398_),
    .A1(_1034_),
    .A2(_1053_));
 sg13g2_o21ai_1 _4856_ (.B1(_1048_),
    .Y(_1399_),
    .A1(_1013_),
    .A2(_1049_));
 sg13g2_o21ai_1 _4857_ (.B1(_1041_),
    .Y(_1400_),
    .A1(_1016_),
    .A2(_1042_));
 sg13g2_o21ai_1 _4858_ (.B1(_1400_),
    .Y(_1401_),
    .A1(_0002_),
    .A2(_1016_));
 sg13g2_a21oi_1 _4859_ (.A1(net444),
    .A2(net390),
    .Y(_1402_),
    .B1(_1040_));
 sg13g2_o21ai_1 _4860_ (.B1(_1402_),
    .Y(_1403_),
    .A1(_0001_),
    .A2(net390));
 sg13g2_and2_1 _4861_ (.A(_1401_),
    .B(_1403_),
    .X(_1404_));
 sg13g2_nor2_1 _4862_ (.A(_0990_),
    .B(_1404_),
    .Y(_1405_));
 sg13g2_xnor2_1 _4863_ (.Y(_1406_),
    .A(_0990_),
    .B(_1404_));
 sg13g2_a21oi_1 _4864_ (.A1(_1044_),
    .A2(_1046_),
    .Y(_1407_),
    .B1(_1406_));
 sg13g2_nand3_1 _4865_ (.B(_1046_),
    .C(_1406_),
    .A(_1044_),
    .Y(_1408_));
 sg13g2_nor2b_1 _4866_ (.A(_1407_),
    .B_N(_1408_),
    .Y(_1409_));
 sg13g2_xnor2_1 _4867_ (.Y(_1410_),
    .A(_1013_),
    .B(_1409_));
 sg13g2_nand2_1 _4868_ (.Y(_1411_),
    .A(_1399_),
    .B(_1410_));
 sg13g2_xnor2_1 _4869_ (.Y(_1412_),
    .A(_1399_),
    .B(_1410_));
 sg13g2_xor2_1 _4870_ (.B(_1412_),
    .A(_1034_),
    .X(_1413_));
 sg13g2_nand2_1 _4871_ (.Y(_1415_),
    .A(_1398_),
    .B(_1413_));
 sg13g2_xnor2_1 _4872_ (.Y(_1416_),
    .A(_1398_),
    .B(_1413_));
 sg13g2_nor2_1 _4873_ (.A(_1055_),
    .B(_1416_),
    .Y(_1417_));
 sg13g2_xor2_1 _4874_ (.B(_1416_),
    .A(_1055_),
    .X(_1418_));
 sg13g2_inv_1 _4875_ (.Y(_1419_),
    .A(_1418_));
 sg13g2_a21o_2 _4876_ (.A2(_1058_),
    .A1(_1397_),
    .B1(_1419_),
    .X(_1420_));
 sg13g2_o21ai_1 _4877_ (.B1(_1411_),
    .Y(_1421_),
    .A1(_1034_),
    .A2(_1412_));
 sg13g2_xnor2_1 _4878_ (.Y(_1422_),
    .A(_1034_),
    .B(_1405_));
 sg13g2_nor2_1 _4879_ (.A(_1012_),
    .B(_1407_),
    .Y(_1423_));
 sg13g2_a21oi_1 _4880_ (.A1(_1012_),
    .A2(_1408_),
    .Y(_1424_),
    .B1(_1423_));
 sg13g2_xnor2_1 _4881_ (.Y(_1425_),
    .A(_1422_),
    .B(_1424_));
 sg13g2_xnor2_1 _4882_ (.Y(_1426_),
    .A(_1421_),
    .B(_1425_));
 sg13g2_xnor2_1 _4883_ (.Y(_1427_),
    .A(_1415_),
    .B(_1426_));
 sg13g2_nor2_2 _4884_ (.A(_1417_),
    .B(_1427_),
    .Y(_1428_));
 sg13g2_and2_2 _4885_ (.A(_1420_),
    .B(_1428_),
    .X(_1429_));
 sg13g2_inv_2 _4886_ (.Y(_1430_),
    .A(_1429_));
 sg13g2_xnor2_1 _4887_ (.Y(_1431_),
    .A(_1376_),
    .B(net72));
 sg13g2_xor2_1 _4888_ (.B(_1369_),
    .A(_1367_),
    .X(_1432_));
 sg13g2_xnor2_1 _4889_ (.Y(_1433_),
    .A(_1363_),
    .B(_1364_));
 sg13g2_a21o_1 _4890_ (.A2(net423),
    .A1(net449),
    .B1(_1360_),
    .X(_1434_));
 sg13g2_and2_1 _4891_ (.A(_1361_),
    .B(_1434_),
    .X(_1436_));
 sg13g2_nor2_2 _4892_ (.A(_0006_),
    .B(net471),
    .Y(_1437_));
 sg13g2_or2_1 _4893_ (.X(_1438_),
    .B(_1437_),
    .A(_1436_));
 sg13g2_xnor2_1 _4894_ (.Y(_1439_),
    .A(_1361_),
    .B(_1362_));
 sg13g2_or2_1 _4895_ (.X(_1440_),
    .B(_1439_),
    .A(_1438_));
 sg13g2_or2_1 _4896_ (.X(_1441_),
    .B(_1440_),
    .A(_1433_));
 sg13g2_and3_1 _4897_ (.X(_1442_),
    .A(_1356_),
    .B(_1357_),
    .C(_1366_));
 sg13g2_nor3_1 _4898_ (.A(_1358_),
    .B(_1367_),
    .C(_1442_),
    .Y(_1443_));
 sg13g2_nor2_1 _4899_ (.A(_1441_),
    .B(_1443_),
    .Y(_1444_));
 sg13g2_nand2_1 _4900_ (.Y(_1445_),
    .A(_1432_),
    .B(_1444_));
 sg13g2_xor2_1 _4901_ (.B(net64),
    .A(_1370_),
    .X(_1446_));
 sg13g2_or2_1 _4902_ (.X(_1447_),
    .B(_1446_),
    .A(_1445_));
 sg13g2_xor2_1 _4903_ (.B(_1375_),
    .A(_1373_),
    .X(_1448_));
 sg13g2_nand2b_1 _4904_ (.Y(_1449_),
    .B(_1448_),
    .A_N(_1447_));
 sg13g2_nand2_1 _4905_ (.Y(_1450_),
    .A(net378),
    .B(_1449_));
 sg13g2_xor2_1 _4906_ (.B(_1450_),
    .A(_1431_),
    .X(_1451_));
 sg13g2_or3_1 _4907_ (.A(_1250_),
    .B(_1382_),
    .C(_1383_),
    .X(_1452_));
 sg13g2_and2_1 _4908_ (.A(_1384_),
    .B(_1452_),
    .X(_1453_));
 sg13g2_nor2b_1 _4909_ (.A(_1286_),
    .B_N(_1288_),
    .Y(_1454_));
 sg13g2_xnor2_1 _4910_ (.Y(_1455_),
    .A(_1378_),
    .B(_1454_));
 sg13g2_nand2b_1 _4911_ (.Y(_1457_),
    .B(_1431_),
    .A_N(_1449_));
 sg13g2_nand2_1 _4912_ (.Y(_1458_),
    .A(net378),
    .B(_1457_));
 sg13g2_xor2_1 _4913_ (.B(_1458_),
    .A(_1455_),
    .X(_1459_));
 sg13g2_nor2b_1 _4914_ (.A(_1457_),
    .B_N(_1455_),
    .Y(_1460_));
 sg13g2_xnor2_1 _4915_ (.Y(_1461_),
    .A(_1251_),
    .B(_1381_));
 sg13g2_nand2b_1 _4916_ (.Y(_1462_),
    .B(_1460_),
    .A_N(_1461_));
 sg13g2_nand3_1 _4917_ (.B(_1428_),
    .C(_1462_),
    .A(_1420_),
    .Y(_1463_));
 sg13g2_xnor2_1 _4918_ (.Y(_1464_),
    .A(_1463_),
    .B(_1453_));
 sg13g2_xor2_1 _4919_ (.B(_1463_),
    .A(_1453_),
    .X(_1465_));
 sg13g2_xnor2_1 _4920_ (.Y(_1466_),
    .A(_1388_),
    .B(_1390_));
 sg13g2_or2_1 _4921_ (.X(_1467_),
    .B(_1462_),
    .A(_1453_));
 sg13g2_xnor2_1 _4922_ (.Y(_1468_),
    .A(_1385_),
    .B(_1386_));
 sg13g2_nor3_1 _4923_ (.A(_1453_),
    .B(_1462_),
    .C(_1468_),
    .Y(_1469_));
 sg13g2_inv_1 _4924_ (.Y(_1470_),
    .A(_1469_));
 sg13g2_nand3_1 _4925_ (.B(_1428_),
    .C(_1470_),
    .A(_1420_),
    .Y(_1471_));
 sg13g2_xnor2_1 _4926_ (.Y(_1472_),
    .A(_1471_),
    .B(_1466_));
 sg13g2_nand3_1 _4927_ (.B(_1428_),
    .C(_1467_),
    .A(_1420_),
    .Y(_1473_));
 sg13g2_xnor2_1 _4928_ (.Y(_1474_),
    .A(_1468_),
    .B(_1473_));
 sg13g2_inv_1 _4929_ (.Y(_1475_),
    .A(_1474_));
 sg13g2_nor2_1 _4930_ (.A(_1472_),
    .B(_1474_),
    .Y(_1476_));
 sg13g2_or3_1 _4931_ (.A(_1464_),
    .B(_1474_),
    .C(_1472_),
    .X(_1478_));
 sg13g2_nor2b_1 _4932_ (.A(_1466_),
    .B_N(_1469_),
    .Y(_1479_));
 sg13g2_xor2_1 _4933_ (.B(_1394_),
    .A(_1097_),
    .X(_1480_));
 sg13g2_nand3b_1 _4934_ (.B(_1469_),
    .C(_1480_),
    .Y(_1481_),
    .A_N(_1466_));
 sg13g2_nand3_1 _4935_ (.B(_1428_),
    .C(_1481_),
    .A(_1420_),
    .Y(_1482_));
 sg13g2_nor2_1 _4936_ (.A(_1479_),
    .B(_1480_),
    .Y(_1483_));
 sg13g2_a21o_1 _4937_ (.A2(_1428_),
    .A1(_1420_),
    .B1(_1480_),
    .X(_1484_));
 sg13g2_o21ai_1 _4938_ (.B1(_1484_),
    .Y(_1485_),
    .A1(_1482_),
    .A2(_1483_));
 sg13g2_nand3_1 _4939_ (.B(_1395_),
    .C(_1396_),
    .A(_1096_),
    .Y(_1486_));
 sg13g2_and2_1 _4940_ (.A(_1397_),
    .B(_1486_),
    .X(_1487_));
 sg13g2_xnor2_1 _4941_ (.Y(_1488_),
    .A(_1482_),
    .B(_1487_));
 sg13g2_and2_1 _4942_ (.A(_1485_),
    .B(_1488_),
    .X(_1489_));
 sg13g2_nand2_1 _4943_ (.Y(_1490_),
    .A(_1478_),
    .B(_1489_));
 sg13g2_o21ai_1 _4944_ (.B1(_1428_),
    .Y(_1491_),
    .A1(_1481_),
    .A2(_1487_));
 sg13g2_nand3_1 _4945_ (.B(_1397_),
    .C(_1419_),
    .A(_1058_),
    .Y(_1492_));
 sg13g2_and3_1 _4946_ (.X(_1493_),
    .A(_1420_),
    .B(_1491_),
    .C(_1492_));
 sg13g2_a21o_2 _4947_ (.A2(_1478_),
    .A1(_1489_),
    .B1(_1493_),
    .X(_1494_));
 sg13g2_and2_1 _4948_ (.A(_1465_),
    .B(_1494_),
    .X(_1495_));
 sg13g2_xnor2_1 _4949_ (.Y(_1496_),
    .A(_1494_),
    .B(_1464_));
 sg13g2_nor2_1 _4950_ (.A(_1430_),
    .B(_1460_),
    .Y(_1497_));
 sg13g2_xnor2_1 _4951_ (.Y(_1499_),
    .A(_1461_),
    .B(_1497_));
 sg13g2_nand3_1 _4952_ (.B(_1475_),
    .C(_1494_),
    .A(_1465_),
    .Y(_1500_));
 sg13g2_xnor2_1 _4953_ (.Y(_1501_),
    .A(_1475_),
    .B(_1495_));
 sg13g2_and2_1 _4954_ (.A(_1496_),
    .B(_1499_),
    .X(_1502_));
 sg13g2_nand2_2 _4955_ (.Y(_1503_),
    .A(_1496_),
    .B(_1499_));
 sg13g2_a21o_1 _4956_ (.A2(_1503_),
    .A1(_1472_),
    .B1(_1501_),
    .X(_1504_));
 sg13g2_and2_1 _4957_ (.A(_1472_),
    .B(_1500_),
    .X(_1505_));
 sg13g2_a22oi_1 _4958_ (.Y(_1506_),
    .B1(_1500_),
    .B2(_1472_),
    .A2(_1495_),
    .A1(_1476_));
 sg13g2_a21o_1 _4959_ (.A2(_1495_),
    .A1(_1476_),
    .B1(_1505_),
    .X(_1507_));
 sg13g2_nand2_1 _4960_ (.Y(_1508_),
    .A(_1478_),
    .B(_1494_));
 sg13g2_xor2_1 _4961_ (.B(_1508_),
    .A(_1485_),
    .X(_1509_));
 sg13g2_a21oi_1 _4962_ (.A1(_1501_),
    .A2(_1506_),
    .Y(_1510_),
    .B1(_1509_));
 sg13g2_a22oi_1 _4963_ (.Y(_1511_),
    .B1(_1504_),
    .B2(_1510_),
    .A2(_1490_),
    .A1(_1488_));
 sg13g2_nand2b_1 _4964_ (.Y(_1512_),
    .B(_1511_),
    .A_N(_1499_));
 sg13g2_nor2b_1 _4965_ (.A(_1511_),
    .B_N(_1499_),
    .Y(_1513_));
 sg13g2_nor2_1 _4966_ (.A(_1503_),
    .B(_1511_),
    .Y(_1514_));
 sg13g2_xnor2_1 _4967_ (.Y(_1515_),
    .A(_1514_),
    .B(_1501_));
 sg13g2_a21oi_1 _4968_ (.A1(_1475_),
    .A2(_1502_),
    .Y(_1516_),
    .B1(_1511_));
 sg13g2_nand2_1 _4969_ (.Y(_1517_),
    .A(_1507_),
    .B(_1516_));
 sg13g2_xnor2_1 _4970_ (.Y(_1518_),
    .A(_1507_),
    .B(_1516_));
 sg13g2_xnor2_1 _4971_ (.Y(_1520_),
    .A(_1511_),
    .B(_1499_));
 sg13g2_nor2b_1 _4972_ (.A(_1459_),
    .B_N(_1496_),
    .Y(_1521_));
 sg13g2_and2_1 _4973_ (.A(_1521_),
    .B(_1520_),
    .X(_1522_));
 sg13g2_nor3_1 _4974_ (.A(_1515_),
    .B(_1518_),
    .C(_1522_),
    .Y(_1523_));
 sg13g2_or3_1 _4975_ (.A(_1515_),
    .B(_1522_),
    .C(_1518_),
    .X(_1524_));
 sg13g2_xor2_1 _4976_ (.B(_1517_),
    .A(_1509_),
    .X(_1525_));
 sg13g2_xnor2_1 _4977_ (.Y(_1526_),
    .A(_1509_),
    .B(_1517_));
 sg13g2_nor2_2 _4978_ (.A(_1523_),
    .B(_1525_),
    .Y(_1527_));
 sg13g2_a21oi_2 _4979_ (.B1(_1459_),
    .Y(_1528_),
    .A2(_1526_),
    .A1(_1524_));
 sg13g2_o21ai_1 _4980_ (.B1(_1512_),
    .Y(_1529_),
    .A1(_1528_),
    .A2(_1513_));
 sg13g2_xor2_1 _4981_ (.B(_1529_),
    .A(_1496_),
    .X(_1530_));
 sg13g2_inv_1 _4982_ (.Y(_1531_),
    .A(_1530_));
 sg13g2_xor2_1 _4983_ (.B(_1527_),
    .A(_1459_),
    .X(_1532_));
 sg13g2_xnor2_1 _4984_ (.Y(_1533_),
    .A(_1459_),
    .B(_1527_));
 sg13g2_nor2b_1 _4985_ (.A(_1451_),
    .B_N(_1520_),
    .Y(_1534_));
 sg13g2_and2_1 _4986_ (.A(_1532_),
    .B(_1534_),
    .X(_1535_));
 sg13g2_a21o_1 _4987_ (.A2(_1526_),
    .A1(_1524_),
    .B1(_1522_),
    .X(_1536_));
 sg13g2_xor2_1 _4988_ (.B(_1536_),
    .A(net56),
    .X(_1537_));
 sg13g2_xnor2_1 _4989_ (.Y(_1538_),
    .A(_1515_),
    .B(_1536_));
 sg13g2_a21oi_1 _4990_ (.A1(_1532_),
    .A2(_1534_),
    .Y(_1539_),
    .B1(_1538_));
 sg13g2_nand2_1 _4991_ (.Y(_1541_),
    .A(_1530_),
    .B(_1539_));
 sg13g2_o21ai_1 _4992_ (.B1(_1518_),
    .Y(_1542_),
    .A1(net56),
    .A2(_1536_));
 sg13g2_a22oi_1 _4993_ (.Y(_1543_),
    .B1(_1542_),
    .B2(_1524_),
    .A2(_1530_),
    .A1(_1539_));
 sg13g2_xnor2_1 _4994_ (.Y(_1544_),
    .A(_1543_),
    .B(_1451_));
 sg13g2_inv_4 _4995_ (.A(_1544_),
    .Y(_1545_));
 sg13g2_nand2_1 _4996_ (.Y(_1546_),
    .A(net378),
    .B(_1447_));
 sg13g2_xor2_1 _4997_ (.B(_1546_),
    .A(_1448_),
    .X(_1547_));
 sg13g2_inv_1 _4998_ (.Y(_1548_),
    .A(_1547_));
 sg13g2_nor3_2 _4999_ (.A(_1451_),
    .B(_1533_),
    .C(_1543_),
    .Y(_1549_));
 sg13g2_or3_1 _5000_ (.A(_1520_),
    .B(_1528_),
    .C(_1549_),
    .X(_1550_));
 sg13g2_o21ai_1 _5001_ (.B1(_1520_),
    .Y(_1551_),
    .A1(_1528_),
    .A2(_1549_));
 sg13g2_nand2_1 _5002_ (.Y(_1552_),
    .A(_1550_),
    .B(_1551_));
 sg13g2_nor3_1 _5003_ (.A(_1531_),
    .B(_1535_),
    .C(_1543_),
    .Y(_1553_));
 sg13g2_o21ai_1 _5004_ (.B1(_1531_),
    .Y(_1554_),
    .A1(_1535_),
    .A2(_1543_));
 sg13g2_nand2b_1 _5005_ (.Y(_1555_),
    .B(_1554_),
    .A_N(_1553_));
 sg13g2_nor2_1 _5006_ (.A(_1533_),
    .B(_1547_),
    .Y(_1556_));
 sg13g2_nand2_1 _5007_ (.Y(_1557_),
    .A(_1545_),
    .B(_1556_));
 sg13g2_a21oi_1 _5008_ (.A1(_1545_),
    .A2(_1556_),
    .Y(_1558_),
    .B1(_1555_));
 sg13g2_a221oi_1 _5009_ (.B2(_1545_),
    .C1(_1555_),
    .B1(_1556_),
    .A1(_1551_),
    .Y(_1559_),
    .A2(_1550_));
 sg13g2_o21ai_1 _5010_ (.B1(_1541_),
    .Y(_1560_),
    .A1(_1537_),
    .A2(_1553_));
 sg13g2_inv_1 _5011_ (.Y(_1562_),
    .A(_1560_));
 sg13g2_nand2b_1 _5012_ (.Y(_1563_),
    .B(_1560_),
    .A_N(_1559_));
 sg13g2_o21ai_1 _5013_ (.B1(_1548_),
    .Y(_1564_),
    .A1(_1562_),
    .A2(_1559_));
 sg13g2_nand3b_1 _5014_ (.B(_1560_),
    .C(_1547_),
    .Y(_1565_),
    .A_N(_1559_));
 sg13g2_nand2_2 _5015_ (.Y(_1566_),
    .A(_1564_),
    .B(_1565_));
 sg13g2_inv_1 _5016_ (.Y(_1567_),
    .A(_1566_));
 sg13g2_nand2_1 _5017_ (.Y(_1568_),
    .A(net378),
    .B(_1445_));
 sg13g2_xor2_1 _5018_ (.B(_1568_),
    .A(_1446_),
    .X(_1569_));
 sg13g2_inv_1 _5019_ (.Y(_1570_),
    .A(_1569_));
 sg13g2_and2_1 _5020_ (.A(_1557_),
    .B(_1563_),
    .X(_1571_));
 sg13g2_nand2_1 _5021_ (.Y(_1573_),
    .A(_1552_),
    .B(_1571_));
 sg13g2_xnor2_1 _5022_ (.Y(_1574_),
    .A(_1552_),
    .B(_1571_));
 sg13g2_xnor2_1 _5023_ (.Y(_1575_),
    .A(_1564_),
    .B(_1545_));
 sg13g2_o21ai_1 _5024_ (.B1(_1533_),
    .Y(_1576_),
    .A1(_1451_),
    .A2(_1543_));
 sg13g2_nor2b_1 _5025_ (.A(_1549_),
    .B_N(_1576_),
    .Y(_1577_));
 sg13g2_o21ai_1 _5026_ (.B1(_1577_),
    .Y(_1578_),
    .A1(_1544_),
    .A2(_1564_));
 sg13g2_or3_1 _5027_ (.A(_1544_),
    .B(_1564_),
    .C(_1577_),
    .X(_1579_));
 sg13g2_and2_1 _5028_ (.A(_1578_),
    .B(_1579_),
    .X(_1580_));
 sg13g2_nand3b_1 _5029_ (.B(_1578_),
    .C(_1579_),
    .Y(_1581_),
    .A_N(_1575_));
 sg13g2_nor2_1 _5030_ (.A(_1566_),
    .B(_1570_),
    .Y(_1582_));
 sg13g2_nand3_1 _5031_ (.B(_1565_),
    .C(_1569_),
    .A(_1564_),
    .Y(_1584_));
 sg13g2_nand3b_1 _5032_ (.B(_1584_),
    .C(_1575_),
    .Y(_1585_),
    .A_N(_1577_));
 sg13g2_a21o_1 _5033_ (.A2(_1581_),
    .A1(_1585_),
    .B1(_1574_),
    .X(_1586_));
 sg13g2_and2_1 _5034_ (.A(_1555_),
    .B(_1573_),
    .X(_1587_));
 sg13g2_a21oi_2 _5035_ (.B1(_1559_),
    .Y(_1588_),
    .A2(_1587_),
    .A1(_1586_));
 sg13g2_a221oi_1 _5036_ (.B2(_1586_),
    .C1(_1570_),
    .B1(_1587_),
    .A1(_1552_),
    .Y(_1589_),
    .A2(_1558_));
 sg13g2_nand2_1 _5037_ (.Y(_1590_),
    .A(_1569_),
    .B(_1588_));
 sg13g2_nand3_1 _5038_ (.B(_1567_),
    .C(_1545_),
    .A(_1589_),
    .Y(_1591_));
 sg13g2_a21o_1 _5039_ (.A2(_1589_),
    .A1(_1567_),
    .B1(_1575_),
    .X(_1592_));
 sg13g2_and2_1 _5040_ (.A(_1591_),
    .B(_1592_),
    .X(_1593_));
 sg13g2_nor2_1 _5041_ (.A(_1569_),
    .B(_1588_),
    .Y(_1595_));
 sg13g2_xnor2_1 _5042_ (.Y(_1596_),
    .A(_1570_),
    .B(_1588_));
 sg13g2_nor2_1 _5043_ (.A(_1430_),
    .B(_1444_),
    .Y(_1597_));
 sg13g2_xnor2_1 _5044_ (.Y(_1598_),
    .A(_1432_),
    .B(_1597_));
 sg13g2_inv_1 _5045_ (.Y(_1599_),
    .A(_1598_));
 sg13g2_nor2_1 _5046_ (.A(_1566_),
    .B(_1598_),
    .Y(_1600_));
 sg13g2_nand2_1 _5047_ (.Y(_1601_),
    .A(_1596_),
    .B(_1600_));
 sg13g2_inv_1 _5048_ (.Y(_1602_),
    .A(_1601_));
 sg13g2_a221oi_1 _5049_ (.B2(_1587_),
    .C1(_1559_),
    .B1(_1586_),
    .A1(_1575_),
    .Y(_1603_),
    .A2(_1582_));
 sg13g2_nand2_1 _5050_ (.Y(_1604_),
    .A(_1580_),
    .B(_1603_));
 sg13g2_xnor2_1 _5051_ (.Y(_1606_),
    .A(_1580_),
    .B(_1603_));
 sg13g2_a221oi_1 _5052_ (.B2(_1600_),
    .C1(_1606_),
    .B1(_1596_),
    .A1(_1592_),
    .Y(_1607_),
    .A2(_1591_));
 sg13g2_xor2_1 _5053_ (.B(_1604_),
    .A(_1574_),
    .X(_1608_));
 sg13g2_xnor2_1 _5054_ (.Y(_1609_),
    .A(_1574_),
    .B(_1604_));
 sg13g2_nor2_2 _5055_ (.A(_1607_),
    .B(_1608_),
    .Y(_1610_));
 sg13g2_nand2b_1 _5056_ (.Y(_1611_),
    .B(_1609_),
    .A_N(_1607_));
 sg13g2_o21ai_1 _5057_ (.B1(_1599_),
    .Y(_1612_),
    .A1(_1608_),
    .A2(_1607_));
 sg13g2_a21oi_2 _5058_ (.B1(_1595_),
    .Y(_1613_),
    .A2(_1590_),
    .A1(_1612_));
 sg13g2_xnor2_1 _5059_ (.Y(_1614_),
    .A(_1613_),
    .B(_1566_));
 sg13g2_nand3b_1 _5060_ (.B(_1609_),
    .C(_1598_),
    .Y(_1615_),
    .A_N(_1607_));
 sg13g2_and2_1 _5061_ (.A(_1612_),
    .B(_1615_),
    .X(_1616_));
 sg13g2_nand2_1 _5062_ (.Y(_1617_),
    .A(net377),
    .B(_1441_));
 sg13g2_xnor2_1 _5063_ (.Y(_1618_),
    .A(_1443_),
    .B(_1617_));
 sg13g2_inv_1 _5064_ (.Y(_1619_),
    .A(_1618_));
 sg13g2_and2_1 _5065_ (.A(_1616_),
    .B(_1619_),
    .X(_1620_));
 sg13g2_nand4_1 _5066_ (.B(_1612_),
    .C(_1615_),
    .A(_1596_),
    .Y(_1621_),
    .D(_1619_));
 sg13g2_nand3b_1 _5067_ (.B(_1601_),
    .C(_1611_),
    .Y(_1622_),
    .A_N(_1593_));
 sg13g2_o21ai_1 _5068_ (.B1(_1593_),
    .Y(_1623_),
    .A1(_1602_),
    .A2(_1610_));
 sg13g2_nand2_1 _5069_ (.Y(_1624_),
    .A(_1622_),
    .B(_1623_));
 sg13g2_nand3_1 _5070_ (.B(_1622_),
    .C(_1623_),
    .A(_1621_),
    .Y(_1625_));
 sg13g2_nor2_1 _5071_ (.A(_1614_),
    .B(_1625_),
    .Y(_1627_));
 sg13g2_a21o_1 _5072_ (.A2(_1622_),
    .A1(_1606_),
    .B1(_1607_),
    .X(_1628_));
 sg13g2_nor2b_2 _5073_ (.A(_1627_),
    .B_N(_1628_),
    .Y(_1629_));
 sg13g2_o21ai_1 _5074_ (.B1(_1628_),
    .Y(_1630_),
    .A1(_1625_),
    .A2(_1614_));
 sg13g2_a22oi_1 _5075_ (.Y(_1631_),
    .B1(_1620_),
    .B2(_1630_),
    .A2(_1611_),
    .A1(_1599_));
 sg13g2_xnor2_1 _5076_ (.Y(_1632_),
    .A(_1596_),
    .B(_1631_));
 sg13g2_nand2_1 _5077_ (.Y(_1633_),
    .A(_1621_),
    .B(_1630_));
 sg13g2_xor2_1 _5078_ (.B(_1633_),
    .A(_1614_),
    .X(_1634_));
 sg13g2_nor2_1 _5079_ (.A(_1618_),
    .B(_1629_),
    .Y(_1635_));
 sg13g2_xnor2_1 _5080_ (.Y(_1636_),
    .A(_1630_),
    .B(_1619_));
 sg13g2_inv_1 _5081_ (.Y(_1638_),
    .A(_1636_));
 sg13g2_nand3_1 _5082_ (.B(_1433_),
    .C(_1440_),
    .A(net377),
    .Y(_1639_));
 sg13g2_a21o_1 _5083_ (.A2(_1440_),
    .A1(net377),
    .B1(_1433_),
    .X(_1640_));
 sg13g2_and2_1 _5084_ (.A(_1639_),
    .B(_1640_),
    .X(_1641_));
 sg13g2_nor2b_1 _5085_ (.A(_1641_),
    .B_N(_1616_),
    .Y(_1642_));
 sg13g2_nor2b_1 _5086_ (.A(_1636_),
    .B_N(_1642_),
    .Y(_1643_));
 sg13g2_nand2b_1 _5087_ (.Y(_1644_),
    .B(_1642_),
    .A_N(_1636_));
 sg13g2_nand3b_1 _5088_ (.B(_1634_),
    .C(_1644_),
    .Y(_1645_),
    .A_N(_1632_));
 sg13g2_o21ai_1 _5089_ (.B1(_1624_),
    .Y(_1646_),
    .A1(_1614_),
    .A2(_1633_));
 sg13g2_nand2b_2 _5090_ (.Y(_1647_),
    .B(_1646_),
    .A_N(_1627_));
 sg13g2_and2_1 _5091_ (.A(_1645_),
    .B(_1647_),
    .X(_1649_));
 sg13g2_nand2_1 _5092_ (.Y(_1650_),
    .A(_1645_),
    .B(_1647_));
 sg13g2_a221oi_1 _5093_ (.B2(_1647_),
    .C1(_1632_),
    .B1(_1645_),
    .A1(_1638_),
    .Y(_1651_),
    .A2(_1642_));
 sg13g2_nor2_1 _5094_ (.A(_1634_),
    .B(_1651_),
    .Y(_1652_));
 sg13g2_or2_1 _5095_ (.X(_1653_),
    .B(_1651_),
    .A(_1634_));
 sg13g2_and2_1 _5096_ (.A(_1645_),
    .B(_1653_),
    .X(_1654_));
 sg13g2_nand2_1 _5097_ (.Y(_1655_),
    .A(_1645_),
    .B(_1653_));
 sg13g2_a21oi_2 _5098_ (.B1(_1641_),
    .Y(_1656_),
    .A2(_1647_),
    .A1(_1645_));
 sg13g2_and3_1 _5099_ (.X(_1657_),
    .A(_1641_),
    .B(_1645_),
    .C(_1647_));
 sg13g2_or2_1 _5100_ (.X(_1658_),
    .B(_1657_),
    .A(_1656_));
 sg13g2_nand2_1 _5101_ (.Y(_1660_),
    .A(net377),
    .B(_1438_));
 sg13g2_xnor2_1 _5102_ (.Y(_1661_),
    .A(_1439_),
    .B(_1660_));
 sg13g2_nor2_1 _5103_ (.A(_1658_),
    .B(_1661_),
    .Y(_1662_));
 sg13g2_a221oi_1 _5104_ (.B2(_1645_),
    .C1(_1636_),
    .B1(_1647_),
    .A1(_1639_),
    .Y(_1663_),
    .A2(_1640_));
 sg13g2_xnor2_1 _5105_ (.Y(_1664_),
    .A(_1636_),
    .B(_1656_));
 sg13g2_nor4_1 _5106_ (.A(_1636_),
    .B(_1656_),
    .C(_1657_),
    .D(_1661_),
    .Y(_1665_));
 sg13g2_or3_1 _5107_ (.A(_1616_),
    .B(_1635_),
    .C(_1663_),
    .X(_1666_));
 sg13g2_o21ai_1 _5108_ (.B1(_1616_),
    .Y(_1667_),
    .A1(_1663_),
    .A2(_1635_));
 sg13g2_and2_1 _5109_ (.A(_1666_),
    .B(_1667_),
    .X(_1668_));
 sg13g2_a21oi_1 _5110_ (.A1(_1666_),
    .A2(_1667_),
    .Y(_1669_),
    .B1(_1665_));
 sg13g2_a21o_1 _5111_ (.A2(_1666_),
    .A1(_1667_),
    .B1(_1665_),
    .X(_1671_));
 sg13g2_o21ai_1 _5112_ (.B1(_1632_),
    .Y(_1672_),
    .A1(_1643_),
    .A2(_1649_));
 sg13g2_and2_1 _5113_ (.A(_1652_),
    .B(_1672_),
    .X(_1673_));
 sg13g2_nand2_1 _5114_ (.Y(_1674_),
    .A(_1669_),
    .B(_1673_));
 sg13g2_a21oi_2 _5115_ (.B1(_1654_),
    .Y(_1675_),
    .A2(_1673_),
    .A1(_1669_));
 sg13g2_nand2b_1 _5116_ (.Y(_1676_),
    .B(_1672_),
    .A_N(_1651_));
 sg13g2_o21ai_1 _5117_ (.B1(_1676_),
    .Y(_1677_),
    .A1(_1671_),
    .A2(_1655_));
 sg13g2_nand2_1 _5118_ (.Y(_1678_),
    .A(net377),
    .B(_1437_));
 sg13g2_xor2_1 _5119_ (.B(_1678_),
    .A(_1436_),
    .X(_1679_));
 sg13g2_inv_1 _5120_ (.Y(_1680_),
    .A(_1679_));
 sg13g2_nor4_1 _5121_ (.A(_1656_),
    .B(_1657_),
    .C(_1661_),
    .D(_1680_),
    .Y(_1681_));
 sg13g2_or2_1 _5122_ (.X(_1682_),
    .B(_1681_),
    .A(_1664_));
 sg13g2_o21ai_1 _5123_ (.B1(_1676_),
    .Y(_1683_),
    .A1(_1668_),
    .A2(_1682_));
 sg13g2_a22oi_1 _5124_ (.Y(_1684_),
    .B1(_1683_),
    .B2(_1675_),
    .A2(_1674_),
    .A1(_1677_));
 sg13g2_nand2_2 _5125_ (.Y(_1685_),
    .A(_1684_),
    .B(_1675_));
 sg13g2_nand2_2 _5126_ (.Y(_1686_),
    .A(net378),
    .B(_1685_));
 sg13g2_o21ai_1 _5127_ (.B1(net378),
    .Y(_1687_),
    .A1(_1650_),
    .A2(_1685_));
 sg13g2_o21ai_1 _5128_ (.B1(_1687_),
    .Y(_1688_),
    .A1(_1430_),
    .A2(_1629_));
 sg13g2_a21oi_1 _5129_ (.A1(net377),
    .A2(_1611_),
    .Y(_1689_),
    .B1(_1688_));
 sg13g2_nand2_1 _5130_ (.Y(_1690_),
    .A(net377),
    .B(_1588_));
 sg13g2_nand2_1 _5131_ (.Y(_1692_),
    .A(_1689_),
    .B(_1690_));
 sg13g2_a21oi_1 _5132_ (.A1(_1429_),
    .A2(_1563_),
    .Y(_1693_),
    .B1(_1692_));
 sg13g2_nor2_1 _5133_ (.A(_1430_),
    .B(_1543_),
    .Y(_1694_));
 sg13g2_nor2b_1 _5134_ (.A(_1694_),
    .B_N(_1693_),
    .Y(_1695_));
 sg13g2_o21ai_1 _5135_ (.B1(net378),
    .Y(_1696_),
    .A1(_1523_),
    .A2(_1525_));
 sg13g2_and2_1 _5136_ (.A(_1695_),
    .B(_1696_),
    .X(_1697_));
 sg13g2_o21ai_1 _5137_ (.B1(_1697_),
    .Y(_1698_),
    .A1(_1430_),
    .A2(_1511_));
 sg13g2_a21o_1 _5138_ (.A2(_1494_),
    .A1(net377),
    .B1(_1698_),
    .X(_1699_));
 sg13g2_nand2_1 _5139_ (.Y(_1700_),
    .A(\pid.integral[12] ),
    .B(net369));
 sg13g2_nor2b_1 _5140_ (.A(_0007_),
    .B_N(net369),
    .Y(_1701_));
 sg13g2_xor2_1 _5141_ (.B(_1698_),
    .A(_1494_),
    .X(_1703_));
 sg13g2_nand2_1 _5142_ (.Y(_1704_),
    .A(\pid.integral[10] ),
    .B(_1703_));
 sg13g2_xnor2_1 _5143_ (.Y(_1705_),
    .A(_1511_),
    .B(_1697_));
 sg13g2_nor2_1 _5144_ (.A(_0008_),
    .B(_1705_),
    .Y(_1706_));
 sg13g2_nand2_1 _5145_ (.Y(_1707_),
    .A(_0008_),
    .B(_1705_));
 sg13g2_nand2b_1 _5146_ (.Y(_1708_),
    .B(_1707_),
    .A_N(_1706_));
 sg13g2_xnor2_1 _5147_ (.Y(_1709_),
    .A(_1527_),
    .B(_1695_));
 sg13g2_inv_1 _5148_ (.Y(_1710_),
    .A(_1709_));
 sg13g2_nand2_1 _5149_ (.Y(_1711_),
    .A(\pid.integral[8] ),
    .B(_1710_));
 sg13g2_xnor2_1 _5150_ (.Y(_1712_),
    .A(_1543_),
    .B(_1693_));
 sg13g2_nor2_1 _5151_ (.A(_0009_),
    .B(_1712_),
    .Y(_1714_));
 sg13g2_xor2_1 _5152_ (.B(_1692_),
    .A(_1563_),
    .X(_1715_));
 sg13g2_nand2_1 _5153_ (.Y(_1716_),
    .A(\pid.integral[6] ),
    .B(_1715_));
 sg13g2_xnor2_1 _5154_ (.Y(_1717_),
    .A(_1588_),
    .B(_1689_));
 sg13g2_nor2b_1 _5155_ (.A(_0010_),
    .B_N(_1717_),
    .Y(_1718_));
 sg13g2_xnor2_1 _5156_ (.Y(_1719_),
    .A(_0010_),
    .B(_1717_));
 sg13g2_xnor2_1 _5157_ (.Y(_1720_),
    .A(_1610_),
    .B(_1688_));
 sg13g2_nand2_1 _5158_ (.Y(_1721_),
    .A(\pid.integral[4] ),
    .B(_1720_));
 sg13g2_xnor2_1 _5159_ (.Y(_1722_),
    .A(_1629_),
    .B(_1687_));
 sg13g2_nor2_1 _5160_ (.A(_0011_),
    .B(_1722_),
    .Y(_1723_));
 sg13g2_xnor2_1 _5161_ (.Y(_1725_),
    .A(_1650_),
    .B(_1686_));
 sg13g2_nand2_1 _5162_ (.Y(_1726_),
    .A(\pid.integral[2] ),
    .B(_1725_));
 sg13g2_o21ai_1 _5163_ (.B1(_1668_),
    .Y(_1727_),
    .A1(_1662_),
    .A2(_1664_));
 sg13g2_nand3b_1 _5164_ (.B(_1661_),
    .C(_1679_),
    .Y(_1728_),
    .A_N(_1658_));
 sg13g2_nand4_1 _5165_ (.B(_1671_),
    .C(_1727_),
    .A(_1654_),
    .Y(_1729_),
    .D(_1728_));
 sg13g2_nand2_1 _5166_ (.Y(_1730_),
    .A(_1684_),
    .B(_1729_));
 sg13g2_a21oi_1 _5167_ (.A1(_1684_),
    .A2(_1729_),
    .Y(_1731_),
    .B1(_1430_));
 sg13g2_xnor2_1 _5168_ (.Y(_1732_),
    .A(_1675_),
    .B(_1731_));
 sg13g2_and2_1 _5169_ (.A(_0953_),
    .B(_1732_),
    .X(_1733_));
 sg13g2_and2_1 _5170_ (.A(\pid.integral[0] ),
    .B(_1730_),
    .X(_1734_));
 sg13g2_or2_1 _5171_ (.X(_1736_),
    .B(_1732_),
    .A(_0953_));
 sg13g2_nand2b_1 _5172_ (.Y(_1737_),
    .B(_1736_),
    .A_N(_1733_));
 sg13g2_a21oi_1 _5173_ (.A1(_1734_),
    .A2(_1736_),
    .Y(_1738_),
    .B1(_1733_));
 sg13g2_xnor2_1 _5174_ (.Y(_1739_),
    .A(_1725_),
    .B(\pid.integral[2] ));
 sg13g2_o21ai_1 _5175_ (.B1(_1726_),
    .Y(_1740_),
    .A1(_1739_),
    .A2(_1738_));
 sg13g2_nand2_1 _5176_ (.Y(_1741_),
    .A(_0011_),
    .B(_1722_));
 sg13g2_nand2b_1 _5177_ (.Y(_1742_),
    .B(_1741_),
    .A_N(_1723_));
 sg13g2_a21oi_2 _5178_ (.B1(_1723_),
    .Y(_1743_),
    .A2(_1740_),
    .A1(_1741_));
 sg13g2_xnor2_1 _5179_ (.Y(_1744_),
    .A(\pid.integral[4] ),
    .B(_1720_));
 sg13g2_o21ai_1 _5180_ (.B1(_1721_),
    .Y(_1745_),
    .A1(_1744_),
    .A2(_1743_));
 sg13g2_a21oi_2 _5181_ (.B1(_1718_),
    .Y(_1747_),
    .A2(_1719_),
    .A1(_1745_));
 sg13g2_nor2_1 _5182_ (.A(\pid.integral[6] ),
    .B(_1715_),
    .Y(_1748_));
 sg13g2_xor2_1 _5183_ (.B(_1715_),
    .A(\pid.integral[6] ),
    .X(_1749_));
 sg13g2_o21ai_1 _5184_ (.B1(_1716_),
    .Y(_1750_),
    .A1(_1748_),
    .A2(_1747_));
 sg13g2_xor2_1 _5185_ (.B(_1712_),
    .A(_0009_),
    .X(_1751_));
 sg13g2_a21oi_2 _5186_ (.B1(_1714_),
    .Y(_1752_),
    .A2(_1750_),
    .A1(_1751_));
 sg13g2_nor2_1 _5187_ (.A(\pid.integral[8] ),
    .B(_1710_),
    .Y(_1753_));
 sg13g2_xnor2_1 _5188_ (.Y(_1754_),
    .A(\pid.integral[8] ),
    .B(_1709_));
 sg13g2_o21ai_1 _5189_ (.B1(_1711_),
    .Y(_1755_),
    .A1(_1753_),
    .A2(_1752_));
 sg13g2_a21oi_2 _5190_ (.B1(_1706_),
    .Y(_1756_),
    .A2(_1707_),
    .A1(_1755_));
 sg13g2_nor2_1 _5191_ (.A(\pid.integral[10] ),
    .B(_1703_),
    .Y(_1758_));
 sg13g2_xor2_1 _5192_ (.B(_1703_),
    .A(\pid.integral[10] ),
    .X(_1759_));
 sg13g2_o21ai_1 _5193_ (.B1(_1704_),
    .Y(_1760_),
    .A1(_1758_),
    .A2(_1756_));
 sg13g2_xnor2_1 _5194_ (.Y(_1761_),
    .A(_0007_),
    .B(net369));
 sg13g2_a21oi_2 _5195_ (.B1(_1701_),
    .Y(_1762_),
    .A2(_1760_),
    .A1(_1761_));
 sg13g2_xor2_1 _5196_ (.B(net369),
    .A(\pid.integral[12] ),
    .X(_1763_));
 sg13g2_inv_1 _5197_ (.Y(_1764_),
    .A(_1763_));
 sg13g2_o21ai_1 _5198_ (.B1(_1700_),
    .Y(_1765_),
    .A1(_1764_),
    .A2(_1762_));
 sg13g2_or2_1 _5199_ (.X(_1766_),
    .B(_1699_),
    .A(\pid.integral[13] ));
 sg13g2_and2_1 _5200_ (.A(\pid.integral[13] ),
    .B(_1699_),
    .X(_1767_));
 sg13g2_xor2_1 _5201_ (.B(net369),
    .A(\pid.integral[13] ),
    .X(_1768_));
 sg13g2_xnor2_1 _5202_ (.Y(_1769_),
    .A(_1768_),
    .B(_1765_));
 sg13g2_o21ai_1 _5203_ (.B1(_0915_),
    .Y(_1770_),
    .A1(_0916_),
    .A2(_1769_));
 sg13g2_or2_1 _5204_ (.X(_1771_),
    .B(net369),
    .A(_0942_));
 sg13g2_xnor2_1 _5205_ (.Y(_1772_),
    .A(_0942_),
    .B(net369));
 sg13g2_nor2_1 _5206_ (.A(_1765_),
    .B(_1767_),
    .Y(_1773_));
 sg13g2_o21ai_1 _5207_ (.B1(_1766_),
    .Y(_1774_),
    .A1(_1765_),
    .A2(_1767_));
 sg13g2_xnor2_1 _5208_ (.Y(_1775_),
    .A(_1772_),
    .B(_1774_));
 sg13g2_xor2_1 _5209_ (.B(_1775_),
    .A(_0917_),
    .X(_1776_));
 sg13g2_nand2_1 _5210_ (.Y(_1777_),
    .A(_1770_),
    .B(_1776_));
 sg13g2_xnor2_1 _5211_ (.Y(_1779_),
    .A(_2604_),
    .B(_0154_));
 sg13g2_xor2_1 _5212_ (.B(_0910_),
    .A(net35),
    .X(_1780_));
 sg13g2_nand2b_1 _5213_ (.Y(_1781_),
    .B(_1779_),
    .A_N(_1780_));
 sg13g2_xor2_1 _5214_ (.B(_1780_),
    .A(_1779_),
    .X(_1782_));
 sg13g2_xnor2_1 _5215_ (.Y(_1783_),
    .A(_1756_),
    .B(_1759_));
 sg13g2_nand2b_1 _5216_ (.Y(_1784_),
    .B(_1783_),
    .A_N(_1782_));
 sg13g2_nand2_1 _5217_ (.Y(_1785_),
    .A(_1781_),
    .B(_1784_));
 sg13g2_o21ai_1 _5218_ (.B1(net48),
    .Y(_1786_),
    .A1(_0910_),
    .A2(_0911_));
 sg13g2_nor2b_2 _5219_ (.A(_0912_),
    .B_N(_1786_),
    .Y(_1787_));
 sg13g2_and2_1 _5220_ (.A(_0155_),
    .B(_1787_),
    .X(_1788_));
 sg13g2_xnor2_1 _5221_ (.Y(_1790_),
    .A(_0155_),
    .B(_1787_));
 sg13g2_xnor2_1 _5222_ (.Y(_1791_),
    .A(_1761_),
    .B(_1760_));
 sg13g2_nor2_1 _5223_ (.A(_1790_),
    .B(_1791_),
    .Y(_1792_));
 sg13g2_xnor2_1 _5224_ (.Y(_1793_),
    .A(_1790_),
    .B(_1791_));
 sg13g2_nor2b_1 _5225_ (.A(_1793_),
    .B_N(_1785_),
    .Y(_1794_));
 sg13g2_xnor2_1 _5226_ (.Y(_1795_),
    .A(_1785_),
    .B(_1793_));
 sg13g2_xor2_1 _5227_ (.B(_0153_),
    .A(_2619_),
    .X(_1796_));
 sg13g2_xor2_1 _5228_ (.B(_0908_),
    .A(_0742_),
    .X(_1797_));
 sg13g2_and2_1 _5229_ (.A(_1796_),
    .B(_1797_),
    .X(_1798_));
 sg13g2_xnor2_1 _5230_ (.Y(_1799_),
    .A(_1708_),
    .B(_1755_));
 sg13g2_xor2_1 _5231_ (.B(_1797_),
    .A(_1796_),
    .X(_1801_));
 sg13g2_a21oi_1 _5232_ (.A1(_1799_),
    .A2(_1801_),
    .Y(_1802_),
    .B1(_1798_));
 sg13g2_xnor2_1 _5233_ (.Y(_1803_),
    .A(_1782_),
    .B(_1783_));
 sg13g2_nor2b_1 _5234_ (.A(_1802_),
    .B_N(_1803_),
    .Y(_1804_));
 sg13g2_nor2b_1 _5235_ (.A(_1803_),
    .B_N(_1802_),
    .Y(_1805_));
 sg13g2_nor2_1 _5236_ (.A(_1804_),
    .B(_1805_),
    .Y(_1806_));
 sg13g2_nor3_1 _5237_ (.A(net374),
    .B(net370),
    .C(_0900_),
    .Y(_1807_));
 sg13g2_nor2_2 _5238_ (.A(_0904_),
    .B(_1807_),
    .Y(_1808_));
 sg13g2_xor2_1 _5239_ (.B(_0149_),
    .A(_2675_),
    .X(_1809_));
 sg13g2_nand2_1 _5240_ (.Y(_1810_),
    .A(_1808_),
    .B(_1809_));
 sg13g2_xor2_1 _5241_ (.B(_1809_),
    .A(_1808_),
    .X(_1812_));
 sg13g2_xnor2_1 _5242_ (.Y(_1813_),
    .A(_1749_),
    .B(_1747_));
 sg13g2_nand2_1 _5243_ (.Y(_1814_),
    .A(_1812_),
    .B(_1813_));
 sg13g2_xnor2_1 _5244_ (.Y(_1815_),
    .A(_2656_),
    .B(_0150_));
 sg13g2_xor2_1 _5245_ (.B(_0906_),
    .A(net34),
    .X(_1816_));
 sg13g2_or2_1 _5246_ (.X(_1817_),
    .B(_1816_),
    .A(_1815_));
 sg13g2_xnor2_1 _5247_ (.Y(_1818_),
    .A(_1815_),
    .B(_1816_));
 sg13g2_xnor2_1 _5248_ (.Y(_1819_),
    .A(_1751_),
    .B(_1750_));
 sg13g2_or2_1 _5249_ (.X(_1820_),
    .B(_1819_),
    .A(_1818_));
 sg13g2_xnor2_1 _5250_ (.Y(_1821_),
    .A(_1818_),
    .B(_1819_));
 sg13g2_a21oi_1 _5251_ (.A1(_1810_),
    .A2(_1814_),
    .Y(_1823_),
    .B1(_1821_));
 sg13g2_xor2_1 _5252_ (.B(_0147_),
    .A(_2696_),
    .X(_1824_));
 sg13g2_xor2_1 _5253_ (.B(_0902_),
    .A(_0806_),
    .X(_1825_));
 sg13g2_xor2_1 _5254_ (.B(_1825_),
    .A(_1824_),
    .X(_1826_));
 sg13g2_xor2_1 _5255_ (.B(_1745_),
    .A(_1719_),
    .X(_1827_));
 sg13g2_nand2_1 _5256_ (.Y(_1828_),
    .A(_1826_),
    .B(_1827_));
 sg13g2_o21ai_1 _5257_ (.B1(_1828_),
    .Y(_1829_),
    .A1(_1824_),
    .A2(_1825_));
 sg13g2_xor2_1 _5258_ (.B(_1813_),
    .A(_1812_),
    .X(_1830_));
 sg13g2_and2_1 _5259_ (.A(_1829_),
    .B(_1830_),
    .X(_1831_));
 sg13g2_xor2_1 _5260_ (.B(_0146_),
    .A(_2709_),
    .X(_1832_));
 sg13g2_xor2_1 _5261_ (.B(_0901_),
    .A(_0830_),
    .X(_1833_));
 sg13g2_nand2_1 _5262_ (.Y(_1834_),
    .A(_1832_),
    .B(_1833_));
 sg13g2_xnor2_1 _5263_ (.Y(_1835_),
    .A(_1832_),
    .B(_1833_));
 sg13g2_xor2_1 _5264_ (.B(_1744_),
    .A(_1743_),
    .X(_1836_));
 sg13g2_nand2b_1 _5265_ (.Y(_1837_),
    .B(_1836_),
    .A_N(_1835_));
 sg13g2_nand2_1 _5266_ (.Y(_1838_),
    .A(_1834_),
    .B(_1837_));
 sg13g2_xnor2_1 _5267_ (.Y(_1839_),
    .A(_1826_),
    .B(_1827_));
 sg13g2_nand2b_1 _5268_ (.Y(_1840_),
    .B(_1838_),
    .A_N(_1839_));
 sg13g2_xnor2_1 _5269_ (.Y(_1841_),
    .A(_0853_),
    .B(_0897_));
 sg13g2_xor2_1 _5270_ (.B(_0145_),
    .A(_0091_),
    .X(_1842_));
 sg13g2_and2_1 _5271_ (.A(_1841_),
    .B(_1842_),
    .X(_1844_));
 sg13g2_xor2_1 _5272_ (.B(_1842_),
    .A(_1841_),
    .X(_1845_));
 sg13g2_xnor2_1 _5273_ (.Y(_1846_),
    .A(_1742_),
    .B(_1740_));
 sg13g2_a21oi_1 _5274_ (.A1(_1845_),
    .A2(_1846_),
    .Y(_1847_),
    .B1(_1844_));
 sg13g2_xnor2_1 _5275_ (.Y(_1848_),
    .A(_1835_),
    .B(_1836_));
 sg13g2_nor2b_1 _5276_ (.A(_1847_),
    .B_N(_1848_),
    .Y(_1849_));
 sg13g2_xnor2_1 _5277_ (.Y(_1850_),
    .A(_0112_),
    .B(_0144_));
 sg13g2_xnor2_1 _5278_ (.Y(_1851_),
    .A(_0874_),
    .B(_0896_));
 sg13g2_nor2_1 _5279_ (.A(_1850_),
    .B(_1851_),
    .Y(_1852_));
 sg13g2_xnor2_1 _5280_ (.Y(_1853_),
    .A(_1850_),
    .B(_1851_));
 sg13g2_xnor2_1 _5281_ (.Y(_1855_),
    .A(_1739_),
    .B(_1738_));
 sg13g2_nor2_1 _5282_ (.A(_1853_),
    .B(_1855_),
    .Y(_1856_));
 sg13g2_nor2_1 _5283_ (.A(_1852_),
    .B(_1856_),
    .Y(_1857_));
 sg13g2_xor2_1 _5284_ (.B(_1846_),
    .A(_1845_),
    .X(_1858_));
 sg13g2_nand2b_1 _5285_ (.Y(_1859_),
    .B(_1858_),
    .A_N(_1857_));
 sg13g2_nor2_1 _5286_ (.A(net373),
    .B(_0143_),
    .Y(_1860_));
 sg13g2_xor2_1 _5287_ (.B(_1860_),
    .A(_0132_),
    .X(_1861_));
 sg13g2_nor2_1 _5288_ (.A(_0870_),
    .B(_0892_),
    .Y(_1862_));
 sg13g2_nand4_1 _5289_ (.B(_0877_),
    .C(_0880_),
    .A(_0858_),
    .Y(_1863_),
    .D(_0883_));
 sg13g2_nand3_1 _5290_ (.B(_1862_),
    .C(_0879_),
    .A(_1863_),
    .Y(_1864_));
 sg13g2_nor2_1 _5291_ (.A(_0883_),
    .B(_0885_),
    .Y(_1866_));
 sg13g2_o21ai_1 _5292_ (.B1(_0888_),
    .Y(_1867_),
    .A1(_0881_),
    .A2(_1866_));
 sg13g2_nor2b_1 _5293_ (.A(_0893_),
    .B_N(_0892_),
    .Y(_1868_));
 sg13g2_nand3b_1 _5294_ (.B(_1867_),
    .C(_1868_),
    .Y(_1869_),
    .A_N(_0879_));
 sg13g2_nor2_1 _5295_ (.A(net374),
    .B(_0893_),
    .Y(_1870_));
 sg13g2_nand3b_1 _5296_ (.B(_1864_),
    .C(_1869_),
    .Y(_1871_),
    .A_N(_0895_));
 sg13g2_nand2_2 _5297_ (.Y(_1872_),
    .A(_0893_),
    .B(_1864_));
 sg13g2_nand3_1 _5298_ (.B(_1869_),
    .C(_1870_),
    .A(_1864_),
    .Y(_1873_));
 sg13g2_o21ai_1 _5299_ (.B1(_1873_),
    .Y(_1874_),
    .A1(_1872_),
    .A2(_0896_));
 sg13g2_xnor2_1 _5300_ (.Y(_1875_),
    .A(_1874_),
    .B(_1861_));
 sg13g2_xnor2_1 _5301_ (.Y(_1877_),
    .A(_1737_),
    .B(_1734_));
 sg13g2_nand2b_1 _5302_ (.Y(_1878_),
    .B(_1877_),
    .A_N(_1875_));
 sg13g2_o21ai_1 _5303_ (.B1(_1878_),
    .Y(_1879_),
    .A1(_1861_),
    .A2(_1874_));
 sg13g2_xnor2_1 _5304_ (.Y(_1880_),
    .A(_1853_),
    .B(_1855_));
 sg13g2_nand2b_1 _5305_ (.Y(_1881_),
    .B(_1879_),
    .A_N(_1880_));
 sg13g2_xor2_1 _5306_ (.B(_1730_),
    .A(net121),
    .X(_1882_));
 sg13g2_xor2_1 _5307_ (.B(_1871_),
    .A(_0143_),
    .X(_1883_));
 sg13g2_nand2_1 _5308_ (.Y(_1884_),
    .A(_1882_),
    .B(_1883_));
 sg13g2_o21ai_1 _5309_ (.B1(_1884_),
    .Y(_1885_),
    .A1(_0143_),
    .A2(_1871_));
 sg13g2_xnor2_1 _5310_ (.Y(_1886_),
    .A(_1875_),
    .B(_1877_));
 sg13g2_nand2_1 _5311_ (.Y(_1888_),
    .A(_1885_),
    .B(_1886_));
 sg13g2_xor2_1 _5312_ (.B(_1879_),
    .A(_1880_),
    .X(_1889_));
 sg13g2_or2_1 _5313_ (.X(_1890_),
    .B(_1888_),
    .A(_1889_));
 sg13g2_xor2_1 _5314_ (.B(_1858_),
    .A(_1857_),
    .X(_1891_));
 sg13g2_a21o_1 _5315_ (.A2(_1881_),
    .A1(_1890_),
    .B1(_1891_),
    .X(_1892_));
 sg13g2_xor2_1 _5316_ (.B(_1848_),
    .A(_1847_),
    .X(_1893_));
 sg13g2_a21oi_2 _5317_ (.B1(_1893_),
    .Y(_1894_),
    .A2(_1859_),
    .A1(_1892_));
 sg13g2_xnor2_1 _5318_ (.Y(_1895_),
    .A(_1838_),
    .B(_1839_));
 sg13g2_o21ai_1 _5319_ (.B1(_1895_),
    .Y(_1896_),
    .A1(_1894_),
    .A2(_1849_));
 sg13g2_xnor2_1 _5320_ (.Y(_1897_),
    .A(_1829_),
    .B(_1830_));
 sg13g2_a21oi_2 _5321_ (.B1(_1897_),
    .Y(_1899_),
    .A2(_1840_),
    .A1(_1896_));
 sg13g2_nand3_1 _5322_ (.B(_1814_),
    .C(_1821_),
    .A(_1810_),
    .Y(_1900_));
 sg13g2_nor2b_1 _5323_ (.A(_1823_),
    .B_N(_1900_),
    .Y(_1901_));
 sg13g2_o21ai_1 _5324_ (.B1(_1901_),
    .Y(_1902_),
    .A1(_1899_),
    .A2(_1831_));
 sg13g2_nor2b_2 _5325_ (.A(_1823_),
    .B_N(_1902_),
    .Y(_1903_));
 sg13g2_xnor2_1 _5326_ (.Y(_1904_),
    .A(_0759_),
    .B(_0907_));
 sg13g2_xnor2_1 _5327_ (.Y(_1905_),
    .A(_2639_),
    .B(_0152_));
 sg13g2_xnor2_1 _5328_ (.Y(_1906_),
    .A(_1754_),
    .B(_1752_));
 sg13g2_xor2_1 _5329_ (.B(_1905_),
    .A(_1904_),
    .X(_1907_));
 sg13g2_and2_1 _5330_ (.A(_1906_),
    .B(_1907_),
    .X(_1908_));
 sg13g2_a21o_1 _5331_ (.A2(_1905_),
    .A1(_1904_),
    .B1(_1908_),
    .X(_1910_));
 sg13g2_xnor2_1 _5332_ (.Y(_1911_),
    .A(_1799_),
    .B(_1801_));
 sg13g2_nor2b_1 _5333_ (.A(_1911_),
    .B_N(_1910_),
    .Y(_1912_));
 sg13g2_xnor2_1 _5334_ (.Y(_1913_),
    .A(_1910_),
    .B(_1911_));
 sg13g2_inv_1 _5335_ (.Y(_1914_),
    .A(_1913_));
 sg13g2_and2_1 _5336_ (.A(_1817_),
    .B(_1820_),
    .X(_1915_));
 sg13g2_xnor2_1 _5337_ (.Y(_1916_),
    .A(_1906_),
    .B(_1907_));
 sg13g2_and2_1 _5338_ (.A(_1915_),
    .B(_1916_),
    .X(_1917_));
 sg13g2_nand2_1 _5339_ (.Y(_1918_),
    .A(_1915_),
    .B(_1916_));
 sg13g2_nor2_1 _5340_ (.A(_1915_),
    .B(_1916_),
    .Y(_1919_));
 sg13g2_nor4_2 _5341_ (.A(_1903_),
    .B(_1914_),
    .C(_1917_),
    .Y(_1921_),
    .D(_1919_));
 sg13g2_nand3_1 _5342_ (.B(_1921_),
    .C(_1806_),
    .A(_1795_),
    .Y(_1922_));
 sg13g2_nand2_1 _5343_ (.Y(_1923_),
    .A(_1913_),
    .B(_1919_));
 sg13g2_nand2b_1 _5344_ (.Y(_1924_),
    .B(_1923_),
    .A_N(_1912_));
 sg13g2_nand3_1 _5345_ (.B(_1806_),
    .C(_1924_),
    .A(_1795_),
    .Y(_1925_));
 sg13g2_a21oi_1 _5346_ (.A1(_1795_),
    .A2(_1804_),
    .Y(_1926_),
    .B1(_1794_));
 sg13g2_nand3_1 _5347_ (.B(_1925_),
    .C(_1926_),
    .A(_1922_),
    .Y(_1927_));
 sg13g2_xnor2_1 _5348_ (.Y(_1928_),
    .A(_1763_),
    .B(_1762_));
 sg13g2_a21oi_1 _5349_ (.A1(_0917_),
    .A2(_1928_),
    .Y(_1929_),
    .B1(_0914_));
 sg13g2_xor2_1 _5350_ (.B(_0917_),
    .A(_1769_),
    .X(_1930_));
 sg13g2_nor2_1 _5351_ (.A(_1929_),
    .B(_1930_),
    .Y(_1932_));
 sg13g2_xor2_1 _5352_ (.B(_1930_),
    .A(_1929_),
    .X(_1933_));
 sg13g2_xor2_1 _5353_ (.B(_1928_),
    .A(_0917_),
    .X(_1934_));
 sg13g2_o21ai_1 _5354_ (.B1(_1934_),
    .Y(_1935_),
    .A1(_1788_),
    .A2(_1792_));
 sg13g2_inv_1 _5355_ (.Y(_1936_),
    .A(_1935_));
 sg13g2_or3_1 _5356_ (.A(_1788_),
    .B(_1792_),
    .C(_1934_),
    .X(_1937_));
 sg13g2_nand3_1 _5357_ (.B(_1935_),
    .C(_1937_),
    .A(_1933_),
    .Y(_1938_));
 sg13g2_nand4_1 _5358_ (.B(_1927_),
    .C(_1935_),
    .A(_1933_),
    .Y(_1939_),
    .D(_1937_));
 sg13g2_a21oi_1 _5359_ (.A1(_1933_),
    .A2(_1936_),
    .Y(_1940_),
    .B1(_1932_));
 sg13g2_xnor2_1 _5360_ (.Y(_1941_),
    .A(_1770_),
    .B(_1776_));
 sg13g2_a21o_1 _5361_ (.A2(_1939_),
    .A1(_1940_),
    .B1(_1941_),
    .X(_1942_));
 sg13g2_nand3_1 _5362_ (.B(net369),
    .C(_1773_),
    .A(_0942_),
    .Y(_1943_));
 sg13g2_o21ai_1 _5363_ (.B1(_1943_),
    .Y(_1944_),
    .A1(_1771_),
    .A2(_1774_));
 sg13g2_xor2_1 _5364_ (.B(_1944_),
    .A(net97),
    .X(_1945_));
 sg13g2_a21oi_1 _5365_ (.A1(_0915_),
    .A2(_1775_),
    .Y(_1946_),
    .B1(_0916_));
 sg13g2_xnor2_1 _5366_ (.Y(_1947_),
    .A(_1945_),
    .B(_1946_));
 sg13g2_and3_1 _5367_ (.X(_1948_),
    .A(_1777_),
    .B(_1942_),
    .C(_1947_));
 sg13g2_a21oi_2 _5368_ (.B1(_1947_),
    .Y(_1949_),
    .A2(_1777_),
    .A1(_1942_));
 sg13g2_or2_1 _5369_ (.X(_1950_),
    .B(_1949_),
    .A(_1948_));
 sg13g2_nand3_1 _5370_ (.B(_1940_),
    .C(_1941_),
    .A(_1939_),
    .Y(_1951_));
 sg13g2_mux2_1 _5371_ (.A0(_1805_),
    .A1(_1804_),
    .S(_1795_),
    .X(_1953_));
 sg13g2_nand2b_1 _5372_ (.Y(_1954_),
    .B(_1953_),
    .A_N(_1924_));
 sg13g2_nand2_1 _5373_ (.Y(_1955_),
    .A(_1925_),
    .B(_1954_));
 sg13g2_o21ai_1 _5374_ (.B1(_1923_),
    .Y(_1956_),
    .A1(_1913_),
    .A2(_1918_));
 sg13g2_nand3_1 _5375_ (.B(_1955_),
    .C(_1956_),
    .A(_1903_),
    .Y(_1957_));
 sg13g2_mux2_1 _5376_ (.A0(_1937_),
    .A1(_1935_),
    .S(_1933_),
    .X(_1958_));
 sg13g2_mux2_1 _5377_ (.A0(_1958_),
    .A1(_1938_),
    .S(_1927_),
    .X(_1959_));
 sg13g2_a221oi_1 _5378_ (.B2(_1922_),
    .C1(_1959_),
    .B1(_1957_),
    .A1(_1951_),
    .Y(_1960_),
    .A2(_1942_));
 sg13g2_or3_1 _5379_ (.A(_1831_),
    .B(_1899_),
    .C(_1901_),
    .X(_1961_));
 sg13g2_nand2_1 _5380_ (.Y(_1962_),
    .A(_1902_),
    .B(_1961_));
 sg13g2_nand3_1 _5381_ (.B(_1896_),
    .C(_1897_),
    .A(_1840_),
    .Y(_1964_));
 sg13g2_nor2b_1 _5382_ (.A(_1899_),
    .B_N(_1964_),
    .Y(_1965_));
 sg13g2_or3_1 _5383_ (.A(_1849_),
    .B(_1894_),
    .C(_1895_),
    .X(_1966_));
 sg13g2_and2_1 _5384_ (.A(_1896_),
    .B(_1966_),
    .X(_1967_));
 sg13g2_nand3_1 _5385_ (.B(_1892_),
    .C(_1893_),
    .A(_1859_),
    .Y(_1968_));
 sg13g2_nor2b_1 _5386_ (.A(_1894_),
    .B_N(_1968_),
    .Y(_1969_));
 sg13g2_nand3_1 _5387_ (.B(_1890_),
    .C(_1891_),
    .A(_1881_),
    .Y(_1970_));
 sg13g2_nand2_1 _5388_ (.Y(_1971_),
    .A(_1892_),
    .B(_1970_));
 sg13g2_inv_1 _5389_ (.Y(_1972_),
    .A(_1971_));
 sg13g2_xnor2_1 _5390_ (.Y(_1973_),
    .A(_1888_),
    .B(_1889_));
 sg13g2_inv_1 _5391_ (.Y(_1975_),
    .A(_1973_));
 sg13g2_xor2_1 _5392_ (.B(_1883_),
    .A(_1882_),
    .X(_1976_));
 sg13g2_xor2_1 _5393_ (.B(_1886_),
    .A(_1885_),
    .X(_1977_));
 sg13g2_or4_1 _5394_ (.A(_1972_),
    .B(_1975_),
    .C(_1976_),
    .D(_1977_),
    .X(_1978_));
 sg13g2_nor4_1 _5395_ (.A(_1965_),
    .B(_1967_),
    .C(_1969_),
    .D(_1978_),
    .Y(_1979_));
 sg13g2_nand3_1 _5396_ (.B(_1962_),
    .C(_1979_),
    .A(_1960_),
    .Y(_1980_));
 sg13g2_nand3_1 _5397_ (.B(_1950_),
    .C(_1980_),
    .A(net451),
    .Y(_1981_));
 sg13g2_o21ai_1 _5398_ (.B1(_1960_),
    .Y(_1982_),
    .A1(_1948_),
    .A2(_1949_));
 sg13g2_and4_1 _5399_ (.A(_1972_),
    .B(_1975_),
    .C(_1976_),
    .D(_1977_),
    .X(_1983_));
 sg13g2_nand4_1 _5400_ (.B(_1967_),
    .C(_1969_),
    .A(_1965_),
    .Y(_1984_),
    .D(_1983_));
 sg13g2_nor2_2 _5401_ (.A(_1962_),
    .B(_1984_),
    .Y(_1986_));
 sg13g2_nor3_2 _5402_ (.A(_1976_),
    .B(_1986_),
    .C(net88),
    .Y(_1987_));
 sg13g2_o21ai_1 _5403_ (.B1(net102),
    .Y(_0058_),
    .A1(_1981_),
    .A2(_1987_));
 sg13g2_nand2b_1 _5404_ (.Y(_1988_),
    .B(net106),
    .A_N(\pid.state[3] ));
 sg13g2_nor3_2 _5405_ (.A(_1977_),
    .B(net88),
    .C(_1986_),
    .Y(_1989_));
 sg13g2_o21ai_1 _5406_ (.B1(net107),
    .Y(_0059_),
    .A1(_1981_),
    .A2(_1989_));
 sg13g2_nand2b_1 _5407_ (.Y(_1990_),
    .B(net108),
    .A_N(net451));
 sg13g2_nor3_2 _5408_ (.A(_1975_),
    .B(net88),
    .C(_1986_),
    .Y(_1991_));
 sg13g2_o21ai_1 _5409_ (.B1(net109),
    .Y(_0060_),
    .A1(_1981_),
    .A2(_1991_));
 sg13g2_nand2b_1 _5410_ (.Y(_1992_),
    .B(net104),
    .A_N(net451));
 sg13g2_nor3_2 _5411_ (.A(net88),
    .B(_1972_),
    .C(_1986_),
    .Y(_1994_));
 sg13g2_o21ai_1 _5412_ (.B1(net105),
    .Y(_0061_),
    .A1(_1981_),
    .A2(_1994_));
 sg13g2_nand2b_1 _5413_ (.Y(_1995_),
    .B(net117),
    .A_N(net451));
 sg13g2_nor2_2 _5414_ (.A(net88),
    .B(_1969_),
    .Y(_1996_));
 sg13g2_o21ai_1 _5415_ (.B1(net118),
    .Y(_0062_),
    .A1(_1996_),
    .A2(_1981_));
 sg13g2_nand2b_1 _5416_ (.Y(_1997_),
    .B(net114),
    .A_N(net451));
 sg13g2_nor2_1 _5417_ (.A(_1967_),
    .B(net88),
    .Y(_1998_));
 sg13g2_o21ai_1 _5418_ (.B1(net115),
    .Y(_0063_),
    .A1(_1981_),
    .A2(_1998_));
 sg13g2_nand2b_1 _5419_ (.Y(_1999_),
    .B(net127),
    .A_N(net451));
 sg13g2_nor2_1 _5420_ (.A(_1965_),
    .B(net88),
    .Y(_2000_));
 sg13g2_o21ai_1 _5421_ (.B1(net128),
    .Y(_0064_),
    .A1(_2000_),
    .A2(_1981_));
 sg13g2_nand2b_1 _5422_ (.Y(_2002_),
    .B(net129),
    .A_N(net451));
 sg13g2_nor2b_1 _5423_ (.A(net88),
    .B_N(_1962_),
    .Y(_2003_));
 sg13g2_o21ai_1 _5424_ (.B1(net130),
    .Y(_0065_),
    .A1(_1981_),
    .A2(_2003_));
 sg13g2_nor2_1 _5425_ (.A(net460),
    .B(net145),
    .Y(_2004_));
 sg13g2_a21oi_1 _5426_ (.A1(net460),
    .A2(_1007_),
    .Y(_0066_),
    .B1(_2004_));
 sg13g2_nor2_1 _5427_ (.A(net460),
    .B(net147),
    .Y(_2005_));
 sg13g2_a21oi_1 _5428_ (.A1(net460),
    .A2(_1050_),
    .Y(_0067_),
    .B1(_2005_));
 sg13g2_nor2_1 _5429_ (.A(net460),
    .B(net148),
    .Y(_2006_));
 sg13g2_a21oi_1 _5430_ (.A1(net460),
    .A2(_1115_),
    .Y(_0068_),
    .B1(_2006_));
 sg13g2_nor2_1 _5431_ (.A(net459),
    .B(net150),
    .Y(_2008_));
 sg13g2_a21oi_1 _5432_ (.A1(net460),
    .A2(_1169_),
    .Y(_0069_),
    .B1(_2008_));
 sg13g2_nor2_1 _5433_ (.A(net458),
    .B(net139),
    .Y(_2009_));
 sg13g2_a21oi_1 _5434_ (.A1(net459),
    .A2(_1201_),
    .Y(_0070_),
    .B1(_2009_));
 sg13g2_nor2_1 _5435_ (.A(net459),
    .B(net144),
    .Y(_2010_));
 sg13g2_a21oi_1 _5436_ (.A1(net458),
    .A2(_1244_),
    .Y(_0071_),
    .B1(_2010_));
 sg13g2_nor2_1 _5437_ (.A(net458),
    .B(net151),
    .Y(_2011_));
 sg13g2_a21oi_1 _5438_ (.A1(net458),
    .A2(_1287_),
    .Y(_0072_),
    .B1(_2011_));
 sg13g2_nor2_1 _5439_ (.A(net458),
    .B(net141),
    .Y(_2012_));
 sg13g2_a21oi_1 _5440_ (.A1(net458),
    .A2(_1319_),
    .Y(_0073_),
    .B1(_2012_));
 sg13g2_nor2_1 _5441_ (.A(net458),
    .B(net143),
    .Y(_2014_));
 sg13g2_a21oi_1 _5442_ (.A1(net458),
    .A2(_1351_),
    .Y(_0074_),
    .B1(_2014_));
 sg13g2_mux2_1 _5443_ (.A0(net121),
    .A1(_1882_),
    .S(net427),
    .X(_0075_));
 sg13g2_mux2_1 _5444_ (.A0(net90),
    .A1(_1877_),
    .S(net427),
    .X(_0076_));
 sg13g2_nor2_1 _5445_ (.A(net103),
    .B(net428),
    .Y(_2015_));
 sg13g2_a21oi_1 _5446_ (.A1(net428),
    .A2(_1855_),
    .Y(_0077_),
    .B1(_2015_));
 sg13g2_mux2_1 _5447_ (.A0(net91),
    .A1(_1846_),
    .S(net428),
    .X(_0078_));
 sg13g2_mux2_1 _5448_ (.A0(net113),
    .A1(_1836_),
    .S(net427),
    .X(_0079_));
 sg13g2_mux2_1 _5449_ (.A0(net93),
    .A1(_1827_),
    .S(net427),
    .X(_0080_));
 sg13g2_mux2_1 _5450_ (.A0(net132),
    .A1(_1813_),
    .S(net427),
    .X(_0081_));
 sg13g2_nor2_1 _5451_ (.A(net89),
    .B(net428),
    .Y(_2017_));
 sg13g2_a21oi_1 _5452_ (.A1(net427),
    .A2(_1819_),
    .Y(_0082_),
    .B1(_2017_));
 sg13g2_mux2_1 _5453_ (.A0(net131),
    .A1(_1906_),
    .S(net429),
    .X(_0083_));
 sg13g2_mux2_1 _5454_ (.A0(net92),
    .A1(_1799_),
    .S(net429),
    .X(_0084_));
 sg13g2_mux2_1 _5455_ (.A0(net125),
    .A1(_1783_),
    .S(net429),
    .X(_0085_));
 sg13g2_nor2_1 _5456_ (.A(net96),
    .B(net429),
    .Y(_2018_));
 sg13g2_a21oi_2 _5457_ (.B1(_2018_),
    .Y(_0086_),
    .A2(net429),
    .A1(_1791_));
 sg13g2_mux2_1 _5458_ (.A0(net112),
    .A1(_1928_),
    .S(net429),
    .X(_0087_));
 sg13g2_nor2_1 _5459_ (.A(net116),
    .B(net429),
    .Y(_2019_));
 sg13g2_a21oi_1 _5460_ (.A1(net429),
    .A2(_1769_),
    .Y(_0088_),
    .B1(_2019_));
 sg13g2_mux2_1 _5461_ (.A0(net94),
    .A1(_1775_),
    .S(net427),
    .X(_0089_));
 sg13g2_mux2_1 _5462_ (.A0(net97),
    .A1(_1945_),
    .S(net427),
    .X(_0090_));
 sg13g2_dfrbp_1 _5463_ (.CLK(clknet_4_8__leaf_clk),
    .RESET_B(net480),
    .D(_0031_),
    .Q_N(_2761_),
    .Q(\pid.Kd[0] ));
 sg13g2_dfrbp_1 _5464_ (.CLK(clknet_4_8__leaf_clk),
    .RESET_B(net480),
    .D(_0032_),
    .Q_N(_0019_),
    .Q(\pid.Kd[1] ));
 sg13g2_dfrbp_1 _5465_ (.CLK(clknet_4_2__leaf_clk),
    .RESET_B(net480),
    .D(_0033_),
    .Q_N(_0018_),
    .Q(\pid.Kd[2] ));
 sg13g2_dfrbp_1 _5466_ (.CLK(clknet_4_2__leaf_clk),
    .RESET_B(net480),
    .D(_0034_),
    .Q_N(_0017_),
    .Q(\pid.Kd[3] ));
 sg13g2_dfrbp_1 _5467_ (.CLK(clknet_4_1__leaf_clk),
    .RESET_B(net477),
    .D(_0035_),
    .Q_N(_0016_),
    .Q(\pid.Kd[4] ));
 sg13g2_dfrbp_1 _5468_ (.CLK(clknet_4_0__leaf_clk),
    .RESET_B(net477),
    .D(_0036_),
    .Q_N(_0015_),
    .Q(\pid.Kd[5] ));
 sg13g2_dfrbp_1 _5469_ (.CLK(clknet_4_0__leaf_clk),
    .RESET_B(net477),
    .D(_0037_),
    .Q_N(_0014_),
    .Q(\pid.Kd[6] ));
 sg13g2_dfrbp_1 _5470_ (.CLK(clknet_4_0__leaf_clk),
    .RESET_B(net477),
    .D(_0038_),
    .Q_N(_0013_),
    .Q(\pid.Kd[7] ));
 sg13g2_dfrbp_1 _5471_ (.CLK(clknet_4_0__leaf_clk),
    .RESET_B(net477),
    .D(_0039_),
    .Q_N(_2760_),
    .Q(\pid.Kd[8] ));
 sg13g2_dfrbp_1 _5472_ (.CLK(clknet_4_3__leaf_clk),
    .RESET_B(net478),
    .D(net33),
    .Q_N(\pid.state[0] ),
    .Q(_0029_));
 sg13g2_dfrbp_1 _5473_ (.CLK(clknet_4_12__leaf_clk),
    .RESET_B(net479),
    .D(net453),
    .Q_N(_2762_),
    .Q(\pid.state[1] ));
 sg13g2_dfrbp_1 _5474_ (.CLK(clknet_4_3__leaf_clk),
    .RESET_B(net476),
    .D(net460),
    .Q_N(_2763_),
    .Q(\pid.state[2] ));
 sg13g2_dfrbp_1 _5475_ (.CLK(clknet_4_11__leaf_clk),
    .RESET_B(net483),
    .D(net124),
    .Q_N(_2759_),
    .Q(\pid.state[3] ));
 sg13g2_dfrbp_1 _5476_ (.CLK(clknet_4_13__leaf_clk),
    .RESET_B(net479),
    .D(_0040_),
    .Q_N(_0006_),
    .Q(\pid.Ki[0] ));
 sg13g2_dfrbp_1 _5477_ (.CLK(clknet_4_12__leaf_clk),
    .RESET_B(net479),
    .D(net99),
    .Q_N(_0003_),
    .Q(\pid.Ki[1] ));
 sg13g2_dfrbp_1 _5478_ (.CLK(clknet_4_7__leaf_clk),
    .RESET_B(net478),
    .D(_0042_),
    .Q_N(_2758_),
    .Q(\pid.Ki[2] ));
 sg13g2_dfrbp_1 _5479_ (.CLK(clknet_4_7__leaf_clk),
    .RESET_B(net478),
    .D(_0043_),
    .Q_N(_2757_),
    .Q(\pid.Ki[3] ));
 sg13g2_dfrbp_1 _5480_ (.CLK(clknet_4_6__leaf_clk),
    .RESET_B(net478),
    .D(_0044_),
    .Q_N(_0005_),
    .Q(\pid.Ki[4] ));
 sg13g2_dfrbp_1 _5481_ (.CLK(clknet_4_7__leaf_clk),
    .RESET_B(net479),
    .D(net137),
    .Q_N(_0004_),
    .Q(\pid.Ki[5] ));
 sg13g2_dfrbp_1 _5482_ (.CLK(clknet_4_7__leaf_clk),
    .RESET_B(net476),
    .D(_0046_),
    .Q_N(_2756_),
    .Q(\pid.Ki[6] ));
 sg13g2_dfrbp_1 _5483_ (.CLK(clknet_4_5__leaf_clk),
    .RESET_B(net477),
    .D(_0047_),
    .Q_N(_0002_),
    .Q(\pid.Ki[7] ));
 sg13g2_dfrbp_1 _5484_ (.CLK(clknet_4_5__leaf_clk),
    .RESET_B(net477),
    .D(_0048_),
    .Q_N(_0001_),
    .Q(\pid.Ki[8] ));
 sg13g2_dfrbp_1 _5485_ (.CLK(clknet_4_8__leaf_clk),
    .RESET_B(net480),
    .D(_0049_),
    .Q_N(_2755_),
    .Q(\pid.prev_error[0] ));
 sg13g2_dfrbp_1 _5486_ (.CLK(clknet_4_6__leaf_clk),
    .RESET_B(net478),
    .D(_0050_),
    .Q_N(_2754_),
    .Q(\pid.prev_error[1] ));
 sg13g2_dfrbp_1 _5487_ (.CLK(clknet_4_6__leaf_clk),
    .RESET_B(net479),
    .D(net120),
    .Q_N(_2753_),
    .Q(\pid.prev_error[2] ));
 sg13g2_dfrbp_1 _5488_ (.CLK(clknet_4_12__leaf_clk),
    .RESET_B(net484),
    .D(_0052_),
    .Q_N(_2752_),
    .Q(\pid.prev_error[3] ));
 sg13g2_dfrbp_1 _5489_ (.CLK(clknet_4_6__leaf_clk),
    .RESET_B(net479),
    .D(_0053_),
    .Q_N(_2751_),
    .Q(\pid.prev_error[4] ));
 sg13g2_dfrbp_1 _5490_ (.CLK(clknet_4_2__leaf_clk),
    .RESET_B(net479),
    .D(_0054_),
    .Q_N(_2750_),
    .Q(\pid.prev_error[5] ));
 sg13g2_dfrbp_1 _5491_ (.CLK(clknet_4_2__leaf_clk),
    .RESET_B(net480),
    .D(_0055_),
    .Q_N(_2749_),
    .Q(\pid.prev_error[6] ));
 sg13g2_dfrbp_1 _5492_ (.CLK(clknet_4_3__leaf_clk),
    .RESET_B(net480),
    .D(_0056_),
    .Q_N(_2748_),
    .Q(\pid.prev_error[7] ));
 sg13g2_dfrbp_1 _5493_ (.CLK(clknet_4_3__leaf_clk),
    .RESET_B(net478),
    .D(_0057_),
    .Q_N(_2747_),
    .Q(\pid.prev_error[8] ));
 sg13g2_dfrbp_1 _5494_ (.CLK(clknet_4_10__leaf_clk),
    .RESET_B(net482),
    .D(_0058_),
    .Q_N(_2746_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _5495_ (.CLK(clknet_4_14__leaf_clk),
    .RESET_B(net483),
    .D(_0059_),
    .Q_N(_2745_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _5496_ (.CLK(clknet_4_10__leaf_clk),
    .RESET_B(net483),
    .D(_0060_),
    .Q_N(_2744_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _5497_ (.CLK(clknet_4_10__leaf_clk),
    .RESET_B(net483),
    .D(_0061_),
    .Q_N(_2743_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _5498_ (.CLK(clknet_4_10__leaf_clk),
    .RESET_B(net483),
    .D(_0062_),
    .Q_N(_2742_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _5499_ (.CLK(clknet_4_11__leaf_clk),
    .RESET_B(net483),
    .D(_0063_),
    .Q_N(_2741_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _5500_ (.CLK(clknet_4_9__leaf_clk),
    .RESET_B(net483),
    .D(_0064_),
    .Q_N(_2740_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _5501_ (.CLK(clknet_4_9__leaf_clk),
    .RESET_B(net483),
    .D(_0065_),
    .Q_N(_2739_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _5502_ (.CLK(clknet_4_1__leaf_clk),
    .RESET_B(net478),
    .D(_0066_),
    .Q_N(_0028_),
    .Q(\pid.Kp[0] ));
 sg13g2_dfrbp_1 _5503_ (.CLK(clknet_4_1__leaf_clk),
    .RESET_B(net478),
    .D(_0067_),
    .Q_N(_0027_),
    .Q(\pid.Kp[1] ));
 sg13g2_dfrbp_1 _5504_ (.CLK(clknet_4_1__leaf_clk),
    .RESET_B(net485),
    .D(_0068_),
    .Q_N(_0026_),
    .Q(\pid.Kp[2] ));
 sg13g2_dfrbp_1 _5505_ (.CLK(clknet_4_4__leaf_clk),
    .RESET_B(net476),
    .D(_0069_),
    .Q_N(_0023_),
    .Q(\pid.Kp[3] ));
 sg13g2_dfrbp_1 _5506_ (.CLK(clknet_4_4__leaf_clk),
    .RESET_B(net476),
    .D(_0070_),
    .Q_N(_0025_),
    .Q(\pid.Kp[4] ));
 sg13g2_dfrbp_1 _5507_ (.CLK(clknet_4_4__leaf_clk),
    .RESET_B(net476),
    .D(_0071_),
    .Q_N(_0024_),
    .Q(\pid.Kp[5] ));
 sg13g2_dfrbp_1 _5508_ (.CLK(clknet_4_4__leaf_clk),
    .RESET_B(net476),
    .D(_0072_),
    .Q_N(_0022_),
    .Q(\pid.Kp[6] ));
 sg13g2_dfrbp_1 _5509_ (.CLK(clknet_4_5__leaf_clk),
    .RESET_B(net476),
    .D(_0073_),
    .Q_N(_0021_),
    .Q(\pid.Kp[7] ));
 sg13g2_dfrbp_1 _5510_ (.CLK(clknet_4_5__leaf_clk),
    .RESET_B(net476),
    .D(_0074_),
    .Q_N(_0020_),
    .Q(\pid.Kp[8] ));
 sg13g2_dfrbp_1 _5511_ (.CLK(clknet_4_14__leaf_clk),
    .RESET_B(net481),
    .D(_0075_),
    .Q_N(_2738_),
    .Q(\pid.integral[0] ));
 sg13g2_dfrbp_1 _5512_ (.CLK(clknet_4_14__leaf_clk),
    .RESET_B(net481),
    .D(_0076_),
    .Q_N(_0012_),
    .Q(\pid.integral[1] ));
 sg13g2_dfrbp_1 _5513_ (.CLK(clknet_4_15__leaf_clk),
    .RESET_B(net481),
    .D(_0077_),
    .Q_N(_2737_),
    .Q(\pid.integral[2] ));
 sg13g2_dfrbp_1 _5514_ (.CLK(clknet_4_14__leaf_clk),
    .RESET_B(net481),
    .D(_0078_),
    .Q_N(_0011_),
    .Q(\pid.integral[3] ));
 sg13g2_dfrbp_1 _5515_ (.CLK(clknet_4_15__leaf_clk),
    .RESET_B(net482),
    .D(_0079_),
    .Q_N(_2736_),
    .Q(\pid.integral[4] ));
 sg13g2_dfrbp_1 _5516_ (.CLK(clknet_4_15__leaf_clk),
    .RESET_B(net482),
    .D(_0080_),
    .Q_N(_0010_),
    .Q(\pid.integral[5] ));
 sg13g2_dfrbp_1 _5517_ (.CLK(clknet_4_15__leaf_clk),
    .RESET_B(net482),
    .D(_0081_),
    .Q_N(_2735_),
    .Q(\pid.integral[6] ));
 sg13g2_dfrbp_1 _5518_ (.CLK(clknet_4_11__leaf_clk),
    .RESET_B(net481),
    .D(_0082_),
    .Q_N(_0009_),
    .Q(\pid.integral[7] ));
 sg13g2_dfrbp_1 _5519_ (.CLK(clknet_4_13__leaf_clk),
    .RESET_B(net481),
    .D(_0083_),
    .Q_N(_2734_),
    .Q(\pid.integral[8] ));
 sg13g2_dfrbp_1 _5520_ (.CLK(clknet_4_13__leaf_clk),
    .RESET_B(net484),
    .D(_0084_),
    .Q_N(_0008_),
    .Q(\pid.integral[9] ));
 sg13g2_dfrbp_1 _5521_ (.CLK(clknet_4_13__leaf_clk),
    .RESET_B(net484),
    .D(_0085_),
    .Q_N(_2733_),
    .Q(\pid.integral[10] ));
 sg13g2_dfrbp_1 _5522_ (.CLK(clknet_4_12__leaf_clk),
    .RESET_B(net484),
    .D(_0086_),
    .Q_N(_0007_),
    .Q(\pid.integral[11] ));
 sg13g2_dfrbp_1 _5523_ (.CLK(clknet_4_8__leaf_clk),
    .RESET_B(net484),
    .D(_0087_),
    .Q_N(_2732_),
    .Q(\pid.integral[12] ));
 sg13g2_dfrbp_1 _5524_ (.CLK(clknet_4_9__leaf_clk),
    .RESET_B(net484),
    .D(_0088_),
    .Q_N(_2731_),
    .Q(\pid.integral[13] ));
 sg13g2_dfrbp_1 _5525_ (.CLK(clknet_4_9__leaf_clk),
    .RESET_B(net481),
    .D(_0089_),
    .Q_N(_2730_),
    .Q(\pid.integral[14] ));
 sg13g2_dfrbp_1 _5526_ (.CLK(clknet_4_11__leaf_clk),
    .RESET_B(net481),
    .D(_0090_),
    .Q_N(_2729_),
    .Q(\pid.integral[15] ));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_pid_controller_18 (.L_LO(net18));
 sg13g2_tielo tt_um_pid_controller_19 (.L_LO(net19));
 sg13g2_tielo tt_um_pid_controller_20 (.L_LO(net20));
 sg13g2_tielo tt_um_pid_controller_21 (.L_LO(net21));
 sg13g2_tielo tt_um_pid_controller_22 (.L_LO(net22));
 sg13g2_tielo tt_um_pid_controller_23 (.L_LO(net23));
 sg13g2_tielo tt_um_pid_controller_24 (.L_LO(net24));
 sg13g2_tielo tt_um_pid_controller_25 (.L_LO(net25));
 sg13g2_tielo tt_um_pid_controller_26 (.L_LO(net26));
 sg13g2_tielo tt_um_pid_controller_27 (.L_LO(net27));
 sg13g2_tielo tt_um_pid_controller_28 (.L_LO(net28));
 sg13g2_tielo tt_um_pid_controller_29 (.L_LO(net29));
 sg13g2_tielo tt_um_pid_controller_30 (.L_LO(net30));
 sg13g2_tielo tt_um_pid_controller_31 (.L_LO(net31));
 sg13g2_tielo tt_um_pid_controller_32 (.L_LO(net32));
 sg13g2_tiehi _5472__33 (.L_HI(net33));
 sg13g2_buf_2 fanout369 (.A(_1699_),
    .X(net369));
 sg13g2_buf_8 fanout370 (.A(_0790_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_2544_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_2543_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_2543_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(net375),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(net376),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_0642_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(net378),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_1429_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_2077_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(net381),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_2084_),
    .X(net381));
 sg13g2_buf_4 fanout382 (.X(net382),
    .A(_2081_));
 sg13g2_buf_1 fanout383 (.A(_2081_),
    .X(net383));
 sg13g2_buf_4 fanout384 (.X(net384),
    .A(_0933_));
 sg13g2_buf_1 fanout385 (.A(_0933_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_2063_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_2063_),
    .X(net387));
 sg13g2_buf_4 fanout388 (.X(net388),
    .A(_2054_));
 sg13g2_buf_2 fanout389 (.A(_2038_),
    .X(net389));
 sg13g2_buf_4 fanout390 (.X(net390),
    .A(net391));
 sg13g2_buf_4 fanout391 (.X(net391),
    .A(_2037_));
 sg13g2_buf_8 fanout392 (.A(net395),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(net395),
    .X(net393));
 sg13g2_buf_8 fanout394 (.A(net395),
    .X(net394));
 sg13g2_buf_4 fanout395 (.X(net395),
    .A(_2035_));
 sg13g2_buf_4 fanout396 (.X(net396),
    .A(_0161_));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(_2055_));
 sg13g2_buf_2 fanout398 (.A(net400),
    .X(net398));
 sg13g2_buf_1 fanout399 (.A(net400),
    .X(net399));
 sg13g2_buf_8 fanout400 (.A(_2026_),
    .X(net400));
 sg13g2_buf_4 fanout401 (.X(net401),
    .A(_2100_));
 sg13g2_buf_8 fanout402 (.A(net403),
    .X(net402));
 sg13g2_buf_4 fanout403 (.X(net403),
    .A(net405));
 sg13g2_buf_4 fanout404 (.X(net404),
    .A(net51));
 sg13g2_buf_8 fanout405 (.A(_2016_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(net407),
    .X(net406));
 sg13g2_buf_4 fanout407 (.X(net407),
    .A(_1931_));
 sg13g2_buf_4 fanout408 (.X(net408),
    .A(net409));
 sg13g2_buf_2 fanout409 (.A(_1931_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(net411),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_2101_),
    .X(net411));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(_1822_));
 sg13g2_buf_2 fanout413 (.A(_1822_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(net415),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_1822_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(net417),
    .X(net416));
 sg13g2_buf_4 fanout417 (.X(net417),
    .A(_1757_));
 sg13g2_buf_4 fanout418 (.X(net418),
    .A(_1746_));
 sg13g2_buf_2 fanout419 (.A(_1746_),
    .X(net419));
 sg13g2_buf_4 fanout420 (.X(net420),
    .A(net424));
 sg13g2_buf_1 fanout421 (.A(net424),
    .X(net421));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(net423));
 sg13g2_buf_2 fanout423 (.A(net424),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_1659_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(net426),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(net430),
    .X(net426));
 sg13g2_buf_4 fanout427 (.X(net427),
    .A(net430));
 sg13g2_buf_1 fanout428 (.A(net430),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(net430),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_1561_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(net432),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(\pid.Kp[8] ),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(net434),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(\pid.Kp[7] ),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(\pid.Kp[6] ),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(net437),
    .X(net436));
 sg13g2_buf_1 fanout437 (.A(\pid.Kp[4] ),
    .X(net437));
 sg13g2_buf_4 fanout438 (.X(net438),
    .A(\pid.Kp[3] ));
 sg13g2_buf_4 fanout439 (.X(net439),
    .A(\pid.Kp[2] ));
 sg13g2_buf_4 fanout440 (.X(net440),
    .A(\pid.Kp[1] ));
 sg13g2_buf_4 fanout441 (.X(net441),
    .A(\pid.Kp[0] ));
 sg13g2_buf_4 fanout442 (.X(net442),
    .A(\pid.Ki[8] ));
 sg13g2_buf_2 fanout443 (.A(\pid.Ki[7] ),
    .X(net443));
 sg13g2_buf_4 fanout444 (.X(net444),
    .A(\pid.Ki[6] ));
 sg13g2_buf_4 fanout445 (.X(net445),
    .A(\pid.Ki[4] ));
 sg13g2_buf_4 fanout446 (.X(net446),
    .A(\pid.Ki[3] ));
 sg13g2_buf_2 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_4 fanout448 (.X(net448),
    .A(\pid.Ki[2] ));
 sg13g2_buf_4 fanout449 (.X(net449),
    .A(\pid.Ki[0] ));
 sg13g2_buf_1 fanout450 (.A(\pid.Ki[0] ),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(\pid.state[3] ),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(net454),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(net454),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(net136),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(net457),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(net457),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(net123),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(net459),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(net133),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(net133),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(net161),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(net162),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(net152),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(net159),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(net156),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(net154),
    .X(net466));
 sg13g2_buf_1 fanout467 (.A(\pid.Kd[2] ),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(net160),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(net140),
    .X(net470));
 sg13g2_buf_4 fanout471 (.X(net471),
    .A(_1594_));
 sg13g2_buf_2 fanout472 (.A(_1594_),
    .X(net472));
 sg13g2_buf_4 fanout473 (.X(net473),
    .A(_1594_));
 sg13g2_buf_2 fanout474 (.A(net3),
    .X(net474));
 sg13g2_buf_16 fanout475 (.X(net475),
    .A(net2));
 sg13g2_buf_4 fanout476 (.X(net476),
    .A(net477));
 sg13g2_buf_4 fanout477 (.X(net477),
    .A(net485));
 sg13g2_buf_4 fanout478 (.X(net478),
    .A(net479));
 sg13g2_buf_4 fanout479 (.X(net479),
    .A(net480));
 sg13g2_buf_4 fanout480 (.X(net480),
    .A(net485));
 sg13g2_buf_4 fanout481 (.X(net481),
    .A(net484));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(net485));
 sg13g2_buf_4 fanout483 (.X(net483),
    .A(net484));
 sg13g2_buf_4 fanout484 (.X(net484),
    .A(net485));
 sg13g2_buf_2 fanout485 (.A(rst_n),
    .X(net485));
 sg13g2_buf_4 input1 (.X(net1),
    .A(ui_in[0]));
 sg13g2_buf_16 input2 (.X(net2),
    .A(ui_in[1]));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[2]));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[3]));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[4]));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[5]));
 sg13g2_buf_4 input7 (.X(net7),
    .A(ui_in[6]));
 sg13g2_buf_4 input8 (.X(net8),
    .A(ui_in[7]));
 sg13g2_buf_4 input9 (.X(net9),
    .A(uio_in[0]));
 sg13g2_buf_2 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_4 input13 (.X(net13),
    .A(uio_in[4]));
 sg13g2_buf_4 input14 (.X(net14),
    .A(uio_in[5]));
 sg13g2_buf_4 input15 (.X(net15),
    .A(uio_in[6]));
 sg13g2_buf_4 input16 (.X(net16),
    .A(uio_in[7]));
 sg13g2_tielo tt_um_pid_controller_17 (.L_LO(net17));
 sg13g2_buf_2 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_2 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_2 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_2 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_2 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_2 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_2 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_2 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_2 clkbuf_4_0__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_0__leaf_clk));
 sg13g2_buf_2 clkbuf_4_1__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_1__leaf_clk));
 sg13g2_buf_2 clkbuf_4_2__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_2__leaf_clk));
 sg13g2_buf_2 clkbuf_4_3__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_3__leaf_clk));
 sg13g2_buf_2 clkbuf_4_4__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_4__leaf_clk));
 sg13g2_buf_2 clkbuf_4_5__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_5__leaf_clk));
 sg13g2_buf_2 clkbuf_4_6__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_6__leaf_clk));
 sg13g2_buf_2 clkbuf_4_7__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_7__leaf_clk));
 sg13g2_buf_2 clkbuf_4_8__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_8__leaf_clk));
 sg13g2_buf_2 clkbuf_4_9__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_9__leaf_clk));
 sg13g2_buf_2 clkbuf_4_10__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_10__leaf_clk));
 sg13g2_buf_2 clkbuf_4_11__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_11__leaf_clk));
 sg13g2_buf_2 clkbuf_4_12__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_12__leaf_clk));
 sg13g2_buf_2 clkbuf_4_13__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_13__leaf_clk));
 sg13g2_buf_2 clkbuf_4_14__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_14__leaf_clk));
 sg13g2_buf_2 clkbuf_4_15__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_15__leaf_clk));
 sg13g2_dlygate4sd1_1 rebuffer1 (.A(_0775_),
    .X(net34));
 sg13g2_dlygate4sd1_1 rebuffer2 (.A(_0722_),
    .X(net35));
 sg13g2_buf_1 rebuffer3 (.A(net67),
    .X(net36));
 sg13g2_buf_2 rebuffer4 (.A(net67),
    .X(net37));
 sg13g2_buf_2 rebuffer5 (.A(net67),
    .X(net38));
 sg13g2_buf_1 rebuffer6 (.A(_0617_),
    .X(net39));
 sg13g2_dlygate4sd1_1 rebuffer7 (.A(_0612_),
    .X(net40));
 sg13g2_buf_2 rebuffer8 (.A(_0524_),
    .X(net41));
 sg13g2_dlygate4sd1_1 rebuffer9 (.A(_0455_),
    .X(net42));
 sg13g2_dlygate4sd1_1 rebuffer10 (.A(_0607_),
    .X(net43));
 sg13g2_dlygate4sd1_1 rebuffer11 (.A(_0741_),
    .X(net44));
 sg13g2_buf_1 rebuffer12 (.A(_0617_),
    .X(net45));
 sg13g2_dlygate4sd1_1 rebuffer13 (.A(_1909_),
    .X(net46));
 sg13g2_dlygate4sd1_1 rebuffer14 (.A(_0519_),
    .X(net47));
 sg13g2_dlygate4sd1_1 rebuffer15 (.A(_0709_),
    .X(net48));
 sg13g2_dlygate4sd1_1 rebuffer16 (.A(_0491_),
    .X(net49));
 sg13g2_dlygate4sd1_1 rebuffer17 (.A(net81),
    .X(net50));
 sg13g2_buf_2 rebuffer18 (.A(net405),
    .X(net51));
 sg13g2_dlygate4sd1_1 rebuffer19 (.A(net51),
    .X(net52));
 sg13g2_buf_1 rebuffer20 (.A(_2034_),
    .X(net53));
 sg13g2_dlygate4sd1_1 rebuffer21 (.A(_2034_),
    .X(net54));
 sg13g2_buf_2 rebuffer22 (.A(_2034_),
    .X(net55));
 sg13g2_dlygate4sd1_1 rebuffer23 (.A(_1515_),
    .X(net56));
 sg13g2_dlygate4sd1_1 rebuffer24 (.A(_0604_),
    .X(net57));
 sg13g2_dlygate4sd1_1 rebuffer25 (.A(_1309_),
    .X(net58));
 sg13g2_dlygate4sd1_1 rebuffer26 (.A(_0486_),
    .X(net59));
 sg13g2_buf_1 rebuffer27 (.A(_2033_),
    .X(net60));
 sg13g2_dlygate4sd1_1 rebuffer28 (.A(_2033_),
    .X(net61));
 sg13g2_dlygate4sd1_1 rebuffer29 (.A(net61),
    .X(net62));
 sg13g2_dlygate4sd1_1 rebuffer30 (.A(_1245_),
    .X(net63));
 sg13g2_dlygate4sd1_1 rebuffer31 (.A(_1371_),
    .X(net64));
 sg13g2_dlygate4sd1_1 rebuffer32 (.A(_1240_),
    .X(net65));
 sg13g2_buf_1 rebuffer33 (.A(_1876_),
    .X(net66));
 sg13g2_buf_8 rebuffer34 (.A(net85),
    .X(net67));
 sg13g2_dlygate4sd1_1 rebuffer35 (.A(_0456_),
    .X(net68));
 sg13g2_buf_1 rebuffer36 (.A(net76),
    .X(net69));
 sg13g2_dlygate4sd1_1 rebuffer37 (.A(_0443_),
    .X(net70));
 sg13g2_dlygate4sd1_1 rebuffer38 (.A(_0406_),
    .X(net71));
 sg13g2_dlygate4sd1_1 rebuffer39 (.A(_1377_),
    .X(net72));
 sg13g2_dlygate4sd1_1 rebuffer40 (.A(_1238_),
    .X(net73));
 sg13g2_dlygate4sd1_1 rebuffer41 (.A(_1193_),
    .X(net74));
 sg13g2_dlygate4sd1_1 rebuffer42 (.A(_1160_),
    .X(net75));
 sg13g2_buf_1 rebuffer43 (.A(net84),
    .X(net76));
 sg13g2_dlygate4sd1_1 rebuffer44 (.A(_1205_),
    .X(net77));
 sg13g2_buf_2 rebuffer45 (.A(_0362_),
    .X(net78));
 sg13g2_dlygate4sd1_1 rebuffer46 (.A(_1162_),
    .X(net79));
 sg13g2_buf_1 rebuffer47 (.A(_2025_),
    .X(net80));
 sg13g2_dlygate4sd3_1 rebuffer48 (.A(_2001_),
    .X(net81));
 sg13g2_dlygate4sd1_1 rebuffer49 (.A(_2001_),
    .X(net82));
 sg13g2_dlygate4sd1_1 rebuffer50 (.A(_1648_),
    .X(net83));
 sg13g2_buf_1 rebuffer51 (.A(_2025_),
    .X(net84));
 sg13g2_buf_2 rebuffer52 (.A(_1876_),
    .X(net85));
 sg13g2_dlygate4sd1_1 rebuffer53 (.A(_1236_),
    .X(net86));
 sg13g2_buf_2 rebuffer54 (.A(_2516_),
    .X(net87));
 sg13g2_buf_8 rebuffer55 (.A(_1982_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold56 (.A(\pid.integral[7] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold57 (.A(\pid.integral[1] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold58 (.A(\pid.integral[3] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold59 (.A(\pid.integral[9] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold60 (.A(\pid.integral[5] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold61 (.A(\pid.integral[14] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold62 (.A(\pid.prev_error[7] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold63 (.A(\pid.integral[11] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold64 (.A(\pid.integral[15] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold65 (.A(\pid.Ki[1] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0041_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold67 (.A(\pid.prev_error[8] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold68 (.A(uo_out[0]),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold69 (.A(_2040_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold70 (.A(\pid.integral[2] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold71 (.A(uo_out[3]),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold72 (.A(_1992_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold73 (.A(uo_out[1]),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold74 (.A(_1988_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold75 (.A(uo_out[2]),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold76 (.A(_1990_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold77 (.A(\pid.prev_error[1] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold78 (.A(\pid.prev_error[4] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold79 (.A(\pid.integral[12] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold80 (.A(\pid.integral[4] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold81 (.A(uo_out[5]),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold82 (.A(_1997_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold83 (.A(\pid.integral[13] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold84 (.A(uo_out[4]),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold85 (.A(_1995_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold86 (.A(\pid.prev_error[2] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0051_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold88 (.A(\pid.integral[0] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold89 (.A(\pid.prev_error[6] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold90 (.A(\pid.state[1] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0000_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold92 (.A(\pid.integral[10] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold93 (.A(\pid.prev_error[3] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold94 (.A(uo_out[6]),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold95 (.A(_1999_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold96 (.A(uo_out[7]),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold97 (.A(_2002_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold98 (.A(\pid.integral[8] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold99 (.A(\pid.integral[6] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold100 (.A(\pid.state[0] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold101 (.A(\pid.prev_error[0] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold102 (.A(\pid.prev_error[5] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold103 (.A(\pid.state[2] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0045_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold105 (.A(\pid.Kd[3] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold106 (.A(net437),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold107 (.A(\pid.Kd[0] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold108 (.A(net434),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold109 (.A(net449),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold110 (.A(net432),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold111 (.A(\pid.Kp[5] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold112 (.A(net441),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold113 (.A(net446),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold114 (.A(net440),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold115 (.A(net439),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold116 (.A(net442),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold117 (.A(net438),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold118 (.A(net435),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold119 (.A(\pid.Kd[6] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold120 (.A(net445),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold121 (.A(\pid.Kd[2] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold122 (.A(net444),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold123 (.A(\pid.Kd[4] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold124 (.A(net448),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold125 (.A(net443),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold126 (.A(\pid.Kd[5] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold127 (.A(\pid.Kd[1] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold128 (.A(\pid.Kd[8] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold129 (.A(\pid.Kd[7] ),
    .X(net162));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_4 FILLER_0_154 ();
 sg13g2_fill_1 FILLER_0_158 ();
 sg13g2_fill_2 FILLER_0_163 ();
 sg13g2_fill_1 FILLER_0_165 ();
 sg13g2_decap_4 FILLER_0_172 ();
 sg13g2_fill_1 FILLER_0_176 ();
 sg13g2_fill_2 FILLER_0_180 ();
 sg13g2_decap_8 FILLER_0_188 ();
 sg13g2_decap_8 FILLER_0_202 ();
 sg13g2_decap_8 FILLER_0_209 ();
 sg13g2_decap_8 FILLER_0_216 ();
 sg13g2_decap_8 FILLER_0_223 ();
 sg13g2_decap_8 FILLER_0_230 ();
 sg13g2_fill_1 FILLER_0_237 ();
 sg13g2_decap_8 FILLER_0_248 ();
 sg13g2_decap_8 FILLER_0_255 ();
 sg13g2_decap_8 FILLER_0_262 ();
 sg13g2_decap_8 FILLER_0_274 ();
 sg13g2_decap_8 FILLER_0_281 ();
 sg13g2_fill_2 FILLER_0_288 ();
 sg13g2_fill_1 FILLER_0_290 ();
 sg13g2_decap_8 FILLER_0_296 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_310 ();
 sg13g2_decap_8 FILLER_0_317 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_4 FILLER_1_133 ();
 sg13g2_fill_1 FILLER_1_137 ();
 sg13g2_fill_1 FILLER_1_171 ();
 sg13g2_fill_1 FILLER_1_188 ();
 sg13g2_fill_1 FILLER_1_201 ();
 sg13g2_fill_2 FILLER_1_214 ();
 sg13g2_fill_1 FILLER_1_216 ();
 sg13g2_fill_2 FILLER_1_230 ();
 sg13g2_fill_1 FILLER_1_232 ();
 sg13g2_decap_4 FILLER_1_254 ();
 sg13g2_fill_1 FILLER_1_258 ();
 sg13g2_fill_2 FILLER_1_279 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_4 FILLER_2_126 ();
 sg13g2_fill_2 FILLER_2_130 ();
 sg13g2_fill_2 FILLER_2_156 ();
 sg13g2_fill_2 FILLER_2_233 ();
 sg13g2_fill_2 FILLER_2_259 ();
 sg13g2_fill_1 FILLER_2_261 ();
 sg13g2_decap_8 FILLER_2_320 ();
 sg13g2_decap_8 FILLER_2_327 ();
 sg13g2_decap_8 FILLER_2_334 ();
 sg13g2_decap_8 FILLER_2_341 ();
 sg13g2_decap_8 FILLER_2_348 ();
 sg13g2_decap_8 FILLER_2_355 ();
 sg13g2_decap_8 FILLER_2_362 ();
 sg13g2_decap_8 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_376 ();
 sg13g2_decap_8 FILLER_2_383 ();
 sg13g2_decap_8 FILLER_2_390 ();
 sg13g2_decap_8 FILLER_2_397 ();
 sg13g2_decap_4 FILLER_2_404 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_fill_1 FILLER_3_126 ();
 sg13g2_fill_2 FILLER_3_160 ();
 sg13g2_fill_1 FILLER_3_196 ();
 sg13g2_fill_1 FILLER_3_297 ();
 sg13g2_decap_8 FILLER_3_314 ();
 sg13g2_decap_8 FILLER_3_321 ();
 sg13g2_decap_8 FILLER_3_328 ();
 sg13g2_decap_8 FILLER_3_335 ();
 sg13g2_decap_8 FILLER_3_342 ();
 sg13g2_decap_8 FILLER_3_349 ();
 sg13g2_decap_8 FILLER_3_356 ();
 sg13g2_decap_8 FILLER_3_363 ();
 sg13g2_decap_8 FILLER_3_370 ();
 sg13g2_decap_8 FILLER_3_377 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_4 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_4 FILLER_4_112 ();
 sg13g2_fill_1 FILLER_4_159 ();
 sg13g2_fill_2 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_170 ();
 sg13g2_fill_2 FILLER_4_184 ();
 sg13g2_decap_8 FILLER_4_198 ();
 sg13g2_decap_8 FILLER_4_205 ();
 sg13g2_fill_2 FILLER_4_212 ();
 sg13g2_decap_4 FILLER_4_235 ();
 sg13g2_fill_1 FILLER_4_239 ();
 sg13g2_decap_8 FILLER_4_248 ();
 sg13g2_decap_8 FILLER_4_255 ();
 sg13g2_decap_4 FILLER_4_262 ();
 sg13g2_decap_8 FILLER_4_275 ();
 sg13g2_decap_8 FILLER_4_282 ();
 sg13g2_decap_4 FILLER_4_289 ();
 sg13g2_decap_4 FILLER_4_297 ();
 sg13g2_fill_2 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_321 ();
 sg13g2_decap_8 FILLER_4_328 ();
 sg13g2_decap_8 FILLER_4_335 ();
 sg13g2_decap_8 FILLER_4_342 ();
 sg13g2_decap_8 FILLER_4_349 ();
 sg13g2_decap_8 FILLER_4_356 ();
 sg13g2_decap_8 FILLER_4_363 ();
 sg13g2_decap_8 FILLER_4_370 ();
 sg13g2_decap_8 FILLER_4_377 ();
 sg13g2_decap_8 FILLER_4_384 ();
 sg13g2_decap_8 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_fill_2 FILLER_5_126 ();
 sg13g2_fill_2 FILLER_5_148 ();
 sg13g2_fill_1 FILLER_5_150 ();
 sg13g2_fill_1 FILLER_5_167 ();
 sg13g2_fill_2 FILLER_5_180 ();
 sg13g2_fill_2 FILLER_5_187 ();
 sg13g2_fill_1 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_194 ();
 sg13g2_decap_8 FILLER_5_201 ();
 sg13g2_decap_8 FILLER_5_208 ();
 sg13g2_decap_8 FILLER_5_215 ();
 sg13g2_decap_8 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_229 ();
 sg13g2_decap_4 FILLER_5_236 ();
 sg13g2_fill_2 FILLER_5_240 ();
 sg13g2_decap_8 FILLER_5_272 ();
 sg13g2_fill_2 FILLER_5_287 ();
 sg13g2_fill_2 FILLER_5_298 ();
 sg13g2_fill_1 FILLER_5_300 ();
 sg13g2_fill_2 FILLER_5_306 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_4 FILLER_6_126 ();
 sg13g2_fill_2 FILLER_6_130 ();
 sg13g2_fill_2 FILLER_6_148 ();
 sg13g2_decap_8 FILLER_6_162 ();
 sg13g2_fill_2 FILLER_6_185 ();
 sg13g2_fill_2 FILLER_6_195 ();
 sg13g2_fill_1 FILLER_6_197 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_4 FILLER_6_217 ();
 sg13g2_fill_1 FILLER_6_230 ();
 sg13g2_fill_2 FILLER_6_275 ();
 sg13g2_fill_1 FILLER_6_282 ();
 sg13g2_fill_2 FILLER_6_291 ();
 sg13g2_decap_8 FILLER_6_317 ();
 sg13g2_decap_8 FILLER_6_324 ();
 sg13g2_decap_8 FILLER_6_331 ();
 sg13g2_decap_8 FILLER_6_338 ();
 sg13g2_decap_8 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_352 ();
 sg13g2_decap_8 FILLER_6_359 ();
 sg13g2_decap_8 FILLER_6_366 ();
 sg13g2_decap_8 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_fill_1 FILLER_7_150 ();
 sg13g2_fill_1 FILLER_7_159 ();
 sg13g2_fill_2 FILLER_7_188 ();
 sg13g2_fill_2 FILLER_7_211 ();
 sg13g2_fill_1 FILLER_7_213 ();
 sg13g2_fill_2 FILLER_7_248 ();
 sg13g2_fill_1 FILLER_7_290 ();
 sg13g2_fill_2 FILLER_7_296 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_4 FILLER_8_119 ();
 sg13g2_fill_2 FILLER_8_123 ();
 sg13g2_fill_2 FILLER_8_146 ();
 sg13g2_decap_8 FILLER_8_156 ();
 sg13g2_decap_4 FILLER_8_163 ();
 sg13g2_fill_1 FILLER_8_167 ();
 sg13g2_decap_4 FILLER_8_189 ();
 sg13g2_fill_1 FILLER_8_193 ();
 sg13g2_fill_2 FILLER_8_262 ();
 sg13g2_fill_1 FILLER_8_264 ();
 sg13g2_decap_4 FILLER_8_269 ();
 sg13g2_fill_1 FILLER_8_273 ();
 sg13g2_fill_2 FILLER_8_281 ();
 sg13g2_decap_8 FILLER_8_311 ();
 sg13g2_decap_8 FILLER_8_318 ();
 sg13g2_decap_8 FILLER_8_325 ();
 sg13g2_decap_8 FILLER_8_332 ();
 sg13g2_decap_8 FILLER_8_339 ();
 sg13g2_decap_8 FILLER_8_346 ();
 sg13g2_decap_8 FILLER_8_353 ();
 sg13g2_decap_8 FILLER_8_360 ();
 sg13g2_decap_8 FILLER_8_367 ();
 sg13g2_decap_8 FILLER_8_374 ();
 sg13g2_decap_8 FILLER_8_381 ();
 sg13g2_decap_8 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_4 FILLER_9_119 ();
 sg13g2_fill_1 FILLER_9_123 ();
 sg13g2_fill_1 FILLER_9_147 ();
 sg13g2_fill_2 FILLER_9_156 ();
 sg13g2_decap_4 FILLER_9_166 ();
 sg13g2_fill_2 FILLER_9_179 ();
 sg13g2_fill_1 FILLER_9_181 ();
 sg13g2_decap_8 FILLER_9_194 ();
 sg13g2_fill_2 FILLER_9_201 ();
 sg13g2_fill_2 FILLER_9_216 ();
 sg13g2_fill_1 FILLER_9_218 ();
 sg13g2_fill_2 FILLER_9_244 ();
 sg13g2_fill_1 FILLER_9_246 ();
 sg13g2_decap_8 FILLER_9_251 ();
 sg13g2_decap_8 FILLER_9_258 ();
 sg13g2_decap_8 FILLER_9_268 ();
 sg13g2_decap_4 FILLER_9_275 ();
 sg13g2_fill_1 FILLER_9_279 ();
 sg13g2_fill_2 FILLER_9_284 ();
 sg13g2_fill_1 FILLER_9_286 ();
 sg13g2_decap_8 FILLER_9_296 ();
 sg13g2_decap_8 FILLER_9_303 ();
 sg13g2_decap_8 FILLER_9_323 ();
 sg13g2_decap_8 FILLER_9_330 ();
 sg13g2_decap_8 FILLER_9_337 ();
 sg13g2_decap_8 FILLER_9_344 ();
 sg13g2_decap_8 FILLER_9_351 ();
 sg13g2_decap_8 FILLER_9_358 ();
 sg13g2_decap_8 FILLER_9_365 ();
 sg13g2_decap_8 FILLER_9_372 ();
 sg13g2_decap_8 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_fill_2 FILLER_10_112 ();
 sg13g2_fill_1 FILLER_10_114 ();
 sg13g2_fill_2 FILLER_10_160 ();
 sg13g2_fill_1 FILLER_10_162 ();
 sg13g2_fill_2 FILLER_10_184 ();
 sg13g2_fill_1 FILLER_10_186 ();
 sg13g2_decap_4 FILLER_10_205 ();
 sg13g2_fill_2 FILLER_10_209 ();
 sg13g2_fill_1 FILLER_10_215 ();
 sg13g2_fill_2 FILLER_10_221 ();
 sg13g2_fill_1 FILLER_10_223 ();
 sg13g2_fill_1 FILLER_10_232 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_fill_2 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_261 ();
 sg13g2_fill_1 FILLER_10_268 ();
 sg13g2_fill_2 FILLER_10_286 ();
 sg13g2_fill_1 FILLER_10_288 ();
 sg13g2_decap_8 FILLER_10_297 ();
 sg13g2_decap_8 FILLER_10_330 ();
 sg13g2_decap_8 FILLER_10_337 ();
 sg13g2_decap_8 FILLER_10_344 ();
 sg13g2_decap_8 FILLER_10_351 ();
 sg13g2_decap_8 FILLER_10_358 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_fill_2 FILLER_11_119 ();
 sg13g2_fill_1 FILLER_11_134 ();
 sg13g2_fill_2 FILLER_11_151 ();
 sg13g2_decap_4 FILLER_11_174 ();
 sg13g2_fill_2 FILLER_11_183 ();
 sg13g2_fill_1 FILLER_11_185 ();
 sg13g2_decap_8 FILLER_11_194 ();
 sg13g2_decap_4 FILLER_11_206 ();
 sg13g2_fill_2 FILLER_11_238 ();
 sg13g2_fill_1 FILLER_11_250 ();
 sg13g2_fill_2 FILLER_11_291 ();
 sg13g2_decap_8 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_325 ();
 sg13g2_decap_8 FILLER_11_332 ();
 sg13g2_decap_8 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_4 FILLER_12_112 ();
 sg13g2_fill_2 FILLER_12_116 ();
 sg13g2_fill_2 FILLER_12_172 ();
 sg13g2_fill_1 FILLER_12_174 ();
 sg13g2_decap_4 FILLER_12_183 ();
 sg13g2_fill_1 FILLER_12_187 ();
 sg13g2_fill_2 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_215 ();
 sg13g2_fill_2 FILLER_12_222 ();
 sg13g2_fill_1 FILLER_12_224 ();
 sg13g2_fill_1 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_314 ();
 sg13g2_decap_8 FILLER_12_321 ();
 sg13g2_decap_8 FILLER_12_328 ();
 sg13g2_decap_8 FILLER_12_335 ();
 sg13g2_decap_8 FILLER_12_342 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_356 ();
 sg13g2_decap_8 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_370 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_4 FILLER_13_112 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_fill_2 FILLER_13_134 ();
 sg13g2_decap_8 FILLER_13_150 ();
 sg13g2_decap_8 FILLER_13_157 ();
 sg13g2_decap_4 FILLER_13_164 ();
 sg13g2_fill_1 FILLER_13_168 ();
 sg13g2_fill_2 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_decap_4 FILLER_13_207 ();
 sg13g2_fill_2 FILLER_13_211 ();
 sg13g2_decap_8 FILLER_13_223 ();
 sg13g2_decap_4 FILLER_13_230 ();
 sg13g2_fill_1 FILLER_13_234 ();
 sg13g2_decap_4 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_300 ();
 sg13g2_decap_8 FILLER_13_307 ();
 sg13g2_decap_8 FILLER_13_314 ();
 sg13g2_decap_8 FILLER_13_321 ();
 sg13g2_decap_8 FILLER_13_328 ();
 sg13g2_decap_8 FILLER_13_335 ();
 sg13g2_decap_8 FILLER_13_342 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_fill_1 FILLER_14_126 ();
 sg13g2_fill_2 FILLER_14_132 ();
 sg13g2_fill_2 FILLER_14_151 ();
 sg13g2_fill_1 FILLER_14_153 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_fill_2 FILLER_14_165 ();
 sg13g2_fill_1 FILLER_14_167 ();
 sg13g2_decap_8 FILLER_14_181 ();
 sg13g2_decap_8 FILLER_14_188 ();
 sg13g2_fill_2 FILLER_14_195 ();
 sg13g2_decap_8 FILLER_14_236 ();
 sg13g2_decap_8 FILLER_14_243 ();
 sg13g2_decap_8 FILLER_14_254 ();
 sg13g2_decap_8 FILLER_14_261 ();
 sg13g2_fill_1 FILLER_14_268 ();
 sg13g2_decap_8 FILLER_14_277 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_decap_4 FILLER_14_291 ();
 sg13g2_fill_1 FILLER_14_295 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_fill_1 FILLER_15_119 ();
 sg13g2_fill_1 FILLER_15_142 ();
 sg13g2_fill_1 FILLER_15_250 ();
 sg13g2_decap_4 FILLER_15_256 ();
 sg13g2_fill_2 FILLER_15_260 ();
 sg13g2_fill_1 FILLER_15_284 ();
 sg13g2_fill_1 FILLER_15_294 ();
 sg13g2_fill_2 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_328 ();
 sg13g2_decap_8 FILLER_15_335 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_decap_8 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_fill_2 FILLER_16_128 ();
 sg13g2_fill_1 FILLER_16_138 ();
 sg13g2_fill_1 FILLER_16_147 ();
 sg13g2_fill_2 FILLER_16_217 ();
 sg13g2_fill_1 FILLER_16_219 ();
 sg13g2_decap_4 FILLER_16_235 ();
 sg13g2_fill_2 FILLER_16_239 ();
 sg13g2_fill_2 FILLER_16_270 ();
 sg13g2_fill_2 FILLER_16_290 ();
 sg13g2_fill_1 FILLER_16_292 ();
 sg13g2_decap_8 FILLER_16_318 ();
 sg13g2_decap_8 FILLER_16_325 ();
 sg13g2_decap_8 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_fill_2 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_121 ();
 sg13g2_fill_1 FILLER_17_138 ();
 sg13g2_fill_2 FILLER_17_144 ();
 sg13g2_fill_1 FILLER_17_146 ();
 sg13g2_fill_2 FILLER_17_151 ();
 sg13g2_decap_4 FILLER_17_188 ();
 sg13g2_fill_1 FILLER_17_192 ();
 sg13g2_fill_1 FILLER_17_198 ();
 sg13g2_fill_2 FILLER_17_264 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_fill_2 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_121 ();
 sg13g2_fill_1 FILLER_18_137 ();
 sg13g2_fill_2 FILLER_18_148 ();
 sg13g2_fill_1 FILLER_18_150 ();
 sg13g2_decap_8 FILLER_18_159 ();
 sg13g2_decap_4 FILLER_18_169 ();
 sg13g2_fill_2 FILLER_18_173 ();
 sg13g2_fill_1 FILLER_18_188 ();
 sg13g2_fill_2 FILLER_18_213 ();
 sg13g2_fill_1 FILLER_18_215 ();
 sg13g2_fill_2 FILLER_18_221 ();
 sg13g2_fill_1 FILLER_18_223 ();
 sg13g2_fill_2 FILLER_18_232 ();
 sg13g2_fill_1 FILLER_18_234 ();
 sg13g2_fill_2 FILLER_18_267 ();
 sg13g2_fill_1 FILLER_18_269 ();
 sg13g2_decap_8 FILLER_18_299 ();
 sg13g2_decap_8 FILLER_18_306 ();
 sg13g2_fill_2 FILLER_18_313 ();
 sg13g2_decap_8 FILLER_18_320 ();
 sg13g2_fill_2 FILLER_18_331 ();
 sg13g2_fill_1 FILLER_18_333 ();
 sg13g2_decap_4 FILLER_18_344 ();
 sg13g2_fill_2 FILLER_18_348 ();
 sg13g2_decap_8 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_fill_2 FILLER_19_147 ();
 sg13g2_fill_1 FILLER_19_149 ();
 sg13g2_fill_1 FILLER_19_159 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_fill_2 FILLER_19_223 ();
 sg13g2_fill_2 FILLER_19_249 ();
 sg13g2_fill_1 FILLER_19_251 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_decap_4 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_293 ();
 sg13g2_fill_2 FILLER_19_300 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_decap_8 FILLER_19_370 ();
 sg13g2_decap_8 FILLER_19_377 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_138 ();
 sg13g2_fill_2 FILLER_20_149 ();
 sg13g2_decap_4 FILLER_20_172 ();
 sg13g2_fill_2 FILLER_20_176 ();
 sg13g2_fill_2 FILLER_20_182 ();
 sg13g2_fill_1 FILLER_20_184 ();
 sg13g2_decap_4 FILLER_20_194 ();
 sg13g2_fill_1 FILLER_20_198 ();
 sg13g2_decap_8 FILLER_20_212 ();
 sg13g2_decap_4 FILLER_20_219 ();
 sg13g2_fill_2 FILLER_20_223 ();
 sg13g2_decap_8 FILLER_20_234 ();
 sg13g2_fill_2 FILLER_20_241 ();
 sg13g2_fill_1 FILLER_20_243 ();
 sg13g2_decap_8 FILLER_20_278 ();
 sg13g2_decap_8 FILLER_20_285 ();
 sg13g2_fill_1 FILLER_20_292 ();
 sg13g2_fill_1 FILLER_20_310 ();
 sg13g2_fill_2 FILLER_20_319 ();
 sg13g2_fill_1 FILLER_20_321 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_fill_2 FILLER_21_162 ();
 sg13g2_fill_2 FILLER_21_174 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_fill_2 FILLER_21_203 ();
 sg13g2_fill_1 FILLER_21_205 ();
 sg13g2_decap_8 FILLER_21_215 ();
 sg13g2_decap_8 FILLER_21_222 ();
 sg13g2_decap_4 FILLER_21_229 ();
 sg13g2_fill_2 FILLER_21_238 ();
 sg13g2_fill_2 FILLER_21_248 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_fill_2 FILLER_21_266 ();
 sg13g2_fill_1 FILLER_21_268 ();
 sg13g2_fill_2 FILLER_21_294 ();
 sg13g2_fill_1 FILLER_21_296 ();
 sg13g2_fill_2 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_350 ();
 sg13g2_fill_1 FILLER_21_363 ();
 sg13g2_decap_8 FILLER_21_377 ();
 sg13g2_decap_8 FILLER_21_384 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_fill_2 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_107 ();
 sg13g2_fill_2 FILLER_22_153 ();
 sg13g2_fill_1 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_4 FILLER_22_196 ();
 sg13g2_fill_2 FILLER_22_221 ();
 sg13g2_fill_1 FILLER_22_223 ();
 sg13g2_fill_1 FILLER_22_233 ();
 sg13g2_fill_1 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_324 ();
 sg13g2_fill_1 FILLER_22_331 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_119 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_decap_4 FILLER_23_149 ();
 sg13g2_fill_2 FILLER_23_153 ();
 sg13g2_decap_8 FILLER_23_167 ();
 sg13g2_decap_8 FILLER_23_174 ();
 sg13g2_decap_8 FILLER_23_181 ();
 sg13g2_fill_2 FILLER_23_188 ();
 sg13g2_decap_4 FILLER_23_194 ();
 sg13g2_fill_2 FILLER_23_198 ();
 sg13g2_decap_4 FILLER_23_205 ();
 sg13g2_fill_1 FILLER_23_209 ();
 sg13g2_fill_2 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_225 ();
 sg13g2_fill_2 FILLER_23_238 ();
 sg13g2_fill_1 FILLER_23_297 ();
 sg13g2_decap_8 FILLER_23_334 ();
 sg13g2_decap_8 FILLER_23_341 ();
 sg13g2_decap_4 FILLER_23_348 ();
 sg13g2_fill_2 FILLER_23_352 ();
 sg13g2_decap_8 FILLER_23_359 ();
 sg13g2_decap_8 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_4 FILLER_24_126 ();
 sg13g2_fill_2 FILLER_24_130 ();
 sg13g2_decap_8 FILLER_24_143 ();
 sg13g2_decap_8 FILLER_24_150 ();
 sg13g2_decap_8 FILLER_24_157 ();
 sg13g2_decap_8 FILLER_24_169 ();
 sg13g2_fill_2 FILLER_24_176 ();
 sg13g2_fill_2 FILLER_24_224 ();
 sg13g2_fill_1 FILLER_24_226 ();
 sg13g2_decap_8 FILLER_24_254 ();
 sg13g2_fill_2 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_326 ();
 sg13g2_decap_4 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_353 ();
 sg13g2_decap_4 FILLER_24_360 ();
 sg13g2_fill_2 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_119 ();
 sg13g2_fill_1 FILLER_25_121 ();
 sg13g2_decap_4 FILLER_25_155 ();
 sg13g2_fill_2 FILLER_25_198 ();
 sg13g2_decap_8 FILLER_25_205 ();
 sg13g2_decap_4 FILLER_25_212 ();
 sg13g2_fill_2 FILLER_25_216 ();
 sg13g2_decap_8 FILLER_25_228 ();
 sg13g2_fill_2 FILLER_25_235 ();
 sg13g2_decap_8 FILLER_25_246 ();
 sg13g2_decap_8 FILLER_25_253 ();
 sg13g2_decap_8 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_267 ();
 sg13g2_fill_2 FILLER_25_281 ();
 sg13g2_fill_1 FILLER_25_283 ();
 sg13g2_decap_8 FILLER_25_288 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_fill_2 FILLER_25_321 ();
 sg13g2_decap_4 FILLER_25_336 ();
 sg13g2_fill_2 FILLER_25_361 ();
 sg13g2_fill_1 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_79 ();
 sg13g2_decap_8 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_95 ();
 sg13g2_decap_8 FILLER_26_102 ();
 sg13g2_decap_8 FILLER_26_109 ();
 sg13g2_fill_2 FILLER_26_116 ();
 sg13g2_fill_1 FILLER_26_139 ();
 sg13g2_fill_1 FILLER_26_162 ();
 sg13g2_decap_8 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_174 ();
 sg13g2_fill_1 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_195 ();
 sg13g2_decap_4 FILLER_26_201 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_215 ();
 sg13g2_decap_8 FILLER_26_222 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_fill_1 FILLER_26_235 ();
 sg13g2_fill_2 FILLER_26_241 ();
 sg13g2_fill_1 FILLER_26_243 ();
 sg13g2_fill_1 FILLER_26_270 ();
 sg13g2_fill_2 FILLER_26_306 ();
 sg13g2_fill_1 FILLER_26_320 ();
 sg13g2_decap_4 FILLER_26_341 ();
 sg13g2_fill_1 FILLER_26_345 ();
 sg13g2_fill_2 FILLER_26_359 ();
 sg13g2_fill_1 FILLER_26_361 ();
 sg13g2_fill_2 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_fill_2 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_65 ();
 sg13g2_fill_1 FILLER_27_79 ();
 sg13g2_decap_8 FILLER_27_96 ();
 sg13g2_decap_8 FILLER_27_103 ();
 sg13g2_decap_8 FILLER_27_110 ();
 sg13g2_fill_2 FILLER_27_146 ();
 sg13g2_decap_4 FILLER_27_174 ();
 sg13g2_fill_1 FILLER_27_178 ();
 sg13g2_fill_2 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_185 ();
 sg13g2_decap_8 FILLER_27_190 ();
 sg13g2_fill_2 FILLER_27_210 ();
 sg13g2_fill_1 FILLER_27_227 ();
 sg13g2_fill_2 FILLER_27_259 ();
 sg13g2_fill_1 FILLER_27_270 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_4 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_60 ();
 sg13g2_fill_1 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_104 ();
 sg13g2_decap_8 FILLER_28_111 ();
 sg13g2_fill_2 FILLER_28_118 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_fill_2 FILLER_28_161 ();
 sg13g2_fill_2 FILLER_28_177 ();
 sg13g2_fill_1 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_decap_4 FILLER_28_209 ();
 sg13g2_fill_2 FILLER_28_213 ();
 sg13g2_decap_4 FILLER_28_233 ();
 sg13g2_fill_1 FILLER_28_250 ();
 sg13g2_fill_1 FILLER_28_281 ();
 sg13g2_fill_2 FILLER_28_290 ();
 sg13g2_fill_2 FILLER_28_338 ();
 sg13g2_fill_1 FILLER_28_340 ();
 sg13g2_fill_2 FILLER_28_349 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_fill_1 FILLER_29_90 ();
 sg13g2_decap_8 FILLER_29_111 ();
 sg13g2_decap_8 FILLER_29_118 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_142 ();
 sg13g2_fill_1 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_178 ();
 sg13g2_decap_4 FILLER_29_192 ();
 sg13g2_fill_1 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_fill_2 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_271 ();
 sg13g2_fill_2 FILLER_29_296 ();
 sg13g2_fill_2 FILLER_29_335 ();
 sg13g2_fill_1 FILLER_29_337 ();
 sg13g2_decap_4 FILLER_29_345 ();
 sg13g2_fill_2 FILLER_29_349 ();
 sg13g2_fill_2 FILLER_29_354 ();
 sg13g2_fill_1 FILLER_29_356 ();
 sg13g2_decap_4 FILLER_29_362 ();
 sg13g2_fill_2 FILLER_29_366 ();
 sg13g2_decap_8 FILLER_29_373 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_4 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_97 ();
 sg13g2_decap_8 FILLER_30_115 ();
 sg13g2_decap_8 FILLER_30_122 ();
 sg13g2_decap_8 FILLER_30_129 ();
 sg13g2_decap_4 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_140 ();
 sg13g2_decap_4 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_decap_4 FILLER_30_197 ();
 sg13g2_fill_1 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_fill_2 FILLER_30_230 ();
 sg13g2_fill_1 FILLER_30_232 ();
 sg13g2_fill_2 FILLER_30_254 ();
 sg13g2_fill_2 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_289 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_fill_2 FILLER_30_334 ();
 sg13g2_fill_1 FILLER_30_349 ();
 sg13g2_fill_1 FILLER_30_358 ();
 sg13g2_fill_2 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_30_386 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_65 ();
 sg13g2_decap_8 FILLER_31_74 ();
 sg13g2_decap_8 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_fill_1 FILLER_31_107 ();
 sg13g2_decap_8 FILLER_31_134 ();
 sg13g2_decap_4 FILLER_31_141 ();
 sg13g2_fill_2 FILLER_31_145 ();
 sg13g2_decap_4 FILLER_31_151 ();
 sg13g2_decap_8 FILLER_31_179 ();
 sg13g2_fill_1 FILLER_31_186 ();
 sg13g2_decap_4 FILLER_31_200 ();
 sg13g2_fill_1 FILLER_31_217 ();
 sg13g2_fill_1 FILLER_31_226 ();
 sg13g2_fill_2 FILLER_31_237 ();
 sg13g2_fill_1 FILLER_31_239 ();
 sg13g2_fill_2 FILLER_31_248 ();
 sg13g2_fill_1 FILLER_31_250 ();
 sg13g2_fill_2 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_262 ();
 sg13g2_fill_2 FILLER_31_340 ();
 sg13g2_decap_4 FILLER_31_350 ();
 sg13g2_fill_1 FILLER_31_354 ();
 sg13g2_fill_2 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_decap_8 FILLER_31_393 ();
 sg13g2_decap_8 FILLER_31_400 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_56 ();
 sg13g2_fill_2 FILLER_32_81 ();
 sg13g2_decap_4 FILLER_32_88 ();
 sg13g2_fill_2 FILLER_32_141 ();
 sg13g2_decap_8 FILLER_32_148 ();
 sg13g2_fill_2 FILLER_32_155 ();
 sg13g2_fill_1 FILLER_32_185 ();
 sg13g2_fill_1 FILLER_32_198 ();
 sg13g2_fill_1 FILLER_32_203 ();
 sg13g2_fill_2 FILLER_32_308 ();
 sg13g2_fill_1 FILLER_32_325 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_fill_1 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_4 FILLER_33_49 ();
 sg13g2_fill_1 FILLER_33_95 ();
 sg13g2_fill_2 FILLER_33_101 ();
 sg13g2_fill_2 FILLER_33_134 ();
 sg13g2_decap_8 FILLER_33_162 ();
 sg13g2_fill_1 FILLER_33_169 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_4 FILLER_33_189 ();
 sg13g2_fill_1 FILLER_33_193 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_fill_2 FILLER_33_217 ();
 sg13g2_fill_1 FILLER_33_219 ();
 sg13g2_fill_1 FILLER_33_233 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_decap_4 FILLER_33_252 ();
 sg13g2_fill_1 FILLER_33_256 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_315 ();
 sg13g2_decap_4 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_348 ();
 sg13g2_decap_8 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_380 ();
 sg13g2_decap_8 FILLER_33_387 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_56 ();
 sg13g2_fill_2 FILLER_34_60 ();
 sg13g2_fill_2 FILLER_34_71 ();
 sg13g2_decap_4 FILLER_34_76 ();
 sg13g2_fill_1 FILLER_34_80 ();
 sg13g2_decap_8 FILLER_34_90 ();
 sg13g2_fill_1 FILLER_34_97 ();
 sg13g2_decap_8 FILLER_34_107 ();
 sg13g2_decap_8 FILLER_34_114 ();
 sg13g2_fill_1 FILLER_34_131 ();
 sg13g2_fill_2 FILLER_34_160 ();
 sg13g2_decap_4 FILLER_34_172 ();
 sg13g2_decap_8 FILLER_34_180 ();
 sg13g2_fill_2 FILLER_34_187 ();
 sg13g2_decap_4 FILLER_34_205 ();
 sg13g2_fill_2 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_decap_8 FILLER_34_254 ();
 sg13g2_fill_2 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_315 ();
 sg13g2_fill_2 FILLER_34_360 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_decap_8 FILLER_34_375 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_fill_2 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_51 ();
 sg13g2_decap_8 FILLER_35_73 ();
 sg13g2_decap_4 FILLER_35_80 ();
 sg13g2_fill_2 FILLER_35_89 ();
 sg13g2_fill_1 FILLER_35_91 ();
 sg13g2_decap_4 FILLER_35_114 ();
 sg13g2_fill_2 FILLER_35_118 ();
 sg13g2_fill_2 FILLER_35_129 ();
 sg13g2_fill_1 FILLER_35_131 ();
 sg13g2_decap_4 FILLER_35_136 ();
 sg13g2_fill_1 FILLER_35_140 ();
 sg13g2_fill_2 FILLER_35_163 ();
 sg13g2_fill_1 FILLER_35_180 ();
 sg13g2_fill_2 FILLER_35_196 ();
 sg13g2_fill_2 FILLER_35_212 ();
 sg13g2_decap_4 FILLER_35_232 ();
 sg13g2_fill_2 FILLER_35_246 ();
 sg13g2_fill_1 FILLER_35_248 ();
 sg13g2_fill_2 FILLER_35_269 ();
 sg13g2_fill_1 FILLER_35_271 ();
 sg13g2_fill_2 FILLER_35_292 ();
 sg13g2_fill_1 FILLER_35_294 ();
 sg13g2_fill_1 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_383 ();
 sg13g2_decap_8 FILLER_35_390 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_44 ();
 sg13g2_decap_4 FILLER_36_76 ();
 sg13g2_fill_1 FILLER_36_80 ();
 sg13g2_fill_1 FILLER_36_93 ();
 sg13g2_fill_2 FILLER_36_102 ();
 sg13g2_fill_1 FILLER_36_104 ();
 sg13g2_fill_2 FILLER_36_109 ();
 sg13g2_decap_8 FILLER_36_137 ();
 sg13g2_decap_4 FILLER_36_144 ();
 sg13g2_fill_2 FILLER_36_148 ();
 sg13g2_fill_1 FILLER_36_153 ();
 sg13g2_fill_2 FILLER_36_160 ();
 sg13g2_fill_1 FILLER_36_162 ();
 sg13g2_fill_1 FILLER_36_167 ();
 sg13g2_fill_1 FILLER_36_195 ();
 sg13g2_fill_2 FILLER_36_276 ();
 sg13g2_fill_1 FILLER_36_278 ();
 sg13g2_fill_2 FILLER_36_318 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_fill_1 FILLER_36_335 ();
 sg13g2_decap_8 FILLER_36_341 ();
 sg13g2_fill_1 FILLER_36_348 ();
 sg13g2_fill_2 FILLER_36_361 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_fill_2 FILLER_37_64 ();
 sg13g2_fill_2 FILLER_37_107 ();
 sg13g2_fill_1 FILLER_37_109 ();
 sg13g2_fill_2 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_135 ();
 sg13g2_decap_8 FILLER_37_145 ();
 sg13g2_fill_1 FILLER_37_152 ();
 sg13g2_fill_2 FILLER_37_165 ();
 sg13g2_fill_2 FILLER_37_200 ();
 sg13g2_decap_4 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_311 ();
 sg13g2_fill_2 FILLER_37_324 ();
 sg13g2_fill_1 FILLER_37_326 ();
 sg13g2_decap_8 FILLER_37_344 ();
 sg13g2_decap_8 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_4 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_85 ();
 sg13g2_fill_1 FILLER_38_87 ();
 sg13g2_fill_2 FILLER_38_155 ();
 sg13g2_fill_1 FILLER_38_157 ();
 sg13g2_fill_2 FILLER_38_193 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_fill_1 FILLER_38_208 ();
 sg13g2_decap_4 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_226 ();
 sg13g2_fill_2 FILLER_38_297 ();
 sg13g2_fill_1 FILLER_38_304 ();
 sg13g2_fill_2 FILLER_38_330 ();
 sg13g2_fill_1 FILLER_38_332 ();
 sg13g2_fill_2 FILLER_38_346 ();
 sg13g2_fill_1 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_367 ();
 sg13g2_decap_4 FILLER_38_374 ();
 sg13g2_fill_2 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_fill_2 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_73 ();
 sg13g2_decap_8 FILLER_39_80 ();
 sg13g2_fill_2 FILLER_39_87 ();
 sg13g2_decap_4 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_115 ();
 sg13g2_decap_4 FILLER_39_122 ();
 sg13g2_fill_1 FILLER_39_130 ();
 sg13g2_decap_8 FILLER_39_158 ();
 sg13g2_decap_8 FILLER_39_165 ();
 sg13g2_fill_1 FILLER_39_184 ();
 sg13g2_decap_8 FILLER_39_194 ();
 sg13g2_decap_8 FILLER_39_201 ();
 sg13g2_fill_1 FILLER_39_208 ();
 sg13g2_decap_4 FILLER_39_235 ();
 sg13g2_decap_4 FILLER_39_243 ();
 sg13g2_fill_1 FILLER_39_247 ();
 sg13g2_fill_2 FILLER_39_276 ();
 sg13g2_fill_1 FILLER_39_278 ();
 sg13g2_fill_1 FILLER_39_303 ();
 sg13g2_decap_8 FILLER_39_330 ();
 sg13g2_fill_1 FILLER_39_337 ();
 sg13g2_decap_4 FILLER_39_376 ();
 sg13g2_fill_2 FILLER_39_380 ();
 sg13g2_decap_8 FILLER_39_395 ();
 sg13g2_decap_8 FILLER_39_402 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_fill_2 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_66 ();
 sg13g2_decap_8 FILLER_40_73 ();
 sg13g2_decap_4 FILLER_40_80 ();
 sg13g2_fill_1 FILLER_40_84 ();
 sg13g2_fill_2 FILLER_40_89 ();
 sg13g2_decap_8 FILLER_40_100 ();
 sg13g2_decap_4 FILLER_40_107 ();
 sg13g2_fill_2 FILLER_40_111 ();
 sg13g2_decap_4 FILLER_40_117 ();
 sg13g2_fill_1 FILLER_40_124 ();
 sg13g2_decap_4 FILLER_40_133 ();
 sg13g2_fill_1 FILLER_40_137 ();
 sg13g2_decap_4 FILLER_40_150 ();
 sg13g2_fill_2 FILLER_40_168 ();
 sg13g2_fill_2 FILLER_40_185 ();
 sg13g2_fill_1 FILLER_40_187 ();
 sg13g2_decap_8 FILLER_40_195 ();
 sg13g2_decap_8 FILLER_40_202 ();
 sg13g2_fill_2 FILLER_40_209 ();
 sg13g2_fill_1 FILLER_40_211 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_fill_1 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_244 ();
 sg13g2_decap_8 FILLER_40_251 ();
 sg13g2_fill_2 FILLER_40_284 ();
 sg13g2_fill_1 FILLER_40_318 ();
 sg13g2_fill_2 FILLER_40_352 ();
 sg13g2_fill_1 FILLER_40_384 ();
 sg13g2_decap_8 FILLER_40_390 ();
 sg13g2_decap_8 FILLER_40_397 ();
 sg13g2_decap_4 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_fill_2 FILLER_41_56 ();
 sg13g2_fill_1 FILLER_41_58 ();
 sg13g2_decap_4 FILLER_41_70 ();
 sg13g2_fill_2 FILLER_41_74 ();
 sg13g2_fill_1 FILLER_41_107 ();
 sg13g2_decap_4 FILLER_41_140 ();
 sg13g2_fill_1 FILLER_41_144 ();
 sg13g2_decap_4 FILLER_41_149 ();
 sg13g2_fill_1 FILLER_41_153 ();
 sg13g2_fill_2 FILLER_41_175 ();
 sg13g2_fill_2 FILLER_41_182 ();
 sg13g2_fill_2 FILLER_41_189 ();
 sg13g2_fill_1 FILLER_41_191 ();
 sg13g2_fill_2 FILLER_41_197 ();
 sg13g2_fill_2 FILLER_41_208 ();
 sg13g2_fill_1 FILLER_41_214 ();
 sg13g2_fill_2 FILLER_41_244 ();
 sg13g2_fill_2 FILLER_41_311 ();
 sg13g2_fill_2 FILLER_41_325 ();
 sg13g2_decap_4 FILLER_41_335 ();
 sg13g2_fill_1 FILLER_41_339 ();
 sg13g2_decap_4 FILLER_41_350 ();
 sg13g2_fill_2 FILLER_41_354 ();
 sg13g2_fill_2 FILLER_41_364 ();
 sg13g2_fill_1 FILLER_41_366 ();
 sg13g2_decap_8 FILLER_41_395 ();
 sg13g2_decap_8 FILLER_41_402 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_fill_1 FILLER_42_49 ();
 sg13g2_fill_1 FILLER_42_99 ();
 sg13g2_fill_2 FILLER_42_112 ();
 sg13g2_fill_1 FILLER_42_114 ();
 sg13g2_fill_2 FILLER_42_141 ();
 sg13g2_fill_1 FILLER_42_143 ();
 sg13g2_fill_2 FILLER_42_149 ();
 sg13g2_fill_1 FILLER_42_151 ();
 sg13g2_fill_2 FILLER_42_156 ();
 sg13g2_fill_2 FILLER_42_167 ();
 sg13g2_fill_1 FILLER_42_169 ();
 sg13g2_decap_8 FILLER_42_186 ();
 sg13g2_fill_2 FILLER_42_193 ();
 sg13g2_fill_1 FILLER_42_210 ();
 sg13g2_fill_2 FILLER_42_247 ();
 sg13g2_fill_1 FILLER_42_286 ();
 sg13g2_fill_2 FILLER_42_299 ();
 sg13g2_decap_8 FILLER_42_304 ();
 sg13g2_decap_8 FILLER_42_311 ();
 sg13g2_decap_4 FILLER_42_318 ();
 sg13g2_fill_2 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_332 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_fill_2 FILLER_42_371 ();
 sg13g2_fill_1 FILLER_42_373 ();
 sg13g2_decap_8 FILLER_42_390 ();
 sg13g2_decap_8 FILLER_42_397 ();
 sg13g2_decap_4 FILLER_42_404 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_4 FILLER_43_42 ();
 sg13g2_fill_1 FILLER_43_46 ();
 sg13g2_fill_2 FILLER_43_73 ();
 sg13g2_fill_2 FILLER_43_93 ();
 sg13g2_fill_1 FILLER_43_99 ();
 sg13g2_fill_1 FILLER_43_130 ();
 sg13g2_decap_4 FILLER_43_137 ();
 sg13g2_fill_2 FILLER_43_153 ();
 sg13g2_fill_2 FILLER_43_299 ();
 sg13g2_fill_1 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_372 ();
 sg13g2_decap_8 FILLER_43_379 ();
 sg13g2_decap_8 FILLER_43_386 ();
 sg13g2_decap_8 FILLER_43_393 ();
 sg13g2_decap_8 FILLER_43_400 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_66 ();
 sg13g2_decap_8 FILLER_44_73 ();
 sg13g2_decap_8 FILLER_44_80 ();
 sg13g2_fill_1 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_101 ();
 sg13g2_fill_1 FILLER_44_108 ();
 sg13g2_decap_8 FILLER_44_113 ();
 sg13g2_decap_8 FILLER_44_120 ();
 sg13g2_decap_8 FILLER_44_146 ();
 sg13g2_fill_1 FILLER_44_153 ();
 sg13g2_decap_8 FILLER_44_171 ();
 sg13g2_decap_8 FILLER_44_178 ();
 sg13g2_decap_8 FILLER_44_185 ();
 sg13g2_fill_2 FILLER_44_230 ();
 sg13g2_fill_2 FILLER_44_258 ();
 sg13g2_fill_1 FILLER_44_260 ();
 sg13g2_decap_4 FILLER_44_269 ();
 sg13g2_fill_1 FILLER_44_278 ();
 sg13g2_decap_4 FILLER_44_283 ();
 sg13g2_fill_1 FILLER_44_287 ();
 sg13g2_fill_2 FILLER_44_327 ();
 sg13g2_decap_8 FILLER_44_383 ();
 sg13g2_decap_8 FILLER_44_390 ();
 sg13g2_decap_8 FILLER_44_397 ();
 sg13g2_decap_4 FILLER_44_404 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_4 FILLER_45_42 ();
 sg13g2_fill_2 FILLER_45_46 ();
 sg13g2_decap_8 FILLER_45_61 ();
 sg13g2_decap_4 FILLER_45_68 ();
 sg13g2_fill_1 FILLER_45_72 ();
 sg13g2_decap_4 FILLER_45_81 ();
 sg13g2_fill_2 FILLER_45_119 ();
 sg13g2_fill_1 FILLER_45_121 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_fill_2 FILLER_45_153 ();
 sg13g2_decap_8 FILLER_45_174 ();
 sg13g2_decap_8 FILLER_45_181 ();
 sg13g2_decap_4 FILLER_45_188 ();
 sg13g2_fill_2 FILLER_45_192 ();
 sg13g2_fill_2 FILLER_45_220 ();
 sg13g2_fill_1 FILLER_45_222 ();
 sg13g2_fill_2 FILLER_45_271 ();
 sg13g2_fill_1 FILLER_45_273 ();
 sg13g2_fill_2 FILLER_45_300 ();
 sg13g2_fill_2 FILLER_45_347 ();
 sg13g2_decap_8 FILLER_45_394 ();
 sg13g2_decap_8 FILLER_45_401 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_fill_1 FILLER_46_42 ();
 sg13g2_fill_2 FILLER_46_63 ();
 sg13g2_fill_2 FILLER_46_73 ();
 sg13g2_fill_2 FILLER_46_83 ();
 sg13g2_fill_1 FILLER_46_114 ();
 sg13g2_decap_8 FILLER_46_137 ();
 sg13g2_decap_8 FILLER_46_144 ();
 sg13g2_fill_1 FILLER_46_151 ();
 sg13g2_fill_1 FILLER_46_160 ();
 sg13g2_fill_2 FILLER_46_174 ();
 sg13g2_fill_2 FILLER_46_181 ();
 sg13g2_decap_4 FILLER_46_196 ();
 sg13g2_fill_1 FILLER_46_221 ();
 sg13g2_decap_4 FILLER_46_260 ();
 sg13g2_fill_2 FILLER_46_264 ();
 sg13g2_decap_4 FILLER_46_286 ();
 sg13g2_fill_2 FILLER_46_290 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_fill_2 FILLER_46_308 ();
 sg13g2_fill_1 FILLER_46_310 ();
 sg13g2_fill_1 FILLER_46_315 ();
 sg13g2_decap_4 FILLER_46_336 ();
 sg13g2_fill_2 FILLER_46_340 ();
 sg13g2_decap_8 FILLER_46_346 ();
 sg13g2_decap_8 FILLER_46_353 ();
 sg13g2_decap_8 FILLER_46_360 ();
 sg13g2_fill_2 FILLER_46_367 ();
 sg13g2_fill_1 FILLER_46_369 ();
 sg13g2_decap_8 FILLER_46_390 ();
 sg13g2_decap_8 FILLER_46_397 ();
 sg13g2_decap_4 FILLER_46_404 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_fill_2 FILLER_47_54 ();
 sg13g2_fill_1 FILLER_47_56 ();
 sg13g2_fill_2 FILLER_47_82 ();
 sg13g2_fill_1 FILLER_47_84 ();
 sg13g2_fill_1 FILLER_47_90 ();
 sg13g2_fill_1 FILLER_47_120 ();
 sg13g2_fill_2 FILLER_47_130 ();
 sg13g2_fill_1 FILLER_47_132 ();
 sg13g2_fill_2 FILLER_47_141 ();
 sg13g2_fill_2 FILLER_47_160 ();
 sg13g2_fill_1 FILLER_47_162 ();
 sg13g2_decap_4 FILLER_47_190 ();
 sg13g2_fill_2 FILLER_47_194 ();
 sg13g2_decap_8 FILLER_47_200 ();
 sg13g2_decap_8 FILLER_47_207 ();
 sg13g2_fill_1 FILLER_47_214 ();
 sg13g2_decap_8 FILLER_47_227 ();
 sg13g2_decap_8 FILLER_47_239 ();
 sg13g2_fill_1 FILLER_47_246 ();
 sg13g2_fill_2 FILLER_47_252 ();
 sg13g2_fill_1 FILLER_47_254 ();
 sg13g2_fill_1 FILLER_47_291 ();
 sg13g2_fill_2 FILLER_47_312 ();
 sg13g2_fill_1 FILLER_47_314 ();
 sg13g2_decap_4 FILLER_47_319 ();
 sg13g2_fill_2 FILLER_47_323 ();
 sg13g2_fill_2 FILLER_47_350 ();
 sg13g2_fill_1 FILLER_47_352 ();
 sg13g2_fill_2 FILLER_47_366 ();
 sg13g2_decap_4 FILLER_47_372 ();
 sg13g2_fill_1 FILLER_47_376 ();
 sg13g2_fill_2 FILLER_47_382 ();
 sg13g2_decap_8 FILLER_47_396 ();
 sg13g2_decap_4 FILLER_47_403 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_fill_1 FILLER_48_49 ();
 sg13g2_fill_2 FILLER_48_95 ();
 sg13g2_fill_1 FILLER_48_97 ();
 sg13g2_decap_8 FILLER_48_103 ();
 sg13g2_decap_8 FILLER_48_110 ();
 sg13g2_fill_1 FILLER_48_117 ();
 sg13g2_fill_2 FILLER_48_123 ();
 sg13g2_fill_1 FILLER_48_125 ();
 sg13g2_fill_1 FILLER_48_136 ();
 sg13g2_fill_2 FILLER_48_158 ();
 sg13g2_fill_1 FILLER_48_160 ();
 sg13g2_fill_1 FILLER_48_200 ();
 sg13g2_fill_1 FILLER_48_206 ();
 sg13g2_decap_8 FILLER_48_234 ();
 sg13g2_fill_1 FILLER_48_241 ();
 sg13g2_decap_8 FILLER_48_250 ();
 sg13g2_decap_4 FILLER_48_257 ();
 sg13g2_fill_1 FILLER_48_261 ();
 sg13g2_fill_1 FILLER_48_275 ();
 sg13g2_fill_2 FILLER_48_290 ();
 sg13g2_fill_1 FILLER_48_292 ();
 sg13g2_decap_4 FILLER_48_326 ();
 sg13g2_fill_2 FILLER_48_330 ();
 sg13g2_fill_2 FILLER_48_406 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_fill_2 FILLER_49_49 ();
 sg13g2_fill_1 FILLER_49_51 ();
 sg13g2_fill_2 FILLER_49_69 ();
 sg13g2_fill_1 FILLER_49_71 ();
 sg13g2_decap_8 FILLER_49_81 ();
 sg13g2_decap_8 FILLER_49_101 ();
 sg13g2_decap_8 FILLER_49_108 ();
 sg13g2_fill_2 FILLER_49_115 ();
 sg13g2_fill_1 FILLER_49_121 ();
 sg13g2_fill_2 FILLER_49_134 ();
 sg13g2_fill_1 FILLER_49_136 ();
 sg13g2_fill_2 FILLER_49_158 ();
 sg13g2_fill_1 FILLER_49_160 ();
 sg13g2_fill_2 FILLER_49_209 ();
 sg13g2_fill_1 FILLER_49_211 ();
 sg13g2_fill_2 FILLER_49_280 ();
 sg13g2_fill_1 FILLER_49_282 ();
 sg13g2_fill_1 FILLER_49_312 ();
 sg13g2_decap_4 FILLER_49_339 ();
 sg13g2_fill_1 FILLER_49_343 ();
 sg13g2_fill_2 FILLER_49_349 ();
 sg13g2_decap_4 FILLER_49_355 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_fill_2 FILLER_49_375 ();
 sg13g2_decap_8 FILLER_49_401 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_fill_2 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_64 ();
 sg13g2_decap_8 FILLER_50_71 ();
 sg13g2_fill_2 FILLER_50_78 ();
 sg13g2_fill_2 FILLER_50_92 ();
 sg13g2_decap_4 FILLER_50_101 ();
 sg13g2_fill_2 FILLER_50_105 ();
 sg13g2_fill_1 FILLER_50_129 ();
 sg13g2_fill_1 FILLER_50_135 ();
 sg13g2_decap_8 FILLER_50_141 ();
 sg13g2_fill_2 FILLER_50_160 ();
 sg13g2_fill_1 FILLER_50_162 ();
 sg13g2_fill_1 FILLER_50_167 ();
 sg13g2_fill_1 FILLER_50_176 ();
 sg13g2_fill_1 FILLER_50_229 ();
 sg13g2_fill_2 FILLER_50_238 ();
 sg13g2_fill_2 FILLER_50_364 ();
 sg13g2_decap_4 FILLER_50_378 ();
 sg13g2_fill_1 FILLER_50_382 ();
 sg13g2_decap_8 FILLER_50_388 ();
 sg13g2_decap_8 FILLER_50_395 ();
 sg13g2_fill_1 FILLER_50_402 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_4 FILLER_51_42 ();
 sg13g2_fill_2 FILLER_51_46 ();
 sg13g2_decap_8 FILLER_51_60 ();
 sg13g2_fill_1 FILLER_51_80 ();
 sg13g2_fill_2 FILLER_51_86 ();
 sg13g2_fill_2 FILLER_51_109 ();
 sg13g2_fill_1 FILLER_51_111 ();
 sg13g2_fill_2 FILLER_51_133 ();
 sg13g2_decap_4 FILLER_51_147 ();
 sg13g2_fill_2 FILLER_51_151 ();
 sg13g2_fill_2 FILLER_51_158 ();
 sg13g2_decap_8 FILLER_51_164 ();
 sg13g2_fill_2 FILLER_51_197 ();
 sg13g2_fill_1 FILLER_51_199 ();
 sg13g2_fill_2 FILLER_51_213 ();
 sg13g2_fill_1 FILLER_51_215 ();
 sg13g2_fill_2 FILLER_51_259 ();
 sg13g2_decap_8 FILLER_51_313 ();
 sg13g2_decap_8 FILLER_51_320 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_fill_2 FILLER_52_49 ();
 sg13g2_fill_1 FILLER_52_61 ();
 sg13g2_fill_1 FILLER_52_91 ();
 sg13g2_decap_4 FILLER_52_95 ();
 sg13g2_fill_1 FILLER_52_99 ();
 sg13g2_decap_4 FILLER_52_105 ();
 sg13g2_fill_1 FILLER_52_109 ();
 sg13g2_decap_8 FILLER_52_127 ();
 sg13g2_fill_1 FILLER_52_134 ();
 sg13g2_fill_2 FILLER_52_144 ();
 sg13g2_fill_1 FILLER_52_146 ();
 sg13g2_decap_4 FILLER_52_171 ();
 sg13g2_decap_8 FILLER_52_182 ();
 sg13g2_decap_4 FILLER_52_189 ();
 sg13g2_decap_8 FILLER_52_203 ();
 sg13g2_fill_2 FILLER_52_222 ();
 sg13g2_fill_2 FILLER_52_247 ();
 sg13g2_fill_1 FILLER_52_249 ();
 sg13g2_decap_8 FILLER_52_272 ();
 sg13g2_decap_8 FILLER_52_279 ();
 sg13g2_decap_4 FILLER_52_286 ();
 sg13g2_fill_2 FILLER_52_290 ();
 sg13g2_fill_2 FILLER_52_305 ();
 sg13g2_fill_1 FILLER_52_307 ();
 sg13g2_fill_2 FILLER_52_330 ();
 sg13g2_fill_1 FILLER_52_332 ();
 sg13g2_decap_4 FILLER_52_338 ();
 sg13g2_fill_2 FILLER_52_366 ();
 sg13g2_fill_1 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_4 FILLER_53_35 ();
 sg13g2_fill_1 FILLER_53_39 ();
 sg13g2_fill_2 FILLER_53_64 ();
 sg13g2_fill_1 FILLER_53_66 ();
 sg13g2_fill_2 FILLER_53_84 ();
 sg13g2_fill_1 FILLER_53_86 ();
 sg13g2_decap_4 FILLER_53_92 ();
 sg13g2_fill_1 FILLER_53_96 ();
 sg13g2_fill_1 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_122 ();
 sg13g2_decap_4 FILLER_53_129 ();
 sg13g2_fill_1 FILLER_53_133 ();
 sg13g2_fill_2 FILLER_53_156 ();
 sg13g2_fill_1 FILLER_53_158 ();
 sg13g2_decap_4 FILLER_53_167 ();
 sg13g2_decap_8 FILLER_53_207 ();
 sg13g2_fill_1 FILLER_53_214 ();
 sg13g2_fill_2 FILLER_53_277 ();
 sg13g2_fill_1 FILLER_53_279 ();
 sg13g2_decap_4 FILLER_53_284 ();
 sg13g2_decap_4 FILLER_53_293 ();
 sg13g2_fill_2 FILLER_53_297 ();
 sg13g2_fill_1 FILLER_53_303 ();
 sg13g2_decap_4 FILLER_53_313 ();
 sg13g2_decap_8 FILLER_53_325 ();
 sg13g2_decap_8 FILLER_53_332 ();
 sg13g2_fill_1 FILLER_53_339 ();
 sg13g2_decap_8 FILLER_53_349 ();
 sg13g2_decap_8 FILLER_53_356 ();
 sg13g2_decap_8 FILLER_53_363 ();
 sg13g2_decap_8 FILLER_53_370 ();
 sg13g2_decap_4 FILLER_53_405 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_4 FILLER_54_42 ();
 sg13g2_fill_1 FILLER_54_57 ();
 sg13g2_fill_1 FILLER_54_68 ();
 sg13g2_fill_2 FILLER_54_79 ();
 sg13g2_fill_1 FILLER_54_81 ();
 sg13g2_decap_8 FILLER_54_115 ();
 sg13g2_fill_1 FILLER_54_122 ();
 sg13g2_decap_8 FILLER_54_144 ();
 sg13g2_decap_8 FILLER_54_151 ();
 sg13g2_fill_1 FILLER_54_173 ();
 sg13g2_decap_8 FILLER_54_273 ();
 sg13g2_decap_8 FILLER_54_280 ();
 sg13g2_fill_1 FILLER_54_287 ();
 sg13g2_fill_1 FILLER_54_360 ();
 sg13g2_decap_8 FILLER_54_366 ();
 sg13g2_fill_1 FILLER_54_373 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_fill_2 FILLER_55_64 ();
 sg13g2_fill_2 FILLER_55_71 ();
 sg13g2_fill_1 FILLER_55_73 ();
 sg13g2_fill_2 FILLER_55_87 ();
 sg13g2_fill_1 FILLER_55_89 ();
 sg13g2_fill_2 FILLER_55_98 ();
 sg13g2_fill_1 FILLER_55_100 ();
 sg13g2_decap_4 FILLER_55_109 ();
 sg13g2_fill_2 FILLER_55_113 ();
 sg13g2_fill_1 FILLER_55_140 ();
 sg13g2_fill_2 FILLER_55_146 ();
 sg13g2_fill_2 FILLER_55_168 ();
 sg13g2_fill_1 FILLER_55_170 ();
 sg13g2_fill_2 FILLER_55_179 ();
 sg13g2_fill_2 FILLER_55_195 ();
 sg13g2_fill_1 FILLER_55_197 ();
 sg13g2_decap_4 FILLER_55_250 ();
 sg13g2_fill_2 FILLER_55_254 ();
 sg13g2_decap_8 FILLER_55_375 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_fill_1 FILLER_56_49 ();
 sg13g2_decap_4 FILLER_56_58 ();
 sg13g2_fill_1 FILLER_56_62 ();
 sg13g2_decap_8 FILLER_56_76 ();
 sg13g2_decap_4 FILLER_56_88 ();
 sg13g2_fill_2 FILLER_56_92 ();
 sg13g2_fill_2 FILLER_56_112 ();
 sg13g2_fill_1 FILLER_56_131 ();
 sg13g2_fill_1 FILLER_56_148 ();
 sg13g2_fill_2 FILLER_56_179 ();
 sg13g2_fill_1 FILLER_56_181 ();
 sg13g2_fill_2 FILLER_56_190 ();
 sg13g2_decap_4 FILLER_56_196 ();
 sg13g2_fill_1 FILLER_56_200 ();
 sg13g2_fill_1 FILLER_56_252 ();
 sg13g2_fill_2 FILLER_56_293 ();
 sg13g2_fill_1 FILLER_56_295 ();
 sg13g2_fill_2 FILLER_56_310 ();
 sg13g2_fill_1 FILLER_56_312 ();
 sg13g2_fill_2 FILLER_56_330 ();
 sg13g2_fill_2 FILLER_56_350 ();
 sg13g2_fill_1 FILLER_56_357 ();
 sg13g2_fill_1 FILLER_56_364 ();
 sg13g2_decap_4 FILLER_56_383 ();
 sg13g2_fill_2 FILLER_56_387 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_4 FILLER_57_70 ();
 sg13g2_fill_1 FILLER_57_74 ();
 sg13g2_fill_1 FILLER_57_90 ();
 sg13g2_fill_1 FILLER_57_103 ();
 sg13g2_decap_4 FILLER_57_112 ();
 sg13g2_fill_2 FILLER_57_116 ();
 sg13g2_fill_2 FILLER_57_130 ();
 sg13g2_fill_2 FILLER_57_151 ();
 sg13g2_fill_1 FILLER_57_153 ();
 sg13g2_decap_8 FILLER_57_167 ();
 sg13g2_decap_8 FILLER_57_183 ();
 sg13g2_decap_8 FILLER_57_190 ();
 sg13g2_decap_8 FILLER_57_197 ();
 sg13g2_decap_8 FILLER_57_204 ();
 sg13g2_decap_8 FILLER_57_211 ();
 sg13g2_decap_8 FILLER_57_218 ();
 sg13g2_decap_8 FILLER_57_225 ();
 sg13g2_decap_8 FILLER_57_232 ();
 sg13g2_decap_8 FILLER_57_239 ();
 sg13g2_decap_4 FILLER_57_246 ();
 sg13g2_fill_2 FILLER_57_273 ();
 sg13g2_fill_1 FILLER_57_275 ();
 sg13g2_fill_2 FILLER_57_288 ();
 sg13g2_fill_2 FILLER_57_295 ();
 sg13g2_decap_4 FILLER_57_308 ();
 sg13g2_decap_8 FILLER_57_332 ();
 sg13g2_decap_8 FILLER_57_339 ();
 sg13g2_decap_4 FILLER_57_346 ();
 sg13g2_fill_1 FILLER_57_350 ();
 sg13g2_decap_8 FILLER_57_401 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_4 FILLER_58_42 ();
 sg13g2_decap_4 FILLER_58_75 ();
 sg13g2_fill_2 FILLER_58_90 ();
 sg13g2_fill_1 FILLER_58_92 ();
 sg13g2_decap_4 FILLER_58_98 ();
 sg13g2_decap_4 FILLER_58_107 ();
 sg13g2_fill_2 FILLER_58_111 ();
 sg13g2_decap_8 FILLER_58_117 ();
 sg13g2_fill_2 FILLER_58_124 ();
 sg13g2_decap_8 FILLER_58_129 ();
 sg13g2_decap_8 FILLER_58_136 ();
 sg13g2_decap_8 FILLER_58_143 ();
 sg13g2_decap_8 FILLER_58_150 ();
 sg13g2_fill_2 FILLER_58_157 ();
 sg13g2_fill_2 FILLER_58_169 ();
 sg13g2_decap_4 FILLER_58_188 ();
 sg13g2_decap_8 FILLER_58_197 ();
 sg13g2_fill_2 FILLER_58_204 ();
 sg13g2_fill_2 FILLER_58_211 ();
 sg13g2_fill_1 FILLER_58_213 ();
 sg13g2_decap_8 FILLER_58_231 ();
 sg13g2_fill_2 FILLER_58_238 ();
 sg13g2_decap_4 FILLER_58_276 ();
 sg13g2_fill_1 FILLER_58_280 ();
 sg13g2_fill_2 FILLER_58_303 ();
 sg13g2_fill_1 FILLER_58_305 ();
 sg13g2_fill_2 FILLER_58_311 ();
 sg13g2_fill_1 FILLER_58_313 ();
 sg13g2_fill_2 FILLER_58_333 ();
 sg13g2_decap_8 FILLER_58_354 ();
 sg13g2_decap_8 FILLER_58_374 ();
 sg13g2_decap_8 FILLER_58_381 ();
 sg13g2_fill_2 FILLER_58_388 ();
 sg13g2_fill_1 FILLER_58_390 ();
 sg13g2_decap_4 FILLER_58_403 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_4 FILLER_59_56 ();
 sg13g2_fill_1 FILLER_59_60 ();
 sg13g2_fill_2 FILLER_59_82 ();
 sg13g2_decap_4 FILLER_59_99 ();
 sg13g2_fill_2 FILLER_59_128 ();
 sg13g2_fill_2 FILLER_59_152 ();
 sg13g2_fill_1 FILLER_59_154 ();
 sg13g2_fill_2 FILLER_59_167 ();
 sg13g2_fill_1 FILLER_59_169 ();
 sg13g2_fill_2 FILLER_59_178 ();
 sg13g2_decap_4 FILLER_59_260 ();
 sg13g2_fill_1 FILLER_59_264 ();
 sg13g2_fill_1 FILLER_59_304 ();
 sg13g2_decap_8 FILLER_59_313 ();
 sg13g2_decap_4 FILLER_59_320 ();
 sg13g2_fill_1 FILLER_59_324 ();
 sg13g2_decap_8 FILLER_59_333 ();
 sg13g2_decap_8 FILLER_59_381 ();
 sg13g2_fill_2 FILLER_59_388 ();
 sg13g2_fill_1 FILLER_59_390 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_fill_1 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_75 ();
 sg13g2_decap_4 FILLER_60_82 ();
 sg13g2_fill_1 FILLER_60_86 ();
 sg13g2_decap_8 FILLER_60_95 ();
 sg13g2_decap_8 FILLER_60_102 ();
 sg13g2_fill_1 FILLER_60_109 ();
 sg13g2_decap_4 FILLER_60_151 ();
 sg13g2_fill_1 FILLER_60_155 ();
 sg13g2_fill_2 FILLER_60_181 ();
 sg13g2_decap_4 FILLER_60_188 ();
 sg13g2_fill_1 FILLER_60_192 ();
 sg13g2_fill_1 FILLER_60_197 ();
 sg13g2_fill_2 FILLER_60_220 ();
 sg13g2_fill_1 FILLER_60_222 ();
 sg13g2_fill_2 FILLER_60_234 ();
 sg13g2_decap_8 FILLER_60_318 ();
 sg13g2_fill_1 FILLER_60_325 ();
 sg13g2_decap_8 FILLER_60_331 ();
 sg13g2_decap_8 FILLER_60_346 ();
 sg13g2_decap_8 FILLER_60_353 ();
 sg13g2_decap_4 FILLER_60_377 ();
 sg13g2_fill_2 FILLER_60_381 ();
 sg13g2_fill_2 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_fill_2 FILLER_61_58 ();
 sg13g2_decap_8 FILLER_61_86 ();
 sg13g2_fill_2 FILLER_61_93 ();
 sg13g2_fill_1 FILLER_61_110 ();
 sg13g2_fill_2 FILLER_61_126 ();
 sg13g2_fill_1 FILLER_61_140 ();
 sg13g2_fill_2 FILLER_61_145 ();
 sg13g2_fill_1 FILLER_61_147 ();
 sg13g2_decap_8 FILLER_61_180 ();
 sg13g2_fill_2 FILLER_61_187 ();
 sg13g2_fill_2 FILLER_61_199 ();
 sg13g2_fill_1 FILLER_61_201 ();
 sg13g2_decap_8 FILLER_61_207 ();
 sg13g2_decap_4 FILLER_61_214 ();
 sg13g2_fill_1 FILLER_61_218 ();
 sg13g2_decap_8 FILLER_61_226 ();
 sg13g2_decap_8 FILLER_61_233 ();
 sg13g2_decap_4 FILLER_61_240 ();
 sg13g2_fill_2 FILLER_61_253 ();
 sg13g2_fill_2 FILLER_61_263 ();
 sg13g2_fill_1 FILLER_61_265 ();
 sg13g2_decap_4 FILLER_61_276 ();
 sg13g2_fill_2 FILLER_61_301 ();
 sg13g2_decap_4 FILLER_61_347 ();
 sg13g2_fill_2 FILLER_61_359 ();
 sg13g2_fill_1 FILLER_61_369 ();
 sg13g2_fill_2 FILLER_61_383 ();
 sg13g2_fill_1 FILLER_61_385 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_4 FILLER_62_35 ();
 sg13g2_fill_2 FILLER_62_39 ();
 sg13g2_fill_2 FILLER_62_74 ();
 sg13g2_decap_8 FILLER_62_81 ();
 sg13g2_decap_4 FILLER_62_88 ();
 sg13g2_decap_4 FILLER_62_100 ();
 sg13g2_fill_2 FILLER_62_104 ();
 sg13g2_decap_8 FILLER_62_115 ();
 sg13g2_decap_8 FILLER_62_122 ();
 sg13g2_decap_8 FILLER_62_129 ();
 sg13g2_decap_8 FILLER_62_136 ();
 sg13g2_fill_2 FILLER_62_143 ();
 sg13g2_fill_1 FILLER_62_165 ();
 sg13g2_fill_2 FILLER_62_179 ();
 sg13g2_fill_2 FILLER_62_194 ();
 sg13g2_fill_1 FILLER_62_196 ();
 sg13g2_decap_4 FILLER_62_211 ();
 sg13g2_decap_4 FILLER_62_237 ();
 sg13g2_fill_2 FILLER_62_250 ();
 sg13g2_fill_1 FILLER_62_252 ();
 sg13g2_fill_2 FILLER_62_307 ();
 sg13g2_fill_2 FILLER_62_321 ();
 sg13g2_fill_1 FILLER_62_339 ();
 sg13g2_fill_1 FILLER_62_368 ();
 sg13g2_fill_1 FILLER_62_377 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_85 ();
 sg13g2_decap_4 FILLER_63_92 ();
 sg13g2_fill_1 FILLER_63_122 ();
 sg13g2_decap_4 FILLER_63_127 ();
 sg13g2_fill_1 FILLER_63_131 ();
 sg13g2_fill_2 FILLER_63_144 ();
 sg13g2_fill_1 FILLER_63_146 ();
 sg13g2_decap_8 FILLER_63_155 ();
 sg13g2_decap_8 FILLER_63_162 ();
 sg13g2_fill_1 FILLER_63_169 ();
 sg13g2_fill_1 FILLER_63_182 ();
 sg13g2_fill_2 FILLER_63_191 ();
 sg13g2_fill_1 FILLER_63_193 ();
 sg13g2_fill_1 FILLER_63_225 ();
 sg13g2_fill_2 FILLER_63_234 ();
 sg13g2_fill_1 FILLER_63_236 ();
 sg13g2_fill_1 FILLER_63_282 ();
 sg13g2_fill_2 FILLER_63_303 ();
 sg13g2_fill_2 FILLER_63_309 ();
 sg13g2_decap_4 FILLER_63_328 ();
 sg13g2_fill_2 FILLER_63_336 ();
 sg13g2_decap_4 FILLER_63_342 ();
 sg13g2_decap_4 FILLER_63_361 ();
 sg13g2_fill_2 FILLER_63_374 ();
 sg13g2_fill_1 FILLER_63_376 ();
 sg13g2_fill_1 FILLER_63_385 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_fill_2 FILLER_64_49 ();
 sg13g2_fill_1 FILLER_64_51 ();
 sg13g2_fill_2 FILLER_64_78 ();
 sg13g2_fill_1 FILLER_64_80 ();
 sg13g2_decap_4 FILLER_64_104 ();
 sg13g2_fill_2 FILLER_64_120 ();
 sg13g2_fill_1 FILLER_64_122 ();
 sg13g2_fill_2 FILLER_64_135 ();
 sg13g2_fill_1 FILLER_64_137 ();
 sg13g2_decap_4 FILLER_64_143 ();
 sg13g2_decap_8 FILLER_64_160 ();
 sg13g2_decap_4 FILLER_64_167 ();
 sg13g2_fill_2 FILLER_64_171 ();
 sg13g2_fill_1 FILLER_64_213 ();
 sg13g2_decap_4 FILLER_64_266 ();
 sg13g2_fill_2 FILLER_64_280 ();
 sg13g2_fill_1 FILLER_64_357 ();
 sg13g2_fill_2 FILLER_64_374 ();
 sg13g2_fill_1 FILLER_64_376 ();
 sg13g2_decap_4 FILLER_64_388 ();
 sg13g2_fill_2 FILLER_64_406 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_fill_2 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_74 ();
 sg13g2_fill_2 FILLER_65_81 ();
 sg13g2_decap_8 FILLER_65_87 ();
 sg13g2_fill_1 FILLER_65_94 ();
 sg13g2_fill_2 FILLER_65_100 ();
 sg13g2_fill_1 FILLER_65_102 ();
 sg13g2_fill_2 FILLER_65_115 ();
 sg13g2_fill_2 FILLER_65_135 ();
 sg13g2_decap_8 FILLER_65_171 ();
 sg13g2_fill_2 FILLER_65_178 ();
 sg13g2_fill_1 FILLER_65_185 ();
 sg13g2_decap_4 FILLER_65_210 ();
 sg13g2_fill_1 FILLER_65_214 ();
 sg13g2_decap_4 FILLER_65_244 ();
 sg13g2_fill_2 FILLER_65_248 ();
 sg13g2_decap_8 FILLER_65_300 ();
 sg13g2_decap_4 FILLER_65_307 ();
 sg13g2_fill_2 FILLER_65_311 ();
 sg13g2_fill_2 FILLER_65_333 ();
 sg13g2_fill_1 FILLER_65_335 ();
 sg13g2_decap_8 FILLER_65_340 ();
 sg13g2_fill_1 FILLER_65_347 ();
 sg13g2_decap_8 FILLER_65_361 ();
 sg13g2_decap_8 FILLER_65_368 ();
 sg13g2_decap_8 FILLER_65_375 ();
 sg13g2_fill_2 FILLER_65_382 ();
 sg13g2_fill_1 FILLER_65_399 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_4 FILLER_66_49 ();
 sg13g2_fill_2 FILLER_66_53 ();
 sg13g2_fill_1 FILLER_66_74 ();
 sg13g2_decap_8 FILLER_66_80 ();
 sg13g2_fill_1 FILLER_66_111 ();
 sg13g2_fill_2 FILLER_66_168 ();
 sg13g2_decap_4 FILLER_66_175 ();
 sg13g2_fill_2 FILLER_66_179 ();
 sg13g2_fill_2 FILLER_66_186 ();
 sg13g2_decap_8 FILLER_66_196 ();
 sg13g2_decap_8 FILLER_66_203 ();
 sg13g2_decap_8 FILLER_66_210 ();
 sg13g2_decap_8 FILLER_66_217 ();
 sg13g2_decap_4 FILLER_66_224 ();
 sg13g2_fill_1 FILLER_66_228 ();
 sg13g2_fill_2 FILLER_66_264 ();
 sg13g2_fill_1 FILLER_66_266 ();
 sg13g2_decap_8 FILLER_66_287 ();
 sg13g2_decap_8 FILLER_66_294 ();
 sg13g2_fill_1 FILLER_66_301 ();
 sg13g2_decap_8 FILLER_66_306 ();
 sg13g2_fill_1 FILLER_66_313 ();
 sg13g2_fill_2 FILLER_66_336 ();
 sg13g2_fill_2 FILLER_66_348 ();
 sg13g2_fill_1 FILLER_66_350 ();
 sg13g2_fill_2 FILLER_66_359 ();
 sg13g2_decap_8 FILLER_66_379 ();
 sg13g2_fill_2 FILLER_66_395 ();
 sg13g2_fill_1 FILLER_66_397 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_4 FILLER_67_49 ();
 sg13g2_fill_1 FILLER_67_53 ();
 sg13g2_decap_4 FILLER_67_92 ();
 sg13g2_fill_1 FILLER_67_96 ();
 sg13g2_decap_8 FILLER_67_116 ();
 sg13g2_decap_4 FILLER_67_123 ();
 sg13g2_fill_2 FILLER_67_127 ();
 sg13g2_fill_1 FILLER_67_133 ();
 sg13g2_decap_4 FILLER_67_138 ();
 sg13g2_decap_4 FILLER_67_146 ();
 sg13g2_fill_1 FILLER_67_150 ();
 sg13g2_fill_2 FILLER_67_155 ();
 sg13g2_fill_1 FILLER_67_157 ();
 sg13g2_decap_4 FILLER_67_163 ();
 sg13g2_fill_1 FILLER_67_167 ();
 sg13g2_decap_4 FILLER_67_176 ();
 sg13g2_fill_2 FILLER_67_188 ();
 sg13g2_fill_1 FILLER_67_195 ();
 sg13g2_decap_8 FILLER_67_208 ();
 sg13g2_fill_2 FILLER_67_215 ();
 sg13g2_fill_1 FILLER_67_217 ();
 sg13g2_fill_2 FILLER_67_238 ();
 sg13g2_fill_1 FILLER_67_295 ();
 sg13g2_fill_1 FILLER_67_328 ();
 sg13g2_fill_2 FILLER_67_344 ();
 sg13g2_fill_2 FILLER_67_361 ();
 sg13g2_fill_1 FILLER_67_363 ();
 sg13g2_fill_2 FILLER_67_380 ();
 sg13g2_fill_1 FILLER_67_402 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_fill_2 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_100 ();
 sg13g2_fill_2 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_130 ();
 sg13g2_fill_1 FILLER_68_137 ();
 sg13g2_decap_4 FILLER_68_142 ();
 sg13g2_fill_1 FILLER_68_146 ();
 sg13g2_fill_2 FILLER_68_152 ();
 sg13g2_fill_1 FILLER_68_154 ();
 sg13g2_decap_4 FILLER_68_164 ();
 sg13g2_fill_2 FILLER_68_168 ();
 sg13g2_fill_2 FILLER_68_200 ();
 sg13g2_fill_1 FILLER_68_202 ();
 sg13g2_fill_1 FILLER_68_212 ();
 sg13g2_decap_8 FILLER_68_314 ();
 sg13g2_fill_2 FILLER_68_321 ();
 sg13g2_fill_1 FILLER_68_323 ();
 sg13g2_fill_2 FILLER_68_336 ();
 sg13g2_decap_4 FILLER_68_342 ();
 sg13g2_fill_2 FILLER_68_346 ();
 sg13g2_decap_4 FILLER_68_356 ();
 sg13g2_fill_1 FILLER_68_360 ();
 sg13g2_fill_2 FILLER_68_366 ();
 sg13g2_decap_8 FILLER_68_378 ();
 sg13g2_fill_1 FILLER_68_394 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_fill_2 FILLER_69_56 ();
 sg13g2_fill_1 FILLER_69_58 ();
 sg13g2_fill_2 FILLER_69_64 ();
 sg13g2_fill_1 FILLER_69_97 ();
 sg13g2_decap_4 FILLER_69_101 ();
 sg13g2_fill_1 FILLER_69_110 ();
 sg13g2_fill_2 FILLER_69_126 ();
 sg13g2_fill_2 FILLER_69_133 ();
 sg13g2_fill_2 FILLER_69_147 ();
 sg13g2_decap_8 FILLER_69_161 ();
 sg13g2_fill_2 FILLER_69_168 ();
 sg13g2_fill_1 FILLER_69_170 ();
 sg13g2_fill_2 FILLER_69_184 ();
 sg13g2_fill_1 FILLER_69_186 ();
 sg13g2_decap_4 FILLER_69_211 ();
 sg13g2_fill_1 FILLER_69_215 ();
 sg13g2_fill_2 FILLER_69_221 ();
 sg13g2_decap_4 FILLER_69_295 ();
 sg13g2_fill_2 FILLER_69_299 ();
 sg13g2_fill_2 FILLER_69_345 ();
 sg13g2_fill_1 FILLER_69_347 ();
 sg13g2_fill_2 FILLER_69_352 ();
 sg13g2_fill_1 FILLER_69_362 ();
 sg13g2_fill_2 FILLER_69_379 ();
 sg13g2_fill_1 FILLER_69_391 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_fill_2 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_71 ();
 sg13g2_decap_8 FILLER_70_78 ();
 sg13g2_fill_2 FILLER_70_85 ();
 sg13g2_fill_1 FILLER_70_87 ();
 sg13g2_fill_2 FILLER_70_92 ();
 sg13g2_fill_1 FILLER_70_99 ();
 sg13g2_fill_1 FILLER_70_104 ();
 sg13g2_fill_2 FILLER_70_139 ();
 sg13g2_fill_2 FILLER_70_144 ();
 sg13g2_decap_8 FILLER_70_170 ();
 sg13g2_fill_1 FILLER_70_177 ();
 sg13g2_decap_4 FILLER_70_190 ();
 sg13g2_fill_2 FILLER_70_199 ();
 sg13g2_fill_1 FILLER_70_201 ();
 sg13g2_fill_2 FILLER_70_225 ();
 sg13g2_fill_1 FILLER_70_227 ();
 sg13g2_fill_1 FILLER_70_280 ();
 sg13g2_decap_4 FILLER_70_320 ();
 sg13g2_fill_1 FILLER_70_324 ();
 sg13g2_fill_2 FILLER_70_333 ();
 sg13g2_fill_1 FILLER_70_335 ();
 sg13g2_fill_2 FILLER_70_343 ();
 sg13g2_fill_1 FILLER_70_345 ();
 sg13g2_fill_2 FILLER_70_358 ();
 sg13g2_decap_8 FILLER_70_372 ();
 sg13g2_decap_4 FILLER_70_379 ();
 sg13g2_fill_1 FILLER_70_383 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_fill_1 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_75 ();
 sg13g2_decap_8 FILLER_71_82 ();
 sg13g2_decap_4 FILLER_71_89 ();
 sg13g2_fill_1 FILLER_71_93 ();
 sg13g2_decap_4 FILLER_71_98 ();
 sg13g2_fill_2 FILLER_71_102 ();
 sg13g2_decap_8 FILLER_71_122 ();
 sg13g2_decap_8 FILLER_71_129 ();
 sg13g2_fill_1 FILLER_71_136 ();
 sg13g2_decap_4 FILLER_71_142 ();
 sg13g2_fill_1 FILLER_71_146 ();
 sg13g2_decap_8 FILLER_71_160 ();
 sg13g2_fill_2 FILLER_71_167 ();
 sg13g2_fill_1 FILLER_71_169 ();
 sg13g2_fill_1 FILLER_71_191 ();
 sg13g2_decap_4 FILLER_71_200 ();
 sg13g2_fill_1 FILLER_71_209 ();
 sg13g2_fill_2 FILLER_71_215 ();
 sg13g2_fill_1 FILLER_71_217 ();
 sg13g2_fill_2 FILLER_71_291 ();
 sg13g2_fill_1 FILLER_71_307 ();
 sg13g2_decap_8 FILLER_71_321 ();
 sg13g2_decap_8 FILLER_71_328 ();
 sg13g2_fill_2 FILLER_71_335 ();
 sg13g2_decap_8 FILLER_71_342 ();
 sg13g2_decap_8 FILLER_71_349 ();
 sg13g2_decap_8 FILLER_71_356 ();
 sg13g2_fill_1 FILLER_71_380 ();
 sg13g2_fill_2 FILLER_71_384 ();
 sg13g2_fill_1 FILLER_71_386 ();
 sg13g2_fill_2 FILLER_71_392 ();
 sg13g2_fill_1 FILLER_71_394 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_fill_1 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_fill_1 FILLER_72_126 ();
 sg13g2_fill_1 FILLER_72_132 ();
 sg13g2_fill_2 FILLER_72_142 ();
 sg13g2_decap_8 FILLER_72_148 ();
 sg13g2_decap_4 FILLER_72_155 ();
 sg13g2_fill_1 FILLER_72_174 ();
 sg13g2_fill_2 FILLER_72_191 ();
 sg13g2_fill_1 FILLER_72_193 ();
 sg13g2_decap_4 FILLER_72_199 ();
 sg13g2_fill_1 FILLER_72_210 ();
 sg13g2_fill_2 FILLER_72_231 ();
 sg13g2_fill_1 FILLER_72_233 ();
 sg13g2_fill_2 FILLER_72_266 ();
 sg13g2_fill_1 FILLER_72_268 ();
 sg13g2_fill_1 FILLER_72_279 ();
 sg13g2_fill_2 FILLER_72_306 ();
 sg13g2_fill_1 FILLER_72_308 ();
 sg13g2_decap_4 FILLER_72_329 ();
 sg13g2_fill_2 FILLER_72_341 ();
 sg13g2_decap_4 FILLER_72_354 ();
 sg13g2_fill_1 FILLER_72_358 ();
 sg13g2_fill_2 FILLER_72_367 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_114 ();
 sg13g2_fill_2 FILLER_73_121 ();
 sg13g2_fill_2 FILLER_73_131 ();
 sg13g2_decap_8 FILLER_73_156 ();
 sg13g2_decap_4 FILLER_73_163 ();
 sg13g2_fill_2 FILLER_73_167 ();
 sg13g2_fill_1 FILLER_73_177 ();
 sg13g2_decap_4 FILLER_73_183 ();
 sg13g2_fill_1 FILLER_73_187 ();
 sg13g2_fill_2 FILLER_73_228 ();
 sg13g2_fill_1 FILLER_73_230 ();
 sg13g2_fill_2 FILLER_73_246 ();
 sg13g2_fill_1 FILLER_73_248 ();
 sg13g2_fill_2 FILLER_73_330 ();
 sg13g2_fill_2 FILLER_73_345 ();
 sg13g2_fill_1 FILLER_73_347 ();
 sg13g2_fill_2 FILLER_73_356 ();
 sg13g2_fill_1 FILLER_73_358 ();
 sg13g2_fill_2 FILLER_73_367 ();
 sg13g2_fill_1 FILLER_73_369 ();
 sg13g2_fill_2 FILLER_73_406 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_4 FILLER_74_56 ();
 sg13g2_fill_1 FILLER_74_60 ();
 sg13g2_fill_1 FILLER_74_95 ();
 sg13g2_fill_1 FILLER_74_104 ();
 sg13g2_fill_2 FILLER_74_145 ();
 sg13g2_fill_2 FILLER_74_153 ();
 sg13g2_decap_8 FILLER_74_170 ();
 sg13g2_fill_1 FILLER_74_177 ();
 sg13g2_fill_2 FILLER_74_190 ();
 sg13g2_fill_1 FILLER_74_192 ();
 sg13g2_decap_4 FILLER_74_211 ();
 sg13g2_fill_2 FILLER_74_215 ();
 sg13g2_decap_8 FILLER_74_221 ();
 sg13g2_fill_2 FILLER_74_228 ();
 sg13g2_fill_1 FILLER_74_240 ();
 sg13g2_fill_2 FILLER_74_267 ();
 sg13g2_fill_1 FILLER_74_269 ();
 sg13g2_fill_2 FILLER_74_279 ();
 sg13g2_fill_2 FILLER_74_353 ();
 sg13g2_decap_8 FILLER_74_367 ();
 sg13g2_fill_1 FILLER_74_377 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_fill_1 FILLER_75_82 ();
 sg13g2_fill_2 FILLER_75_89 ();
 sg13g2_fill_1 FILLER_75_91 ();
 sg13g2_fill_2 FILLER_75_137 ();
 sg13g2_decap_8 FILLER_75_179 ();
 sg13g2_decap_4 FILLER_75_186 ();
 sg13g2_fill_1 FILLER_75_190 ();
 sg13g2_fill_1 FILLER_75_199 ();
 sg13g2_fill_2 FILLER_75_216 ();
 sg13g2_fill_2 FILLER_75_226 ();
 sg13g2_fill_2 FILLER_75_246 ();
 sg13g2_fill_1 FILLER_75_248 ();
 sg13g2_fill_2 FILLER_75_305 ();
 sg13g2_fill_1 FILLER_75_307 ();
 sg13g2_fill_1 FILLER_75_318 ();
 sg13g2_fill_2 FILLER_75_339 ();
 sg13g2_fill_1 FILLER_75_341 ();
 sg13g2_fill_2 FILLER_75_363 ();
 sg13g2_fill_1 FILLER_75_370 ();
 sg13g2_fill_2 FILLER_75_388 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_4 FILLER_76_77 ();
 sg13g2_fill_1 FILLER_76_95 ();
 sg13g2_fill_1 FILLER_76_101 ();
 sg13g2_fill_1 FILLER_76_128 ();
 sg13g2_fill_1 FILLER_76_201 ();
 sg13g2_fill_2 FILLER_76_226 ();
 sg13g2_fill_2 FILLER_76_263 ();
 sg13g2_fill_2 FILLER_76_343 ();
 sg13g2_fill_1 FILLER_76_345 ();
 sg13g2_fill_2 FILLER_76_377 ();
 sg13g2_fill_2 FILLER_76_391 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_fill_2 FILLER_77_84 ();
 sg13g2_fill_1 FILLER_77_90 ();
 sg13g2_fill_2 FILLER_77_130 ();
 sg13g2_fill_1 FILLER_77_146 ();
 sg13g2_fill_1 FILLER_77_154 ();
 sg13g2_fill_1 FILLER_77_179 ();
 sg13g2_fill_2 FILLER_77_278 ();
 sg13g2_fill_1 FILLER_77_394 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_4 FILLER_78_77 ();
 sg13g2_fill_1 FILLER_78_94 ();
 sg13g2_fill_2 FILLER_78_165 ();
 sg13g2_fill_1 FILLER_78_167 ();
 sg13g2_decap_8 FILLER_78_186 ();
 sg13g2_fill_1 FILLER_78_217 ();
 sg13g2_fill_1 FILLER_78_263 ();
 sg13g2_fill_2 FILLER_78_315 ();
 sg13g2_fill_1 FILLER_78_331 ();
 sg13g2_fill_1 FILLER_78_350 ();
 sg13g2_fill_2 FILLER_78_381 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_4 FILLER_79_84 ();
 sg13g2_fill_1 FILLER_79_88 ();
 sg13g2_fill_2 FILLER_79_98 ();
 sg13g2_fill_1 FILLER_79_100 ();
 sg13g2_decap_4 FILLER_79_114 ();
 sg13g2_fill_2 FILLER_79_118 ();
 sg13g2_fill_2 FILLER_79_135 ();
 sg13g2_fill_1 FILLER_79_137 ();
 sg13g2_fill_1 FILLER_79_142 ();
 sg13g2_fill_2 FILLER_79_153 ();
 sg13g2_decap_4 FILLER_79_165 ();
 sg13g2_decap_8 FILLER_79_179 ();
 sg13g2_decap_8 FILLER_79_186 ();
 sg13g2_decap_8 FILLER_79_193 ();
 sg13g2_decap_4 FILLER_79_200 ();
 sg13g2_fill_1 FILLER_79_225 ();
 sg13g2_fill_2 FILLER_79_249 ();
 sg13g2_fill_2 FILLER_79_316 ();
 sg13g2_fill_1 FILLER_79_318 ();
 sg13g2_fill_1 FILLER_79_325 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_fill_2 FILLER_80_109 ();
 sg13g2_fill_1 FILLER_80_111 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_4 FILLER_80_208 ();
 sg13g2_fill_2 FILLER_80_212 ();
 sg13g2_decap_4 FILLER_80_218 ();
 sg13g2_fill_2 FILLER_80_338 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_399 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net25;
 assign uio_out[1] = net26;
 assign uio_out[2] = net27;
 assign uio_out[3] = net28;
 assign uio_out[4] = net29;
 assign uio_out[5] = net30;
 assign uio_out[6] = net31;
 assign uio_out[7] = net32;
endmodule

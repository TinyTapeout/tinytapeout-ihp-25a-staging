module tt_um_vga_cbtest (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire clknet_0_clk;
 wire hsync;
 wire \pix_x[0] ;
 wire \pix_x[1] ;
 wire \pix_x[2] ;
 wire \pix_x[3] ;
 wire \pix_x[4] ;
 wire \pix_x[5] ;
 wire \pix_x[6] ;
 wire \pix_x[7] ;
 wire \pix_x[8] ;
 wire \pix_x[9] ;
 wire \pix_y[0] ;
 wire \pix_y[1] ;
 wire \pix_y[2] ;
 wire \pix_y[3] ;
 wire \pix_y[4] ;
 wire \pix_y[5] ;
 wire \pix_y[6] ;
 wire \pix_y[7] ;
 wire \pix_y[8] ;
 wire \pix_y[9] ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire \vga_sync_gen.vsync ;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net1;
 wire net2;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;

 sg13g2_inv_1 _0502_ (.Y(_0419_),
    .A(net67));
 sg13g2_inv_1 _0503_ (.Y(_0420_),
    .A(\pix_y[6] ));
 sg13g2_inv_1 _0504_ (.Y(_0421_),
    .A(\pix_y[5] ));
 sg13g2_inv_1 _0505_ (.Y(_0422_),
    .A(net234));
 sg13g2_inv_2 _0506_ (.Y(_0423_),
    .A(net238));
 sg13g2_inv_2 _0507_ (.Y(_0424_),
    .A(net230));
 sg13g2_inv_2 _0508_ (.Y(_0425_),
    .A(net226));
 sg13g2_inv_1 _0509_ (.Y(_0426_),
    .A(\pix_y[4] ));
 sg13g2_inv_1 _0510_ (.Y(_0427_),
    .A(net1));
 sg13g2_inv_1 _0511_ (.Y(_0428_),
    .A(net250));
 sg13g2_inv_1 _0512_ (.Y(_0429_),
    .A(net254));
 sg13g2_inv_1 _0513_ (.Y(_0430_),
    .A(net245));
 sg13g2_inv_2 _0514_ (.Y(_0431_),
    .A(net240));
 sg13g2_nor2_2 _0515_ (.A(net229),
    .B(_0425_),
    .Y(_0432_));
 sg13g2_inv_1 _0516_ (.Y(_0433_),
    .A(_0432_));
 sg13g2_nand2_1 _0517_ (.Y(_0434_),
    .A(net233),
    .B(_0432_));
 sg13g2_nor2b_2 _0518_ (.A(net237),
    .B_N(net233),
    .Y(_0435_));
 sg13g2_nand2b_2 _0519_ (.Y(_0436_),
    .B(net233),
    .A_N(net237));
 sg13g2_nand3_1 _0520_ (.B(_0424_),
    .C(net221),
    .A(net224),
    .Y(_0437_));
 sg13g2_nand2_2 _0521_ (.Y(_0438_),
    .A(\pix_y[5] ),
    .B(\pix_y[4] ));
 sg13g2_nor2b_1 _0522_ (.A(net61),
    .B_N(\pix_y[7] ),
    .Y(_0439_));
 sg13g2_nand3_1 _0523_ (.B(\pix_y[6] ),
    .C(_0439_),
    .A(\pix_y[8] ),
    .Y(_0440_));
 sg13g2_nand2b_1 _0524_ (.Y(_0441_),
    .B(_0438_),
    .A_N(_0440_));
 sg13g2_a221oi_1 _0525_ (.B2(net46),
    .C1(_0441_),
    .B1(_0437_),
    .A1(net224),
    .Y(_0001_),
    .A2(_0434_));
 sg13g2_nor2b_1 _0526_ (.A(net240),
    .B_N(net252),
    .Y(_0442_));
 sg13g2_nand2b_2 _0527_ (.Y(_0443_),
    .B(net252),
    .A_N(net241));
 sg13g2_nor2b_1 _0528_ (.A(net240),
    .B_N(net249),
    .Y(_0444_));
 sg13g2_nand2b_2 _0529_ (.Y(_0445_),
    .B(net249),
    .A_N(net240));
 sg13g2_or2_1 _0530_ (.X(_0446_),
    .B(net253),
    .A(net248));
 sg13g2_nor2b_1 _0531_ (.A(net247),
    .B_N(net242),
    .Y(_0447_));
 sg13g2_nand2b_2 _0532_ (.Y(_0448_),
    .B(net239),
    .A_N(net250));
 sg13g2_nor2b_1 _0533_ (.A(net253),
    .B_N(net243),
    .Y(_0449_));
 sg13g2_nand2b_2 _0534_ (.Y(_0450_),
    .B(net241),
    .A_N(net252));
 sg13g2_nor4_2 _0535_ (.A(net219),
    .B(net217),
    .C(net214),
    .Y(_0451_),
    .D(_0449_));
 sg13g2_nand3b_1 _0536_ (.B(\pix_x[9] ),
    .C(net63),
    .Y(_0452_),
    .A_N(net58));
 sg13g2_nor2_1 _0537_ (.A(_0451_),
    .B(net64),
    .Y(_0000_));
 sg13g2_and2_1 _0538_ (.A(net66),
    .B(net48),
    .X(_0453_));
 sg13g2_and3_2 _0539_ (.X(_0454_),
    .A(net257),
    .B(net51),
    .C(_0453_));
 sg13g2_nor2_2 _0540_ (.A(net249),
    .B(_0443_),
    .Y(_0455_));
 sg13g2_nor2b_1 _0541_ (.A(net78),
    .B_N(\pix_x[8] ),
    .Y(_0456_));
 sg13g2_nand4_1 _0542_ (.B(_0454_),
    .C(_0455_),
    .A(\pix_x[9] ),
    .Y(_0457_),
    .D(_0456_));
 sg13g2_and2_1 _0543_ (.A(net1),
    .B(_0457_),
    .X(_0037_));
 sg13g2_nand2_2 _0544_ (.Y(_0038_),
    .A(net1),
    .B(_0457_));
 sg13g2_and2_1 _0545_ (.A(net45),
    .B(net197),
    .X(_0012_));
 sg13g2_nor2_1 _0546_ (.A(\pix_x[0] ),
    .B(net48),
    .Y(_0039_));
 sg13g2_nor3_1 _0547_ (.A(_0427_),
    .B(_0453_),
    .C(net49),
    .Y(_0013_));
 sg13g2_o21ai_1 _0548_ (.B1(net1),
    .Y(_0040_),
    .A1(net51),
    .A2(_0453_));
 sg13g2_a21oi_1 _0549_ (.A1(net51),
    .A2(_0453_),
    .Y(_0014_),
    .B1(_0040_));
 sg13g2_a21oi_1 _0550_ (.A1(net51),
    .A2(_0453_),
    .Y(_0041_),
    .B1(net257));
 sg13g2_nor3_1 _0551_ (.A(_0427_),
    .B(_0454_),
    .C(_0041_),
    .Y(_0015_));
 sg13g2_xor2_1 _0552_ (.B(_0454_),
    .A(net71),
    .X(_0042_));
 sg13g2_nor2_1 _0553_ (.A(_0038_),
    .B(_0042_),
    .Y(_0016_));
 sg13g2_and2_1 _0554_ (.A(net251),
    .B(net255),
    .X(_0043_));
 sg13g2_nand2_2 _0555_ (.Y(_0044_),
    .A(net251),
    .B(net256));
 sg13g2_and3_1 _0556_ (.X(_0045_),
    .A(net247),
    .B(net253),
    .C(_0454_));
 sg13g2_a21oi_1 _0557_ (.A1(net253),
    .A2(_0454_),
    .Y(_0046_),
    .B1(net247));
 sg13g2_nor3_1 _0558_ (.A(_0038_),
    .B(_0045_),
    .C(_0046_),
    .Y(_0017_));
 sg13g2_and2_1 _0559_ (.A(net242),
    .B(_0045_),
    .X(_0047_));
 sg13g2_nor2_1 _0560_ (.A(net242),
    .B(_0045_),
    .Y(_0048_));
 sg13g2_nor3_1 _0561_ (.A(_0038_),
    .B(_0047_),
    .C(_0048_),
    .Y(_0018_));
 sg13g2_nor2b_1 _0562_ (.A(net65),
    .B_N(_0045_),
    .Y(_0049_));
 sg13g2_o21ai_1 _0563_ (.B1(net197),
    .Y(_0050_),
    .A1(net63),
    .A2(_0049_));
 sg13g2_a21oi_1 _0564_ (.A1(net63),
    .A2(_0049_),
    .Y(_0019_),
    .B1(_0050_));
 sg13g2_a21oi_1 _0565_ (.A1(\pix_x[7] ),
    .A2(_0047_),
    .Y(_0051_),
    .B1(net58));
 sg13g2_and3_1 _0566_ (.X(_0052_),
    .A(net63),
    .B(net58),
    .C(_0047_));
 sg13g2_nor3_1 _0567_ (.A(_0038_),
    .B(net59),
    .C(_0052_),
    .Y(_0020_));
 sg13g2_a21oi_1 _0568_ (.A1(net74),
    .A2(_0052_),
    .Y(_0053_),
    .B1(_0038_));
 sg13g2_o21ai_1 _0569_ (.B1(_0053_),
    .Y(_0054_),
    .A1(net74),
    .A2(_0052_));
 sg13g2_inv_1 _0570_ (.Y(_0021_),
    .A(_0054_));
 sg13g2_nor2_1 _0571_ (.A(net232),
    .B(net236),
    .Y(_0055_));
 sg13g2_nand2_2 _0572_ (.Y(_0056_),
    .A(_0422_),
    .B(_0423_));
 sg13g2_nor2_1 _0573_ (.A(net224),
    .B(\pix_y[4] ),
    .Y(_0057_));
 sg13g2_nor2_2 _0574_ (.A(_0424_),
    .B(_0425_),
    .Y(_0058_));
 sg13g2_nand2_2 _0575_ (.Y(_0059_),
    .A(net229),
    .B(net226));
 sg13g2_nor3_1 _0576_ (.A(\pix_y[8] ),
    .B(\pix_y[7] ),
    .C(\pix_y[6] ),
    .Y(_0060_));
 sg13g2_nand4_1 _0577_ (.B(_0057_),
    .C(_0058_),
    .A(\pix_y[9] ),
    .Y(_0061_),
    .D(_0060_));
 sg13g2_o21ai_1 _0578_ (.B1(net1),
    .Y(_0062_),
    .A1(_0056_),
    .A2(_0061_));
 sg13g2_or2_2 _0579_ (.X(_0063_),
    .B(_0062_),
    .A(_0457_));
 sg13g2_inv_1 _0580_ (.Y(_0064_),
    .A(_0063_));
 sg13g2_a22oi_1 _0581_ (.Y(_0065_),
    .B1(_0064_),
    .B2(net56),
    .A2(_0037_),
    .A1(net238));
 sg13g2_inv_1 _0582_ (.Y(_0022_),
    .A(net57));
 sg13g2_nor2_1 _0583_ (.A(net235),
    .B(_0423_),
    .Y(_0066_));
 sg13g2_nand2b_1 _0584_ (.Y(_0067_),
    .B(net236),
    .A_N(net232));
 sg13g2_nand2_2 _0585_ (.Y(_0068_),
    .A(net220),
    .B(net210));
 sg13g2_nand2_1 _0586_ (.Y(_0069_),
    .A(_0064_),
    .B(_0068_));
 sg13g2_o21ai_1 _0587_ (.B1(_0069_),
    .Y(_0023_),
    .A1(net223),
    .A2(_0038_));
 sg13g2_nand2_1 _0588_ (.Y(_0070_),
    .A(net228),
    .B(net197));
 sg13g2_and2_1 _0589_ (.A(net232),
    .B(net236),
    .X(_0071_));
 sg13g2_nand2_1 _0590_ (.Y(_0072_),
    .A(net233),
    .B(net237));
 sg13g2_xnor2_1 _0591_ (.Y(_0073_),
    .A(net228),
    .B(net208));
 sg13g2_o21ai_1 _0592_ (.B1(_0070_),
    .Y(_0024_),
    .A1(_0063_),
    .A2(_0073_));
 sg13g2_nand2_1 _0593_ (.Y(_0074_),
    .A(net226),
    .B(net197));
 sg13g2_nor2_1 _0594_ (.A(net70),
    .B(net207),
    .Y(_0075_));
 sg13g2_xnor2_1 _0595_ (.Y(_0076_),
    .A(net226),
    .B(_0075_));
 sg13g2_o21ai_1 _0596_ (.B1(_0074_),
    .Y(_0025_),
    .A1(_0063_),
    .A2(_0076_));
 sg13g2_and2_1 _0597_ (.A(_0038_),
    .B(_0062_),
    .X(_0077_));
 sg13g2_nor3_1 _0598_ (.A(net197),
    .B(_0059_),
    .C(net207),
    .Y(_0078_));
 sg13g2_xnor2_1 _0599_ (.Y(_0079_),
    .A(net77),
    .B(_0078_));
 sg13g2_nor2_1 _0600_ (.A(_0077_),
    .B(_0079_),
    .Y(_0026_));
 sg13g2_nand2_1 _0601_ (.Y(_0080_),
    .A(net224),
    .B(net197));
 sg13g2_nor3_1 _0602_ (.A(net72),
    .B(_0059_),
    .C(net207),
    .Y(_0081_));
 sg13g2_xnor2_1 _0603_ (.Y(_0082_),
    .A(net224),
    .B(_0081_));
 sg13g2_o21ai_1 _0604_ (.B1(_0080_),
    .Y(_0027_),
    .A1(_0063_),
    .A2(_0082_));
 sg13g2_nor4_2 _0605_ (.A(_0438_),
    .B(net197),
    .C(_0059_),
    .Y(_0083_),
    .D(net207));
 sg13g2_xnor2_1 _0606_ (.Y(_0084_),
    .A(net75),
    .B(_0083_));
 sg13g2_nor2_1 _0607_ (.A(_0077_),
    .B(net76),
    .Y(_0028_));
 sg13g2_nand2_1 _0608_ (.Y(_0085_),
    .A(net69),
    .B(net197));
 sg13g2_nor4_1 _0609_ (.A(net53),
    .B(_0438_),
    .C(_0059_),
    .D(net207),
    .Y(_0086_));
 sg13g2_xnor2_1 _0610_ (.Y(_0087_),
    .A(net69),
    .B(_0086_));
 sg13g2_o21ai_1 _0611_ (.B1(_0085_),
    .Y(_0029_),
    .A1(_0063_),
    .A2(_0087_));
 sg13g2_nand3_1 _0612_ (.B(\pix_y[6] ),
    .C(_0083_),
    .A(\pix_y[7] ),
    .Y(_0088_));
 sg13g2_or2_1 _0613_ (.X(_0089_),
    .B(_0088_),
    .A(_0419_));
 sg13g2_nor2b_1 _0614_ (.A(_0077_),
    .B_N(_0089_),
    .Y(_0090_));
 sg13g2_nand2b_1 _0615_ (.Y(_0091_),
    .B(_0089_),
    .A_N(_0077_));
 sg13g2_a21oi_1 _0616_ (.A1(_0419_),
    .A2(_0088_),
    .Y(_0030_),
    .B1(_0091_));
 sg13g2_nor2_1 _0617_ (.A(_0440_),
    .B(_0062_),
    .Y(_0092_));
 sg13g2_a22oi_1 _0618_ (.Y(_0093_),
    .B1(_0092_),
    .B2(_0083_),
    .A2(_0090_),
    .A1(net61));
 sg13g2_inv_1 _0619_ (.Y(_0031_),
    .A(net62));
 sg13g2_nor2_1 _0620_ (.A(net252),
    .B(net258),
    .Y(_0094_));
 sg13g2_nor2_2 _0621_ (.A(net247),
    .B(\pix_x[3] ),
    .Y(_0095_));
 sg13g2_a21oi_1 _0622_ (.A1(net253),
    .A2(net257),
    .Y(_0096_),
    .B1(net247));
 sg13g2_o21ai_1 _0623_ (.B1(net242),
    .Y(_0097_),
    .A1(_0094_),
    .A2(_0096_));
 sg13g2_nor2_2 _0624_ (.A(net245),
    .B(net239),
    .Y(_0098_));
 sg13g2_or2_2 _0625_ (.X(_0099_),
    .B(net244),
    .A(net245));
 sg13g2_nor2_2 _0626_ (.A(_0044_),
    .B(_0099_),
    .Y(_0100_));
 sg13g2_nand3b_1 _0627_ (.B(net234),
    .C(_0097_),
    .Y(_0101_),
    .A_N(_0100_));
 sg13g2_nor2b_2 _0628_ (.A(net257),
    .B_N(net248),
    .Y(_0102_));
 sg13g2_nor2_1 _0629_ (.A(_0431_),
    .B(_0096_),
    .Y(_0103_));
 sg13g2_nand2_1 _0630_ (.Y(_0104_),
    .A(net247),
    .B(net257));
 sg13g2_a21oi_1 _0631_ (.A1(net248),
    .A2(net257),
    .Y(_0105_),
    .B1(net242));
 sg13g2_nor3_1 _0632_ (.A(net238),
    .B(net248),
    .C(_0429_),
    .Y(_0106_));
 sg13g2_or3_1 _0633_ (.A(_0103_),
    .B(_0105_),
    .C(_0106_),
    .X(_0107_));
 sg13g2_a22oi_1 _0634_ (.Y(_0108_),
    .B1(_0107_),
    .B2(net223),
    .A2(_0102_),
    .A1(_0435_));
 sg13g2_a21oi_1 _0635_ (.A1(_0101_),
    .A2(_0108_),
    .Y(_0109_),
    .B1(_0059_));
 sg13g2_nor2b_2 _0636_ (.A(net251),
    .B_N(net255),
    .Y(_0110_));
 sg13g2_nand2b_2 _0637_ (.Y(_0111_),
    .B(net255),
    .A_N(net251));
 sg13g2_nand3b_1 _0638_ (.B(net258),
    .C(net249),
    .Y(_0112_),
    .A_N(net252));
 sg13g2_nand2_1 _0639_ (.Y(_0113_),
    .A(_0431_),
    .B(_0112_));
 sg13g2_nand2b_1 _0640_ (.Y(_0114_),
    .B(net240),
    .A_N(net246));
 sg13g2_o21ai_1 _0641_ (.B1(net244),
    .Y(_0115_),
    .A1(_0430_),
    .A2(net203));
 sg13g2_a21oi_1 _0642_ (.A1(_0113_),
    .A2(_0115_),
    .Y(_0116_),
    .B1(_0056_));
 sg13g2_nor2_2 _0643_ (.A(_0099_),
    .B(_0111_),
    .Y(_0117_));
 sg13g2_nand2_1 _0644_ (.Y(_0118_),
    .A(_0098_),
    .B(net204));
 sg13g2_nor2_2 _0645_ (.A(net216),
    .B(net203),
    .Y(_0119_));
 sg13g2_nand2_1 _0646_ (.Y(_0120_),
    .A(net217),
    .B(net204));
 sg13g2_o21ai_1 _0647_ (.B1(net238),
    .Y(_0121_),
    .A1(_0445_),
    .A2(_0111_));
 sg13g2_nor2b_1 _0648_ (.A(net247),
    .B_N(net257),
    .Y(_0122_));
 sg13g2_nor2_1 _0649_ (.A(_0448_),
    .B(net203),
    .Y(_0123_));
 sg13g2_nand2_1 _0650_ (.Y(_0124_),
    .A(net214),
    .B(net204));
 sg13g2_nor2_1 _0651_ (.A(_0121_),
    .B(_0123_),
    .Y(_0125_));
 sg13g2_nor2_2 _0652_ (.A(net210),
    .B(_0119_),
    .Y(_0126_));
 sg13g2_a221oi_1 _0653_ (.B2(_0126_),
    .C1(net229),
    .B1(_0124_),
    .A1(net233),
    .Y(_0127_),
    .A2(_0118_));
 sg13g2_nand2b_1 _0654_ (.Y(_0128_),
    .B(_0127_),
    .A_N(_0116_));
 sg13g2_nand2b_1 _0655_ (.Y(_0129_),
    .B(net246),
    .A_N(net258));
 sg13g2_and2_2 _0656_ (.A(net245),
    .B(net239),
    .X(_0130_));
 sg13g2_nand2_2 _0657_ (.Y(_0131_),
    .A(net246),
    .B(net241));
 sg13g2_nor2_2 _0658_ (.A(_0450_),
    .B(_0129_),
    .Y(_0132_));
 sg13g2_nand2_1 _0659_ (.Y(_0133_),
    .A(net205),
    .B(_0130_));
 sg13g2_nor2_1 _0660_ (.A(net220),
    .B(_0132_),
    .Y(_0134_));
 sg13g2_o21ai_1 _0661_ (.B1(net228),
    .Y(_0135_),
    .A1(_0068_),
    .A2(_0119_));
 sg13g2_a221oi_1 _0662_ (.B2(_0118_),
    .C1(_0135_),
    .B1(_0134_),
    .A1(_0126_),
    .Y(_0136_),
    .A2(_0133_));
 sg13g2_nor2_1 _0663_ (.A(net225),
    .B(_0136_),
    .Y(_0137_));
 sg13g2_a22oi_1 _0664_ (.Y(_0138_),
    .B1(_0122_),
    .B2(_0423_),
    .A2(_0446_),
    .A1(net242));
 sg13g2_nand3_1 _0665_ (.B(_0113_),
    .C(_0138_),
    .A(net234),
    .Y(_0139_));
 sg13g2_a221oi_1 _0666_ (.B2(net198),
    .C1(_0433_),
    .B1(_0132_),
    .A1(net223),
    .Y(_0140_),
    .A2(_0117_));
 sg13g2_a221oi_1 _0667_ (.B2(_0140_),
    .C1(_0109_),
    .B1(_0139_),
    .A1(_0128_),
    .Y(_0141_),
    .A2(_0137_));
 sg13g2_nor2_1 _0668_ (.A(\pix_y[4] ),
    .B(_0141_),
    .Y(_0142_));
 sg13g2_nand2_1 _0669_ (.Y(_0143_),
    .A(\pix_y[6] ),
    .B(net46));
 sg13g2_nor2b_2 _0670_ (.A(net255),
    .B_N(net251),
    .Y(_0144_));
 sg13g2_nand2b_1 _0671_ (.Y(_0145_),
    .B(net253),
    .A_N(net258));
 sg13g2_xnor2_1 _0672_ (.Y(_0146_),
    .A(net251),
    .B(net255));
 sg13g2_xor2_1 _0673_ (.B(net255),
    .A(net251),
    .X(_0147_));
 sg13g2_nand3_1 _0674_ (.B(net214),
    .C(_0147_),
    .A(net236),
    .Y(_0148_));
 sg13g2_nor2_2 _0675_ (.A(net254),
    .B(_0445_),
    .Y(_0149_));
 sg13g2_nor2_2 _0676_ (.A(net255),
    .B(_0448_),
    .Y(_0150_));
 sg13g2_a21oi_1 _0677_ (.A1(net254),
    .A2(_0150_),
    .Y(_0151_),
    .B1(_0149_));
 sg13g2_a21o_1 _0678_ (.A2(_0150_),
    .A1(net254),
    .B1(_0149_),
    .X(_0152_));
 sg13g2_nand2_1 _0679_ (.Y(_0153_),
    .A(net233),
    .B(_0124_));
 sg13g2_a21oi_1 _0680_ (.A1(_0148_),
    .A2(_0152_),
    .Y(_0154_),
    .B1(_0153_));
 sg13g2_a22oi_1 _0681_ (.Y(_0155_),
    .B1(_0147_),
    .B2(net214),
    .A2(_0095_),
    .A1(net219));
 sg13g2_nor2_2 _0682_ (.A(net243),
    .B(_0104_),
    .Y(_0156_));
 sg13g2_nor2_1 _0683_ (.A(_0150_),
    .B(_0156_),
    .Y(_0157_));
 sg13g2_a221oi_1 _0684_ (.B2(net212),
    .C1(_0154_),
    .B1(_0157_),
    .A1(_0126_),
    .Y(_0158_),
    .A2(_0155_));
 sg13g2_nor2_2 _0685_ (.A(_0010_),
    .B(net233),
    .Y(_0159_));
 sg13g2_nand2b_2 _0686_ (.Y(_0160_),
    .B(net245),
    .A_N(_0009_));
 sg13g2_nor2_2 _0687_ (.A(net203),
    .B(_0160_),
    .Y(_0161_));
 sg13g2_nand2_1 _0688_ (.Y(_0162_),
    .A(_0159_),
    .B(_0161_));
 sg13g2_nand3_1 _0689_ (.B(net212),
    .C(_0119_),
    .A(net225),
    .Y(_0163_));
 sg13g2_a22oi_1 _0690_ (.Y(_0164_),
    .B1(_0163_),
    .B2(net228),
    .A2(_0162_),
    .A1(_0432_));
 sg13g2_o21ai_1 _0691_ (.B1(_0164_),
    .Y(_0165_),
    .A1(net225),
    .A2(_0158_));
 sg13g2_a21o_1 _0692_ (.A2(_0165_),
    .A1(\pix_y[4] ),
    .B1(_0143_),
    .X(_0166_));
 sg13g2_nor2_1 _0693_ (.A(_0110_),
    .B(net202),
    .Y(_0167_));
 sg13g2_nand2_1 _0694_ (.Y(_0168_),
    .A(net203),
    .B(_0130_));
 sg13g2_nor2_2 _0695_ (.A(net202),
    .B(_0147_),
    .Y(_0169_));
 sg13g2_a22oi_1 _0696_ (.Y(_0170_),
    .B1(_0130_),
    .B2(_0146_),
    .A2(net204),
    .A1(net217));
 sg13g2_nand2b_1 _0697_ (.Y(_0171_),
    .B(net232),
    .A_N(_0170_));
 sg13g2_nor2_1 _0698_ (.A(net216),
    .B(net200),
    .Y(_0172_));
 sg13g2_o21ai_1 _0699_ (.B1(net211),
    .Y(_0173_),
    .A1(_0132_),
    .A2(_0172_));
 sg13g2_o21ai_1 _0700_ (.B1(net198),
    .Y(_0174_),
    .A1(_0117_),
    .A2(_0169_));
 sg13g2_nand3_1 _0701_ (.B(_0173_),
    .C(_0174_),
    .A(_0171_),
    .Y(_0175_));
 sg13g2_o21ai_1 _0702_ (.B1(net244),
    .Y(_0176_),
    .A1(net250),
    .A2(_0146_));
 sg13g2_a22oi_1 _0703_ (.Y(_0177_),
    .B1(_0176_),
    .B2(net233),
    .A2(_0159_),
    .A1(_0115_));
 sg13g2_a21oi_1 _0704_ (.A1(_0430_),
    .A2(_0144_),
    .Y(_0178_),
    .B1(net239));
 sg13g2_nand2_1 _0705_ (.Y(_0179_),
    .A(net229),
    .B(_0425_));
 sg13g2_nor3_1 _0706_ (.A(_0177_),
    .B(_0178_),
    .C(_0179_),
    .Y(_0180_));
 sg13g2_nand3_1 _0707_ (.B(net246),
    .C(net240),
    .A(net252),
    .Y(_0181_));
 sg13g2_nand2_1 _0708_ (.Y(_0182_),
    .A(_0130_),
    .B(_0144_));
 sg13g2_a21oi_1 _0709_ (.A1(net216),
    .A2(net202),
    .Y(_0183_),
    .B1(net200));
 sg13g2_a22oi_1 _0710_ (.Y(_0184_),
    .B1(_0183_),
    .B2(net198),
    .A2(_0132_),
    .A1(net208));
 sg13g2_nand3_1 _0711_ (.B(net211),
    .C(_0147_),
    .A(net214),
    .Y(_0185_));
 sg13g2_o21ai_1 _0712_ (.B1(net221),
    .Y(_0186_),
    .A1(_0150_),
    .A2(_0172_));
 sg13g2_nand3_1 _0713_ (.B(_0185_),
    .C(_0186_),
    .A(_0184_),
    .Y(_0187_));
 sg13g2_a21oi_1 _0714_ (.A1(_0432_),
    .A2(_0187_),
    .Y(_0188_),
    .B1(_0180_));
 sg13g2_nor2_1 _0715_ (.A(_0010_),
    .B(net223),
    .Y(_0189_));
 sg13g2_nor3_1 _0716_ (.A(net250),
    .B(_0009_),
    .C(net200),
    .Y(_0190_));
 sg13g2_a221oi_1 _0717_ (.B2(_0159_),
    .C1(_0425_),
    .B1(_0190_),
    .A1(_0100_),
    .Y(_0191_),
    .A2(_0189_));
 sg13g2_a21oi_1 _0718_ (.A1(net212),
    .A2(_0100_),
    .Y(_0192_),
    .B1(net225));
 sg13g2_nor4_1 _0719_ (.A(_0426_),
    .B(_0007_),
    .C(_0191_),
    .D(_0192_),
    .Y(_0193_));
 sg13g2_nor2_1 _0720_ (.A(net236),
    .B(_0117_),
    .Y(_0194_));
 sg13g2_a22oi_1 _0721_ (.Y(_0195_),
    .B1(_0098_),
    .B2(net204),
    .A2(_0095_),
    .A1(net239));
 sg13g2_a221oi_1 _0722_ (.B2(net236),
    .C1(net232),
    .B1(_0195_),
    .A1(_0168_),
    .Y(_0196_),
    .A2(_0194_));
 sg13g2_o21ai_1 _0723_ (.B1(net221),
    .Y(_0197_),
    .A1(_0119_),
    .A2(_0150_));
 sg13g2_nor3_1 _0724_ (.A(net206),
    .B(net200),
    .C(_0160_),
    .Y(_0198_));
 sg13g2_nand3b_1 _0725_ (.B(net225),
    .C(_0197_),
    .Y(_0199_),
    .A_N(_0198_));
 sg13g2_o21ai_1 _0726_ (.B1(net211),
    .Y(_0200_),
    .A1(_0117_),
    .A2(_0169_));
 sg13g2_nor3_1 _0727_ (.A(net211),
    .B(_0147_),
    .C(_0160_),
    .Y(_0201_));
 sg13g2_nor2_1 _0728_ (.A(net225),
    .B(_0201_),
    .Y(_0202_));
 sg13g2_a21oi_1 _0729_ (.A1(_0200_),
    .A2(_0202_),
    .Y(_0203_),
    .B1(net228));
 sg13g2_o21ai_1 _0730_ (.B1(_0203_),
    .Y(_0204_),
    .A1(_0196_),
    .A2(_0199_));
 sg13g2_a21oi_1 _0731_ (.A1(_0120_),
    .A2(_0182_),
    .Y(_0205_),
    .B1(net232));
 sg13g2_o21ai_1 _0732_ (.B1(net232),
    .Y(_0206_),
    .A1(net236),
    .A2(_0117_));
 sg13g2_a21oi_1 _0733_ (.A1(_0182_),
    .A2(_0206_),
    .Y(_0207_),
    .B1(_0125_));
 sg13g2_o21ai_1 _0734_ (.B1(_0058_),
    .Y(_0208_),
    .A1(_0205_),
    .A2(_0207_));
 sg13g2_a21oi_1 _0735_ (.A1(net217),
    .A2(net205),
    .Y(_0209_),
    .B1(net232));
 sg13g2_o21ai_1 _0736_ (.B1(_0209_),
    .Y(_0210_),
    .A1(net236),
    .A2(_0170_));
 sg13g2_nand2b_1 _0737_ (.Y(_0211_),
    .B(_0133_),
    .A_N(_0210_));
 sg13g2_a221oi_1 _0738_ (.B2(net208),
    .C1(_0179_),
    .B1(_0195_),
    .A1(_0120_),
    .Y(_0212_),
    .A2(_0134_));
 sg13g2_a21oi_1 _0739_ (.A1(_0211_),
    .A2(_0212_),
    .Y(_0213_),
    .B1(_0438_));
 sg13g2_nand3_1 _0740_ (.B(_0208_),
    .C(_0213_),
    .A(_0204_),
    .Y(_0214_));
 sg13g2_a21oi_1 _0741_ (.A1(_0058_),
    .A2(_0175_),
    .Y(_0215_),
    .B1(\pix_y[4] ));
 sg13g2_o21ai_1 _0742_ (.B1(_0420_),
    .Y(_0216_),
    .A1(net224),
    .A2(_0193_));
 sg13g2_a21oi_1 _0743_ (.A1(_0188_),
    .A2(_0215_),
    .Y(_0217_),
    .B1(_0216_));
 sg13g2_nand2_1 _0744_ (.Y(_0218_),
    .A(_0214_),
    .B(_0217_));
 sg13g2_o21ai_1 _0745_ (.B1(_0218_),
    .Y(_0219_),
    .A1(_0142_),
    .A2(_0166_));
 sg13g2_nand2b_1 _0746_ (.Y(_0220_),
    .B(_0003_),
    .A_N(net249));
 sg13g2_nand2_1 _0747_ (.Y(_0221_),
    .A(net249),
    .B(net205));
 sg13g2_mux2_1 _0748_ (.A0(_0003_),
    .A1(net205),
    .S(net249),
    .X(_0222_));
 sg13g2_and2_1 _0749_ (.A(net240),
    .B(_0222_),
    .X(_0223_));
 sg13g2_a221oi_1 _0750_ (.B2(net240),
    .C1(_0121_),
    .B1(_0222_),
    .A1(net258),
    .Y(_0224_),
    .A2(_0455_));
 sg13g2_nand3b_1 _0751_ (.B(net241),
    .C(_0003_),
    .Y(_0225_),
    .A_N(net252));
 sg13g2_nand2_2 _0752_ (.Y(_0226_),
    .A(_0181_),
    .B(_0225_));
 sg13g2_nor3_1 _0753_ (.A(\pix_y[0] ),
    .B(_0117_),
    .C(_0226_),
    .Y(_0227_));
 sg13g2_or3_1 _0754_ (.A(net234),
    .B(_0224_),
    .C(_0227_),
    .X(_0228_));
 sg13g2_nor2_1 _0755_ (.A(net215),
    .B(_0146_),
    .Y(_0229_));
 sg13g2_a21oi_1 _0756_ (.A1(_0112_),
    .A2(_0220_),
    .Y(_0230_),
    .B1(_0431_));
 sg13g2_or2_1 _0757_ (.X(_0231_),
    .B(_0230_),
    .A(_0229_));
 sg13g2_nand3_1 _0758_ (.B(net203),
    .C(net201),
    .A(_0447_),
    .Y(_0232_));
 sg13g2_nand3b_1 _0759_ (.B(_0112_),
    .C(_0232_),
    .Y(_0233_),
    .A_N(_0455_));
 sg13g2_a221oi_1 _0760_ (.B2(net209),
    .C1(_0424_),
    .B1(_0233_),
    .A1(net222),
    .Y(_0234_),
    .A2(_0231_));
 sg13g2_a22oi_1 _0761_ (.Y(_0235_),
    .B1(net201),
    .B2(net214),
    .A2(_0095_),
    .A1(_0442_));
 sg13g2_a21o_1 _0762_ (.A2(_0235_),
    .A1(_0112_),
    .B1(net210),
    .X(_0236_));
 sg13g2_a21o_1 _0763_ (.A2(net215),
    .A1(_0443_),
    .B1(_0102_),
    .X(_0237_));
 sg13g2_nand2_1 _0764_ (.Y(_0238_),
    .A(_0449_),
    .B(_0104_));
 sg13g2_o21ai_1 _0765_ (.B1(_0237_),
    .Y(_0239_),
    .A1(_0095_),
    .A2(_0238_));
 sg13g2_a21oi_2 _0766_ (.B1(_0144_),
    .Y(_0240_),
    .A2(net215),
    .A1(_0443_));
 sg13g2_nand2b_1 _0767_ (.Y(_0241_),
    .B(_0004_),
    .A_N(net247));
 sg13g2_a21oi_1 _0768_ (.A1(_0221_),
    .A2(_0241_),
    .Y(_0242_),
    .B1(_0431_));
 sg13g2_o21ai_1 _0769_ (.B1(net209),
    .Y(_0243_),
    .A1(_0240_),
    .A2(_0242_));
 sg13g2_a21oi_1 _0770_ (.A1(_0112_),
    .A2(_0241_),
    .Y(_0244_),
    .B1(_0431_));
 sg13g2_nand2b_1 _0771_ (.Y(_0245_),
    .B(net252),
    .A_N(_0003_));
 sg13g2_o21ai_1 _0772_ (.B1(_0245_),
    .Y(_0246_),
    .A1(net219),
    .A2(net218));
 sg13g2_nand2b_1 _0773_ (.Y(_0247_),
    .B(_0246_),
    .A_N(_0244_));
 sg13g2_a22oi_1 _0774_ (.Y(_0248_),
    .B1(_0247_),
    .B2(net222),
    .A2(_0239_),
    .A1(net213));
 sg13g2_nand4_1 _0775_ (.B(_0236_),
    .C(_0243_),
    .A(_0424_),
    .Y(_0249_),
    .D(_0248_));
 sg13g2_a21oi_1 _0776_ (.A1(_0228_),
    .A2(_0234_),
    .Y(_0250_),
    .B1(net227));
 sg13g2_o21ai_1 _0777_ (.B1(net213),
    .Y(_0251_),
    .A1(_0240_),
    .A2(_0244_));
 sg13g2_o21ai_1 _0778_ (.B1(net239),
    .Y(_0252_),
    .A1(net245),
    .A2(net205));
 sg13g2_o21ai_1 _0779_ (.B1(net202),
    .Y(_0253_),
    .A1(net258),
    .A2(_0450_));
 sg13g2_a21oi_1 _0780_ (.A1(_0423_),
    .A2(_0105_),
    .Y(_0254_),
    .B1(net223));
 sg13g2_o21ai_1 _0781_ (.B1(_0254_),
    .Y(_0255_),
    .A1(_0240_),
    .A2(_0253_));
 sg13g2_a21o_1 _0782_ (.A2(_0237_),
    .A1(_0131_),
    .B1(net210),
    .X(_0256_));
 sg13g2_nand4_1 _0783_ (.B(_0251_),
    .C(_0255_),
    .A(net230),
    .Y(_0257_),
    .D(_0256_));
 sg13g2_o21ai_1 _0784_ (.B1(net213),
    .Y(_0258_),
    .A1(_0149_),
    .A2(_0150_));
 sg13g2_nor2_1 _0785_ (.A(_0436_),
    .B(_0131_),
    .Y(_0259_));
 sg13g2_a21oi_1 _0786_ (.A1(_0443_),
    .A2(_0450_),
    .Y(_0260_),
    .B1(net258));
 sg13g2_o21ai_1 _0787_ (.B1(net199),
    .Y(_0261_),
    .A1(_0156_),
    .A2(_0260_));
 sg13g2_a22oi_1 _0788_ (.Y(_0262_),
    .B1(_0259_),
    .B2(net200),
    .A2(_0156_),
    .A1(net234));
 sg13g2_a21oi_1 _0789_ (.A1(net209),
    .A2(_0244_),
    .Y(_0263_),
    .B1(net230));
 sg13g2_nand4_1 _0790_ (.B(_0261_),
    .C(_0262_),
    .A(_0258_),
    .Y(_0264_),
    .D(_0263_));
 sg13g2_and3_1 _0791_ (.X(_0265_),
    .A(net227),
    .B(_0257_),
    .C(_0264_));
 sg13g2_a21o_1 _0792_ (.A2(_0250_),
    .A1(_0249_),
    .B1(_0265_),
    .X(_0266_));
 sg13g2_nand2b_1 _0793_ (.Y(_0267_),
    .B(_0115_),
    .A_N(_0178_));
 sg13g2_o21ai_1 _0794_ (.B1(net221),
    .Y(_0268_),
    .A1(net251),
    .A2(net216));
 sg13g2_o21ai_1 _0795_ (.B1(_0268_),
    .Y(_0269_),
    .A1(net210),
    .A2(_0156_));
 sg13g2_nand2_1 _0796_ (.Y(_0270_),
    .A(net256),
    .B(net214));
 sg13g2_nand3_1 _0797_ (.B(_0099_),
    .C(_0270_),
    .A(net198),
    .Y(_0271_));
 sg13g2_nor2_1 _0798_ (.A(_0429_),
    .B(net215),
    .Y(_0272_));
 sg13g2_nor2_1 _0799_ (.A(net220),
    .B(_0272_),
    .Y(_0273_));
 sg13g2_o21ai_1 _0800_ (.B1(net212),
    .Y(_0274_),
    .A1(_0099_),
    .A2(_0110_));
 sg13g2_a22oi_1 _0801_ (.Y(_0275_),
    .B1(net200),
    .B2(net214),
    .A2(net203),
    .A1(_0098_));
 sg13g2_and2_1 _0802_ (.A(net212),
    .B(_0275_),
    .X(_0276_));
 sg13g2_a221oi_1 _0803_ (.B2(_0098_),
    .C1(net206),
    .B1(_0147_),
    .A1(net204),
    .Y(_0277_),
    .A2(_0130_));
 sg13g2_nor4_1 _0804_ (.A(net228),
    .B(_0273_),
    .C(_0276_),
    .D(_0277_),
    .Y(_0278_));
 sg13g2_a21o_1 _0805_ (.A2(_0176_),
    .A1(_0113_),
    .B1(net206),
    .X(_0279_));
 sg13g2_a221oi_1 _0806_ (.B2(_0133_),
    .C1(_0424_),
    .B1(_0269_),
    .A1(net211),
    .Y(_0280_),
    .A2(_0267_));
 sg13g2_a221oi_1 _0807_ (.B2(_0280_),
    .C1(net225),
    .B1(_0279_),
    .A1(_0271_),
    .Y(_0281_),
    .A2(_0278_));
 sg13g2_a22oi_1 _0808_ (.Y(_0282_),
    .B1(_0161_),
    .B2(net211),
    .A2(_0100_),
    .A1(net221));
 sg13g2_nand2_1 _0809_ (.Y(_0283_),
    .A(_0058_),
    .B(_0282_));
 sg13g2_nor4_2 _0810_ (.A(net238),
    .B(net250),
    .C(net256),
    .Y(_0284_),
    .D(_0009_));
 sg13g2_nor4_1 _0811_ (.A(net250),
    .B(_0009_),
    .C(_0146_),
    .D(_0284_),
    .Y(_0285_));
 sg13g2_a21oi_1 _0812_ (.A1(_0429_),
    .A2(_0284_),
    .Y(_0286_),
    .B1(net235));
 sg13g2_nor2b_1 _0813_ (.A(_0285_),
    .B_N(_0286_),
    .Y(_0287_));
 sg13g2_o21ai_1 _0814_ (.B1(net208),
    .Y(_0288_),
    .A1(_0099_),
    .A2(net200));
 sg13g2_o21ai_1 _0815_ (.B1(_0288_),
    .Y(_0289_),
    .A1(net220),
    .A2(_0161_));
 sg13g2_o21ai_1 _0816_ (.B1(_0432_),
    .Y(_0290_),
    .A1(_0287_),
    .A2(_0289_));
 sg13g2_nand4_1 _0817_ (.B(_0002_),
    .C(_0283_),
    .A(\pix_y[5] ),
    .Y(_0291_),
    .D(_0290_));
 sg13g2_nor2_1 _0818_ (.A(net224),
    .B(_0426_),
    .Y(_0292_));
 sg13g2_nor2_1 _0819_ (.A(net255),
    .B(net216),
    .Y(_0293_));
 sg13g2_a21oi_1 _0820_ (.A1(_0431_),
    .A2(_0102_),
    .Y(_0294_),
    .B1(net234));
 sg13g2_nand2_1 _0821_ (.Y(_0295_),
    .A(net218),
    .B(_0043_));
 sg13g2_a21oi_1 _0822_ (.A1(net234),
    .A2(_0295_),
    .Y(_0296_),
    .B1(_0294_));
 sg13g2_o21ai_1 _0823_ (.B1(net238),
    .Y(_0297_),
    .A1(_0223_),
    .A2(_0296_));
 sg13g2_a22oi_1 _0824_ (.Y(_0298_),
    .B1(_0122_),
    .B2(net219),
    .A2(net218),
    .A1(_0004_));
 sg13g2_a21o_1 _0825_ (.A2(_0298_),
    .A1(_0270_),
    .B1(_0056_),
    .X(_0299_));
 sg13g2_o21ai_1 _0826_ (.B1(_0435_),
    .Y(_0300_),
    .A1(_0455_),
    .A2(_0150_));
 sg13g2_and3_1 _0827_ (.X(_0301_),
    .A(net231),
    .B(_0299_),
    .C(_0300_));
 sg13g2_nor2_1 _0828_ (.A(net216),
    .B(_0144_),
    .Y(_0302_));
 sg13g2_nor2_1 _0829_ (.A(_0043_),
    .B(net202),
    .Y(_0303_));
 sg13g2_nand2_1 _0830_ (.Y(_0304_),
    .A(_0044_),
    .B(_0130_));
 sg13g2_a22oi_1 _0831_ (.Y(_0305_),
    .B1(net201),
    .B2(net218),
    .A2(_0095_),
    .A1(_0442_));
 sg13g2_nand2_1 _0832_ (.Y(_0306_),
    .A(_0304_),
    .B(_0305_));
 sg13g2_o21ai_1 _0833_ (.B1(_0306_),
    .Y(_0307_),
    .A1(net199),
    .A2(_0294_));
 sg13g2_nor2_1 _0834_ (.A(net220),
    .B(_0298_),
    .Y(_0308_));
 sg13g2_a21oi_1 _0835_ (.A1(net246),
    .A2(net205),
    .Y(_0309_),
    .B1(net223));
 sg13g2_a221oi_1 _0836_ (.B2(_0309_),
    .C1(net230),
    .B1(_0253_),
    .A1(net209),
    .Y(_0310_),
    .A2(_0149_));
 sg13g2_nor2b_1 _0837_ (.A(_0308_),
    .B_N(_0310_),
    .Y(_0311_));
 sg13g2_a221oi_1 _0838_ (.B2(_0311_),
    .C1(net227),
    .B1(_0307_),
    .A1(_0297_),
    .Y(_0312_),
    .A2(_0301_));
 sg13g2_o21ai_1 _0839_ (.B1(net221),
    .Y(_0313_),
    .A1(_0169_),
    .A2(_0293_));
 sg13g2_nand2_1 _0840_ (.Y(_0314_),
    .A(net215),
    .B(_0181_));
 sg13g2_nand3_1 _0841_ (.B(net201),
    .C(_0314_),
    .A(net209),
    .Y(_0315_));
 sg13g2_o21ai_1 _0842_ (.B1(net198),
    .Y(_0316_),
    .A1(_0123_),
    .A2(_0156_));
 sg13g2_a21o_1 _0843_ (.A2(_0295_),
    .A1(_0182_),
    .B1(_0056_),
    .X(_0317_));
 sg13g2_nand4_1 _0844_ (.B(_0315_),
    .C(_0316_),
    .A(_0313_),
    .Y(_0318_),
    .D(_0317_));
 sg13g2_nor2_1 _0845_ (.A(net205),
    .B(net202),
    .Y(_0319_));
 sg13g2_nor3_1 _0846_ (.A(_0043_),
    .B(net205),
    .C(net202),
    .Y(_0320_));
 sg13g2_nor2_1 _0847_ (.A(net216),
    .B(net204),
    .Y(_0321_));
 sg13g2_o21ai_1 _0848_ (.B1(net198),
    .Y(_0322_),
    .A1(_0320_),
    .A2(_0321_));
 sg13g2_o21ai_1 _0849_ (.B1(net208),
    .Y(_0323_),
    .A1(_0150_),
    .A2(_0156_));
 sg13g2_o21ai_1 _0850_ (.B1(_0146_),
    .Y(_0324_),
    .A1(net219),
    .A2(net217));
 sg13g2_a21o_1 _0851_ (.A2(_0324_),
    .A1(_0182_),
    .B1(net220),
    .X(_0325_));
 sg13g2_nand2b_1 _0852_ (.Y(_0326_),
    .B(net211),
    .A_N(_0195_));
 sg13g2_nand4_1 _0853_ (.B(_0323_),
    .C(_0325_),
    .A(_0322_),
    .Y(_0327_),
    .D(_0326_));
 sg13g2_a22oi_1 _0854_ (.Y(_0328_),
    .B1(_0327_),
    .B2(_0058_),
    .A2(_0318_),
    .A1(_0432_));
 sg13g2_nand2b_1 _0855_ (.Y(_0329_),
    .B(_0328_),
    .A_N(_0312_));
 sg13g2_o21ai_1 _0856_ (.B1(\pix_y[6] ),
    .Y(_0330_),
    .A1(_0281_),
    .A2(_0291_));
 sg13g2_a221oi_1 _0857_ (.B2(_0329_),
    .C1(_0330_),
    .B1(_0292_),
    .A1(_0057_),
    .Y(_0331_),
    .A2(_0266_));
 sg13g2_a21oi_1 _0858_ (.A1(_0246_),
    .A2(_0252_),
    .Y(_0332_),
    .B1(net206));
 sg13g2_a22oi_1 _0859_ (.Y(_0333_),
    .B1(net203),
    .B2(_0130_),
    .A2(_0095_),
    .A1(net219));
 sg13g2_a21o_1 _0860_ (.A2(_0333_),
    .A1(_0120_),
    .B1(_0056_),
    .X(_0334_));
 sg13g2_a21oi_1 _0861_ (.A1(net245),
    .A2(net200),
    .Y(_0335_),
    .B1(net239));
 sg13g2_o21ai_1 _0862_ (.B1(net222),
    .Y(_0336_),
    .A1(_0167_),
    .A2(_0335_));
 sg13g2_or2_1 _0863_ (.X(_0337_),
    .B(_0246_),
    .A(_0067_));
 sg13g2_a21oi_1 _0864_ (.A1(_0181_),
    .A2(_0225_),
    .Y(_0338_),
    .B1(net210));
 sg13g2_nand2_1 _0865_ (.Y(_0339_),
    .A(net199),
    .B(_0226_));
 sg13g2_nor3_1 _0866_ (.A(_0423_),
    .B(net249),
    .C(_0443_),
    .Y(_0340_));
 sg13g2_nor3_1 _0867_ (.A(net223),
    .B(_0110_),
    .C(net202),
    .Y(_0341_));
 sg13g2_nor3_1 _0868_ (.A(net215),
    .B(_0043_),
    .C(net208),
    .Y(_0342_));
 sg13g2_a21oi_1 _0869_ (.A1(net215),
    .A2(_0114_),
    .Y(_0343_),
    .B1(_0111_));
 sg13g2_or2_1 _0870_ (.X(_0344_),
    .B(_0332_),
    .A(net230));
 sg13g2_nand4_1 _0871_ (.B(_0336_),
    .C(_0337_),
    .A(_0334_),
    .Y(_0345_),
    .D(_0339_));
 sg13g2_nor4_1 _0872_ (.A(_0424_),
    .B(_0340_),
    .C(_0341_),
    .D(_0342_),
    .Y(_0346_));
 sg13g2_a221oi_1 _0873_ (.B2(net209),
    .C1(_0338_),
    .B1(_0343_),
    .A1(net213),
    .Y(_0347_),
    .A2(_0253_));
 sg13g2_a21oi_1 _0874_ (.A1(_0346_),
    .A2(_0347_),
    .Y(_0348_),
    .B1(net227));
 sg13g2_o21ai_1 _0875_ (.B1(_0348_),
    .Y(_0349_),
    .A1(_0344_),
    .A2(_0345_));
 sg13g2_a21o_1 _0876_ (.A2(_0246_),
    .A1(_0097_),
    .B1(net220),
    .X(_0350_));
 sg13g2_a21oi_1 _0877_ (.A1(net248),
    .A2(net253),
    .Y(_0351_),
    .B1(net242));
 sg13g2_a22oi_1 _0878_ (.Y(_0352_),
    .B1(_0351_),
    .B2(_0446_),
    .A2(_0095_),
    .A1(net242));
 sg13g2_nand2b_1 _0879_ (.Y(_0353_),
    .B(net208),
    .A_N(_0352_));
 sg13g2_nand2b_1 _0880_ (.Y(_0354_),
    .B(net198),
    .A_N(_0195_));
 sg13g2_nand4_1 _0881_ (.B(_0350_),
    .C(_0353_),
    .A(_0334_),
    .Y(_0355_),
    .D(_0354_));
 sg13g2_a22oi_1 _0882_ (.Y(_0356_),
    .B1(net217),
    .B2(_0147_),
    .A2(net219),
    .A1(_0428_));
 sg13g2_or2_1 _0883_ (.X(_0357_),
    .B(_0229_),
    .A(_0455_));
 sg13g2_a21o_1 _0884_ (.A2(_0356_),
    .A1(_0124_),
    .B1(net206),
    .X(_0358_));
 sg13g2_a21o_1 _0885_ (.A2(_0305_),
    .A1(_0304_),
    .B1(_0056_),
    .X(_0359_));
 sg13g2_o21ai_1 _0886_ (.B1(_0435_),
    .Y(_0360_),
    .A1(_0156_),
    .A2(_0319_));
 sg13g2_o21ai_1 _0887_ (.B1(_0431_),
    .Y(_0361_),
    .A1(_0094_),
    .A2(_0096_));
 sg13g2_nand2_1 _0888_ (.Y(_0362_),
    .A(net257),
    .B(_0004_));
 sg13g2_nand3_1 _0889_ (.B(_0129_),
    .C(_0362_),
    .A(net243),
    .Y(_0363_));
 sg13g2_nand3_1 _0890_ (.B(_0361_),
    .C(_0363_),
    .A(net199),
    .Y(_0364_));
 sg13g2_nand4_1 _0891_ (.B(_0359_),
    .C(_0360_),
    .A(_0358_),
    .Y(_0365_),
    .D(_0364_));
 sg13g2_a22oi_1 _0892_ (.Y(_0366_),
    .B1(_0365_),
    .B2(_0058_),
    .A2(_0355_),
    .A1(_0432_));
 sg13g2_a21oi_1 _0893_ (.A1(_0349_),
    .A2(_0366_),
    .Y(_0367_),
    .B1(_0438_));
 sg13g2_o21ai_1 _0894_ (.B1(net222),
    .Y(_0368_),
    .A1(_0223_),
    .A2(_0357_));
 sg13g2_o21ai_1 _0895_ (.B1(net199),
    .Y(_0369_),
    .A1(_0223_),
    .A2(_0272_));
 sg13g2_nand2b_1 _0896_ (.Y(_0370_),
    .B(net219),
    .A_N(_0095_));
 sg13g2_a21oi_1 _0897_ (.A1(_0304_),
    .A2(_0370_),
    .Y(_0371_),
    .B1(_0056_));
 sg13g2_nor3_1 _0898_ (.A(net230),
    .B(_0332_),
    .C(_0371_),
    .Y(_0372_));
 sg13g2_and3_1 _0899_ (.X(_0373_),
    .A(_0368_),
    .B(_0369_),
    .C(_0372_));
 sg13g2_a21oi_1 _0900_ (.A1(net216),
    .A2(_0168_),
    .Y(_0374_),
    .B1(net210));
 sg13g2_a21oi_1 _0901_ (.A1(net217),
    .A2(_0044_),
    .Y(_0375_),
    .B1(_0167_));
 sg13g2_o21ai_1 _0902_ (.B1(net228),
    .Y(_0376_),
    .A1(net206),
    .A2(_0375_));
 sg13g2_a21oi_1 _0903_ (.A1(_0443_),
    .A2(net215),
    .Y(_0377_),
    .B1(_0146_));
 sg13g2_o21ai_1 _0904_ (.B1(net221),
    .Y(_0378_),
    .A1(_0169_),
    .A2(_0377_));
 sg13g2_a21oi_1 _0905_ (.A1(net245),
    .A2(_0044_),
    .Y(_0379_),
    .B1(net239));
 sg13g2_o21ai_1 _0906_ (.B1(net213),
    .Y(_0380_),
    .A1(_0226_),
    .A2(_0379_));
 sg13g2_nand2_1 _0907_ (.Y(_0381_),
    .A(_0378_),
    .B(_0380_));
 sg13g2_nor3_1 _0908_ (.A(_0374_),
    .B(_0376_),
    .C(_0381_),
    .Y(_0382_));
 sg13g2_o21ai_1 _0909_ (.B1(net225),
    .Y(_0383_),
    .A1(_0373_),
    .A2(_0382_));
 sg13g2_o21ai_1 _0910_ (.B1(net199),
    .Y(_0384_),
    .A1(_0240_),
    .A2(_0319_));
 sg13g2_nor2_1 _0911_ (.A(_0044_),
    .B(net206),
    .Y(_0385_));
 sg13g2_a221oi_1 _0912_ (.B2(_0114_),
    .C1(net230),
    .B1(_0385_),
    .A1(net223),
    .Y(_0386_),
    .A2(_0284_));
 sg13g2_o21ai_1 _0913_ (.B1(net221),
    .Y(_0387_),
    .A1(_0302_),
    .A2(_0320_));
 sg13g2_nand3_1 _0914_ (.B(_0386_),
    .C(_0387_),
    .A(_0384_),
    .Y(_0388_));
 sg13g2_o21ai_1 _0915_ (.B1(net234),
    .Y(_0389_),
    .A1(_0229_),
    .A2(_0303_));
 sg13g2_o21ai_1 _0916_ (.B1(_0068_),
    .Y(_0390_),
    .A1(_0130_),
    .A2(_0293_));
 sg13g2_nand3_1 _0917_ (.B(_0044_),
    .C(net211),
    .A(net217),
    .Y(_0391_));
 sg13g2_nand4_1 _0918_ (.B(_0389_),
    .C(_0390_),
    .A(net230),
    .Y(_0392_),
    .D(_0391_));
 sg13g2_a21oi_1 _0919_ (.A1(_0388_),
    .A2(_0392_),
    .Y(_0393_),
    .B1(net227));
 sg13g2_nor3_1 _0920_ (.A(_0421_),
    .B(\pix_y[4] ),
    .C(_0393_),
    .Y(_0394_));
 sg13g2_o21ai_1 _0921_ (.B1(net213),
    .Y(_0395_),
    .A1(_0103_),
    .A2(_0351_));
 sg13g2_nor2_1 _0922_ (.A(net210),
    .B(_0161_),
    .Y(_0396_));
 sg13g2_a221oi_1 _0923_ (.B2(net208),
    .C1(_0396_),
    .B1(_0275_),
    .A1(net222),
    .Y(_0397_),
    .A2(_0267_));
 sg13g2_a21oi_1 _0924_ (.A1(_0395_),
    .A2(_0397_),
    .Y(_0398_),
    .B1(_0433_));
 sg13g2_o21ai_1 _0925_ (.B1(_0274_),
    .Y(_0399_),
    .A1(net220),
    .A2(_0161_));
 sg13g2_nor2_1 _0926_ (.A(net206),
    .B(_0100_),
    .Y(_0400_));
 sg13g2_o21ai_1 _0927_ (.B1(_0400_),
    .Y(_0401_),
    .A1(_0448_),
    .A2(_0044_));
 sg13g2_a21oi_1 _0928_ (.A1(net198),
    .A2(_0151_),
    .Y(_0402_),
    .B1(_0399_));
 sg13g2_a21oi_1 _0929_ (.A1(_0401_),
    .A2(_0402_),
    .Y(_0403_),
    .B1(_0059_));
 sg13g2_nor2_1 _0930_ (.A(net237),
    .B(_0100_),
    .Y(_0404_));
 sg13g2_nor4_1 _0931_ (.A(_0424_),
    .B(net222),
    .C(_0126_),
    .D(_0404_),
    .Y(_0405_));
 sg13g2_o21ai_1 _0932_ (.B1(_0405_),
    .Y(_0406_),
    .A1(_0153_),
    .A2(_0156_));
 sg13g2_nand2_1 _0933_ (.Y(_0407_),
    .A(net204),
    .B(_0259_));
 sg13g2_o21ai_1 _0934_ (.B1(_0100_),
    .Y(_0408_),
    .A1(net222),
    .A2(_0159_));
 sg13g2_a21o_1 _0935_ (.A2(_0408_),
    .A1(_0407_),
    .B1(net228),
    .X(_0409_));
 sg13g2_nand3_1 _0936_ (.B(_0406_),
    .C(_0409_),
    .A(_0425_),
    .Y(_0410_));
 sg13g2_nor4_1 _0937_ (.A(net224),
    .B(_0426_),
    .C(_0398_),
    .D(_0403_),
    .Y(_0411_));
 sg13g2_a221oi_1 _0938_ (.B2(_0411_),
    .C1(_0367_),
    .B1(_0410_),
    .A1(_0383_),
    .Y(_0412_),
    .A2(_0394_));
 sg13g2_a21oi_1 _0939_ (.A1(_0420_),
    .A2(_0412_),
    .Y(_0413_),
    .B1(_0331_));
 sg13g2_nand2_1 _0940_ (.Y(_0414_),
    .A(_0439_),
    .B(net79));
 sg13g2_nor4_2 _0941_ (.A(net74),
    .B(net67),
    .C(_0427_),
    .Y(_0415_),
    .D(_0414_));
 sg13g2_nand2_1 _0942_ (.Y(_0416_),
    .A(_0219_),
    .B(_0415_));
 sg13g2_inv_1 _0943_ (.Y(_0034_),
    .A(_0416_));
 sg13g2_nand2_1 _0944_ (.Y(_0417_),
    .A(_0413_),
    .B(_0415_));
 sg13g2_inv_1 _0945_ (.Y(_0033_),
    .A(_0417_));
 sg13g2_a22oi_1 _0946_ (.Y(_0032_),
    .B1(_0416_),
    .B2(_0417_),
    .A2(_0413_),
    .A1(_0219_));
 sg13g2_nor2_1 _0947_ (.A(_0219_),
    .B(_0417_),
    .Y(_0035_));
 sg13g2_a21oi_1 _0948_ (.A1(net53),
    .A2(_0412_),
    .Y(_0418_),
    .B1(_0331_));
 sg13g2_nor2_1 _0949_ (.A(_0416_),
    .B(net54),
    .Y(_0036_));
 sg13g2_dfrbp_1 _0950_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net28),
    .D(_0012_),
    .Q_N(_0011_),
    .Q(\pix_x[0] ));
 sg13g2_dfrbp_1 _0951_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net42),
    .D(net50),
    .Q_N(_0472_),
    .Q(\pix_x[1] ));
 sg13g2_dfrbp_1 _0952_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net41),
    .D(net52),
    .Q_N(_0471_),
    .Q(\pix_x[2] ));
 sg13g2_dfrbp_1 _0953_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net40),
    .D(_0015_),
    .Q_N(_0003_),
    .Q(\pix_x[3] ));
 sg13g2_dfrbp_1 _0954_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net38),
    .D(_0016_),
    .Q_N(_0004_),
    .Q(\pix_x[4] ));
 sg13g2_dfrbp_1 _0955_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net37),
    .D(_0017_),
    .Q_N(_0008_),
    .Q(\pix_x[5] ));
 sg13g2_dfrbp_1 _0956_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net36),
    .D(_0018_),
    .Q_N(_0009_),
    .Q(\pix_x[6] ));
 sg13g2_dfrbp_1 _0957_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net35),
    .D(_0019_),
    .Q_N(_0470_),
    .Q(\pix_x[7] ));
 sg13g2_dfrbp_1 _0958_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net34),
    .D(net60),
    .Q_N(_0469_),
    .Q(\pix_x[8] ));
 sg13g2_dfrbp_1 _0959_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net39),
    .D(_0021_),
    .Q_N(_0473_),
    .Q(\pix_x[9] ));
 sg13g2_dfrbp_1 _0960_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net33),
    .D(_0000_),
    .Q_N(_0468_),
    .Q(hsync));
 sg13g2_dfrbp_1 _0961_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net32),
    .D(_0022_),
    .Q_N(_0010_),
    .Q(\pix_y[0] ));
 sg13g2_dfrbp_1 _0962_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net30),
    .D(_0023_),
    .Q_N(_0467_),
    .Q(\pix_y[1] ));
 sg13g2_dfrbp_1 _0963_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net27),
    .D(_0024_),
    .Q_N(_0007_),
    .Q(\pix_y[2] ));
 sg13g2_dfrbp_1 _0964_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net25),
    .D(_0025_),
    .Q_N(_0466_),
    .Q(\pix_y[3] ));
 sg13g2_dfrbp_1 _0965_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net23),
    .D(_0026_),
    .Q_N(_0002_),
    .Q(\pix_y[4] ));
 sg13g2_dfrbp_1 _0966_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net21),
    .D(net73),
    .Q_N(_0005_),
    .Q(\pix_y[5] ));
 sg13g2_dfrbp_1 _0967_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net19),
    .D(_0028_),
    .Q_N(_0006_),
    .Q(\pix_y[6] ));
 sg13g2_dfrbp_1 _0968_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net44),
    .D(_0029_),
    .Q_N(_0465_),
    .Q(\pix_y[7] ));
 sg13g2_dfrbp_1 _0969_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net31),
    .D(net68),
    .Q_N(_0464_),
    .Q(\pix_y[8] ));
 sg13g2_dfrbp_1 _0970_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net24),
    .D(_0031_),
    .Q_N(_0474_),
    .Q(\pix_y[9] ));
 sg13g2_dfrbp_1 _0971_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net26),
    .D(net47),
    .Q_N(_0463_),
    .Q(\vga_sync_gen.vsync ));
 sg13g2_dfrbp_1 _0972_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net22),
    .D(_0032_),
    .Q_N(_0462_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _0973_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net20),
    .D(_0033_),
    .Q_N(_0461_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _0974_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net18),
    .D(_0034_),
    .Q_N(_0460_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _0975_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net43),
    .D(_0035_),
    .Q_N(_0459_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _0976_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net29),
    .D(net55),
    .Q_N(_0458_),
    .Q(uo_out[5]));
 sg13g2_tiehi _0967__19 (.L_HI(net19));
 sg13g2_tiehi _0973__20 (.L_HI(net20));
 sg13g2_tiehi _0966__21 (.L_HI(net21));
 sg13g2_tiehi _0972__22 (.L_HI(net22));
 sg13g2_tiehi _0965__23 (.L_HI(net23));
 sg13g2_tiehi _0970__24 (.L_HI(net24));
 sg13g2_tiehi _0964__25 (.L_HI(net25));
 sg13g2_tiehi _0971__26 (.L_HI(net26));
 sg13g2_tiehi _0963__27 (.L_HI(net27));
 sg13g2_tiehi _0950__28 (.L_HI(net28));
 sg13g2_tiehi _0976__29 (.L_HI(net29));
 sg13g2_tiehi _0962__30 (.L_HI(net30));
 sg13g2_tiehi _0969__31 (.L_HI(net31));
 sg13g2_tiehi _0961__32 (.L_HI(net32));
 sg13g2_tiehi _0960__33 (.L_HI(net33));
 sg13g2_tiehi _0958__34 (.L_HI(net34));
 sg13g2_tiehi _0957__35 (.L_HI(net35));
 sg13g2_tiehi _0956__36 (.L_HI(net36));
 sg13g2_tiehi _0955__37 (.L_HI(net37));
 sg13g2_tiehi _0954__38 (.L_HI(net38));
 sg13g2_tiehi _0959__39 (.L_HI(net39));
 sg13g2_tiehi _0953__40 (.L_HI(net40));
 sg13g2_tiehi _0952__41 (.L_HI(net41));
 sg13g2_tiehi _0951__42 (.L_HI(net42));
 sg13g2_tiehi _0975__43 (.L_HI(net43));
 sg13g2_tiehi _0968__44 (.L_HI(net44));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_vga_cbtest_3 (.L_LO(net3));
 sg13g2_tielo tt_um_vga_cbtest_4 (.L_LO(net4));
 sg13g2_tielo tt_um_vga_cbtest_5 (.L_LO(net5));
 sg13g2_tielo tt_um_vga_cbtest_6 (.L_LO(net6));
 sg13g2_tielo tt_um_vga_cbtest_7 (.L_LO(net7));
 sg13g2_tielo tt_um_vga_cbtest_8 (.L_LO(net8));
 sg13g2_tielo tt_um_vga_cbtest_9 (.L_LO(net9));
 sg13g2_tielo tt_um_vga_cbtest_10 (.L_LO(net10));
 sg13g2_tielo tt_um_vga_cbtest_11 (.L_LO(net11));
 sg13g2_tielo tt_um_vga_cbtest_12 (.L_LO(net12));
 sg13g2_tielo tt_um_vga_cbtest_13 (.L_LO(net13));
 sg13g2_tielo tt_um_vga_cbtest_14 (.L_LO(net14));
 sg13g2_tielo tt_um_vga_cbtest_15 (.L_LO(net15));
 sg13g2_tielo tt_um_vga_cbtest_16 (.L_LO(net16));
 sg13g2_tielo tt_um_vga_cbtest_17 (.L_LO(net17));
 sg13g2_tiehi _0974__18 (.L_HI(net18));
 sg13g2_buf_1 _1020_ (.A(uo_out[4]),
    .X(uo_out[0]));
 sg13g2_buf_1 _1021_ (.A(\vga_sync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1022_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout197 (.X(net197),
    .A(_0037_));
 sg13g2_buf_4 fanout198 (.X(net198),
    .A(_0066_));
 sg13g2_buf_2 fanout199 (.A(_0066_),
    .X(net199));
 sg13g2_buf_4 fanout200 (.X(net200),
    .A(_0145_));
 sg13g2_buf_1 fanout201 (.A(_0145_),
    .X(net201));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(_0131_));
 sg13g2_buf_4 fanout203 (.X(net203),
    .A(_0111_));
 sg13g2_buf_2 fanout204 (.A(_0110_),
    .X(net204));
 sg13g2_buf_4 fanout205 (.X(net205),
    .A(_0094_));
 sg13g2_buf_2 fanout206 (.A(_0072_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_0072_),
    .X(net207));
 sg13g2_buf_4 fanout208 (.X(net208),
    .A(_0071_));
 sg13g2_buf_2 fanout209 (.A(_0071_),
    .X(net209));
 sg13g2_buf_4 fanout210 (.X(net210),
    .A(_0067_));
 sg13g2_buf_2 fanout211 (.A(net213),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(net213),
    .X(net212));
 sg13g2_buf_4 fanout213 (.X(net213),
    .A(_0055_));
 sg13g2_buf_4 fanout214 (.X(net214),
    .A(_0447_));
 sg13g2_buf_2 fanout215 (.A(_0445_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_0445_),
    .X(net216));
 sg13g2_buf_4 fanout217 (.X(net217),
    .A(_0444_));
 sg13g2_buf_2 fanout218 (.A(_0444_),
    .X(net218));
 sg13g2_buf_4 fanout219 (.X(net219),
    .A(_0442_));
 sg13g2_buf_4 fanout220 (.X(net220),
    .A(_0436_));
 sg13g2_buf_4 fanout221 (.X(net221),
    .A(net222));
 sg13g2_buf_4 fanout222 (.X(net222),
    .A(_0435_));
 sg13g2_buf_4 fanout223 (.X(net223),
    .A(_0422_));
 sg13g2_buf_2 fanout224 (.A(\pix_y[5] ),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(net227),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(net227),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(\pix_y[3] ),
    .X(net227));
 sg13g2_buf_4 fanout228 (.X(net228),
    .A(net231));
 sg13g2_buf_2 fanout229 (.A(net231),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(net231),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(net80),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(net235),
    .X(net232));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(net235));
 sg13g2_buf_2 fanout234 (.A(net235),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(\pix_y[1] ),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(net238),
    .X(net236));
 sg13g2_buf_1 fanout237 (.A(net238),
    .X(net237));
 sg13g2_buf_4 fanout238 (.X(net238),
    .A(\pix_y[0] ));
 sg13g2_buf_2 fanout239 (.A(net244),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net243),
    .X(net240));
 sg13g2_buf_1 fanout241 (.A(net243),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(net243),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(net244),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(\pix_x[6] ),
    .X(net244));
 sg13g2_buf_4 fanout245 (.X(net245),
    .A(_0008_));
 sg13g2_buf_2 fanout246 (.A(_0008_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(net248),
    .X(net247));
 sg13g2_buf_1 fanout248 (.A(net250),
    .X(net248));
 sg13g2_buf_4 fanout249 (.X(net249),
    .A(net250));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(\pix_x[5] ));
 sg13g2_buf_2 fanout251 (.A(net254),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(net253),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(net254),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(\pix_x[4] ),
    .X(net254));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(net256));
 sg13g2_buf_2 fanout256 (.A(\pix_x[3] ),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(net258),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(\pix_x[3] ),
    .X(net258));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_tielo tt_um_vga_cbtest_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0011_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0005_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0001_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold4 (.A(\pix_x[1] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0039_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0013_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold7 (.A(\pix_x[2] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0014_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0006_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0418_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0036_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0010_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0065_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold14 (.A(\pix_x[8] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0051_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0020_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold17 (.A(\pix_y[9] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0093_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold19 (.A(\pix_x[7] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0452_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0009_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold22 (.A(\pix_x[0] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold23 (.A(\pix_y[8] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0030_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold25 (.A(\pix_y[7] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0007_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0004_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0002_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0027_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold30 (.A(\pix_x[9] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold31 (.A(\pix_y[6] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0084_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold33 (.A(\pix_y[4] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold34 (.A(\pix_x[7] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0456_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold36 (.A(\pix_y[2] ),
    .X(net80));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_4 FILLER_16_280 ();
 sg13g2_fill_1 FILLER_16_284 ();
 sg13g2_decap_8 FILLER_16_290 ();
 sg13g2_decap_8 FILLER_16_297 ();
 sg13g2_decap_8 FILLER_16_304 ();
 sg13g2_decap_8 FILLER_16_311 ();
 sg13g2_decap_8 FILLER_16_318 ();
 sg13g2_decap_8 FILLER_16_325 ();
 sg13g2_decap_8 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_4 FILLER_17_224 ();
 sg13g2_decap_4 FILLER_17_235 ();
 sg13g2_fill_2 FILLER_17_239 ();
 sg13g2_fill_2 FILLER_17_245 ();
 sg13g2_decap_4 FILLER_17_251 ();
 sg13g2_fill_1 FILLER_17_255 ();
 sg13g2_decap_8 FILLER_17_263 ();
 sg13g2_decap_8 FILLER_17_270 ();
 sg13g2_fill_2 FILLER_17_277 ();
 sg13g2_fill_1 FILLER_17_279 ();
 sg13g2_decap_8 FILLER_17_296 ();
 sg13g2_fill_2 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_317 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_331 ();
 sg13g2_decap_8 FILLER_17_338 ();
 sg13g2_decap_8 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_4 FILLER_18_196 ();
 sg13g2_fill_1 FILLER_18_200 ();
 sg13g2_fill_1 FILLER_18_206 ();
 sg13g2_decap_4 FILLER_18_211 ();
 sg13g2_fill_2 FILLER_18_215 ();
 sg13g2_fill_1 FILLER_18_243 ();
 sg13g2_fill_1 FILLER_18_248 ();
 sg13g2_fill_2 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_266 ();
 sg13g2_decap_4 FILLER_18_272 ();
 sg13g2_fill_1 FILLER_18_276 ();
 sg13g2_decap_4 FILLER_18_292 ();
 sg13g2_fill_2 FILLER_18_296 ();
 sg13g2_fill_2 FILLER_18_317 ();
 sg13g2_fill_1 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_4 FILLER_19_161 ();
 sg13g2_fill_1 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_198 ();
 sg13g2_decap_8 FILLER_19_227 ();
 sg13g2_fill_1 FILLER_19_234 ();
 sg13g2_decap_8 FILLER_19_256 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_fill_2 FILLER_19_288 ();
 sg13g2_fill_1 FILLER_19_290 ();
 sg13g2_fill_2 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_303 ();
 sg13g2_fill_2 FILLER_19_309 ();
 sg13g2_decap_4 FILLER_19_331 ();
 sg13g2_fill_1 FILLER_19_335 ();
 sg13g2_fill_1 FILLER_19_341 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_fill_2 FILLER_20_179 ();
 sg13g2_decap_4 FILLER_20_191 ();
 sg13g2_fill_1 FILLER_20_195 ();
 sg13g2_fill_1 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_207 ();
 sg13g2_fill_1 FILLER_20_209 ();
 sg13g2_decap_4 FILLER_20_214 ();
 sg13g2_fill_1 FILLER_20_218 ();
 sg13g2_decap_4 FILLER_20_224 ();
 sg13g2_fill_2 FILLER_20_228 ();
 sg13g2_fill_2 FILLER_20_234 ();
 sg13g2_fill_1 FILLER_20_236 ();
 sg13g2_fill_2 FILLER_20_266 ();
 sg13g2_fill_1 FILLER_20_268 ();
 sg13g2_decap_4 FILLER_20_279 ();
 sg13g2_decap_4 FILLER_20_289 ();
 sg13g2_decap_4 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_fill_1 FILLER_21_177 ();
 sg13g2_fill_2 FILLER_21_186 ();
 sg13g2_fill_1 FILLER_21_188 ();
 sg13g2_fill_2 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_226 ();
 sg13g2_fill_1 FILLER_21_233 ();
 sg13g2_decap_4 FILLER_21_253 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_fill_2 FILLER_21_300 ();
 sg13g2_fill_1 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_fill_2 FILLER_21_336 ();
 sg13g2_fill_1 FILLER_21_338 ();
 sg13g2_fill_2 FILLER_21_344 ();
 sg13g2_fill_1 FILLER_21_346 ();
 sg13g2_decap_4 FILLER_21_358 ();
 sg13g2_fill_2 FILLER_21_362 ();
 sg13g2_fill_2 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_fill_1 FILLER_22_154 ();
 sg13g2_fill_1 FILLER_22_182 ();
 sg13g2_fill_2 FILLER_22_188 ();
 sg13g2_fill_2 FILLER_22_195 ();
 sg13g2_fill_1 FILLER_22_197 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_4 FILLER_22_210 ();
 sg13g2_fill_1 FILLER_22_214 ();
 sg13g2_decap_4 FILLER_22_225 ();
 sg13g2_fill_2 FILLER_22_229 ();
 sg13g2_fill_1 FILLER_22_260 ();
 sg13g2_decap_4 FILLER_22_275 ();
 sg13g2_fill_1 FILLER_22_279 ();
 sg13g2_decap_8 FILLER_22_306 ();
 sg13g2_fill_2 FILLER_22_313 ();
 sg13g2_fill_1 FILLER_22_315 ();
 sg13g2_decap_4 FILLER_22_329 ();
 sg13g2_fill_1 FILLER_22_333 ();
 sg13g2_decap_4 FILLER_22_339 ();
 sg13g2_fill_2 FILLER_22_352 ();
 sg13g2_fill_1 FILLER_22_354 ();
 sg13g2_fill_2 FILLER_22_367 ();
 sg13g2_fill_1 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_388 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_4 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_194 ();
 sg13g2_fill_2 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_213 ();
 sg13g2_fill_2 FILLER_23_221 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_230 ();
 sg13g2_fill_2 FILLER_23_250 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_fill_1 FILLER_23_282 ();
 sg13g2_decap_8 FILLER_23_304 ();
 sg13g2_fill_1 FILLER_23_311 ();
 sg13g2_fill_2 FILLER_23_317 ();
 sg13g2_decap_4 FILLER_23_324 ();
 sg13g2_fill_2 FILLER_23_341 ();
 sg13g2_fill_1 FILLER_23_343 ();
 sg13g2_fill_2 FILLER_23_359 ();
 sg13g2_fill_1 FILLER_23_361 ();
 sg13g2_fill_2 FILLER_23_372 ();
 sg13g2_fill_1 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_4 FILLER_24_161 ();
 sg13g2_fill_1 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_193 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_4 FILLER_24_245 ();
 sg13g2_fill_2 FILLER_24_249 ();
 sg13g2_decap_4 FILLER_24_256 ();
 sg13g2_fill_2 FILLER_24_266 ();
 sg13g2_fill_1 FILLER_24_268 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_fill_2 FILLER_24_280 ();
 sg13g2_fill_1 FILLER_24_282 ();
 sg13g2_fill_2 FILLER_24_300 ();
 sg13g2_fill_1 FILLER_24_327 ();
 sg13g2_fill_2 FILLER_24_365 ();
 sg13g2_fill_1 FILLER_24_367 ();
 sg13g2_fill_1 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_4 FILLER_25_154 ();
 sg13g2_fill_1 FILLER_25_158 ();
 sg13g2_decap_4 FILLER_25_167 ();
 sg13g2_decap_4 FILLER_25_190 ();
 sg13g2_fill_1 FILLER_25_209 ();
 sg13g2_decap_8 FILLER_25_216 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_fill_2 FILLER_25_230 ();
 sg13g2_decap_4 FILLER_25_238 ();
 sg13g2_fill_2 FILLER_25_255 ();
 sg13g2_fill_1 FILLER_25_257 ();
 sg13g2_fill_2 FILLER_25_264 ();
 sg13g2_fill_1 FILLER_25_288 ();
 sg13g2_fill_2 FILLER_25_294 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_fill_2 FILLER_25_311 ();
 sg13g2_fill_1 FILLER_25_330 ();
 sg13g2_fill_2 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_344 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_fill_1 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_decap_4 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_decap_4 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_260 ();
 sg13g2_decap_8 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_278 ();
 sg13g2_fill_2 FILLER_26_284 ();
 sg13g2_fill_1 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_fill_2 FILLER_26_319 ();
 sg13g2_decap_4 FILLER_26_326 ();
 sg13g2_decap_4 FILLER_26_334 ();
 sg13g2_fill_2 FILLER_26_338 ();
 sg13g2_decap_4 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_154 ();
 sg13g2_fill_2 FILLER_27_180 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_decap_4 FILLER_27_192 ();
 sg13g2_fill_2 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_fill_2 FILLER_27_217 ();
 sg13g2_fill_2 FILLER_27_224 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_fill_2 FILLER_27_254 ();
 sg13g2_fill_1 FILLER_27_256 ();
 sg13g2_fill_1 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_fill_1 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_297 ();
 sg13g2_fill_2 FILLER_27_304 ();
 sg13g2_fill_1 FILLER_27_306 ();
 sg13g2_fill_2 FILLER_27_345 ();
 sg13g2_fill_2 FILLER_27_352 ();
 sg13g2_fill_1 FILLER_27_354 ();
 sg13g2_fill_2 FILLER_27_360 ();
 sg13g2_fill_1 FILLER_27_362 ();
 sg13g2_decap_8 FILLER_27_369 ();
 sg13g2_fill_1 FILLER_27_376 ();
 sg13g2_fill_2 FILLER_27_387 ();
 sg13g2_fill_1 FILLER_27_389 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_4 FILLER_28_154 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_decap_4 FILLER_28_173 ();
 sg13g2_fill_2 FILLER_28_183 ();
 sg13g2_fill_1 FILLER_28_185 ();
 sg13g2_decap_4 FILLER_28_198 ();
 sg13g2_fill_1 FILLER_28_217 ();
 sg13g2_fill_1 FILLER_28_231 ();
 sg13g2_decap_4 FILLER_28_247 ();
 sg13g2_fill_2 FILLER_28_269 ();
 sg13g2_fill_1 FILLER_28_271 ();
 sg13g2_fill_1 FILLER_28_278 ();
 sg13g2_fill_2 FILLER_28_290 ();
 sg13g2_fill_1 FILLER_28_292 ();
 sg13g2_fill_2 FILLER_28_307 ();
 sg13g2_fill_2 FILLER_28_321 ();
 sg13g2_fill_1 FILLER_28_333 ();
 sg13g2_decap_8 FILLER_28_346 ();
 sg13g2_fill_2 FILLER_28_353 ();
 sg13g2_decap_8 FILLER_28_370 ();
 sg13g2_fill_1 FILLER_28_377 ();
 sg13g2_decap_4 FILLER_28_383 ();
 sg13g2_fill_2 FILLER_28_387 ();
 sg13g2_decap_4 FILLER_28_393 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_154 ();
 sg13g2_fill_1 FILLER_29_172 ();
 sg13g2_fill_2 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_191 ();
 sg13g2_decap_8 FILLER_29_202 ();
 sg13g2_decap_8 FILLER_29_209 ();
 sg13g2_fill_1 FILLER_29_216 ();
 sg13g2_decap_8 FILLER_29_230 ();
 sg13g2_decap_8 FILLER_29_237 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_fill_2 FILLER_29_277 ();
 sg13g2_decap_4 FILLER_29_291 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_decap_8 FILLER_29_312 ();
 sg13g2_decap_4 FILLER_29_319 ();
 sg13g2_decap_4 FILLER_29_328 ();
 sg13g2_fill_1 FILLER_29_332 ();
 sg13g2_decap_4 FILLER_29_337 ();
 sg13g2_fill_1 FILLER_29_348 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_4 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_decap_8 FILLER_30_156 ();
 sg13g2_fill_1 FILLER_30_168 ();
 sg13g2_fill_2 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_176 ();
 sg13g2_fill_2 FILLER_30_182 ();
 sg13g2_fill_2 FILLER_30_233 ();
 sg13g2_fill_1 FILLER_30_235 ();
 sg13g2_decap_4 FILLER_30_265 ();
 sg13g2_fill_1 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_2 FILLER_30_380 ();
 sg13g2_decap_8 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_decap_4 FILLER_31_211 ();
 sg13g2_fill_1 FILLER_31_215 ();
 sg13g2_fill_1 FILLER_31_231 ();
 sg13g2_decap_4 FILLER_31_237 ();
 sg13g2_decap_8 FILLER_31_251 ();
 sg13g2_decap_4 FILLER_31_258 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_4 FILLER_31_273 ();
 sg13g2_fill_1 FILLER_31_308 ();
 sg13g2_decap_4 FILLER_31_317 ();
 sg13g2_fill_2 FILLER_31_321 ();
 sg13g2_fill_2 FILLER_31_342 ();
 sg13g2_fill_1 FILLER_31_361 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_4 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_188 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_decap_4 FILLER_32_314 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_fill_2 FILLER_32_333 ();
 sg13g2_fill_1 FILLER_32_335 ();
 sg13g2_decap_8 FILLER_32_398 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_fill_1 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_152 ();
 sg13g2_decap_4 FILLER_33_159 ();
 sg13g2_decap_8 FILLER_33_235 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_fill_2 FILLER_33_251 ();
 sg13g2_decap_8 FILLER_33_258 ();
 sg13g2_fill_2 FILLER_33_265 ();
 sg13g2_fill_2 FILLER_33_282 ();
 sg13g2_fill_2 FILLER_33_307 ();
 sg13g2_fill_1 FILLER_33_321 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_fill_1 FILLER_34_161 ();
 sg13g2_fill_2 FILLER_34_183 ();
 sg13g2_fill_1 FILLER_34_264 ();
 sg13g2_fill_2 FILLER_34_304 ();
 sg13g2_decap_4 FILLER_34_313 ();
 sg13g2_fill_2 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_fill_2 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_182 ();
 sg13g2_fill_1 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_208 ();
 sg13g2_fill_1 FILLER_35_226 ();
 sg13g2_fill_2 FILLER_35_253 ();
 sg13g2_decap_4 FILLER_35_259 ();
 sg13g2_fill_2 FILLER_35_263 ();
 sg13g2_fill_2 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_273 ();
 sg13g2_fill_2 FILLER_35_352 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_decap_8 FILLER_36_171 ();
 sg13g2_fill_1 FILLER_36_178 ();
 sg13g2_fill_2 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_266 ();
 sg13g2_fill_2 FILLER_36_290 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_fill_2 FILLER_36_326 ();
 sg13g2_fill_2 FILLER_36_337 ();
 sg13g2_fill_2 FILLER_36_362 ();
 sg13g2_fill_1 FILLER_36_364 ();
 sg13g2_fill_2 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_fill_1 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_202 ();
 sg13g2_fill_1 FILLER_37_212 ();
 sg13g2_fill_2 FILLER_37_239 ();
 sg13g2_fill_2 FILLER_37_249 ();
 sg13g2_fill_1 FILLER_37_251 ();
 sg13g2_decap_8 FILLER_37_307 ();
 sg13g2_decap_8 FILLER_37_356 ();
 sg13g2_fill_2 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_369 ();
 sg13g2_decap_8 FILLER_37_376 ();
 sg13g2_decap_8 FILLER_37_383 ();
 sg13g2_decap_8 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_fill_2 FILLER_38_220 ();
 sg13g2_fill_1 FILLER_38_222 ();
 sg13g2_decap_4 FILLER_38_227 ();
 sg13g2_fill_2 FILLER_38_231 ();
 sg13g2_decap_4 FILLER_38_267 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_decap_4 FILLER_38_277 ();
 sg13g2_fill_2 FILLER_38_281 ();
 sg13g2_decap_8 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_fill_2 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_326 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_352 ();
 sg13g2_decap_8 FILLER_38_359 ();
 sg13g2_decap_8 FILLER_38_366 ();
 sg13g2_fill_2 FILLER_38_373 ();
 sg13g2_fill_1 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
endmodule

module tt_um_ephrenm_tsal (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire \top_instance.adc_data[0] ;
 wire \top_instance.adc_data[10] ;
 wire \top_instance.adc_data[11] ;
 wire \top_instance.adc_data[1] ;
 wire \top_instance.adc_data[2] ;
 wire \top_instance.adc_data[3] ;
 wire \top_instance.adc_data[4] ;
 wire \top_instance.adc_data[5] ;
 wire \top_instance.adc_data[6] ;
 wire \top_instance.adc_data[7] ;
 wire \top_instance.adc_data[8] ;
 wire \top_instance.adc_data[9] ;
 wire \top_instance.adc_inst.bit_counter[0] ;
 wire \top_instance.adc_inst.bit_counter[1] ;
 wire \top_instance.adc_inst.bit_counter[2] ;
 wire \top_instance.adc_inst.bit_counter[3] ;
 wire \top_instance.adc_inst.bit_counter[4] ;
 wire \top_instance.adc_inst.bit_counter[5] ;
 wire \top_instance.adc_inst.clk_counter[0] ;
 wire \top_instance.adc_inst.clk_counter[1] ;
 wire \top_instance.adc_inst.clk_counter[2] ;
 wire \top_instance.adc_inst.clk_counter[3] ;
 wire \top_instance.adc_inst.clk_counter[4] ;
 wire \top_instance.adc_inst.clk_counter[5] ;
 wire \top_instance.adc_inst.clk_counter[6] ;
 wire \top_instance.adc_inst.clk_counter[7] ;
 wire \top_instance.adc_inst.clk_counter[8] ;
 wire \top_instance.adc_inst.clk_counter[9] ;
 wire \top_instance.adc_inst.cs ;
 wire \top_instance.adc_inst.data_in_reg ;
 wire \top_instance.adc_inst.data_ready ;
 wire \top_instance.adc_inst.sclk ;
 wire \top_instance.comparator_inst.comp_reg[0] ;
 wire \top_instance.comparator_inst.comp_reg[1] ;
 wire \top_instance.comparator_inst.comp_reg[2] ;
 wire \top_instance.comparator_inst.comp_reg[3] ;
 wire \top_instance.comparator_inst.comp_reg[4] ;
 wire \top_instance.comparator_inst.comp_reg[5] ;
 wire \top_instance.comparator_inst.comp_reg[6] ;
 wire \top_instance.comparator_inst.comp_reg[7] ;
 wire \top_instance.comparator_inst.green_enable ;
 wire \top_instance.comparator_inst.in[0] ;
 wire \top_instance.comparator_inst.in[1] ;
 wire \top_instance.comparator_inst.in[2] ;
 wire \top_instance.comparator_inst.in[3] ;
 wire \top_instance.comparator_inst.in[4] ;
 wire \top_instance.comparator_inst.in[5] ;
 wire \top_instance.comparator_inst.in[6] ;
 wire \top_instance.comparator_inst.in[7] ;
 wire \top_instance.comparator_inst.input_reg[0] ;
 wire \top_instance.comparator_inst.input_reg[1] ;
 wire \top_instance.comparator_inst.input_reg[2] ;
 wire \top_instance.comparator_inst.input_reg[3] ;
 wire \top_instance.comparator_inst.input_reg[4] ;
 wire \top_instance.comparator_inst.input_reg[5] ;
 wire \top_instance.comparator_inst.input_reg[6] ;
 wire \top_instance.comparator_inst.input_reg[7] ;
 wire \top_instance.comparator_inst.red_enable ;
 wire \top_instance.green_led ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[0] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[10] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[11] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[12] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[13] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[14] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[15] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[16] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[17] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[18] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[19] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[1] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[20] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[21] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[22] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[23] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[2] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[3] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[4] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[5] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[6] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[7] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[8] ;
 wire \top_instance.pulse_generator_inst.red_ctrl_counter[9] ;
 wire \top_instance.pulse_generator_inst.red_led ;
 wire net131;
 wire net11;
 wire net12;
 wire clknet_0_clk;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;

 sg13g2_inv_1 _418_ (.Y(_082_),
    .A(net233));
 sg13g2_inv_1 _419_ (.Y(_083_),
    .A(net141));
 sg13g2_inv_1 _420_ (.Y(_084_),
    .A(\top_instance.comparator_inst.input_reg[6] ));
 sg13g2_inv_1 _421_ (.Y(_085_),
    .A(net145));
 sg13g2_inv_1 _422_ (.Y(_086_),
    .A(\top_instance.comparator_inst.input_reg[5] ));
 sg13g2_inv_1 _423_ (.Y(_087_),
    .A(net137));
 sg13g2_inv_1 _424_ (.Y(_088_),
    .A(\top_instance.comparator_inst.input_reg[4] ));
 sg13g2_inv_1 _425_ (.Y(_089_),
    .A(net143));
 sg13g2_inv_1 _426_ (.Y(_090_),
    .A(net149));
 sg13g2_inv_1 _427_ (.Y(_091_),
    .A(\top_instance.comparator_inst.input_reg[2] ));
 sg13g2_inv_1 _428_ (.Y(_092_),
    .A(net139));
 sg13g2_inv_1 _429_ (.Y(_093_),
    .A(net133));
 sg13g2_inv_1 _430_ (.Y(_094_),
    .A(net135));
 sg13g2_inv_1 _431_ (.Y(_095_),
    .A(net170));
 sg13g2_inv_1 _432_ (.Y(_096_),
    .A(net167));
 sg13g2_inv_1 _433_ (.Y(_097_),
    .A(\top_instance.pulse_generator_inst.red_ctrl_counter[15] ));
 sg13g2_inv_2 _434_ (.Y(_098_),
    .A(net243));
 sg13g2_inv_1 _435_ (.Y(_099_),
    .A(net227));
 sg13g2_inv_1 _436_ (.Y(_100_),
    .A(net153));
 sg13g2_inv_1 _437_ (.Y(_101_),
    .A(net237));
 sg13g2_inv_1 _438_ (.Y(_102_),
    .A(net57));
 sg13g2_inv_1 _439_ (.Y(_103_),
    .A(\top_instance.adc_data[11] ));
 sg13g2_inv_1 _440_ (.Y(_104_),
    .A(\top_instance.adc_data[10] ));
 sg13g2_inv_1 _441_ (.Y(_105_),
    .A(\top_instance.comparator_inst.comp_reg[5] ));
 sg13g2_inv_1 _442_ (.Y(_106_),
    .A(\top_instance.adc_data[9] ));
 sg13g2_inv_1 _443_ (.Y(_107_),
    .A(\top_instance.adc_data[8] ));
 sg13g2_inv_1 _444_ (.Y(_108_),
    .A(\top_instance.adc_data[7] ));
 sg13g2_inv_1 _445_ (.Y(_109_),
    .A(\top_instance.adc_data[6] ));
 sg13g2_inv_1 _446_ (.Y(_110_),
    .A(\top_instance.adc_data[5] ));
 sg13g2_inv_1 _447_ (.Y(_111_),
    .A(\top_instance.adc_data[4] ));
 sg13g2_inv_1 _448_ (.Y(_112_),
    .A(net67));
 sg13g2_inv_1 _449_ (.Y(_113_),
    .A(_006_));
 sg13g2_nand2b_1 _450_ (.Y(_114_),
    .B(\top_instance.comparator_inst.comp_reg[3] ),
    .A_N(\top_instance.comparator_inst.input_reg[3] ));
 sg13g2_nand2b_1 _451_ (.Y(_115_),
    .B(\top_instance.comparator_inst.input_reg[1] ),
    .A_N(\top_instance.comparator_inst.comp_reg[1] ));
 sg13g2_nand2b_1 _452_ (.Y(_116_),
    .B(\top_instance.comparator_inst.input_reg[0] ),
    .A_N(\top_instance.comparator_inst.comp_reg[0] ));
 sg13g2_nor2b_1 _453_ (.A(\top_instance.comparator_inst.input_reg[1] ),
    .B_N(\top_instance.comparator_inst.comp_reg[1] ),
    .Y(_117_));
 sg13g2_a221oi_1 _454_ (.B2(_116_),
    .C1(_117_),
    .B1(_115_),
    .A1(_091_),
    .Y(_118_),
    .A2(\top_instance.comparator_inst.comp_reg[2] ));
 sg13g2_nand2b_1 _455_ (.Y(_119_),
    .B(\top_instance.comparator_inst.input_reg[3] ),
    .A_N(\top_instance.comparator_inst.comp_reg[3] ));
 sg13g2_o21ai_1 _456_ (.B1(_119_),
    .Y(_120_),
    .A1(_091_),
    .A2(\top_instance.comparator_inst.comp_reg[2] ));
 sg13g2_o21ai_1 _457_ (.B1(_114_),
    .Y(_121_),
    .A1(_118_),
    .A2(_120_));
 sg13g2_o21ai_1 _458_ (.B1(_121_),
    .Y(_122_),
    .A1(_088_),
    .A2(\top_instance.comparator_inst.comp_reg[4] ));
 sg13g2_a22oi_1 _459_ (.Y(_123_),
    .B1(\top_instance.comparator_inst.comp_reg[4] ),
    .B2(_088_),
    .A2(\top_instance.comparator_inst.comp_reg[5] ),
    .A1(_086_));
 sg13g2_a22oi_1 _460_ (.Y(_124_),
    .B1(_122_),
    .B2(_123_),
    .A2(_105_),
    .A1(\top_instance.comparator_inst.input_reg[5] ));
 sg13g2_a21oi_1 _461_ (.A1(_084_),
    .A2(net203),
    .Y(_125_),
    .B1(_124_));
 sg13g2_nand2b_1 _462_ (.Y(_126_),
    .B(\top_instance.comparator_inst.input_reg[6] ),
    .A_N(\top_instance.comparator_inst.comp_reg[6] ));
 sg13g2_o21ai_1 _463_ (.B1(_126_),
    .Y(_127_),
    .A1(_082_),
    .A2(net183));
 sg13g2_nor2_1 _464_ (.A(_125_),
    .B(_127_),
    .Y(_128_));
 sg13g2_a21oi_1 _465_ (.A1(_082_),
    .A2(net183),
    .Y(_002_),
    .B1(_128_));
 sg13g2_a21o_1 _466_ (.A2(net183),
    .A1(_082_),
    .B1(_128_),
    .X(_000_));
 sg13g2_and2_1 _467_ (.A(net70),
    .B(net132),
    .X(_008_));
 sg13g2_nor3_1 _468_ (.A(net179),
    .B(net232),
    .C(net248),
    .Y(_129_));
 sg13g2_nor4_2 _469_ (.A(net179),
    .B(\top_instance.adc_inst.clk_counter[1] ),
    .C(net195),
    .Y(_130_),
    .D(\top_instance.adc_inst.clk_counter[2] ));
 sg13g2_nand2b_1 _470_ (.Y(_131_),
    .B(_130_),
    .A_N(net209));
 sg13g2_nor2_1 _471_ (.A(\top_instance.adc_inst.clk_counter[4] ),
    .B(\top_instance.adc_inst.clk_counter[5] ),
    .Y(_132_));
 sg13g2_nor2_1 _472_ (.A(\top_instance.adc_inst.clk_counter[7] ),
    .B(\top_instance.adc_inst.clk_counter[6] ),
    .Y(_133_));
 sg13g2_and3_1 _473_ (.X(_134_),
    .A(_130_),
    .B(_132_),
    .C(_133_));
 sg13g2_nor2_1 _474_ (.A(net219),
    .B(\top_instance.adc_inst.clk_counter[8] ),
    .Y(_135_));
 sg13g2_nand2_2 _475_ (.Y(_136_),
    .A(_134_),
    .B(_135_));
 sg13g2_nand2_2 _476_ (.Y(_137_),
    .A(net69),
    .B(_136_));
 sg13g2_xnor2_1 _477_ (.Y(_138_),
    .A(net209),
    .B(_130_));
 sg13g2_nor2_1 _478_ (.A(_137_),
    .B(net210),
    .Y(_009_));
 sg13g2_and3_1 _479_ (.X(_139_),
    .A(net236),
    .B(\top_instance.pulse_generator_inst.red_ctrl_counter[4] ),
    .C(\top_instance.pulse_generator_inst.red_ctrl_counter[3] ));
 sg13g2_nand4_1 _480_ (.B(\top_instance.pulse_generator_inst.red_ctrl_counter[2] ),
    .C(\top_instance.pulse_generator_inst.red_ctrl_counter[1] ),
    .A(\top_instance.pulse_generator_inst.red_ctrl_counter[3] ),
    .Y(_140_),
    .D(\top_instance.pulse_generator_inst.red_ctrl_counter[0] ));
 sg13g2_nand4_1 _481_ (.B(\top_instance.pulse_generator_inst.red_ctrl_counter[18] ),
    .C(net190),
    .A(net156),
    .Y(_141_),
    .D(net167));
 sg13g2_nor2_1 _482_ (.A(_140_),
    .B(_141_),
    .Y(_142_));
 sg13g2_nor4_1 _483_ (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[15] ),
    .B(_098_),
    .C(\top_instance.pulse_generator_inst.red_ctrl_counter[13] ),
    .D(\top_instance.pulse_generator_inst.red_ctrl_counter[12] ),
    .Y(_143_));
 sg13g2_nor3_1 _484_ (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[23] ),
    .B(\top_instance.pulse_generator_inst.red_ctrl_counter[22] ),
    .C(\top_instance.pulse_generator_inst.red_ctrl_counter[21] ),
    .Y(_144_));
 sg13g2_nand2b_1 _485_ (.Y(_145_),
    .B(\top_instance.pulse_generator_inst.red_ctrl_counter[4] ),
    .A_N(\top_instance.pulse_generator_inst.red_ctrl_counter[7] ));
 sg13g2_nand2b_1 _486_ (.Y(_146_),
    .B(\top_instance.pulse_generator_inst.red_ctrl_counter[5] ),
    .A_N(\top_instance.pulse_generator_inst.red_ctrl_counter[6] ));
 sg13g2_or4_1 _487_ (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[11] ),
    .B(\top_instance.pulse_generator_inst.red_ctrl_counter[10] ),
    .C(_100_),
    .D(\top_instance.pulse_generator_inst.red_ctrl_counter[8] ),
    .X(_147_));
 sg13g2_nor4_1 _488_ (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[20] ),
    .B(_145_),
    .C(_146_),
    .D(_147_),
    .Y(_148_));
 sg13g2_nand4_1 _489_ (.B(_143_),
    .C(_144_),
    .A(_142_),
    .Y(_149_),
    .D(_148_));
 sg13g2_inv_1 _490_ (.Y(_150_),
    .A(_149_));
 sg13g2_o21ai_1 _491_ (.B1(\top_instance.comparator_inst.red_enable ),
    .Y(_151_),
    .A1(\top_instance.pulse_generator_inst.red_led ),
    .A2(_150_));
 sg13g2_o21ai_1 _492_ (.B1(net68),
    .Y(_152_),
    .A1(net151),
    .A2(_149_));
 sg13g2_nor2_1 _493_ (.A(_151_),
    .B(_152_),
    .Y(_010_));
 sg13g2_nand3_1 _494_ (.B(_130_),
    .C(_132_),
    .A(net245),
    .Y(_153_));
 sg13g2_xor2_1 _495_ (.B(_153_),
    .A(net207),
    .X(_154_));
 sg13g2_nor2_1 _496_ (.A(_137_),
    .B(net208),
    .Y(_011_));
 sg13g2_nand2_1 _497_ (.Y(_155_),
    .A(net161),
    .B(_134_));
 sg13g2_or2_1 _498_ (.X(_156_),
    .B(_134_),
    .A(net161));
 sg13g2_a21oi_1 _499_ (.A1(net162),
    .A2(_156_),
    .Y(_012_),
    .B1(_137_));
 sg13g2_xor2_1 _500_ (.B(_155_),
    .A(net219),
    .X(_157_));
 sg13g2_nor2_1 _501_ (.A(_137_),
    .B(_157_),
    .Y(_013_));
 sg13g2_and2_1 _502_ (.A(net69),
    .B(net9),
    .X(_014_));
 sg13g2_o21ai_1 _503_ (.B1(net72),
    .Y(_158_),
    .A1(net60),
    .A2(net200));
 sg13g2_a21oi_1 _504_ (.A1(net59),
    .A2(_111_),
    .Y(_015_),
    .B1(_158_));
 sg13g2_o21ai_1 _505_ (.B1(net72),
    .Y(_159_),
    .A1(net60),
    .A2(net194));
 sg13g2_a21oi_1 _506_ (.A1(net59),
    .A2(_110_),
    .Y(_016_),
    .B1(_159_));
 sg13g2_o21ai_1 _507_ (.B1(net72),
    .Y(_160_),
    .A1(net59),
    .A2(net216));
 sg13g2_a21oi_1 _508_ (.A1(net59),
    .A2(_109_),
    .Y(_017_),
    .B1(_160_));
 sg13g2_o21ai_1 _509_ (.B1(net72),
    .Y(_161_),
    .A1(net59),
    .A2(net206));
 sg13g2_a21oi_1 _510_ (.A1(net59),
    .A2(_108_),
    .Y(_018_),
    .B1(_161_));
 sg13g2_o21ai_1 _511_ (.B1(net73),
    .Y(_162_),
    .A1(net61),
    .A2(net215));
 sg13g2_a21oi_1 _512_ (.A1(net61),
    .A2(_107_),
    .Y(_019_),
    .B1(_162_));
 sg13g2_o21ai_1 _513_ (.B1(net73),
    .Y(_163_),
    .A1(net61),
    .A2(net218));
 sg13g2_a21oi_1 _514_ (.A1(net61),
    .A2(_106_),
    .Y(_020_),
    .B1(_163_));
 sg13g2_o21ai_1 _515_ (.B1(net73),
    .Y(_164_),
    .A1(net62),
    .A2(net203));
 sg13g2_a21oi_1 _516_ (.A1(net62),
    .A2(_104_),
    .Y(_021_),
    .B1(net204));
 sg13g2_o21ai_1 _517_ (.B1(net69),
    .Y(_165_),
    .A1(net62),
    .A2(net183));
 sg13g2_a21oi_1 _518_ (.A1(net62),
    .A2(_103_),
    .Y(_022_),
    .B1(_165_));
 sg13g2_and2_1 _519_ (.A(net69),
    .B(\top_instance.adc_inst.data_in_reg ),
    .X(_023_));
 sg13g2_and2_1 _520_ (.A(net69),
    .B(\top_instance.adc_data[0] ),
    .X(_024_));
 sg13g2_and2_1 _521_ (.A(net70),
    .B(\top_instance.adc_data[1] ),
    .X(_025_));
 sg13g2_and2_1 _522_ (.A(net70),
    .B(\top_instance.adc_data[2] ),
    .X(_026_));
 sg13g2_and2_1 _523_ (.A(net73),
    .B(\top_instance.adc_data[3] ),
    .X(_027_));
 sg13g2_nor2_1 _524_ (.A(_111_),
    .B(net66),
    .Y(_028_));
 sg13g2_nor2_1 _525_ (.A(_110_),
    .B(net66),
    .Y(_029_));
 sg13g2_nor2_1 _526_ (.A(_109_),
    .B(net65),
    .Y(_030_));
 sg13g2_nor2_1 _527_ (.A(_108_),
    .B(net65),
    .Y(_031_));
 sg13g2_nor2_1 _528_ (.A(_107_),
    .B(net65),
    .Y(_032_));
 sg13g2_nor2_1 _529_ (.A(_106_),
    .B(net65),
    .Y(_033_));
 sg13g2_nor2_1 _530_ (.A(_104_),
    .B(net65),
    .Y(_034_));
 sg13g2_or2_1 _531_ (.X(_166_),
    .B(\top_instance.adc_inst.bit_counter[0] ),
    .A(\top_instance.adc_inst.bit_counter[1] ));
 sg13g2_nor4_2 _532_ (.A(\top_instance.adc_inst.bit_counter[3] ),
    .B(net177),
    .C(\top_instance.adc_inst.bit_counter[1] ),
    .Y(_167_),
    .D(\top_instance.adc_inst.bit_counter[0] ));
 sg13g2_nor2b_1 _533_ (.A(\top_instance.adc_inst.bit_counter[4] ),
    .B_N(_167_),
    .Y(_168_));
 sg13g2_nor2b_1 _534_ (.A(net165),
    .B_N(_168_),
    .Y(_169_));
 sg13g2_or2_2 _535_ (.X(_170_),
    .B(_169_),
    .A(_136_));
 sg13g2_a21o_1 _536_ (.A2(_169_),
    .A1(net213),
    .B1(_136_),
    .X(_171_));
 sg13g2_nor2_1 _537_ (.A(net220),
    .B(_170_),
    .Y(_172_));
 sg13g2_a21oi_1 _538_ (.A1(net220),
    .A2(_171_),
    .Y(_173_),
    .B1(_172_));
 sg13g2_nor2_1 _539_ (.A(net64),
    .B(_173_),
    .Y(_035_));
 sg13g2_a21oi_1 _540_ (.A1(net235),
    .A2(_172_),
    .Y(_174_),
    .B1(net64));
 sg13g2_o21ai_1 _541_ (.B1(_174_),
    .Y(_175_),
    .A1(net235),
    .A2(_172_));
 sg13g2_inv_1 _542_ (.Y(_036_),
    .A(_175_));
 sg13g2_and2_1 _543_ (.A(net67),
    .B(_171_),
    .X(_176_));
 sg13g2_nand2_1 _544_ (.Y(_177_),
    .A(net67),
    .B(_171_));
 sg13g2_or2_1 _545_ (.X(_178_),
    .B(_166_),
    .A(_113_));
 sg13g2_nand2_1 _546_ (.Y(_179_),
    .A(_113_),
    .B(_166_));
 sg13g2_a21oi_1 _547_ (.A1(_178_),
    .A2(_179_),
    .Y(_180_),
    .B1(_170_));
 sg13g2_a22oi_1 _548_ (.Y(_181_),
    .B1(_180_),
    .B2(net67),
    .A2(_176_),
    .A1(net177));
 sg13g2_inv_1 _549_ (.Y(_037_),
    .A(net178));
 sg13g2_xor2_1 _550_ (.B(_178_),
    .A(net217),
    .X(_182_));
 sg13g2_nor2_1 _551_ (.A(_170_),
    .B(_182_),
    .Y(_183_));
 sg13g2_a22oi_1 _552_ (.Y(_184_),
    .B1(_183_),
    .B2(net67),
    .A2(_176_),
    .A1(net217));
 sg13g2_inv_1 _553_ (.Y(_038_),
    .A(_184_));
 sg13g2_xnor2_1 _554_ (.Y(_185_),
    .A(net201),
    .B(_167_));
 sg13g2_nor3_1 _555_ (.A(net64),
    .B(_170_),
    .C(_185_),
    .Y(_186_));
 sg13g2_a21o_1 _556_ (.A2(_176_),
    .A1(net201),
    .B1(_186_),
    .X(_039_));
 sg13g2_nand3_1 _557_ (.B(_135_),
    .C(_168_),
    .A(_134_),
    .Y(_187_));
 sg13g2_nand2b_1 _558_ (.Y(_188_),
    .B(_169_),
    .A_N(_136_));
 sg13g2_inv_1 _559_ (.Y(_189_),
    .A(_188_));
 sg13g2_nor2_1 _560_ (.A(net213),
    .B(_188_),
    .Y(_190_));
 sg13g2_a21oi_1 _561_ (.A1(net165),
    .A2(_187_),
    .Y(_191_),
    .B1(_190_));
 sg13g2_nor2_1 _562_ (.A(net64),
    .B(net166),
    .Y(_040_));
 sg13g2_nor2_1 _563_ (.A(net64),
    .B(net179),
    .Y(_041_));
 sg13g2_xor2_1 _564_ (.B(net232),
    .A(net179),
    .X(_192_));
 sg13g2_nor2_1 _565_ (.A(net64),
    .B(_192_),
    .Y(_042_));
 sg13g2_o21ai_1 _566_ (.B1(net248),
    .Y(_193_),
    .A1(net179),
    .A2(net232));
 sg13g2_nor2b_1 _567_ (.A(_129_),
    .B_N(_193_),
    .Y(_194_));
 sg13g2_nor2_1 _568_ (.A(net64),
    .B(_194_),
    .Y(_043_));
 sg13g2_xnor2_1 _569_ (.Y(_195_),
    .A(net195),
    .B(_129_));
 sg13g2_nor2_1 _570_ (.A(_177_),
    .B(net196),
    .Y(_044_));
 sg13g2_xnor2_1 _571_ (.Y(_196_),
    .A(net239),
    .B(_131_));
 sg13g2_o21ai_1 _572_ (.B1(net240),
    .Y(_197_),
    .A1(net230),
    .A2(_188_));
 sg13g2_nor2_1 _573_ (.A(net64),
    .B(_197_),
    .Y(_045_));
 sg13g2_a21o_1 _574_ (.A2(_132_),
    .A1(_130_),
    .B1(net245),
    .X(_198_));
 sg13g2_and2_1 _575_ (.A(net246),
    .B(_198_),
    .X(_199_));
 sg13g2_a21oi_1 _576_ (.A1(_136_),
    .A2(_199_),
    .Y(_046_),
    .B1(_177_));
 sg13g2_nor2_1 _577_ (.A(net230),
    .B(_189_),
    .Y(_200_));
 sg13g2_o21ai_1 _578_ (.B1(net69),
    .Y(_047_),
    .A1(_190_),
    .A2(_200_));
 sg13g2_o21ai_1 _579_ (.B1(net69),
    .Y(_201_),
    .A1(net62),
    .A2(_189_));
 sg13g2_nor2_1 _580_ (.A(_190_),
    .B(_201_),
    .Y(_048_));
 sg13g2_o21ai_1 _581_ (.B1(net69),
    .Y(_202_),
    .A1(net147),
    .A2(_170_));
 sg13g2_a21oi_1 _582_ (.A1(_102_),
    .A2(_170_),
    .Y(_049_),
    .B1(_202_));
 sg13g2_o21ai_1 _583_ (.B1(net67),
    .Y(_203_),
    .A1(\top_instance.comparator_inst.red_enable ),
    .A2(net192));
 sg13g2_a21oi_1 _584_ (.A1(\top_instance.comparator_inst.red_enable ),
    .A2(net192),
    .Y(_050_),
    .B1(_203_));
 sg13g2_a21oi_1 _585_ (.A1(\top_instance.comparator_inst.red_enable ),
    .A2(\top_instance.pulse_generator_inst.red_ctrl_counter[0] ),
    .Y(_204_),
    .B1(net172));
 sg13g2_nand3_1 _586_ (.B(net172),
    .C(\top_instance.pulse_generator_inst.red_ctrl_counter[0] ),
    .A(\top_instance.comparator_inst.red_enable ),
    .Y(_205_));
 sg13g2_nand2_1 _587_ (.Y(_206_),
    .A(net68),
    .B(_205_));
 sg13g2_nor2_1 _588_ (.A(net173),
    .B(_206_),
    .Y(_051_));
 sg13g2_nor2b_1 _589_ (.A(net188),
    .B_N(_205_),
    .Y(_207_));
 sg13g2_and4_2 _590_ (.A(\top_instance.comparator_inst.red_enable ),
    .B(net188),
    .C(net172),
    .D(\top_instance.pulse_generator_inst.red_ctrl_counter[0] ),
    .X(_208_));
 sg13g2_nor3_1 _591_ (.A(net65),
    .B(net189),
    .C(_208_),
    .Y(_052_));
 sg13g2_o21ai_1 _592_ (.B1(net67),
    .Y(_209_),
    .A1(net198),
    .A2(_208_));
 sg13g2_a21oi_1 _593_ (.A1(net198),
    .A2(_208_),
    .Y(_053_),
    .B1(_209_));
 sg13g2_a21oi_1 _594_ (.A1(\top_instance.pulse_generator_inst.red_ctrl_counter[3] ),
    .A2(_208_),
    .Y(_210_),
    .B1(net185));
 sg13g2_and3_1 _595_ (.X(_211_),
    .A(net185),
    .B(net198),
    .C(_208_));
 sg13g2_nor3_1 _596_ (.A(net66),
    .B(net186),
    .C(_211_),
    .Y(_054_));
 sg13g2_and2_1 _597_ (.A(_139_),
    .B(_208_),
    .X(_212_));
 sg13g2_o21ai_1 _598_ (.B1(net67),
    .Y(_213_),
    .A1(net236),
    .A2(_211_));
 sg13g2_nor2_1 _599_ (.A(_212_),
    .B(_213_),
    .Y(_055_));
 sg13g2_a21o_2 _600_ (.A2(_150_),
    .A1(\top_instance.comparator_inst.red_enable ),
    .B1(net65),
    .X(_214_));
 sg13g2_xnor2_1 _601_ (.Y(_215_),
    .A(net223),
    .B(_212_));
 sg13g2_nor2_1 _602_ (.A(_214_),
    .B(_215_),
    .Y(_056_));
 sg13g2_a21oi_1 _603_ (.A1(\top_instance.pulse_generator_inst.red_ctrl_counter[6] ),
    .A2(_212_),
    .Y(_216_),
    .B1(net163));
 sg13g2_nand4_1 _604_ (.B(net223),
    .C(_139_),
    .A(net163),
    .Y(_217_),
    .D(_208_));
 sg13g2_inv_1 _605_ (.Y(_218_),
    .A(_217_));
 sg13g2_nor3_1 _606_ (.A(net66),
    .B(net164),
    .C(_218_),
    .Y(_057_));
 sg13g2_o21ai_1 _607_ (.B1(net68),
    .Y(_219_),
    .A1(_101_),
    .A2(_217_));
 sg13g2_a21oi_1 _608_ (.A1(_101_),
    .A2(_217_),
    .Y(_058_),
    .B1(_219_));
 sg13g2_a21oi_1 _609_ (.A1(\top_instance.pulse_generator_inst.red_ctrl_counter[8] ),
    .A2(_218_),
    .Y(_220_),
    .B1(net153));
 sg13g2_nor3_1 _610_ (.A(_100_),
    .B(_101_),
    .C(_217_),
    .Y(_221_));
 sg13g2_nor3_1 _611_ (.A(_214_),
    .B(net154),
    .C(_221_),
    .Y(_059_));
 sg13g2_nor4_2 _612_ (.A(_099_),
    .B(_100_),
    .C(_101_),
    .Y(_222_),
    .D(_217_));
 sg13g2_o21ai_1 _613_ (.B1(net68),
    .Y(_223_),
    .A1(net227),
    .A2(_221_));
 sg13g2_nor2_1 _614_ (.A(_222_),
    .B(net228),
    .Y(_060_));
 sg13g2_nor2_1 _615_ (.A(net211),
    .B(_222_),
    .Y(_224_));
 sg13g2_and2_1 _616_ (.A(net211),
    .B(_222_),
    .X(_225_));
 sg13g2_nor3_1 _617_ (.A(net65),
    .B(net212),
    .C(_225_),
    .Y(_061_));
 sg13g2_o21ai_1 _618_ (.B1(net74),
    .Y(_226_),
    .A1(net175),
    .A2(_225_));
 sg13g2_a21oi_1 _619_ (.A1(net175),
    .A2(_225_),
    .Y(_062_),
    .B1(_226_));
 sg13g2_a21oi_1 _620_ (.A1(\top_instance.pulse_generator_inst.red_ctrl_counter[12] ),
    .A2(_225_),
    .Y(_227_),
    .B1(net159));
 sg13g2_nand4_1 _621_ (.B(net249),
    .C(net211),
    .A(net159),
    .Y(_228_),
    .D(_222_));
 sg13g2_nand2_1 _622_ (.Y(_229_),
    .A(net74),
    .B(_228_));
 sg13g2_nor2_1 _623_ (.A(net160),
    .B(_229_),
    .Y(_063_));
 sg13g2_and2_1 _624_ (.A(_098_),
    .B(_228_),
    .X(_230_));
 sg13g2_nor2_1 _625_ (.A(_098_),
    .B(_228_),
    .Y(_231_));
 sg13g2_nor3_1 _626_ (.A(_214_),
    .B(net244),
    .C(_231_),
    .Y(_064_));
 sg13g2_xnor2_1 _627_ (.Y(_232_),
    .A(net221),
    .B(_231_));
 sg13g2_nor2_1 _628_ (.A(net66),
    .B(net222),
    .Y(_065_));
 sg13g2_a21oi_1 _629_ (.A1(\top_instance.pulse_generator_inst.red_ctrl_counter[15] ),
    .A2(_231_),
    .Y(_233_),
    .B1(net167));
 sg13g2_nor4_2 _630_ (.A(_096_),
    .B(_097_),
    .C(_098_),
    .Y(_234_),
    .D(_228_));
 sg13g2_nor3_1 _631_ (.A(_214_),
    .B(net168),
    .C(_234_),
    .Y(_066_));
 sg13g2_nor2_1 _632_ (.A(net190),
    .B(_234_),
    .Y(_235_));
 sg13g2_and2_1 _633_ (.A(net190),
    .B(_234_),
    .X(_236_));
 sg13g2_nor3_1 _634_ (.A(_214_),
    .B(net191),
    .C(_236_),
    .Y(_067_));
 sg13g2_nor2_1 _635_ (.A(net226),
    .B(_236_),
    .Y(_237_));
 sg13g2_and2_1 _636_ (.A(net226),
    .B(_236_),
    .X(_238_));
 sg13g2_nor3_1 _637_ (.A(_214_),
    .B(_237_),
    .C(_238_),
    .Y(_068_));
 sg13g2_a21oi_1 _638_ (.A1(\top_instance.pulse_generator_inst.red_ctrl_counter[18] ),
    .A2(_236_),
    .Y(_239_),
    .B1(net156));
 sg13g2_nor4_2 _639_ (.A(_097_),
    .B(_098_),
    .C(_141_),
    .Y(_240_),
    .D(_228_));
 sg13g2_nor3_1 _640_ (.A(_214_),
    .B(net157),
    .C(_240_),
    .Y(_069_));
 sg13g2_o21ai_1 _641_ (.B1(net74),
    .Y(_241_),
    .A1(net224),
    .A2(_240_));
 sg13g2_a21oi_1 _642_ (.A1(net224),
    .A2(_240_),
    .Y(_070_),
    .B1(_241_));
 sg13g2_a21oi_1 _643_ (.A1(\top_instance.pulse_generator_inst.red_ctrl_counter[20] ),
    .A2(_240_),
    .Y(_242_),
    .B1(net180));
 sg13g2_nand3_1 _644_ (.B(net224),
    .C(_240_),
    .A(net180),
    .Y(_243_));
 sg13g2_nand2_1 _645_ (.Y(_244_),
    .A(net74),
    .B(_243_));
 sg13g2_nor2_1 _646_ (.A(net181),
    .B(_244_),
    .Y(_071_));
 sg13g2_nand2b_1 _647_ (.Y(_245_),
    .B(_243_),
    .A_N(net241));
 sg13g2_nand4_1 _648_ (.B(net180),
    .C(\top_instance.pulse_generator_inst.red_ctrl_counter[20] ),
    .A(net241),
    .Y(_246_),
    .D(_240_));
 sg13g2_and3_1 _649_ (.X(_072_),
    .A(net74),
    .B(_245_),
    .C(_246_));
 sg13g2_o21ai_1 _650_ (.B1(net74),
    .Y(_247_),
    .A1(_095_),
    .A2(_246_));
 sg13g2_a21oi_1 _651_ (.A1(_095_),
    .A2(_246_),
    .Y(_073_),
    .B1(_247_));
 sg13g2_o21ai_1 _652_ (.B1(net72),
    .Y(_248_),
    .A1(net63),
    .A2(\top_instance.comparator_inst.input_reg[0] ));
 sg13g2_a21oi_1 _653_ (.A1(net63),
    .A2(_094_),
    .Y(_074_),
    .B1(_248_));
 sg13g2_o21ai_1 _654_ (.B1(net72),
    .Y(_249_),
    .A1(net59),
    .A2(\top_instance.comparator_inst.input_reg[1] ));
 sg13g2_a21oi_1 _655_ (.A1(net59),
    .A2(_093_),
    .Y(_075_),
    .B1(_249_));
 sg13g2_o21ai_1 _656_ (.B1(net72),
    .Y(_250_),
    .A1(net60),
    .A2(\top_instance.comparator_inst.input_reg[2] ));
 sg13g2_a21oi_1 _657_ (.A1(net60),
    .A2(_092_),
    .Y(_076_),
    .B1(_250_));
 sg13g2_o21ai_1 _658_ (.B1(net73),
    .Y(_251_),
    .A1(net63),
    .A2(\top_instance.comparator_inst.input_reg[3] ));
 sg13g2_a21oi_1 _659_ (.A1(net60),
    .A2(_090_),
    .Y(_077_),
    .B1(_251_));
 sg13g2_o21ai_1 _660_ (.B1(net72),
    .Y(_252_),
    .A1(net60),
    .A2(\top_instance.comparator_inst.input_reg[4] ));
 sg13g2_a21oi_1 _661_ (.A1(net60),
    .A2(_089_),
    .Y(_078_),
    .B1(_252_));
 sg13g2_o21ai_1 _662_ (.B1(net73),
    .Y(_253_),
    .A1(net61),
    .A2(\top_instance.comparator_inst.input_reg[5] ));
 sg13g2_a21oi_1 _663_ (.A1(net61),
    .A2(_087_),
    .Y(_079_),
    .B1(_253_));
 sg13g2_o21ai_1 _664_ (.B1(net73),
    .Y(_254_),
    .A1(net62),
    .A2(\top_instance.comparator_inst.input_reg[6] ));
 sg13g2_a21oi_1 _665_ (.A1(net61),
    .A2(_085_),
    .Y(_080_),
    .B1(_254_));
 sg13g2_o21ai_1 _666_ (.B1(net70),
    .Y(_255_),
    .A1(\top_instance.comparator_inst.input_reg[7] ),
    .A2(net62));
 sg13g2_a21oi_1 _667_ (.A1(_083_),
    .A2(net62),
    .Y(_081_),
    .B1(_255_));
 sg13g2_dfrbp_1 _668_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net43),
    .D(_008_),
    .Q_N(_324_),
    .Q(\top_instance.green_led ));
 sg13g2_dfrbp_1 _669_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net37),
    .D(_009_),
    .Q_N(_323_),
    .Q(\top_instance.adc_inst.clk_counter[4] ));
 sg13g2_dfrbp_1 _670_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net36),
    .D(net152),
    .Q_N(_003_),
    .Q(\top_instance.pulse_generator_inst.red_led ));
 sg13g2_dfrbp_1 _671_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net34),
    .D(_011_),
    .Q_N(_322_),
    .Q(\top_instance.adc_inst.clk_counter[7] ));
 sg13g2_dfrbp_1 _672_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net33),
    .D(_012_),
    .Q_N(_007_),
    .Q(\top_instance.adc_inst.clk_counter[8] ));
 sg13g2_dfrbp_1 _673_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net32),
    .D(_013_),
    .Q_N(_321_),
    .Q(\top_instance.adc_inst.clk_counter[9] ));
 sg13g2_dfrbp_1 _674_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net31),
    .D(_014_),
    .Q_N(_320_),
    .Q(\top_instance.adc_inst.data_in_reg ));
 sg13g2_dfrbp_1 _675_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net30),
    .D(_015_),
    .Q_N(_319_),
    .Q(\top_instance.comparator_inst.comp_reg[0] ));
 sg13g2_dfrbp_1 _676_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net28),
    .D(_016_),
    .Q_N(_318_),
    .Q(\top_instance.comparator_inst.comp_reg[1] ));
 sg13g2_dfrbp_1 _677_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net128),
    .D(_017_),
    .Q_N(_317_),
    .Q(\top_instance.comparator_inst.comp_reg[2] ));
 sg13g2_dfrbp_1 _678_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net126),
    .D(_018_),
    .Q_N(_316_),
    .Q(\top_instance.comparator_inst.comp_reg[3] ));
 sg13g2_dfrbp_1 _679_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net124),
    .D(_019_),
    .Q_N(_315_),
    .Q(\top_instance.comparator_inst.comp_reg[4] ));
 sg13g2_dfrbp_1 _680_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net122),
    .D(_020_),
    .Q_N(_314_),
    .Q(\top_instance.comparator_inst.comp_reg[5] ));
 sg13g2_dfrbp_1 _681_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net120),
    .D(net205),
    .Q_N(_313_),
    .Q(\top_instance.comparator_inst.comp_reg[6] ));
 sg13g2_dfrbp_1 _682_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net44),
    .D(_022_),
    .Q_N(_325_),
    .Q(\top_instance.comparator_inst.comp_reg[7] ));
 sg13g2_dfrbp_1 _683_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net90),
    .D(net234),
    .Q_N(_326_),
    .Q(\top_instance.comparator_inst.red_enable ));
 sg13g2_dfrbp_1 _684_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net118),
    .D(net184),
    .Q_N(_312_),
    .Q(\top_instance.comparator_inst.green_enable ));
 sg13g2_dfrbp_1 _685_ (.CLK(net57),
    .RESET_B(net116),
    .D(_023_),
    .Q_N(_311_),
    .Q(\top_instance.adc_data[0] ));
 sg13g2_dfrbp_1 _686_ (.CLK(net57),
    .RESET_B(net115),
    .D(_024_),
    .Q_N(_310_),
    .Q(\top_instance.adc_data[1] ));
 sg13g2_dfrbp_1 _687_ (.CLK(net57),
    .RESET_B(net114),
    .D(_025_),
    .Q_N(_309_),
    .Q(\top_instance.adc_data[2] ));
 sg13g2_dfrbp_1 _688_ (.CLK(net58),
    .RESET_B(net113),
    .D(_026_),
    .Q_N(_308_),
    .Q(\top_instance.adc_data[3] ));
 sg13g2_dfrbp_1 _689_ (.CLK(net58),
    .RESET_B(net112),
    .D(_027_),
    .Q_N(_307_),
    .Q(\top_instance.adc_data[4] ));
 sg13g2_dfrbp_1 _690_ (.CLK(net58),
    .RESET_B(net111),
    .D(_028_),
    .Q_N(_306_),
    .Q(\top_instance.adc_data[5] ));
 sg13g2_dfrbp_1 _691_ (.CLK(net58),
    .RESET_B(net110),
    .D(_029_),
    .Q_N(_305_),
    .Q(\top_instance.adc_data[6] ));
 sg13g2_dfrbp_1 _692_ (.CLK(net58),
    .RESET_B(net109),
    .D(_030_),
    .Q_N(_304_),
    .Q(\top_instance.adc_data[7] ));
 sg13g2_dfrbp_1 _693_ (.CLK(net58),
    .RESET_B(net108),
    .D(_031_),
    .Q_N(_303_),
    .Q(\top_instance.adc_data[8] ));
 sg13g2_dfrbp_1 _694_ (.CLK(net57),
    .RESET_B(net107),
    .D(_032_),
    .Q_N(_302_),
    .Q(\top_instance.adc_data[9] ));
 sg13g2_dfrbp_1 _695_ (.CLK(net57),
    .RESET_B(net106),
    .D(_033_),
    .Q_N(_301_),
    .Q(\top_instance.adc_data[10] ));
 sg13g2_dfrbp_1 _696_ (.CLK(net57),
    .RESET_B(net105),
    .D(_034_),
    .Q_N(_300_),
    .Q(\top_instance.adc_data[11] ));
 sg13g2_dfrbp_1 _697_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net104),
    .D(_035_),
    .Q_N(_299_),
    .Q(\top_instance.adc_inst.bit_counter[0] ));
 sg13g2_dfrbp_1 _698_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net102),
    .D(_036_),
    .Q_N(_298_),
    .Q(\top_instance.adc_inst.bit_counter[1] ));
 sg13g2_dfrbp_1 _699_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net100),
    .D(_037_),
    .Q_N(_006_),
    .Q(\top_instance.adc_inst.bit_counter[2] ));
 sg13g2_dfrbp_1 _700_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net98),
    .D(_038_),
    .Q_N(_297_),
    .Q(\top_instance.adc_inst.bit_counter[3] ));
 sg13g2_dfrbp_1 _701_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net88),
    .D(net202),
    .Q_N(_296_),
    .Q(\top_instance.adc_inst.bit_counter[4] ));
 sg13g2_dfrbp_1 _702_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net86),
    .D(_040_),
    .Q_N(_295_),
    .Q(\top_instance.adc_inst.bit_counter[5] ));
 sg13g2_dfrbp_1 _703_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net84),
    .D(_041_),
    .Q_N(_294_),
    .Q(\top_instance.adc_inst.clk_counter[0] ));
 sg13g2_dfrbp_1 _704_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net83),
    .D(_042_),
    .Q_N(_293_),
    .Q(\top_instance.adc_inst.clk_counter[1] ));
 sg13g2_dfrbp_1 _705_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net82),
    .D(_043_),
    .Q_N(_292_),
    .Q(\top_instance.adc_inst.clk_counter[2] ));
 sg13g2_dfrbp_1 _706_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net81),
    .D(net197),
    .Q_N(_291_),
    .Q(\top_instance.adc_inst.clk_counter[3] ));
 sg13g2_dfrbp_1 _707_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net80),
    .D(_045_),
    .Q_N(_290_),
    .Q(\top_instance.adc_inst.clk_counter[5] ));
 sg13g2_dfrbp_1 _708_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net79),
    .D(net247),
    .Q_N(_005_),
    .Q(\top_instance.adc_inst.clk_counter[6] ));
 sg13g2_dfrbp_1 _709_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net78),
    .D(_047_),
    .Q_N(_004_),
    .Q(\top_instance.adc_inst.cs ));
 sg13g2_dfrbp_1 _710_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net76),
    .D(net214),
    .Q_N(_289_),
    .Q(\top_instance.adc_inst.data_ready ));
 sg13g2_dfrbp_1 _711_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net91),
    .D(net148),
    .Q_N(_001_),
    .Q(\top_instance.adc_inst.sclk ));
 sg13g2_dfrbp_1 _712_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net92),
    .D(net1),
    .Q_N(_327_),
    .Q(\top_instance.comparator_inst.in[0] ));
 sg13g2_dfrbp_1 _713_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net93),
    .D(net2),
    .Q_N(_328_),
    .Q(\top_instance.comparator_inst.in[1] ));
 sg13g2_dfrbp_1 _714_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net94),
    .D(net3),
    .Q_N(_329_),
    .Q(\top_instance.comparator_inst.in[2] ));
 sg13g2_dfrbp_1 _715_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net95),
    .D(net4),
    .Q_N(_330_),
    .Q(\top_instance.comparator_inst.in[3] ));
 sg13g2_dfrbp_1 _716_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net96),
    .D(net5),
    .Q_N(_331_),
    .Q(\top_instance.comparator_inst.in[4] ));
 sg13g2_dfrbp_1 _717_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net97),
    .D(net6),
    .Q_N(_332_),
    .Q(\top_instance.comparator_inst.in[5] ));
 sg13g2_dfrbp_1 _718_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net53),
    .D(net7),
    .Q_N(_333_),
    .Q(\top_instance.comparator_inst.in[6] ));
 sg13g2_dfrbp_1 _719_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net56),
    .D(net8),
    .Q_N(_288_),
    .Q(\top_instance.comparator_inst.in[7] ));
 sg13g2_dfrbp_1 _720_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net54),
    .D(net193),
    .Q_N(_287_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[0] ));
 sg13g2_dfrbp_1 _721_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net52),
    .D(net174),
    .Q_N(_286_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[1] ));
 sg13g2_dfrbp_1 _722_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net50),
    .D(_052_),
    .Q_N(_285_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[2] ));
 sg13g2_dfrbp_1 _723_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net48),
    .D(net199),
    .Q_N(_284_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[3] ));
 sg13g2_dfrbp_1 _724_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net46),
    .D(net187),
    .Q_N(_283_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[4] ));
 sg13g2_dfrbp_1 _725_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net42),
    .D(_055_),
    .Q_N(_282_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[5] ));
 sg13g2_dfrbp_1 _726_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net40),
    .D(_056_),
    .Q_N(_281_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[6] ));
 sg13g2_dfrbp_1 _727_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net38),
    .D(_057_),
    .Q_N(_280_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[7] ));
 sg13g2_dfrbp_1 _728_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net29),
    .D(net238),
    .Q_N(_279_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[8] ));
 sg13g2_dfrbp_1 _729_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net127),
    .D(net155),
    .Q_N(_278_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[9] ));
 sg13g2_dfrbp_1 _730_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net123),
    .D(net229),
    .Q_N(_277_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[10] ));
 sg13g2_dfrbp_1 _731_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net119),
    .D(_061_),
    .Q_N(_276_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[11] ));
 sg13g2_dfrbp_1 _732_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net103),
    .D(net176),
    .Q_N(_275_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[12] ));
 sg13g2_dfrbp_1 _733_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net99),
    .D(_063_),
    .Q_N(_274_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[13] ));
 sg13g2_dfrbp_1 _734_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net87),
    .D(_064_),
    .Q_N(_273_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[14] ));
 sg13g2_dfrbp_1 _735_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net77),
    .D(_065_),
    .Q_N(_272_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[15] ));
 sg13g2_dfrbp_1 _736_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net55),
    .D(net169),
    .Q_N(_271_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[16] ));
 sg13g2_dfrbp_1 _737_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net51),
    .D(_067_),
    .Q_N(_270_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[17] ));
 sg13g2_dfrbp_1 _738_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net47),
    .D(_068_),
    .Q_N(_269_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[18] ));
 sg13g2_dfrbp_1 _739_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net41),
    .D(net158),
    .Q_N(_268_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[19] ));
 sg13g2_dfrbp_1 _740_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net35),
    .D(net225),
    .Q_N(_267_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[20] ));
 sg13g2_dfrbp_1 _741_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net125),
    .D(net182),
    .Q_N(_266_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[21] ));
 sg13g2_dfrbp_1 _742_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net117),
    .D(net242),
    .Q_N(_265_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[22] ));
 sg13g2_dfrbp_1 _743_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net89),
    .D(net171),
    .Q_N(_264_),
    .Q(\top_instance.pulse_generator_inst.red_ctrl_counter[23] ));
 sg13g2_dfrbp_1 _744_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net75),
    .D(net136),
    .Q_N(_263_),
    .Q(\top_instance.comparator_inst.input_reg[0] ));
 sg13g2_dfrbp_1 _745_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net49),
    .D(net134),
    .Q_N(_262_),
    .Q(\top_instance.comparator_inst.input_reg[1] ));
 sg13g2_dfrbp_1 _746_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net39),
    .D(net140),
    .Q_N(_261_),
    .Q(\top_instance.comparator_inst.input_reg[2] ));
 sg13g2_dfrbp_1 _747_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net121),
    .D(net150),
    .Q_N(_260_),
    .Q(\top_instance.comparator_inst.input_reg[3] ));
 sg13g2_dfrbp_1 _748_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net85),
    .D(net144),
    .Q_N(_259_),
    .Q(\top_instance.comparator_inst.input_reg[4] ));
 sg13g2_dfrbp_1 _749_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net45),
    .D(net138),
    .Q_N(_258_),
    .Q(\top_instance.comparator_inst.input_reg[5] ));
 sg13g2_dfrbp_1 _750_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net101),
    .D(net146),
    .Q_N(_257_),
    .Q(\top_instance.comparator_inst.input_reg[6] ));
 sg13g2_dfrbp_1 _751_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net129),
    .D(net142),
    .Q_N(_256_),
    .Q(\top_instance.comparator_inst.input_reg[7] ));
 sg13g2_tiehi _728__29 (.L_HI(net29));
 sg13g2_tiehi _675__30 (.L_HI(net30));
 sg13g2_tiehi _674__31 (.L_HI(net31));
 sg13g2_tiehi _673__32 (.L_HI(net32));
 sg13g2_tiehi _672__33 (.L_HI(net33));
 sg13g2_tiehi _671__34 (.L_HI(net34));
 sg13g2_tiehi _740__35 (.L_HI(net35));
 sg13g2_tiehi _670__36 (.L_HI(net36));
 sg13g2_tiehi _669__37 (.L_HI(net37));
 sg13g2_tiehi _727__38 (.L_HI(net38));
 sg13g2_tiehi _746__39 (.L_HI(net39));
 sg13g2_tiehi _726__40 (.L_HI(net40));
 sg13g2_tiehi _739__41 (.L_HI(net41));
 sg13g2_tiehi _725__42 (.L_HI(net42));
 sg13g2_tiehi _668__43 (.L_HI(net43));
 sg13g2_tiehi _682__44 (.L_HI(net44));
 sg13g2_tiehi _749__45 (.L_HI(net45));
 sg13g2_tiehi _724__46 (.L_HI(net46));
 sg13g2_tiehi _738__47 (.L_HI(net47));
 sg13g2_tiehi _723__48 (.L_HI(net48));
 sg13g2_tiehi _745__49 (.L_HI(net49));
 sg13g2_tiehi _722__50 (.L_HI(net50));
 sg13g2_tiehi _737__51 (.L_HI(net51));
 sg13g2_tiehi _721__52 (.L_HI(net52));
 sg13g2_tiehi _718__53 (.L_HI(net53));
 sg13g2_tiehi _720__54 (.L_HI(net54));
 sg13g2_tiehi _736__55 (.L_HI(net55));
 sg13g2_tiehi _719__56 (.L_HI(net56));
 sg13g2_tiehi _744__57 (.L_HI(net75));
 sg13g2_tiehi _710__58 (.L_HI(net76));
 sg13g2_tiehi _735__59 (.L_HI(net77));
 sg13g2_tiehi _709__60 (.L_HI(net78));
 sg13g2_tiehi _708__61 (.L_HI(net79));
 sg13g2_tiehi _707__62 (.L_HI(net80));
 sg13g2_tiehi _706__63 (.L_HI(net81));
 sg13g2_tiehi _705__64 (.L_HI(net82));
 sg13g2_tiehi _704__65 (.L_HI(net83));
 sg13g2_tiehi _703__66 (.L_HI(net84));
 sg13g2_tiehi _748__67 (.L_HI(net85));
 sg13g2_tiehi _702__68 (.L_HI(net86));
 sg13g2_tiehi _734__69 (.L_HI(net87));
 sg13g2_tiehi _701__70 (.L_HI(net88));
 sg13g2_tiehi _743__71 (.L_HI(net89));
 sg13g2_tiehi _683__72 (.L_HI(net90));
 sg13g2_tiehi _711__73 (.L_HI(net91));
 sg13g2_tiehi _712__74 (.L_HI(net92));
 sg13g2_tiehi _713__75 (.L_HI(net93));
 sg13g2_tiehi _714__76 (.L_HI(net94));
 sg13g2_tiehi _715__77 (.L_HI(net95));
 sg13g2_tiehi _716__78 (.L_HI(net96));
 sg13g2_tiehi _717__79 (.L_HI(net97));
 sg13g2_tiehi _700__80 (.L_HI(net98));
 sg13g2_tiehi _733__81 (.L_HI(net99));
 sg13g2_tiehi _699__82 (.L_HI(net100));
 sg13g2_tiehi _750__83 (.L_HI(net101));
 sg13g2_tiehi _698__84 (.L_HI(net102));
 sg13g2_tiehi _732__85 (.L_HI(net103));
 sg13g2_tiehi _697__86 (.L_HI(net104));
 sg13g2_tiehi _696__87 (.L_HI(net105));
 sg13g2_tiehi _695__88 (.L_HI(net106));
 sg13g2_tiehi _694__89 (.L_HI(net107));
 sg13g2_tiehi _693__90 (.L_HI(net108));
 sg13g2_tiehi _692__91 (.L_HI(net109));
 sg13g2_tiehi _691__92 (.L_HI(net110));
 sg13g2_tiehi _690__93 (.L_HI(net111));
 sg13g2_tiehi _689__94 (.L_HI(net112));
 sg13g2_tiehi _688__95 (.L_HI(net113));
 sg13g2_tiehi _687__96 (.L_HI(net114));
 sg13g2_tiehi _686__97 (.L_HI(net115));
 sg13g2_tiehi _685__98 (.L_HI(net116));
 sg13g2_tiehi _742__99 (.L_HI(net117));
 sg13g2_tiehi _684__100 (.L_HI(net118));
 sg13g2_tiehi _731__101 (.L_HI(net119));
 sg13g2_tiehi _681__102 (.L_HI(net120));
 sg13g2_tiehi _747__103 (.L_HI(net121));
 sg13g2_tiehi _680__104 (.L_HI(net122));
 sg13g2_tiehi _730__105 (.L_HI(net123));
 sg13g2_tiehi _679__106 (.L_HI(net124));
 sg13g2_tiehi _741__107 (.L_HI(net125));
 sg13g2_tiehi _678__108 (.L_HI(net126));
 sg13g2_tiehi _729__109 (.L_HI(net127));
 sg13g2_tiehi _677__110 (.L_HI(net128));
 sg13g2_tiehi _751__111 (.L_HI(net129));
 sg13g2_tiehi tt_um_ephrenm_tsal_112 (.L_HI(net130));
 sg13g2_tiehi tt_um_ephrenm_tsal_113 (.L_HI(net131));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_ephrenm_tsal_11 (.L_LO(net11));
 sg13g2_tielo tt_um_ephrenm_tsal_12 (.L_LO(net12));
 sg13g2_tielo tt_um_ephrenm_tsal_13 (.L_LO(net13));
 sg13g2_tielo tt_um_ephrenm_tsal_14 (.L_LO(net14));
 sg13g2_tielo tt_um_ephrenm_tsal_15 (.L_LO(net15));
 sg13g2_tielo tt_um_ephrenm_tsal_16 (.L_LO(net16));
 sg13g2_tielo tt_um_ephrenm_tsal_17 (.L_LO(net17));
 sg13g2_tielo tt_um_ephrenm_tsal_18 (.L_LO(net18));
 sg13g2_tielo tt_um_ephrenm_tsal_19 (.L_LO(net19));
 sg13g2_tielo tt_um_ephrenm_tsal_20 (.L_LO(net20));
 sg13g2_tielo tt_um_ephrenm_tsal_21 (.L_LO(net21));
 sg13g2_tielo tt_um_ephrenm_tsal_22 (.L_LO(net22));
 sg13g2_tielo tt_um_ephrenm_tsal_23 (.L_LO(net23));
 sg13g2_tielo tt_um_ephrenm_tsal_24 (.L_LO(net24));
 sg13g2_tielo tt_um_ephrenm_tsal_25 (.L_LO(net25));
 sg13g2_tielo tt_um_ephrenm_tsal_26 (.L_LO(net26));
 sg13g2_tielo tt_um_ephrenm_tsal_27 (.L_LO(net27));
 sg13g2_tiehi _676__28 (.L_HI(net28));
 sg13g2_buf_1 _856_ (.A(\top_instance.adc_inst.cs ),
    .X(uio_out[0]));
 sg13g2_buf_1 _857_ (.A(net57),
    .X(uio_out[3]));
 sg13g2_buf_1 _858_ (.A(\top_instance.green_led ),
    .X(uo_out[0]));
 sg13g2_buf_1 _859_ (.A(\top_instance.pulse_generator_inst.red_led ),
    .X(uo_out[1]));
 sg13g2_buf_2 fanout57 (.A(\top_instance.adc_inst.sclk ),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(\top_instance.adc_inst.sclk ),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(net60),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(net61),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(net63),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(net231),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(net250),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(net66),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(net66),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_112_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(net71),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(net71),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(net71),
    .X(net69));
 sg13g2_buf_1 fanout70 (.A(net71),
    .X(net70));
 sg13g2_buf_1 fanout71 (.A(rst_n),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(net73),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(rst_n),
    .X(net74));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_tielo tt_um_ephrenm_tsal_10 (.L_LO(net10));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\top_instance.comparator_inst.green_enable ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold2 (.A(\top_instance.comparator_inst.in[1] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold3 (.A(_075_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold4 (.A(\top_instance.comparator_inst.in[0] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold5 (.A(_074_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold6 (.A(\top_instance.comparator_inst.in[5] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold7 (.A(_079_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold8 (.A(\top_instance.comparator_inst.in[2] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold9 (.A(_076_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold10 (.A(\top_instance.comparator_inst.in[7] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold11 (.A(_081_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold12 (.A(\top_instance.comparator_inst.in[4] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold13 (.A(_078_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold14 (.A(\top_instance.comparator_inst.in[6] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold15 (.A(_080_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold16 (.A(_001_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold17 (.A(_049_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold18 (.A(\top_instance.comparator_inst.in[3] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold19 (.A(_077_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold20 (.A(_003_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold21 (.A(_010_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold22 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[9] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold23 (.A(_220_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold24 (.A(_059_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold25 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[19] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold26 (.A(_239_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold27 (.A(_069_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold28 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[13] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold29 (.A(_227_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold30 (.A(_007_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold31 (.A(_155_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold32 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[7] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold33 (.A(_216_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold34 (.A(\top_instance.adc_inst.bit_counter[5] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold35 (.A(_191_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold36 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[16] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold37 (.A(_233_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold38 (.A(_066_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold39 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[23] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold40 (.A(_073_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold41 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[1] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold42 (.A(_204_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold43 (.A(_051_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold44 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[12] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold45 (.A(_062_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold46 (.A(\top_instance.adc_inst.bit_counter[2] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold47 (.A(_181_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold48 (.A(\top_instance.adc_inst.clk_counter[0] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold49 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[21] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold50 (.A(_242_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold51 (.A(_071_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold52 (.A(\top_instance.comparator_inst.comp_reg[7] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold53 (.A(_002_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold54 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[4] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold55 (.A(_210_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold56 (.A(_054_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold57 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[2] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold58 (.A(_207_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold59 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[17] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold60 (.A(_235_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold61 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[0] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold62 (.A(_050_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold63 (.A(\top_instance.comparator_inst.comp_reg[1] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold64 (.A(\top_instance.adc_inst.clk_counter[3] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold65 (.A(_195_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold66 (.A(_044_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold67 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[3] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold68 (.A(_053_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold69 (.A(\top_instance.comparator_inst.comp_reg[0] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold70 (.A(\top_instance.adc_inst.bit_counter[4] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold71 (.A(_039_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold72 (.A(\top_instance.comparator_inst.comp_reg[6] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold73 (.A(_164_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold74 (.A(_021_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold75 (.A(\top_instance.comparator_inst.comp_reg[3] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold76 (.A(\top_instance.adc_inst.clk_counter[7] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold77 (.A(_154_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold78 (.A(\top_instance.adc_inst.clk_counter[4] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold79 (.A(_138_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold80 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[11] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold81 (.A(_224_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold82 (.A(_004_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold83 (.A(_048_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold84 (.A(\top_instance.comparator_inst.comp_reg[4] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold85 (.A(\top_instance.comparator_inst.comp_reg[2] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold86 (.A(\top_instance.adc_inst.bit_counter[3] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold87 (.A(\top_instance.comparator_inst.comp_reg[5] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold88 (.A(\top_instance.adc_inst.clk_counter[9] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold89 (.A(\top_instance.adc_inst.bit_counter[0] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold90 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[15] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold91 (.A(_232_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold92 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[6] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold93 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[20] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold94 (.A(_070_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold95 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[18] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold96 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[10] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold97 (.A(_223_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold98 (.A(_060_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold99 (.A(\top_instance.adc_inst.cs ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold100 (.A(\top_instance.adc_inst.data_ready ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold101 (.A(\top_instance.adc_inst.clk_counter[1] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold102 (.A(\top_instance.comparator_inst.input_reg[7] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold103 (.A(_000_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold104 (.A(\top_instance.adc_inst.bit_counter[1] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold105 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[5] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold106 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[8] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold107 (.A(_058_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold108 (.A(\top_instance.adc_inst.clk_counter[5] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold109 (.A(_196_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold110 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[22] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold111 (.A(_072_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold112 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[14] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold113 (.A(_230_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold114 (.A(_005_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold115 (.A(_153_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold116 (.A(_046_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold117 (.A(\top_instance.adc_inst.clk_counter[2] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold118 (.A(\top_instance.pulse_generator_inst.red_ctrl_counter[12] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold119 (.A(\top_instance.adc_inst.data_ready ),
    .X(net250));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_fill_2 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_4 FILLER_18_245 ();
 sg13g2_fill_2 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_fill_1 FILLER_18_263 ();
 sg13g2_decap_4 FILLER_18_277 ();
 sg13g2_fill_2 FILLER_18_281 ();
 sg13g2_fill_1 FILLER_18_287 ();
 sg13g2_decap_4 FILLER_18_296 ();
 sg13g2_fill_2 FILLER_18_304 ();
 sg13g2_fill_1 FILLER_18_306 ();
 sg13g2_decap_8 FILLER_18_310 ();
 sg13g2_decap_8 FILLER_18_317 ();
 sg13g2_decap_8 FILLER_18_324 ();
 sg13g2_decap_8 FILLER_18_331 ();
 sg13g2_decap_8 FILLER_18_338 ();
 sg13g2_decap_8 FILLER_18_345 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_359 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_decap_8 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_fill_2 FILLER_19_239 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_fill_1 FILLER_19_325 ();
 sg13g2_decap_8 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_decap_4 FILLER_19_344 ();
 sg13g2_fill_1 FILLER_19_348 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_4 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_227 ();
 sg13g2_fill_2 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_345 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_decap_8 FILLER_20_379 ();
 sg13g2_decap_8 FILLER_20_386 ();
 sg13g2_decap_8 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_175 ();
 sg13g2_fill_1 FILLER_21_202 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_fill_2 FILLER_21_239 ();
 sg13g2_fill_1 FILLER_21_241 ();
 sg13g2_fill_1 FILLER_21_268 ();
 sg13g2_fill_2 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_fill_1 FILLER_22_182 ();
 sg13g2_fill_2 FILLER_22_200 ();
 sg13g2_fill_1 FILLER_22_211 ();
 sg13g2_decap_4 FILLER_22_234 ();
 sg13g2_fill_1 FILLER_22_238 ();
 sg13g2_fill_2 FILLER_22_266 ();
 sg13g2_fill_2 FILLER_22_274 ();
 sg13g2_fill_1 FILLER_22_276 ();
 sg13g2_fill_2 FILLER_22_303 ();
 sg13g2_fill_2 FILLER_22_317 ();
 sg13g2_fill_2 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_4 FILLER_23_168 ();
 sg13g2_fill_2 FILLER_23_172 ();
 sg13g2_fill_2 FILLER_23_200 ();
 sg13g2_fill_1 FILLER_23_244 ();
 sg13g2_fill_1 FILLER_23_261 ();
 sg13g2_fill_1 FILLER_23_278 ();
 sg13g2_fill_2 FILLER_23_331 ();
 sg13g2_fill_1 FILLER_23_333 ();
 sg13g2_fill_1 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_380 ();
 sg13g2_decap_8 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_fill_2 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_4 FILLER_24_147 ();
 sg13g2_fill_1 FILLER_24_151 ();
 sg13g2_decap_8 FILLER_24_156 ();
 sg13g2_decap_8 FILLER_24_163 ();
 sg13g2_fill_1 FILLER_24_170 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_fill_2 FILLER_24_327 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_fill_2 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_90 ();
 sg13g2_decap_8 FILLER_25_97 ();
 sg13g2_decap_4 FILLER_25_104 ();
 sg13g2_fill_2 FILLER_25_125 ();
 sg13g2_fill_1 FILLER_25_141 ();
 sg13g2_fill_2 FILLER_25_198 ();
 sg13g2_fill_1 FILLER_25_205 ();
 sg13g2_fill_2 FILLER_25_257 ();
 sg13g2_fill_2 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_321 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_decap_8 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_4 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_67 ();
 sg13g2_fill_2 FILLER_26_72 ();
 sg13g2_fill_1 FILLER_26_74 ();
 sg13g2_fill_1 FILLER_26_79 ();
 sg13g2_fill_1 FILLER_26_89 ();
 sg13g2_fill_2 FILLER_26_145 ();
 sg13g2_fill_1 FILLER_26_147 ();
 sg13g2_fill_1 FILLER_26_166 ();
 sg13g2_fill_2 FILLER_26_171 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_decap_4 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_183 ();
 sg13g2_fill_2 FILLER_26_210 ();
 sg13g2_fill_1 FILLER_26_226 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_fill_2 FILLER_26_297 ();
 sg13g2_fill_2 FILLER_26_325 ();
 sg13g2_fill_2 FILLER_26_334 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_90 ();
 sg13g2_fill_1 FILLER_27_145 ();
 sg13g2_fill_1 FILLER_27_168 ();
 sg13g2_fill_2 FILLER_27_189 ();
 sg13g2_fill_2 FILLER_27_246 ();
 sg13g2_fill_2 FILLER_27_298 ();
 sg13g2_fill_1 FILLER_27_309 ();
 sg13g2_fill_2 FILLER_27_319 ();
 sg13g2_decap_8 FILLER_27_361 ();
 sg13g2_decap_8 FILLER_27_368 ();
 sg13g2_decap_8 FILLER_27_375 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_94 ();
 sg13g2_fill_1 FILLER_28_96 ();
 sg13g2_fill_1 FILLER_28_126 ();
 sg13g2_fill_2 FILLER_28_141 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_fill_1 FILLER_28_183 ();
 sg13g2_fill_2 FILLER_28_193 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_309 ();
 sg13g2_fill_1 FILLER_28_314 ();
 sg13g2_decap_8 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_4 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_67 ();
 sg13g2_decap_4 FILLER_29_81 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_139 ();
 sg13g2_fill_1 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_173 ();
 sg13g2_fill_2 FILLER_29_211 ();
 sg13g2_fill_1 FILLER_29_213 ();
 sg13g2_fill_2 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_254 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_267 ();
 sg13g2_fill_2 FILLER_29_282 ();
 sg13g2_fill_1 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_316 ();
 sg13g2_fill_2 FILLER_29_347 ();
 sg13g2_fill_1 FILLER_29_349 ();
 sg13g2_fill_2 FILLER_29_376 ();
 sg13g2_fill_2 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_1 FILLER_30_145 ();
 sg13g2_fill_2 FILLER_30_155 ();
 sg13g2_fill_1 FILLER_30_157 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_decap_4 FILLER_30_197 ();
 sg13g2_decap_8 FILLER_30_205 ();
 sg13g2_decap_4 FILLER_30_212 ();
 sg13g2_decap_4 FILLER_30_294 ();
 sg13g2_fill_2 FILLER_30_298 ();
 sg13g2_fill_1 FILLER_30_304 ();
 sg13g2_decap_8 FILLER_30_309 ();
 sg13g2_fill_2 FILLER_30_327 ();
 sg13g2_fill_1 FILLER_30_337 ();
 sg13g2_decap_4 FILLER_30_346 ();
 sg13g2_fill_1 FILLER_30_350 ();
 sg13g2_fill_2 FILLER_30_356 ();
 sg13g2_fill_2 FILLER_30_367 ();
 sg13g2_fill_1 FILLER_30_369 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_175 ();
 sg13g2_decap_4 FILLER_31_180 ();
 sg13g2_fill_1 FILLER_31_184 ();
 sg13g2_decap_4 FILLER_31_221 ();
 sg13g2_fill_2 FILLER_31_225 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_fill_2 FILLER_31_245 ();
 sg13g2_fill_2 FILLER_31_263 ();
 sg13g2_fill_1 FILLER_31_265 ();
 sg13g2_decap_4 FILLER_31_270 ();
 sg13g2_fill_2 FILLER_31_274 ();
 sg13g2_fill_1 FILLER_31_283 ();
 sg13g2_fill_2 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_338 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_4 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_60 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_107 ();
 sg13g2_fill_1 FILLER_32_132 ();
 sg13g2_fill_2 FILLER_32_191 ();
 sg13g2_fill_2 FILLER_32_198 ();
 sg13g2_fill_2 FILLER_32_209 ();
 sg13g2_fill_1 FILLER_32_211 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_fill_1 FILLER_32_235 ();
 sg13g2_fill_2 FILLER_32_292 ();
 sg13g2_fill_2 FILLER_32_302 ();
 sg13g2_decap_8 FILLER_32_307 ();
 sg13g2_fill_2 FILLER_32_314 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_decap_4 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_325 ();
 sg13g2_fill_2 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_fill_2 FILLER_33_70 ();
 sg13g2_decap_4 FILLER_33_76 ();
 sg13g2_fill_2 FILLER_33_80 ();
 sg13g2_fill_2 FILLER_33_180 ();
 sg13g2_fill_1 FILLER_33_182 ();
 sg13g2_decap_4 FILLER_33_240 ();
 sg13g2_fill_2 FILLER_33_252 ();
 sg13g2_fill_1 FILLER_33_254 ();
 sg13g2_fill_2 FILLER_33_267 ();
 sg13g2_fill_1 FILLER_33_278 ();
 sg13g2_fill_1 FILLER_33_284 ();
 sg13g2_decap_4 FILLER_33_289 ();
 sg13g2_fill_2 FILLER_33_293 ();
 sg13g2_fill_2 FILLER_33_326 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_79 ();
 sg13g2_fill_1 FILLER_34_133 ();
 sg13g2_fill_2 FILLER_34_160 ();
 sg13g2_fill_2 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_199 ();
 sg13g2_fill_1 FILLER_34_215 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_230 ();
 sg13g2_fill_1 FILLER_34_273 ();
 sg13g2_fill_2 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_353 ();
 sg13g2_fill_2 FILLER_34_369 ();
 sg13g2_fill_2 FILLER_34_381 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_4 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_88 ();
 sg13g2_fill_2 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_290 ();
 sg13g2_fill_2 FILLER_35_297 ();
 sg13g2_fill_1 FILLER_35_299 ();
 sg13g2_fill_2 FILLER_35_314 ();
 sg13g2_fill_1 FILLER_35_346 ();
 sg13g2_fill_1 FILLER_35_383 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_fill_2 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_114 ();
 sg13g2_fill_2 FILLER_36_139 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_fill_2 FILLER_36_182 ();
 sg13g2_fill_1 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_fill_1 FILLER_36_212 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_105 ();
 sg13g2_fill_1 FILLER_37_107 ();
 sg13g2_decap_8 FILLER_37_128 ();
 sg13g2_fill_2 FILLER_37_135 ();
 sg13g2_decap_4 FILLER_37_144 ();
 sg13g2_fill_1 FILLER_37_148 ();
 sg13g2_decap_8 FILLER_37_157 ();
 sg13g2_decap_8 FILLER_37_164 ();
 sg13g2_decap_8 FILLER_37_171 ();
 sg13g2_decap_8 FILLER_37_178 ();
 sg13g2_decap_8 FILLER_37_185 ();
 sg13g2_decap_8 FILLER_37_192 ();
 sg13g2_decap_8 FILLER_37_202 ();
 sg13g2_decap_4 FILLER_37_209 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_fill_1 FILLER_37_297 ();
 sg13g2_fill_1 FILLER_37_322 ();
 sg13g2_fill_1 FILLER_37_332 ();
 sg13g2_fill_1 FILLER_37_360 ();
 sg13g2_fill_1 FILLER_37_387 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_155 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_179 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_decap_4 FILLER_38_220 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_233 ();
 sg13g2_decap_8 FILLER_38_240 ();
 sg13g2_decap_8 FILLER_38_251 ();
 sg13g2_fill_2 FILLER_38_258 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_fill_1 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_380 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net130;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net131;
 assign uio_oe[4] = net12;
 assign uio_oe[5] = net13;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net15;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
 assign uio_out[4] = net18;
 assign uio_out[5] = net19;
 assign uio_out[6] = net20;
 assign uio_out[7] = net21;
 assign uo_out[2] = net22;
 assign uo_out[3] = net23;
 assign uo_out[4] = net24;
 assign uo_out[5] = net25;
 assign uo_out[6] = net26;
 assign uo_out[7] = net27;
endmodule

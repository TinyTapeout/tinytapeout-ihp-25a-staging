module tt_um_alif (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire \lif1.adapt_threshold[0] ;
 wire \lif1.adapt_threshold[1] ;
 wire \lif1.adapt_threshold[2] ;
 wire \lif1.adapt_threshold[3] ;
 wire \lif1.adapt_threshold[4] ;
 wire \lif1.adapt_threshold[5] ;
 wire \lif1.adapt_threshold[6] ;
 wire \lif1.adapt_threshold[7] ;
 wire \lif1.spike ;
 wire \lif1.spike_counter[0] ;
 wire \lif1.spike_counter[1] ;
 wire \lif1.spike_counter[2] ;
 wire \lif1.spike_counter[3] ;
 wire \lif1.spike_counter[4] ;
 wire \lif1.spike_counter[5] ;
 wire \lif1.spike_counter[6] ;
 wire \lif1.spike_counter[7] ;
 wire \lif2.adapt_threshold[0] ;
 wire \lif2.adapt_threshold[1] ;
 wire \lif2.adapt_threshold[2] ;
 wire \lif2.adapt_threshold[3] ;
 wire \lif2.adapt_threshold[4] ;
 wire \lif2.adapt_threshold[5] ;
 wire \lif2.adapt_threshold[6] ;
 wire \lif2.adapt_threshold[7] ;
 wire \lif2.spike ;
 wire \lif2.spike_counter[0] ;
 wire \lif2.spike_counter[1] ;
 wire \lif2.spike_counter[2] ;
 wire \lif2.spike_counter[3] ;
 wire \lif2.spike_counter[4] ;
 wire \lif2.spike_counter[5] ;
 wire \lif2.spike_counter[6] ;
 wire \lif2.spike_counter[7] ;
 wire \lif2.state[0] ;
 wire \lif2.state[1] ;
 wire \lif2.state[2] ;
 wire \lif2.state[3] ;
 wire \lif2.state[4] ;
 wire \lif2.state[5] ;
 wire \lif2.state[6] ;
 wire \lif2.state[7] ;
 wire \lif3.adapt_threshold[0] ;
 wire \lif3.adapt_threshold[1] ;
 wire \lif3.adapt_threshold[2] ;
 wire \lif3.adapt_threshold[3] ;
 wire \lif3.adapt_threshold[4] ;
 wire \lif3.adapt_threshold[5] ;
 wire \lif3.adapt_threshold[6] ;
 wire \lif3.adapt_threshold[7] ;
 wire \lif3.spike ;
 wire \lif3.spike_counter[0] ;
 wire \lif3.spike_counter[1] ;
 wire \lif3.spike_counter[2] ;
 wire \lif3.spike_counter[3] ;
 wire \lif3.spike_counter[4] ;
 wire \lif3.spike_counter[5] ;
 wire \lif3.spike_counter[6] ;
 wire \lif3.spike_counter[7] ;
 wire \lif3.state[0] ;
 wire \lif3.state[1] ;
 wire \lif3.state[2] ;
 wire \lif3.state[3] ;
 wire \lif3.state[4] ;
 wire \lif3.state[5] ;
 wire \lif3.state[6] ;
 wire \lif3.state[7] ;
 wire clknet_0_clk;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;

 sg13g2_inv_1 _0877_ (.Y(_0094_),
    .A(\lif2.adapt_threshold[7] ));
 sg13g2_inv_1 _0878_ (.Y(_0095_),
    .A(\lif2.adapt_threshold[6] ));
 sg13g2_inv_1 _0879_ (.Y(_0096_),
    .A(\lif2.adapt_threshold[5] ));
 sg13g2_inv_1 _0880_ (.Y(_0097_),
    .A(\lif2.adapt_threshold[4] ));
 sg13g2_inv_1 _0881_ (.Y(_0098_),
    .A(net202));
 sg13g2_inv_1 _0882_ (.Y(_0099_),
    .A(\lif1.adapt_threshold[7] ));
 sg13g2_inv_1 _0883_ (.Y(_0100_),
    .A(\lif1.adapt_threshold[5] ));
 sg13g2_inv_1 _0884_ (.Y(_0101_),
    .A(\lif1.adapt_threshold[4] ));
 sg13g2_inv_1 _0885_ (.Y(_0102_),
    .A(\lif1.adapt_threshold[3] ));
 sg13g2_inv_1 _0886_ (.Y(_0103_),
    .A(net207));
 sg13g2_inv_1 _0887_ (.Y(_0104_),
    .A(net208));
 sg13g2_inv_1 _0888_ (.Y(_0105_),
    .A(\lif3.adapt_threshold[6] ));
 sg13g2_inv_1 _0889_ (.Y(_0106_),
    .A(\lif3.adapt_threshold[5] ));
 sg13g2_inv_1 _0890_ (.Y(_0107_),
    .A(\lif3.adapt_threshold[4] ));
 sg13g2_inv_1 _0891_ (.Y(_0108_),
    .A(\lif3.adapt_threshold[3] ));
 sg13g2_inv_1 _0892_ (.Y(_0109_),
    .A(\lif3.adapt_threshold[2] ));
 sg13g2_inv_1 _0893_ (.Y(_0110_),
    .A(\lif3.adapt_threshold[1] ));
 sg13g2_inv_1 _0894_ (.Y(_0111_),
    .A(uo_out[1]));
 sg13g2_inv_1 _0895_ (.Y(_0112_),
    .A(uo_out[2]));
 sg13g2_inv_1 _0896_ (.Y(_0113_),
    .A(uo_out[7]));
 sg13g2_inv_1 _0897_ (.Y(_0114_),
    .A(uo_out[6]));
 sg13g2_inv_1 _0898_ (.Y(_0115_),
    .A(\lif3.state[2] ));
 sg13g2_inv_1 _0899_ (.Y(_0116_),
    .A(\lif3.spike_counter[5] ));
 sg13g2_inv_1 _0900_ (.Y(_0117_),
    .A(\lif2.state[1] ));
 sg13g2_inv_1 _0901_ (.Y(_0118_),
    .A(\lif2.state[3] ));
 sg13g2_inv_1 _0902_ (.Y(_0119_),
    .A(net92));
 sg13g2_inv_1 _0903_ (.Y(_0120_),
    .A(\lif2.state[7] ));
 sg13g2_inv_2 _0904_ (.Y(_0121_),
    .A(\lif2.state[6] ));
 sg13g2_inv_1 _0905_ (.Y(_0122_),
    .A(net91));
 sg13g2_inv_1 _0906_ (.Y(_0123_),
    .A(\lif2.state[4] ));
 sg13g2_inv_1 _0907_ (.Y(_0124_),
    .A(\lif3.state[7] ));
 sg13g2_inv_1 _0908_ (.Y(_0125_),
    .A(net99));
 sg13g2_inv_1 _0909_ (.Y(_0126_),
    .A(\lif3.state[5] ));
 sg13g2_inv_1 _0910_ (.Y(_0127_),
    .A(\lif3.state[4] ));
 sg13g2_inv_1 _0911_ (.Y(_0128_),
    .A(\lif3.state[3] ));
 sg13g2_inv_1 _0912_ (.Y(_0129_),
    .A(\lif3.state[1] ));
 sg13g2_inv_1 _0913_ (.Y(_0130_),
    .A(\lif3.state[0] ));
 sg13g2_inv_1 _0914_ (.Y(_0131_),
    .A(\lif2.spike_counter[6] ));
 sg13g2_inv_1 _0915_ (.Y(_0132_),
    .A(\lif1.spike_counter[5] ));
 sg13g2_inv_1 _0916_ (.Y(_0133_),
    .A(net106));
 sg13g2_inv_1 _0917_ (.Y(_0134_),
    .A(net8));
 sg13g2_inv_1 _0918_ (.Y(_0135_),
    .A(net7));
 sg13g2_inv_1 _0919_ (.Y(_0136_),
    .A(net120));
 sg13g2_nand2b_1 _0920_ (.Y(_0137_),
    .B(uo_out[6]),
    .A_N(\lif1.adapt_threshold[6] ));
 sg13g2_nor2_1 _0921_ (.A(_0100_),
    .B(uo_out[5]),
    .Y(_0138_));
 sg13g2_o21ai_1 _0922_ (.B1(\lif1.adapt_threshold[0] ),
    .Y(_0139_),
    .A1(\lif1.adapt_threshold[1] ),
    .A2(_0111_));
 sg13g2_a22oi_1 _0923_ (.Y(_0140_),
    .B1(_0112_),
    .B2(\lif1.adapt_threshold[2] ),
    .A2(_0111_),
    .A1(\lif1.adapt_threshold[1] ));
 sg13g2_o21ai_1 _0924_ (.B1(_0140_),
    .Y(_0141_),
    .A1(uo_out[0]),
    .A2(_0139_));
 sg13g2_a22oi_1 _0925_ (.Y(_0142_),
    .B1(uo_out[2]),
    .B2(_0103_),
    .A2(net97),
    .A1(_0102_));
 sg13g2_nand2b_1 _0926_ (.Y(_0143_),
    .B(\lif1.adapt_threshold[3] ),
    .A_N(net97));
 sg13g2_o21ai_1 _0927_ (.B1(_0143_),
    .Y(_0144_),
    .A1(_0101_),
    .A2(uo_out[4]));
 sg13g2_a21oi_1 _0928_ (.A1(_0141_),
    .A2(_0142_),
    .Y(_0145_),
    .B1(_0144_));
 sg13g2_a221oi_1 _0929_ (.B2(_0101_),
    .C1(_0145_),
    .B1(uo_out[4]),
    .A1(_0100_),
    .Y(_0146_),
    .A2(uo_out[5]));
 sg13g2_o21ai_1 _0930_ (.B1(_0137_),
    .Y(_0147_),
    .A1(_0138_),
    .A2(_0146_));
 sg13g2_a22oi_1 _0931_ (.Y(_0148_),
    .B1(_0114_),
    .B2(\lif1.adapt_threshold[6] ),
    .A2(_0113_),
    .A1(\lif1.adapt_threshold[7] ));
 sg13g2_a22oi_1 _0932_ (.Y(_0149_),
    .B1(_0147_),
    .B2(_0148_),
    .A2(uo_out[7]),
    .A1(_0099_));
 sg13g2_inv_1 _0933_ (.Y(\lif1.spike ),
    .A(_0149_));
 sg13g2_nor2b_1 _0934_ (.A(\lif2.state[0] ),
    .B_N(\lif2.adapt_threshold[0] ),
    .Y(_0150_));
 sg13g2_o21ai_1 _0935_ (.B1(_0150_),
    .Y(_0151_),
    .A1(\lif2.adapt_threshold[1] ),
    .A2(_0117_));
 sg13g2_a22oi_1 _0936_ (.Y(_0152_),
    .B1(_0119_),
    .B2(\lif2.adapt_threshold[2] ),
    .A2(_0117_),
    .A1(\lif2.adapt_threshold[1] ));
 sg13g2_nor2_1 _0937_ (.A(\lif2.adapt_threshold[3] ),
    .B(_0118_),
    .Y(_0153_));
 sg13g2_a221oi_1 _0938_ (.B2(_0152_),
    .C1(_0153_),
    .B1(_0151_),
    .A1(_0098_),
    .Y(_0154_),
    .A2(net92));
 sg13g2_a221oi_1 _0939_ (.B2(\lif2.adapt_threshold[4] ),
    .C1(_0154_),
    .B1(_0123_),
    .A1(\lif2.adapt_threshold[3] ),
    .Y(_0155_),
    .A2(_0118_));
 sg13g2_a221oi_1 _0940_ (.B2(_0097_),
    .C1(_0155_),
    .B1(\lif2.state[4] ),
    .A1(_0096_),
    .Y(_0156_),
    .A2(net91));
 sg13g2_a221oi_1 _0941_ (.B2(\lif2.adapt_threshold[5] ),
    .C1(_0156_),
    .B1(_0122_),
    .A1(\lif2.adapt_threshold[6] ),
    .Y(_0157_),
    .A2(_0121_));
 sg13g2_a221oi_1 _0942_ (.B2(_0095_),
    .C1(_0157_),
    .B1(\lif2.state[6] ),
    .A1(_0094_),
    .Y(_0158_),
    .A2(\lif2.state[7] ));
 sg13g2_a21oi_1 _0943_ (.A1(\lif2.adapt_threshold[7] ),
    .A2(_0120_),
    .Y(\lif2.spike ),
    .B1(_0158_));
 sg13g2_a22oi_1 _0944_ (.Y(_0159_),
    .B1(_0130_),
    .B2(\lif3.adapt_threshold[0] ),
    .A2(_0129_),
    .A1(\lif3.adapt_threshold[1] ));
 sg13g2_a221oi_1 _0945_ (.B2(_0110_),
    .C1(_0159_),
    .B1(\lif3.state[1] ),
    .A1(_0109_),
    .Y(_0160_),
    .A2(\lif3.state[2] ));
 sg13g2_a221oi_1 _0946_ (.B2(\lif3.adapt_threshold[3] ),
    .C1(_0160_),
    .B1(_0128_),
    .A1(\lif3.adapt_threshold[2] ),
    .Y(_0161_),
    .A2(_0115_));
 sg13g2_a221oi_1 _0947_ (.B2(_0108_),
    .C1(_0161_),
    .B1(\lif3.state[3] ),
    .A1(_0107_),
    .Y(_0162_),
    .A2(\lif3.state[4] ));
 sg13g2_a221oi_1 _0948_ (.B2(\lif3.adapt_threshold[4] ),
    .C1(_0162_),
    .B1(_0127_),
    .A1(\lif3.adapt_threshold[5] ),
    .Y(_0163_),
    .A2(_0126_));
 sg13g2_a221oi_1 _0949_ (.B2(_0106_),
    .C1(_0163_),
    .B1(net100),
    .A1(_0105_),
    .Y(_0164_),
    .A2(net99));
 sg13g2_a221oi_1 _0950_ (.B2(\lif3.adapt_threshold[6] ),
    .C1(_0164_),
    .B1(_0125_),
    .A1(\lif3.adapt_threshold[7] ),
    .Y(_0165_),
    .A2(_0124_));
 sg13g2_a21oi_2 _0951_ (.B1(_0165_),
    .Y(_0166_),
    .A2(\lif3.state[7] ),
    .A1(_0104_));
 sg13g2_inv_1 _0952_ (.Y(\lif3.spike ),
    .A(_0166_));
 sg13g2_nor2_1 _0953_ (.A(\lif3.spike_counter[4] ),
    .B(\lif3.spike_counter[3] ),
    .Y(_0167_));
 sg13g2_a21oi_1 _0954_ (.A1(\lif3.spike_counter[2] ),
    .A2(\lif3.spike_counter[1] ),
    .Y(_0168_),
    .B1(\lif3.spike_counter[6] ));
 sg13g2_nand4_1 _0955_ (.B(_0004_),
    .C(_0167_),
    .A(_0116_),
    .Y(_0169_),
    .D(_0168_));
 sg13g2_nand2_1 _0956_ (.Y(_0170_),
    .A(\lif3.adapt_threshold[1] ),
    .B(\lif3.adapt_threshold[0] ));
 sg13g2_nor2_1 _0957_ (.A(\lif3.adapt_threshold[3] ),
    .B(\lif3.adapt_threshold[2] ),
    .Y(_0171_));
 sg13g2_nand2_1 _0958_ (.Y(_0172_),
    .A(\lif3.adapt_threshold[5] ),
    .B(\lif3.adapt_threshold[4] ));
 sg13g2_a21oi_1 _0959_ (.A1(_0170_),
    .A2(_0171_),
    .Y(_0173_),
    .B1(_0172_));
 sg13g2_nand2_1 _0960_ (.Y(_0174_),
    .A(_0104_),
    .B(_0105_));
 sg13g2_o21ai_1 _0961_ (.B1(_0169_),
    .Y(_0175_),
    .A1(_0173_),
    .A2(_0174_));
 sg13g2_nand2_1 _0962_ (.Y(_0176_),
    .A(_0109_),
    .B(_0110_));
 sg13g2_nand3_1 _0963_ (.B(\lif3.adapt_threshold[3] ),
    .C(_0176_),
    .A(_0107_),
    .Y(_0177_));
 sg13g2_a21oi_1 _0964_ (.A1(_0013_),
    .A2(_0177_),
    .Y(_0178_),
    .B1(_0106_));
 sg13g2_nor2_1 _0965_ (.A(\lif3.adapt_threshold[6] ),
    .B(_0178_),
    .Y(_0179_));
 sg13g2_nor2_1 _0966_ (.A(_0104_),
    .B(_0179_),
    .Y(_0180_));
 sg13g2_o21ai_1 _0967_ (.B1(net90),
    .Y(_0181_),
    .A1(_0166_),
    .A2(_0180_));
 sg13g2_inv_1 _0968_ (.Y(_0182_),
    .A(_0181_));
 sg13g2_mux2_1 _0969_ (.A0(\lif3.spike_counter[3] ),
    .A1(_0003_),
    .S(_0175_),
    .X(_0183_));
 sg13g2_nand2b_1 _0970_ (.Y(_0184_),
    .B(net150),
    .A_N(_0183_));
 sg13g2_xnor2_1 _0971_ (.Y(_0185_),
    .A(net150),
    .B(_0183_));
 sg13g2_o21ai_1 _0972_ (.B1(net107),
    .Y(_0186_),
    .A1(\lif3.adapt_threshold[0] ),
    .A2(_0181_));
 sg13g2_a21oi_1 _0973_ (.A1(_0181_),
    .A2(net151),
    .Y(_0022_),
    .B1(_0186_));
 sg13g2_nand2_1 _0974_ (.Y(_0187_),
    .A(net147),
    .B(\lif3.spike_counter[3] ));
 sg13g2_nand2b_1 _0975_ (.Y(_0188_),
    .B(_0187_),
    .A_N(_0167_));
 sg13g2_nor2_2 _0976_ (.A(\lif3.state[2] ),
    .B(\lif3.state[3] ),
    .Y(_0189_));
 sg13g2_nand2_2 _0977_ (.Y(_0190_),
    .A(\lif3.state[2] ),
    .B(\lif3.state[3] ));
 sg13g2_xor2_1 _0978_ (.B(\lif3.state[3] ),
    .A(\lif3.state[2] ),
    .X(_0191_));
 sg13g2_nand2b_1 _0979_ (.Y(_0192_),
    .B(_0190_),
    .A_N(_0189_));
 sg13g2_mux2_1 _0980_ (.A0(_0188_),
    .A1(_0192_),
    .S(_0175_),
    .X(_0193_));
 sg13g2_and2_1 _0981_ (.A(\lif3.adapt_threshold[1] ),
    .B(_0193_),
    .X(_0194_));
 sg13g2_xnor2_1 _0982_ (.Y(_0195_),
    .A(_0110_),
    .B(_0193_));
 sg13g2_xnor2_1 _0983_ (.Y(_0196_),
    .A(_0184_),
    .B(_0195_));
 sg13g2_a21oi_1 _0984_ (.A1(net175),
    .A2(_0182_),
    .Y(_0197_),
    .B1(net103));
 sg13g2_o21ai_1 _0985_ (.B1(_0197_),
    .Y(_0023_),
    .A1(_0182_),
    .A2(_0196_));
 sg13g2_a21oi_1 _0986_ (.A1(_0184_),
    .A2(_0195_),
    .Y(_0198_),
    .B1(_0194_));
 sg13g2_nand3_1 _0987_ (.B(\lif3.spike_counter[4] ),
    .C(\lif3.spike_counter[3] ),
    .A(net153),
    .Y(_0199_));
 sg13g2_xnor2_1 _0988_ (.Y(_0200_),
    .A(_0116_),
    .B(_0187_));
 sg13g2_nand2_1 _0989_ (.Y(_0201_),
    .A(_0127_),
    .B(_0189_));
 sg13g2_o21ai_1 _0990_ (.B1(\lif3.state[4] ),
    .Y(_0202_),
    .A1(\lif3.state[2] ),
    .A2(\lif3.state[3] ));
 sg13g2_nand2_1 _0991_ (.Y(_0203_),
    .A(_0201_),
    .B(_0202_));
 sg13g2_mux2_1 _0992_ (.A0(_0200_),
    .A1(_0203_),
    .S(net90),
    .X(_0204_));
 sg13g2_xnor2_1 _0993_ (.Y(_0205_),
    .A(_0015_),
    .B(_0204_));
 sg13g2_inv_1 _0994_ (.Y(_0206_),
    .A(_0205_));
 sg13g2_xnor2_1 _0995_ (.Y(_0207_),
    .A(_0198_),
    .B(_0206_));
 sg13g2_o21ai_1 _0996_ (.B1(net107),
    .Y(_0208_),
    .A1(net189),
    .A2(_0181_));
 sg13g2_a21oi_1 _0997_ (.A1(_0181_),
    .A2(_0207_),
    .Y(_0024_),
    .B1(_0208_));
 sg13g2_nand2_1 _0998_ (.Y(_0209_),
    .A(\lif3.adapt_threshold[2] ),
    .B(_0204_));
 sg13g2_o21ai_1 _0999_ (.B1(_0209_),
    .Y(_0210_),
    .A1(_0198_),
    .A2(_0206_));
 sg13g2_xnor2_1 _1000_ (.Y(_0211_),
    .A(_0014_),
    .B(_0199_));
 sg13g2_nand3_1 _1001_ (.B(_0127_),
    .C(_0189_),
    .A(_0126_),
    .Y(_0212_));
 sg13g2_nand2_1 _1002_ (.Y(_0213_),
    .A(\lif3.state[5] ),
    .B(_0201_));
 sg13g2_nand3_1 _1003_ (.B(_0212_),
    .C(_0213_),
    .A(net90),
    .Y(_0214_));
 sg13g2_o21ai_1 _1004_ (.B1(_0214_),
    .Y(_0215_),
    .A1(net90),
    .A2(_0211_));
 sg13g2_nor2_1 _1005_ (.A(_0016_),
    .B(_0215_),
    .Y(_0216_));
 sg13g2_nand2_1 _1006_ (.Y(_0217_),
    .A(_0016_),
    .B(_0215_));
 sg13g2_nand2b_1 _1007_ (.Y(_0218_),
    .B(_0217_),
    .A_N(_0216_));
 sg13g2_xor2_1 _1008_ (.B(_0218_),
    .A(_0210_),
    .X(_0219_));
 sg13g2_a21oi_1 _1009_ (.A1(net176),
    .A2(_0182_),
    .Y(_0220_),
    .B1(net103));
 sg13g2_o21ai_1 _1010_ (.B1(_0220_),
    .Y(_0025_),
    .A1(net83),
    .A2(_0219_));
 sg13g2_a21oi_1 _1011_ (.A1(_0210_),
    .A2(_0217_),
    .Y(_0221_),
    .B1(_0216_));
 sg13g2_nand4_1 _1012_ (.B(\lif3.spike_counter[5] ),
    .C(\lif3.spike_counter[4] ),
    .A(\lif3.spike_counter[6] ),
    .Y(_0222_),
    .D(\lif3.spike_counter[3] ));
 sg13g2_xnor2_1 _1013_ (.Y(_0223_),
    .A(_0004_),
    .B(_0222_));
 sg13g2_nor2_1 _1014_ (.A(net90),
    .B(_0223_),
    .Y(_0224_));
 sg13g2_nand2b_1 _1015_ (.Y(_0225_),
    .B(_0125_),
    .A_N(_0212_));
 sg13g2_xnor2_1 _1016_ (.Y(_0226_),
    .A(_0125_),
    .B(_0212_));
 sg13g2_a21oi_1 _1017_ (.A1(net90),
    .A2(_0226_),
    .Y(_0227_),
    .B1(_0224_));
 sg13g2_xor2_1 _1018_ (.B(_0227_),
    .A(_0013_),
    .X(_0228_));
 sg13g2_xnor2_1 _1019_ (.Y(_0229_),
    .A(_0221_),
    .B(_0228_));
 sg13g2_a21oi_1 _1020_ (.A1(net173),
    .A2(net83),
    .Y(_0230_),
    .B1(net103));
 sg13g2_o21ai_1 _1021_ (.B1(_0230_),
    .Y(_0026_),
    .A1(net83),
    .A2(_0229_));
 sg13g2_nor2_1 _1022_ (.A(\lif3.state[7] ),
    .B(net99),
    .Y(_0231_));
 sg13g2_o21ai_1 _1023_ (.B1(net90),
    .Y(_0232_),
    .A1(\lif3.state[7] ),
    .A2(_0225_));
 sg13g2_a21o_1 _1024_ (.A2(_0225_),
    .A1(\lif3.state[7] ),
    .B1(_0232_),
    .X(_0233_));
 sg13g2_or3_1 _1025_ (.A(_0004_),
    .B(net90),
    .C(_0222_),
    .X(_0234_));
 sg13g2_nand3_1 _1026_ (.B(_0233_),
    .C(_0234_),
    .A(\lif3.adapt_threshold[5] ),
    .Y(_0235_));
 sg13g2_a21o_1 _1027_ (.A2(_0234_),
    .A1(_0233_),
    .B1(\lif3.adapt_threshold[5] ),
    .X(_0236_));
 sg13g2_nand2_1 _1028_ (.Y(_0237_),
    .A(_0235_),
    .B(_0236_));
 sg13g2_nand2_1 _1029_ (.Y(_0238_),
    .A(\lif3.adapt_threshold[4] ),
    .B(_0227_));
 sg13g2_o21ai_1 _1030_ (.B1(_0238_),
    .Y(_0239_),
    .A1(_0221_),
    .A2(_0228_));
 sg13g2_xor2_1 _1031_ (.B(_0239_),
    .A(_0237_),
    .X(_0240_));
 sg13g2_a21oi_1 _1032_ (.A1(net191),
    .A2(net83),
    .Y(_0241_),
    .B1(net104));
 sg13g2_o21ai_1 _1033_ (.B1(_0241_),
    .Y(_0027_),
    .A1(net83),
    .A2(_0240_));
 sg13g2_xnor2_1 _1034_ (.Y(_0242_),
    .A(\lif3.adapt_threshold[6] ),
    .B(_0232_));
 sg13g2_nand2_1 _1035_ (.Y(_0243_),
    .A(_0236_),
    .B(_0239_));
 sg13g2_a21oi_1 _1036_ (.A1(_0235_),
    .A2(_0243_),
    .Y(_0244_),
    .B1(_0242_));
 sg13g2_nand3_1 _1037_ (.B(_0242_),
    .C(_0243_),
    .A(_0235_),
    .Y(_0245_));
 sg13g2_nand2_1 _1038_ (.Y(_0246_),
    .A(_0181_),
    .B(_0245_));
 sg13g2_a21oi_1 _1039_ (.A1(net194),
    .A2(net83),
    .Y(_0247_),
    .B1(net104));
 sg13g2_o21ai_1 _1040_ (.B1(_0247_),
    .Y(_0028_),
    .A1(_0244_),
    .A2(_0246_));
 sg13g2_a21oi_1 _1041_ (.A1(\lif3.adapt_threshold[6] ),
    .A2(_0232_),
    .Y(_0248_),
    .B1(_0244_));
 sg13g2_xnor2_1 _1042_ (.Y(_0249_),
    .A(net178),
    .B(_0232_));
 sg13g2_xnor2_1 _1043_ (.Y(_0250_),
    .A(_0248_),
    .B(_0249_));
 sg13g2_a21oi_1 _1044_ (.A1(net178),
    .A2(net83),
    .Y(_0251_),
    .B1(net104));
 sg13g2_o21ai_1 _1045_ (.B1(_0251_),
    .Y(_0029_),
    .A1(net83),
    .A2(_0250_));
 sg13g2_nand2_1 _1046_ (.Y(_0252_),
    .A(\lif3.state[7] ),
    .B(net99));
 sg13g2_a21oi_1 _1047_ (.A1(net100),
    .A2(_0252_),
    .Y(_0253_),
    .B1(_0231_));
 sg13g2_nor2_1 _1048_ (.A(_0126_),
    .B(_0127_),
    .Y(_0254_));
 sg13g2_xor2_1 _1049_ (.B(\lif3.state[4] ),
    .A(net100),
    .X(_0255_));
 sg13g2_a21oi_1 _1050_ (.A1(\lif3.state[6] ),
    .A2(_0255_),
    .Y(_0256_),
    .B1(_0254_));
 sg13g2_xor2_1 _1051_ (.B(net100),
    .A(net99),
    .X(_0257_));
 sg13g2_xnor2_1 _1052_ (.Y(_0258_),
    .A(\lif3.state[7] ),
    .B(_0257_));
 sg13g2_and2_1 _1053_ (.A(_0256_),
    .B(_0258_),
    .X(_0259_));
 sg13g2_or2_1 _1054_ (.X(_0260_),
    .B(_0258_),
    .A(_0256_));
 sg13g2_xnor2_1 _1055_ (.Y(_0261_),
    .A(net99),
    .B(_0255_));
 sg13g2_nor2_1 _1056_ (.A(_0127_),
    .B(_0128_),
    .Y(_0262_));
 sg13g2_xor2_1 _1057_ (.B(\lif3.state[3] ),
    .A(\lif3.state[4] ),
    .X(_0263_));
 sg13g2_a21oi_1 _1058_ (.A1(net100),
    .A2(_0263_),
    .Y(_0264_),
    .B1(_0262_));
 sg13g2_nor2_1 _1059_ (.A(_0261_),
    .B(_0264_),
    .Y(_0265_));
 sg13g2_xnor2_1 _1060_ (.Y(_0266_),
    .A(net100),
    .B(_0263_));
 sg13g2_a21o_1 _1061_ (.A2(_0202_),
    .A1(_0190_),
    .B1(_0266_),
    .X(_0267_));
 sg13g2_nand3_1 _1062_ (.B(_0202_),
    .C(_0266_),
    .A(_0190_),
    .Y(_0268_));
 sg13g2_inv_1 _1063_ (.Y(_0269_),
    .A(_0268_));
 sg13g2_a21oi_1 _1064_ (.A1(_0129_),
    .A2(_0190_),
    .Y(_0270_),
    .B1(_0189_));
 sg13g2_xnor2_1 _1065_ (.Y(_0271_),
    .A(\lif3.state[4] ),
    .B(_0191_));
 sg13g2_nor2b_1 _1066_ (.A(_0271_),
    .B_N(_0270_),
    .Y(_0272_));
 sg13g2_nand3_1 _1067_ (.B(\lif3.state[3] ),
    .C(\lif3.state[1] ),
    .A(\lif3.state[2] ),
    .Y(_0273_));
 sg13g2_nor2_1 _1068_ (.A(\lif3.state[2] ),
    .B(\lif3.state[1] ),
    .Y(_0274_));
 sg13g2_nand2_1 _1069_ (.Y(_0275_),
    .A(_0128_),
    .B(\lif3.state[0] ));
 sg13g2_o21ai_1 _1070_ (.B1(_0273_),
    .Y(_0276_),
    .A1(_0274_),
    .A2(_0275_));
 sg13g2_xnor2_1 _1071_ (.Y(_0277_),
    .A(_0270_),
    .B(_0271_));
 sg13g2_a21oi_2 _1072_ (.B1(_0272_),
    .Y(_0278_),
    .A2(_0277_),
    .A1(_0276_));
 sg13g2_o21ai_1 _1073_ (.B1(_0267_),
    .Y(_0279_),
    .A1(_0269_),
    .A2(_0278_));
 sg13g2_xnor2_1 _1074_ (.Y(_0280_),
    .A(_0261_),
    .B(_0264_));
 sg13g2_inv_1 _1075_ (.Y(_0281_),
    .A(_0280_));
 sg13g2_a21oi_2 _1076_ (.B1(_0265_),
    .Y(_0282_),
    .A2(_0281_),
    .A1(_0279_));
 sg13g2_nor2b_1 _1077_ (.A(_0259_),
    .B_N(_0260_),
    .Y(_0283_));
 sg13g2_a21oi_2 _1078_ (.B1(_0259_),
    .Y(_0284_),
    .A2(_0282_),
    .A1(_0260_));
 sg13g2_xnor2_1 _1079_ (.Y(_0285_),
    .A(_0253_),
    .B(_0284_));
 sg13g2_nand2b_1 _1080_ (.Y(_0286_),
    .B(net7),
    .A_N(_0285_));
 sg13g2_a21o_1 _1081_ (.A2(_0252_),
    .A1(net100),
    .B1(_0284_),
    .X(_0287_));
 sg13g2_nor4_1 _1082_ (.A(_0124_),
    .B(net99),
    .C(net100),
    .D(_0284_),
    .Y(_0288_));
 sg13g2_a21oi_1 _1083_ (.A1(net99),
    .A2(_0287_),
    .Y(_0289_),
    .B1(_0288_));
 sg13g2_nand2b_1 _1084_ (.Y(_0290_),
    .B(net8),
    .A_N(_0289_));
 sg13g2_xnor2_1 _1085_ (.Y(_0291_),
    .A(net8),
    .B(_0289_));
 sg13g2_nand2b_1 _1086_ (.Y(_0292_),
    .B(_0291_),
    .A_N(_0286_));
 sg13g2_xor2_1 _1087_ (.B(_0291_),
    .A(_0286_),
    .X(_0293_));
 sg13g2_xnor2_1 _1088_ (.Y(_0294_),
    .A(_0282_),
    .B(_0283_));
 sg13g2_and2_1 _1089_ (.A(net6),
    .B(_0294_),
    .X(_0295_));
 sg13g2_xnor2_1 _1090_ (.Y(_0296_),
    .A(net7),
    .B(_0285_));
 sg13g2_nor2_1 _1091_ (.A(_0295_),
    .B(_0296_),
    .Y(_0297_));
 sg13g2_nand2_1 _1092_ (.Y(_0298_),
    .A(_0295_),
    .B(_0296_));
 sg13g2_xnor2_1 _1093_ (.Y(_0299_),
    .A(_0279_),
    .B(_0280_));
 sg13g2_nor2_1 _1094_ (.A(net5),
    .B(_0299_),
    .Y(_0300_));
 sg13g2_xnor2_1 _1095_ (.Y(_0301_),
    .A(net6),
    .B(_0294_));
 sg13g2_nor2_1 _1096_ (.A(_0300_),
    .B(_0301_),
    .Y(_0302_));
 sg13g2_nand2_1 _1097_ (.Y(_0303_),
    .A(_0267_),
    .B(_0268_));
 sg13g2_xor2_1 _1098_ (.B(_0303_),
    .A(_0278_),
    .X(_0304_));
 sg13g2_nand2_1 _1099_ (.Y(_0305_),
    .A(net4),
    .B(_0304_));
 sg13g2_xnor2_1 _1100_ (.Y(_0306_),
    .A(net5),
    .B(_0299_));
 sg13g2_nand2b_1 _1101_ (.Y(_0307_),
    .B(_0306_),
    .A_N(_0305_));
 sg13g2_xnor2_1 _1102_ (.Y(_0308_),
    .A(_0276_),
    .B(_0277_));
 sg13g2_nor2b_1 _1103_ (.A(net3),
    .B_N(_0308_),
    .Y(_0309_));
 sg13g2_xor2_1 _1104_ (.B(_0304_),
    .A(net4),
    .X(_0310_));
 sg13g2_nor2b_1 _1105_ (.A(_0309_),
    .B_N(_0310_),
    .Y(_0311_));
 sg13g2_nor2_1 _1106_ (.A(\lif3.state[0] ),
    .B(_0274_),
    .Y(_0312_));
 sg13g2_xnor2_1 _1107_ (.Y(_0313_),
    .A(_0128_),
    .B(_0312_));
 sg13g2_nand2_1 _1108_ (.Y(_0314_),
    .A(net2),
    .B(_0313_));
 sg13g2_xor2_1 _1109_ (.B(_0308_),
    .A(net3),
    .X(_0315_));
 sg13g2_nor2b_1 _1110_ (.A(_0314_),
    .B_N(_0315_),
    .Y(_0316_));
 sg13g2_xnor2_1 _1111_ (.Y(_0317_),
    .A(_0309_),
    .B(_0310_));
 sg13g2_a21oi_1 _1112_ (.A1(_0316_),
    .A2(_0317_),
    .Y(_0318_),
    .B1(_0311_));
 sg13g2_xor2_1 _1113_ (.B(_0306_),
    .A(_0305_),
    .X(_0319_));
 sg13g2_o21ai_1 _1114_ (.B1(_0307_),
    .Y(_0320_),
    .A1(_0318_),
    .A2(_0319_));
 sg13g2_xor2_1 _1115_ (.B(_0301_),
    .A(_0300_),
    .X(_0321_));
 sg13g2_a21oi_1 _1116_ (.A1(_0320_),
    .A2(_0321_),
    .Y(_0322_),
    .B1(_0302_));
 sg13g2_nor2b_1 _1117_ (.A(_0297_),
    .B_N(_0298_),
    .Y(_0323_));
 sg13g2_a21o_1 _1118_ (.A2(_0322_),
    .A1(_0298_),
    .B1(_0297_),
    .X(_0324_));
 sg13g2_o21ai_1 _1119_ (.B1(_0292_),
    .Y(_0325_),
    .A1(_0293_),
    .A2(_0324_));
 sg13g2_nor2_1 _1120_ (.A(_0257_),
    .B(_0284_),
    .Y(_0326_));
 sg13g2_nor2_1 _1121_ (.A(_0124_),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_nor2_1 _1122_ (.A(net9),
    .B(_0327_),
    .Y(_0328_));
 sg13g2_nand2_1 _1123_ (.Y(_0329_),
    .A(_0290_),
    .B(_0328_));
 sg13g2_nor2_1 _1124_ (.A(_0290_),
    .B(_0328_),
    .Y(_0330_));
 sg13g2_a221oi_1 _1125_ (.B2(_0325_),
    .C1(_0330_),
    .B1(_0329_),
    .A1(net9),
    .Y(_0331_),
    .A2(_0327_));
 sg13g2_xnor2_1 _1126_ (.Y(_0332_),
    .A(net2),
    .B(_0313_));
 sg13g2_a21oi_1 _1127_ (.A1(_0331_),
    .A2(_0332_),
    .Y(_0030_),
    .B1(net104));
 sg13g2_xor2_1 _1128_ (.B(_0315_),
    .A(_0314_),
    .X(_0333_));
 sg13g2_a21oi_1 _1129_ (.A1(_0331_),
    .A2(_0333_),
    .Y(_0031_),
    .B1(net104));
 sg13g2_xnor2_1 _1130_ (.Y(_0334_),
    .A(_0316_),
    .B(_0317_));
 sg13g2_a21oi_1 _1131_ (.A1(_0331_),
    .A2(_0334_),
    .Y(_0032_),
    .B1(net103));
 sg13g2_xnor2_1 _1132_ (.Y(_0335_),
    .A(_0318_),
    .B(_0319_));
 sg13g2_a21oi_1 _1133_ (.A1(_0331_),
    .A2(_0335_),
    .Y(_0033_),
    .B1(net103));
 sg13g2_xnor2_1 _1134_ (.Y(_0336_),
    .A(_0320_),
    .B(_0321_));
 sg13g2_a21oi_1 _1135_ (.A1(_0331_),
    .A2(_0336_),
    .Y(_0034_),
    .B1(net103));
 sg13g2_xor2_1 _1136_ (.B(_0323_),
    .A(_0322_),
    .X(_0337_));
 sg13g2_a21oi_1 _1137_ (.A1(_0331_),
    .A2(_0337_),
    .Y(_0035_),
    .B1(net103));
 sg13g2_xnor2_1 _1138_ (.Y(_0338_),
    .A(_0293_),
    .B(_0324_));
 sg13g2_a21oi_1 _1139_ (.A1(_0331_),
    .A2(_0338_),
    .Y(_0036_),
    .B1(net103));
 sg13g2_nor2_1 _1140_ (.A(_0325_),
    .B(_0329_),
    .Y(_0339_));
 sg13g2_nor2_1 _1141_ (.A(net104),
    .B(_0339_),
    .Y(_0037_));
 sg13g2_nand2_2 _1142_ (.Y(_0340_),
    .A(net107),
    .B(_0166_));
 sg13g2_and3_1 _1143_ (.X(_0038_),
    .A(net107),
    .B(net121),
    .C(_0166_));
 sg13g2_xnor2_1 _1144_ (.Y(_0341_),
    .A(\lif3.spike_counter[1] ),
    .B(net161));
 sg13g2_nor2_1 _1145_ (.A(_0340_),
    .B(net162),
    .Y(_0039_));
 sg13g2_and3_1 _1146_ (.X(_0342_),
    .A(net126),
    .B(\lif3.spike_counter[1] ),
    .C(net161));
 sg13g2_nand3_1 _1147_ (.B(\lif3.spike_counter[1] ),
    .C(net209),
    .A(net126),
    .Y(_0343_));
 sg13g2_a21oi_1 _1148_ (.A1(\lif3.spike_counter[1] ),
    .A2(\lif3.spike_counter[0] ),
    .Y(_0344_),
    .B1(net126));
 sg13g2_nor3_1 _1149_ (.A(_0340_),
    .B(_0342_),
    .C(net127),
    .Y(_0040_));
 sg13g2_xnor2_1 _1150_ (.Y(_0345_),
    .A(net187),
    .B(_0342_));
 sg13g2_nor2_1 _1151_ (.A(_0340_),
    .B(net188),
    .Y(_0041_));
 sg13g2_a21oi_1 _1152_ (.A1(\lif3.spike_counter[3] ),
    .A2(_0342_),
    .Y(_0346_),
    .B1(net147));
 sg13g2_nor2_1 _1153_ (.A(_0187_),
    .B(_0343_),
    .Y(_0347_));
 sg13g2_nor3_1 _1154_ (.A(_0340_),
    .B(net148),
    .C(_0347_),
    .Y(_0042_));
 sg13g2_nor2_1 _1155_ (.A(_0199_),
    .B(_0343_),
    .Y(_0348_));
 sg13g2_nor2_1 _1156_ (.A(net153),
    .B(_0347_),
    .Y(_0349_));
 sg13g2_nor3_1 _1157_ (.A(_0340_),
    .B(_0348_),
    .C(net154),
    .Y(_0043_));
 sg13g2_xnor2_1 _1158_ (.Y(_0350_),
    .A(net155),
    .B(_0348_));
 sg13g2_nor2_1 _1159_ (.A(_0340_),
    .B(net156),
    .Y(_0044_));
 sg13g2_nor3_1 _1160_ (.A(_0014_),
    .B(_0199_),
    .C(_0343_),
    .Y(_0351_));
 sg13g2_xnor2_1 _1161_ (.Y(_0352_),
    .A(net129),
    .B(_0351_));
 sg13g2_nor2_1 _1162_ (.A(_0340_),
    .B(net130),
    .Y(_0045_));
 sg13g2_nor2_1 _1163_ (.A(\lif1.spike_counter[4] ),
    .B(\lif1.spike_counter[3] ),
    .Y(_0353_));
 sg13g2_a21oi_1 _1164_ (.A1(\lif1.spike_counter[2] ),
    .A2(\lif1.spike_counter[1] ),
    .Y(_0354_),
    .B1(\lif1.spike_counter[6] ));
 sg13g2_nand4_1 _1165_ (.B(_0010_),
    .C(_0353_),
    .A(_0132_),
    .Y(_0355_),
    .D(_0354_));
 sg13g2_nand2_1 _1166_ (.Y(_0356_),
    .A(\lif1.adapt_threshold[1] ),
    .B(\lif1.adapt_threshold[0] ));
 sg13g2_nor2_1 _1167_ (.A(\lif1.adapt_threshold[3] ),
    .B(\lif1.adapt_threshold[2] ),
    .Y(_0357_));
 sg13g2_nand2_1 _1168_ (.Y(_0358_),
    .A(\lif1.adapt_threshold[5] ),
    .B(\lif1.adapt_threshold[4] ));
 sg13g2_a21oi_1 _1169_ (.A1(_0356_),
    .A2(_0357_),
    .Y(_0359_),
    .B1(_0358_));
 sg13g2_or2_1 _1170_ (.X(_0360_),
    .B(\lif1.adapt_threshold[6] ),
    .A(\lif1.adapt_threshold[7] ));
 sg13g2_o21ai_1 _1171_ (.B1(_0355_),
    .Y(_0361_),
    .A1(_0359_),
    .A2(_0360_));
 sg13g2_inv_1 _1172_ (.Y(_0362_),
    .A(_0361_));
 sg13g2_or2_1 _1173_ (.X(_0363_),
    .B(\lif1.adapt_threshold[1] ),
    .A(\lif1.adapt_threshold[2] ));
 sg13g2_nand3_1 _1174_ (.B(\lif1.adapt_threshold[3] ),
    .C(_0363_),
    .A(_0101_),
    .Y(_0364_));
 sg13g2_a21oi_1 _1175_ (.A1(_0011_),
    .A2(_0364_),
    .Y(_0365_),
    .B1(_0100_));
 sg13g2_o21ai_1 _1176_ (.B1(\lif1.adapt_threshold[7] ),
    .Y(_0366_),
    .A1(\lif1.adapt_threshold[6] ),
    .A2(_0365_));
 sg13g2_a21oi_1 _1177_ (.A1(\lif1.spike ),
    .A2(_0366_),
    .Y(_0367_),
    .B1(_0362_));
 sg13g2_mux2_1 _1178_ (.A0(\lif1.spike_counter[3] ),
    .A1(_0009_),
    .S(net89),
    .X(_0368_));
 sg13g2_nand2b_1 _1179_ (.Y(_0369_),
    .B(_0008_),
    .A_N(_0368_));
 sg13g2_xor2_1 _1180_ (.B(_0368_),
    .A(_0008_),
    .X(_0370_));
 sg13g2_mux2_1 _1181_ (.A0(_0370_),
    .A1(net205),
    .S(net87),
    .X(_0371_));
 sg13g2_and2_1 _1182_ (.A(net106),
    .B(net206),
    .X(_0046_));
 sg13g2_nand2_1 _1183_ (.Y(_0372_),
    .A(\lif1.spike_counter[4] ),
    .B(\lif1.spike_counter[3] ));
 sg13g2_nand2b_1 _1184_ (.Y(_0373_),
    .B(_0372_),
    .A_N(_0353_));
 sg13g2_nor2_2 _1185_ (.A(net97),
    .B(uo_out[2]),
    .Y(_0374_));
 sg13g2_xnor2_1 _1186_ (.Y(_0375_),
    .A(net97),
    .B(uo_out[2]));
 sg13g2_mux2_1 _1187_ (.A0(_0373_),
    .A1(_0375_),
    .S(net89),
    .X(_0376_));
 sg13g2_nand2_1 _1188_ (.Y(_0377_),
    .A(\lif1.adapt_threshold[1] ),
    .B(_0376_));
 sg13g2_xnor2_1 _1189_ (.Y(_0378_),
    .A(\lif1.adapt_threshold[1] ),
    .B(_0376_));
 sg13g2_nand2b_1 _1190_ (.Y(_0379_),
    .B(_0369_),
    .A_N(_0378_));
 sg13g2_xor2_1 _1191_ (.B(_0378_),
    .A(_0369_),
    .X(_0380_));
 sg13g2_a21oi_1 _1192_ (.A1(net199),
    .A2(net87),
    .Y(_0381_),
    .B1(net101));
 sg13g2_o21ai_1 _1193_ (.B1(_0381_),
    .Y(_0047_),
    .A1(net87),
    .A2(_0380_));
 sg13g2_nand3_1 _1194_ (.B(\lif1.spike_counter[4] ),
    .C(\lif1.spike_counter[3] ),
    .A(\lif1.spike_counter[5] ),
    .Y(_0382_));
 sg13g2_xnor2_1 _1195_ (.Y(_0383_),
    .A(_0132_),
    .B(_0372_));
 sg13g2_nor2_1 _1196_ (.A(net89),
    .B(_0383_),
    .Y(_0384_));
 sg13g2_nor3_1 _1197_ (.A(net97),
    .B(uo_out[2]),
    .C(uo_out[4]),
    .Y(_0385_));
 sg13g2_xnor2_1 _1198_ (.Y(_0386_),
    .A(uo_out[4]),
    .B(_0374_));
 sg13g2_a21oi_1 _1199_ (.A1(_0361_),
    .A2(_0386_),
    .Y(_0387_),
    .B1(_0384_));
 sg13g2_xor2_1 _1200_ (.B(_0387_),
    .A(_0017_),
    .X(_0388_));
 sg13g2_nand3_1 _1201_ (.B(_0379_),
    .C(_0388_),
    .A(_0377_),
    .Y(_0389_));
 sg13g2_a21o_1 _1202_ (.A2(_0379_),
    .A1(_0377_),
    .B1(_0388_),
    .X(_0390_));
 sg13g2_a21oi_1 _1203_ (.A1(_0389_),
    .A2(_0390_),
    .Y(_0391_),
    .B1(net87));
 sg13g2_a21oi_1 _1204_ (.A1(_0103_),
    .A2(net87),
    .Y(_0392_),
    .B1(_0391_));
 sg13g2_and2_1 _1205_ (.A(net106),
    .B(_0392_),
    .X(_0048_));
 sg13g2_nand2_1 _1206_ (.Y(_0393_),
    .A(\lif1.adapt_threshold[2] ),
    .B(_0387_));
 sg13g2_nand4_1 _1207_ (.B(\lif1.spike_counter[5] ),
    .C(\lif1.spike_counter[4] ),
    .A(\lif1.spike_counter[6] ),
    .Y(_0394_),
    .D(\lif1.spike_counter[3] ));
 sg13g2_xor2_1 _1208_ (.B(_0382_),
    .A(\lif1.spike_counter[6] ),
    .X(_0395_));
 sg13g2_nor2b_1 _1209_ (.A(uo_out[5]),
    .B_N(_0385_),
    .Y(_0396_));
 sg13g2_xnor2_1 _1210_ (.Y(_0397_),
    .A(uo_out[5]),
    .B(_0385_));
 sg13g2_nand2_1 _1211_ (.Y(_0398_),
    .A(net89),
    .B(_0397_));
 sg13g2_o21ai_1 _1212_ (.B1(_0398_),
    .Y(_0399_),
    .A1(net89),
    .A2(_0395_));
 sg13g2_or2_1 _1213_ (.X(_0400_),
    .B(_0399_),
    .A(_0018_));
 sg13g2_xnor2_1 _1214_ (.Y(_0401_),
    .A(_0018_),
    .B(_0399_));
 sg13g2_a21o_1 _1215_ (.A2(_0393_),
    .A1(_0390_),
    .B1(_0401_),
    .X(_0402_));
 sg13g2_nand3_1 _1216_ (.B(_0393_),
    .C(_0401_),
    .A(_0390_),
    .Y(_0403_));
 sg13g2_nand2_1 _1217_ (.Y(_0404_),
    .A(_0402_),
    .B(_0403_));
 sg13g2_a21oi_1 _1218_ (.A1(net184),
    .A2(net86),
    .Y(_0405_),
    .B1(net101));
 sg13g2_o21ai_1 _1219_ (.B1(_0405_),
    .Y(_0049_),
    .A1(net86),
    .A2(_0404_));
 sg13g2_or2_1 _1220_ (.X(_0406_),
    .B(net94),
    .A(uo_out[6]));
 sg13g2_nand2_1 _1221_ (.Y(_0407_),
    .A(_0114_),
    .B(_0396_));
 sg13g2_xnor2_1 _1222_ (.Y(_0408_),
    .A(_0114_),
    .B(_0396_));
 sg13g2_a21oi_1 _1223_ (.A1(_0010_),
    .A2(_0394_),
    .Y(_0409_),
    .B1(net89));
 sg13g2_o21ai_1 _1224_ (.B1(_0409_),
    .Y(_0410_),
    .A1(_0010_),
    .A2(_0394_));
 sg13g2_o21ai_1 _1225_ (.B1(_0410_),
    .Y(_0411_),
    .A1(_0362_),
    .A2(_0408_));
 sg13g2_xnor2_1 _1226_ (.Y(_0412_),
    .A(_0011_),
    .B(_0411_));
 sg13g2_a21oi_1 _1227_ (.A1(_0400_),
    .A2(_0402_),
    .Y(_0413_),
    .B1(_0412_));
 sg13g2_nand3_1 _1228_ (.B(_0402_),
    .C(_0412_),
    .A(_0400_),
    .Y(_0414_));
 sg13g2_nand2b_1 _1229_ (.Y(_0415_),
    .B(_0414_),
    .A_N(_0413_));
 sg13g2_a21oi_1 _1230_ (.A1(net163),
    .A2(net86),
    .Y(_0416_),
    .B1(net101));
 sg13g2_o21ai_1 _1231_ (.B1(_0416_),
    .Y(_0050_),
    .A1(net86),
    .A2(_0415_));
 sg13g2_nor2_1 _1232_ (.A(_0101_),
    .B(_0411_),
    .Y(_0417_));
 sg13g2_nor2_1 _1233_ (.A(_0413_),
    .B(_0417_),
    .Y(_0418_));
 sg13g2_or3_1 _1234_ (.A(_0010_),
    .B(net89),
    .C(_0394_),
    .X(_0419_));
 sg13g2_nor2_1 _1235_ (.A(uo_out[7]),
    .B(uo_out[6]),
    .Y(_0420_));
 sg13g2_o21ai_1 _1236_ (.B1(net89),
    .Y(_0421_),
    .A1(uo_out[7]),
    .A2(_0407_));
 sg13g2_a21o_1 _1237_ (.A2(_0407_),
    .A1(uo_out[7]),
    .B1(_0421_),
    .X(_0422_));
 sg13g2_a21oi_1 _1238_ (.A1(_0419_),
    .A2(_0422_),
    .Y(_0423_),
    .B1(\lif1.adapt_threshold[5] ));
 sg13g2_inv_1 _1239_ (.Y(_0424_),
    .A(_0423_));
 sg13g2_nand3_1 _1240_ (.B(_0419_),
    .C(_0422_),
    .A(net170),
    .Y(_0425_));
 sg13g2_nand2_1 _1241_ (.Y(_0426_),
    .A(_0424_),
    .B(_0425_));
 sg13g2_xnor2_1 _1242_ (.Y(_0427_),
    .A(_0418_),
    .B(_0426_));
 sg13g2_a21oi_1 _1243_ (.A1(net170),
    .A2(net86),
    .Y(_0428_),
    .B1(net101));
 sg13g2_o21ai_1 _1244_ (.B1(_0428_),
    .Y(_0051_),
    .A1(net86),
    .A2(_0427_));
 sg13g2_xnor2_1 _1245_ (.Y(_0429_),
    .A(\lif1.adapt_threshold[6] ),
    .B(_0421_));
 sg13g2_o21ai_1 _1246_ (.B1(_0424_),
    .Y(_0430_),
    .A1(_0413_),
    .A2(_0417_));
 sg13g2_a21oi_1 _1247_ (.A1(_0425_),
    .A2(_0430_),
    .Y(_0431_),
    .B1(_0429_));
 sg13g2_nand3_1 _1248_ (.B(_0429_),
    .C(_0430_),
    .A(_0425_),
    .Y(_0432_));
 sg13g2_nand2b_1 _1249_ (.Y(_0433_),
    .B(_0432_),
    .A_N(_0431_));
 sg13g2_a21oi_1 _1250_ (.A1(net204),
    .A2(net87),
    .Y(_0434_),
    .B1(net101));
 sg13g2_o21ai_1 _1251_ (.B1(_0434_),
    .Y(_0052_),
    .A1(net86),
    .A2(_0433_));
 sg13g2_a21oi_1 _1252_ (.A1(\lif1.adapt_threshold[6] ),
    .A2(_0421_),
    .Y(_0435_),
    .B1(_0431_));
 sg13g2_xnor2_1 _1253_ (.Y(_0436_),
    .A(\lif1.adapt_threshold[7] ),
    .B(_0421_));
 sg13g2_xnor2_1 _1254_ (.Y(_0437_),
    .A(_0435_),
    .B(_0436_));
 sg13g2_a21oi_1 _1255_ (.A1(net195),
    .A2(net87),
    .Y(_0438_),
    .B1(net101));
 sg13g2_o21ai_1 _1256_ (.B1(_0438_),
    .Y(_0053_),
    .A1(net86),
    .A2(_0437_));
 sg13g2_and2_1 _1257_ (.A(uo_out[6]),
    .B(net94),
    .X(_0439_));
 sg13g2_xor2_1 _1258_ (.B(net94),
    .A(uo_out[6]),
    .X(_0440_));
 sg13g2_a21oi_1 _1259_ (.A1(uo_out[4]),
    .A2(_0406_),
    .Y(_0441_),
    .B1(_0439_));
 sg13g2_xor2_1 _1260_ (.B(uo_out[6]),
    .A(uo_out[7]),
    .X(_0442_));
 sg13g2_xnor2_1 _1261_ (.Y(_0443_),
    .A(net94),
    .B(_0442_));
 sg13g2_nor2_1 _1262_ (.A(_0441_),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_nand2_1 _1263_ (.Y(_0445_),
    .A(_0441_),
    .B(_0443_));
 sg13g2_xnor2_1 _1264_ (.Y(_0446_),
    .A(net95),
    .B(_0440_));
 sg13g2_and2_1 _1265_ (.A(uo_out[5]),
    .B(net95),
    .X(_0447_));
 sg13g2_xor2_1 _1266_ (.B(net95),
    .A(uo_out[5]),
    .X(_0448_));
 sg13g2_a21oi_1 _1267_ (.A1(uo_out[3]),
    .A2(_0448_),
    .Y(_0449_),
    .B1(_0447_));
 sg13g2_nor2_1 _1268_ (.A(_0446_),
    .B(_0449_),
    .Y(_0450_));
 sg13g2_inv_1 _1269_ (.Y(_0451_),
    .A(_0450_));
 sg13g2_and2_1 _1270_ (.A(uo_out[3]),
    .B(uo_out[4]),
    .X(_0452_));
 sg13g2_xor2_1 _1271_ (.B(uo_out[4]),
    .A(net97),
    .X(_0453_));
 sg13g2_a21o_1 _1272_ (.A2(_0453_),
    .A1(net98),
    .B1(_0452_),
    .X(_0454_));
 sg13g2_xnor2_1 _1273_ (.Y(_0455_),
    .A(uo_out[3]),
    .B(_0448_));
 sg13g2_inv_1 _1274_ (.Y(_0456_),
    .A(_0455_));
 sg13g2_nor2_2 _1275_ (.A(_0454_),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_xnor2_1 _1276_ (.Y(_0458_),
    .A(net98),
    .B(_0453_));
 sg13g2_a21oi_1 _1277_ (.A1(uo_out[3]),
    .A2(net98),
    .Y(_0459_),
    .B1(uo_out[1]));
 sg13g2_nor3_1 _1278_ (.A(_0374_),
    .B(_0458_),
    .C(_0459_),
    .Y(_0460_));
 sg13g2_nand3_1 _1279_ (.B(uo_out[3]),
    .C(uo_out[2]),
    .A(uo_out[1]),
    .Y(_0461_));
 sg13g2_nor2_1 _1280_ (.A(uo_out[1]),
    .B(uo_out[2]),
    .Y(_0462_));
 sg13g2_nand2b_1 _1281_ (.Y(_0463_),
    .B(uo_out[0]),
    .A_N(uo_out[3]));
 sg13g2_o21ai_1 _1282_ (.B1(_0461_),
    .Y(_0464_),
    .A1(_0462_),
    .A2(_0463_));
 sg13g2_o21ai_1 _1283_ (.B1(_0458_),
    .Y(_0465_),
    .A1(_0374_),
    .A2(_0459_));
 sg13g2_nor2b_1 _1284_ (.A(_0460_),
    .B_N(_0465_),
    .Y(_0466_));
 sg13g2_a21oi_1 _1285_ (.A1(_0464_),
    .A2(_0465_),
    .Y(_0467_),
    .B1(_0460_));
 sg13g2_a221oi_1 _1286_ (.B2(_0465_),
    .C1(_0460_),
    .B1(_0464_),
    .A1(_0454_),
    .Y(_0468_),
    .A2(_0456_));
 sg13g2_xnor2_1 _1287_ (.Y(_0469_),
    .A(_0446_),
    .B(_0449_));
 sg13g2_or3_1 _1288_ (.A(_0457_),
    .B(_0468_),
    .C(_0469_),
    .X(_0470_));
 sg13g2_nand2b_2 _1289_ (.Y(_0471_),
    .B(_0445_),
    .A_N(_0444_));
 sg13g2_nor4_2 _1290_ (.A(_0457_),
    .B(_0468_),
    .C(_0469_),
    .Y(_0472_),
    .D(_0471_));
 sg13g2_or4_1 _1291_ (.A(_0457_),
    .B(_0468_),
    .C(_0469_),
    .D(_0471_),
    .X(_0473_));
 sg13g2_a21oi_1 _1292_ (.A1(_0445_),
    .A2(_0450_),
    .Y(_0474_),
    .B1(_0444_));
 sg13g2_a21o_1 _1293_ (.A2(_0450_),
    .A1(_0445_),
    .B1(_0444_),
    .X(_0475_));
 sg13g2_nor3_1 _1294_ (.A(_0406_),
    .B(_0472_),
    .C(_0475_),
    .Y(_0476_));
 sg13g2_nor2_1 _1295_ (.A(_0113_),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_nor2_1 _1296_ (.A(uo_out[7]),
    .B(_0439_),
    .Y(_0478_));
 sg13g2_o21ai_1 _1297_ (.B1(uo_out[6]),
    .Y(_0479_),
    .A1(_0472_),
    .A2(_0475_));
 sg13g2_o21ai_1 _1298_ (.B1(_0479_),
    .Y(_0480_),
    .A1(_0477_),
    .A2(_0478_));
 sg13g2_and2_1 _1299_ (.A(net8),
    .B(_0480_),
    .X(_0481_));
 sg13g2_nor3_1 _1300_ (.A(net9),
    .B(_0477_),
    .C(_0481_),
    .Y(_0482_));
 sg13g2_a21oi_1 _1301_ (.A1(uo_out[5]),
    .A2(_0442_),
    .Y(_0483_),
    .B1(_0420_));
 sg13g2_nand3_1 _1302_ (.B(_0474_),
    .C(_0483_),
    .A(_0473_),
    .Y(_0484_));
 sg13g2_a21o_1 _1303_ (.A2(_0474_),
    .A1(_0473_),
    .B1(_0483_),
    .X(_0485_));
 sg13g2_a21oi_2 _1304_ (.B1(_0135_),
    .Y(_0486_),
    .A2(_0485_),
    .A1(_0484_));
 sg13g2_xnor2_1 _1305_ (.Y(_0487_),
    .A(_0134_),
    .B(_0480_));
 sg13g2_and2_1 _1306_ (.A(_0486_),
    .B(_0487_),
    .X(_0488_));
 sg13g2_xor2_1 _1307_ (.B(_0487_),
    .A(_0486_),
    .X(_0489_));
 sg13g2_a21o_1 _1308_ (.A2(_0470_),
    .A1(_0451_),
    .B1(_0471_),
    .X(_0490_));
 sg13g2_nand3_1 _1309_ (.B(_0470_),
    .C(_0471_),
    .A(_0451_),
    .Y(_0491_));
 sg13g2_and3_1 _1310_ (.X(_0492_),
    .A(net6),
    .B(_0490_),
    .C(_0491_));
 sg13g2_nand3_1 _1311_ (.B(_0490_),
    .C(_0491_),
    .A(net6),
    .Y(_0493_));
 sg13g2_and3_1 _1312_ (.X(_0494_),
    .A(_0135_),
    .B(_0484_),
    .C(_0485_));
 sg13g2_nor3_1 _1313_ (.A(_0486_),
    .B(_0493_),
    .C(_0494_),
    .Y(_0495_));
 sg13g2_or3_1 _1314_ (.A(_0486_),
    .B(_0493_),
    .C(_0494_),
    .X(_0496_));
 sg13g2_o21ai_1 _1315_ (.B1(_0493_),
    .Y(_0497_),
    .A1(_0486_),
    .A2(_0494_));
 sg13g2_o21ai_1 _1316_ (.B1(_0469_),
    .Y(_0498_),
    .A1(_0457_),
    .A2(_0468_));
 sg13g2_and2_1 _1317_ (.A(_0470_),
    .B(_0498_),
    .X(_0499_));
 sg13g2_nor2_1 _1318_ (.A(net5),
    .B(_0499_),
    .Y(_0500_));
 sg13g2_a21oi_1 _1319_ (.A1(_0490_),
    .A2(_0491_),
    .Y(_0501_),
    .B1(net6));
 sg13g2_nor3_1 _1320_ (.A(_0492_),
    .B(_0500_),
    .C(_0501_),
    .Y(_0502_));
 sg13g2_or3_1 _1321_ (.A(_0492_),
    .B(_0500_),
    .C(_0501_),
    .X(_0503_));
 sg13g2_xnor2_1 _1322_ (.Y(_0504_),
    .A(_0454_),
    .B(_0455_));
 sg13g2_xnor2_1 _1323_ (.Y(_0505_),
    .A(_0467_),
    .B(_0504_));
 sg13g2_nand2_1 _1324_ (.Y(_0506_),
    .A(net4),
    .B(_0505_));
 sg13g2_xnor2_1 _1325_ (.Y(_0507_),
    .A(net5),
    .B(_0499_));
 sg13g2_nor2b_1 _1326_ (.A(_0506_),
    .B_N(_0507_),
    .Y(_0508_));
 sg13g2_xnor2_1 _1327_ (.Y(_0509_),
    .A(_0464_),
    .B(_0466_));
 sg13g2_nor2b_1 _1328_ (.A(net3),
    .B_N(_0509_),
    .Y(_0510_));
 sg13g2_xor2_1 _1329_ (.B(_0505_),
    .A(net4),
    .X(_0511_));
 sg13g2_nand2b_1 _1330_ (.Y(_0512_),
    .B(_0511_),
    .A_N(_0510_));
 sg13g2_nor2_1 _1331_ (.A(uo_out[0]),
    .B(_0462_),
    .Y(_0513_));
 sg13g2_xnor2_1 _1332_ (.Y(_0514_),
    .A(uo_out[3]),
    .B(_0513_));
 sg13g2_nor2b_1 _1333_ (.A(net2),
    .B_N(_0514_),
    .Y(_0515_));
 sg13g2_xor2_1 _1334_ (.B(_0509_),
    .A(net3),
    .X(_0516_));
 sg13g2_nand2b_1 _1335_ (.Y(_0517_),
    .B(_0516_),
    .A_N(_0515_));
 sg13g2_nor2b_1 _1336_ (.A(_0511_),
    .B_N(_0510_),
    .Y(_0518_));
 sg13g2_xnor2_1 _1337_ (.Y(_0519_),
    .A(_0510_),
    .B(_0511_));
 sg13g2_o21ai_1 _1338_ (.B1(_0512_),
    .Y(_0520_),
    .A1(_0517_),
    .A2(_0518_));
 sg13g2_nand2b_1 _1339_ (.Y(_0521_),
    .B(_0506_),
    .A_N(_0507_));
 sg13g2_nand2b_1 _1340_ (.Y(_0522_),
    .B(_0521_),
    .A_N(_0508_));
 sg13g2_a21oi_2 _1341_ (.B1(_0508_),
    .Y(_0523_),
    .A2(_0521_),
    .A1(_0520_));
 sg13g2_o21ai_1 _1342_ (.B1(_0500_),
    .Y(_0524_),
    .A1(_0492_),
    .A2(_0501_));
 sg13g2_and2_1 _1343_ (.A(_0503_),
    .B(_0524_),
    .X(_0525_));
 sg13g2_nor2b_1 _1344_ (.A(_0523_),
    .B_N(_0525_),
    .Y(_0526_));
 sg13g2_nor2_1 _1345_ (.A(_0502_),
    .B(_0526_),
    .Y(_0527_));
 sg13g2_o21ai_1 _1346_ (.B1(_0497_),
    .Y(_0528_),
    .A1(_0495_),
    .A2(_0502_));
 sg13g2_nand2_1 _1347_ (.Y(_0529_),
    .A(_0496_),
    .B(_0497_));
 sg13g2_nand4_1 _1348_ (.B(_0497_),
    .C(_0503_),
    .A(_0496_),
    .Y(_0530_),
    .D(_0524_));
 sg13g2_o21ai_1 _1349_ (.B1(_0528_),
    .Y(_0531_),
    .A1(_0523_),
    .A2(_0530_));
 sg13g2_a21oi_1 _1350_ (.A1(_0489_),
    .A2(_0531_),
    .Y(_0532_),
    .B1(_0488_));
 sg13g2_nand2_1 _1351_ (.Y(_0533_),
    .A(net9),
    .B(_0477_));
 sg13g2_o21ai_1 _1352_ (.B1(_0481_),
    .Y(_0534_),
    .A1(net9),
    .A2(_0477_));
 sg13g2_and2_1 _1353_ (.A(_0533_),
    .B(_0534_),
    .X(_0535_));
 sg13g2_a21oi_2 _1354_ (.B1(_0482_),
    .Y(_0536_),
    .A2(_0535_),
    .A1(_0532_));
 sg13g2_xor2_1 _1355_ (.B(_0514_),
    .A(net2),
    .X(_0537_));
 sg13g2_o21ai_1 _1356_ (.B1(net1),
    .Y(_0538_),
    .A1(_0536_),
    .A2(_0537_));
 sg13g2_inv_1 _1357_ (.Y(_0054_),
    .A(_0538_));
 sg13g2_xnor2_1 _1358_ (.Y(_0539_),
    .A(_0515_),
    .B(_0516_));
 sg13g2_o21ai_1 _1359_ (.B1(net1),
    .Y(_0540_),
    .A1(_0536_),
    .A2(_0539_));
 sg13g2_inv_1 _1360_ (.Y(_0055_),
    .A(_0540_));
 sg13g2_xnor2_1 _1361_ (.Y(_0541_),
    .A(_0517_),
    .B(_0519_));
 sg13g2_o21ai_1 _1362_ (.B1(net106),
    .Y(_0542_),
    .A1(_0536_),
    .A2(_0541_));
 sg13g2_inv_1 _1363_ (.Y(_0056_),
    .A(_0542_));
 sg13g2_xnor2_1 _1364_ (.Y(_0543_),
    .A(_0520_),
    .B(_0522_));
 sg13g2_o21ai_1 _1365_ (.B1(net107),
    .Y(_0544_),
    .A1(_0536_),
    .A2(_0543_));
 sg13g2_inv_1 _1366_ (.Y(_0057_),
    .A(_0544_));
 sg13g2_xnor2_1 _1367_ (.Y(_0545_),
    .A(_0523_),
    .B(_0525_));
 sg13g2_o21ai_1 _1368_ (.B1(net107),
    .Y(_0546_),
    .A1(_0536_),
    .A2(_0545_));
 sg13g2_inv_1 _1369_ (.Y(_0058_),
    .A(_0546_));
 sg13g2_xor2_1 _1370_ (.B(_0529_),
    .A(_0527_),
    .X(_0547_));
 sg13g2_o21ai_1 _1371_ (.B1(net107),
    .Y(_0548_),
    .A1(_0536_),
    .A2(_0547_));
 sg13g2_inv_1 _1372_ (.Y(_0059_),
    .A(_0548_));
 sg13g2_xor2_1 _1373_ (.B(_0531_),
    .A(_0489_),
    .X(_0549_));
 sg13g2_o21ai_1 _1374_ (.B1(net106),
    .Y(_0550_),
    .A1(_0536_),
    .A2(_0549_));
 sg13g2_inv_1 _1375_ (.Y(_0060_),
    .A(_0550_));
 sg13g2_a21oi_1 _1376_ (.A1(_0482_),
    .A2(_0532_),
    .Y(_0061_),
    .B1(net101));
 sg13g2_nand2_2 _1377_ (.Y(_0551_),
    .A(net106),
    .B(_0149_));
 sg13g2_and3_1 _1378_ (.X(_0062_),
    .A(net106),
    .B(net122),
    .C(_0149_));
 sg13g2_xnor2_1 _1379_ (.Y(_0552_),
    .A(\lif1.spike_counter[1] ),
    .B(net165));
 sg13g2_nor2_1 _1380_ (.A(_0551_),
    .B(net166),
    .Y(_0063_));
 sg13g2_and3_1 _1381_ (.X(_0553_),
    .A(net137),
    .B(\lif1.spike_counter[1] ),
    .C(net165));
 sg13g2_nand3_1 _1382_ (.B(\lif1.spike_counter[1] ),
    .C(net165),
    .A(net137),
    .Y(_0554_));
 sg13g2_a21oi_1 _1383_ (.A1(\lif1.spike_counter[1] ),
    .A2(\lif1.spike_counter[0] ),
    .Y(_0555_),
    .B1(net137));
 sg13g2_nor3_1 _1384_ (.A(_0551_),
    .B(_0553_),
    .C(net138),
    .Y(_0064_));
 sg13g2_xnor2_1 _1385_ (.Y(_0556_),
    .A(net192),
    .B(_0553_));
 sg13g2_nor2_1 _1386_ (.A(_0551_),
    .B(net193),
    .Y(_0065_));
 sg13g2_a21oi_1 _1387_ (.A1(\lif1.spike_counter[3] ),
    .A2(_0553_),
    .Y(_0557_),
    .B1(net159));
 sg13g2_nor2_1 _1388_ (.A(_0372_),
    .B(_0554_),
    .Y(_0558_));
 sg13g2_nor3_1 _1389_ (.A(_0551_),
    .B(net160),
    .C(_0558_),
    .Y(_0066_));
 sg13g2_xnor2_1 _1390_ (.Y(_0559_),
    .A(net171),
    .B(_0558_));
 sg13g2_nor2_1 _1391_ (.A(_0551_),
    .B(net172),
    .Y(_0067_));
 sg13g2_nor2_1 _1392_ (.A(_0394_),
    .B(_0554_),
    .Y(_0560_));
 sg13g2_a21oi_1 _1393_ (.A1(\lif1.spike_counter[5] ),
    .A2(_0558_),
    .Y(_0561_),
    .B1(net145));
 sg13g2_nor3_1 _1394_ (.A(_0551_),
    .B(_0560_),
    .C(net146),
    .Y(_0068_));
 sg13g2_xnor2_1 _1395_ (.Y(_0562_),
    .A(net131),
    .B(_0560_));
 sg13g2_nor2_1 _1396_ (.A(_0551_),
    .B(net132),
    .Y(_0069_));
 sg13g2_nor2_1 _1397_ (.A(\lif2.spike_counter[4] ),
    .B(\lif2.spike_counter[3] ),
    .Y(_0563_));
 sg13g2_a21oi_1 _1398_ (.A1(\lif2.spike_counter[2] ),
    .A2(\lif2.spike_counter[1] ),
    .Y(_0564_),
    .B1(\lif2.spike_counter[5] ));
 sg13g2_nand4_1 _1399_ (.B(_0007_),
    .C(_0563_),
    .A(_0131_),
    .Y(_0565_),
    .D(_0564_));
 sg13g2_nand2_1 _1400_ (.Y(_0566_),
    .A(\lif2.adapt_threshold[1] ),
    .B(\lif2.adapt_threshold[0] ));
 sg13g2_nor2_1 _1401_ (.A(\lif2.adapt_threshold[3] ),
    .B(\lif2.adapt_threshold[2] ),
    .Y(_0567_));
 sg13g2_nand2_1 _1402_ (.Y(_0568_),
    .A(\lif2.adapt_threshold[5] ),
    .B(\lif2.adapt_threshold[4] ));
 sg13g2_a21oi_1 _1403_ (.A1(_0566_),
    .A2(_0567_),
    .Y(_0569_),
    .B1(_0568_));
 sg13g2_nand2_1 _1404_ (.Y(_0570_),
    .A(_0094_),
    .B(_0095_));
 sg13g2_o21ai_1 _1405_ (.B1(_0565_),
    .Y(_0571_),
    .A1(_0569_),
    .A2(_0570_));
 sg13g2_or2_1 _1406_ (.X(_0572_),
    .B(\lif2.adapt_threshold[1] ),
    .A(\lif2.adapt_threshold[2] ));
 sg13g2_nand3_1 _1407_ (.B(\lif2.adapt_threshold[3] ),
    .C(_0572_),
    .A(_0097_),
    .Y(_0573_));
 sg13g2_a21oi_1 _1408_ (.A1(_0012_),
    .A2(_0573_),
    .Y(_0574_),
    .B1(_0096_));
 sg13g2_o21ai_1 _1409_ (.B1(\lif2.adapt_threshold[7] ),
    .Y(_0575_),
    .A1(\lif2.adapt_threshold[6] ),
    .A2(_0574_));
 sg13g2_nand2_1 _1410_ (.Y(_0576_),
    .A(\lif2.spike ),
    .B(_0575_));
 sg13g2_and2_1 _1411_ (.A(net88),
    .B(_0576_),
    .X(_0577_));
 sg13g2_mux2_1 _1412_ (.A0(\lif2.spike_counter[3] ),
    .A1(_0006_),
    .S(_0571_),
    .X(_0578_));
 sg13g2_nand2b_1 _1413_ (.Y(_0579_),
    .B(_0005_),
    .A_N(_0578_));
 sg13g2_xor2_1 _1414_ (.B(_0578_),
    .A(_0005_),
    .X(_0580_));
 sg13g2_nor2_1 _1415_ (.A(net85),
    .B(_0580_),
    .Y(_0581_));
 sg13g2_nor2b_1 _1416_ (.A(net133),
    .B_N(net85),
    .Y(_0582_));
 sg13g2_nor3_1 _1417_ (.A(net105),
    .B(_0581_),
    .C(_0582_),
    .Y(_0070_));
 sg13g2_nand2_1 _1418_ (.Y(_0583_),
    .A(net143),
    .B(\lif2.spike_counter[3] ));
 sg13g2_nand2b_1 _1419_ (.Y(_0584_),
    .B(_0583_),
    .A_N(_0563_));
 sg13g2_nor2_2 _1420_ (.A(\lif2.state[3] ),
    .B(net92),
    .Y(_0585_));
 sg13g2_nand2_1 _1421_ (.Y(_0586_),
    .A(\lif2.state[3] ),
    .B(net92));
 sg13g2_nand2b_1 _1422_ (.Y(_0587_),
    .B(_0586_),
    .A_N(_0585_));
 sg13g2_mux2_1 _1423_ (.A0(_0584_),
    .A1(_0587_),
    .S(_0571_),
    .X(_0588_));
 sg13g2_and2_1 _1424_ (.A(\lif2.adapt_threshold[1] ),
    .B(_0588_),
    .X(_0589_));
 sg13g2_xor2_1 _1425_ (.B(_0588_),
    .A(\lif2.adapt_threshold[1] ),
    .X(_0590_));
 sg13g2_xnor2_1 _1426_ (.Y(_0591_),
    .A(_0579_),
    .B(_0590_));
 sg13g2_a21oi_1 _1427_ (.A1(net197),
    .A2(net85),
    .Y(_0592_),
    .B1(net105));
 sg13g2_o21ai_1 _1428_ (.B1(_0592_),
    .Y(_0071_),
    .A1(net85),
    .A2(_0591_));
 sg13g2_a21oi_1 _1429_ (.A1(_0579_),
    .A2(_0590_),
    .Y(_0593_),
    .B1(_0589_));
 sg13g2_nand3_1 _1430_ (.B(\lif2.spike_counter[4] ),
    .C(\lif2.spike_counter[3] ),
    .A(\lif2.spike_counter[5] ),
    .Y(_0594_));
 sg13g2_xor2_1 _1431_ (.B(_0583_),
    .A(\lif2.spike_counter[5] ),
    .X(_0595_));
 sg13g2_nand2_1 _1432_ (.Y(_0596_),
    .A(_0123_),
    .B(_0585_));
 sg13g2_o21ai_1 _1433_ (.B1(\lif2.state[4] ),
    .Y(_0597_),
    .A1(\lif2.state[3] ),
    .A2(net92));
 sg13g2_nand2_1 _1434_ (.Y(_0598_),
    .A(_0596_),
    .B(_0597_));
 sg13g2_mux2_1 _1435_ (.A0(_0595_),
    .A1(_0598_),
    .S(net88),
    .X(_0599_));
 sg13g2_xor2_1 _1436_ (.B(_0599_),
    .A(_0000_),
    .X(_0600_));
 sg13g2_xnor2_1 _1437_ (.Y(_0601_),
    .A(_0593_),
    .B(_0600_));
 sg13g2_mux2_1 _1438_ (.A0(_0601_),
    .A1(_0098_),
    .S(net85),
    .X(_0602_));
 sg13g2_nor2_1 _1439_ (.A(net102),
    .B(net203),
    .Y(_0072_));
 sg13g2_nand2_1 _1440_ (.Y(_0603_),
    .A(\lif2.adapt_threshold[2] ),
    .B(_0599_));
 sg13g2_o21ai_1 _1441_ (.B1(_0603_),
    .Y(_0604_),
    .A1(_0593_),
    .A2(_0600_));
 sg13g2_or2_1 _1442_ (.X(_0605_),
    .B(_0594_),
    .A(_0131_));
 sg13g2_xnor2_1 _1443_ (.Y(_0606_),
    .A(_0131_),
    .B(_0594_));
 sg13g2_nor2_1 _1444_ (.A(net91),
    .B(_0596_),
    .Y(_0607_));
 sg13g2_xnor2_1 _1445_ (.Y(_0608_),
    .A(_0122_),
    .B(_0596_));
 sg13g2_nand2_1 _1446_ (.Y(_0609_),
    .A(net88),
    .B(_0608_));
 sg13g2_o21ai_1 _1447_ (.B1(_0609_),
    .Y(_0610_),
    .A1(net88),
    .A2(_0606_));
 sg13g2_nor2_1 _1448_ (.A(_0001_),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_xnor2_1 _1449_ (.Y(_0612_),
    .A(_0001_),
    .B(_0610_));
 sg13g2_inv_1 _1450_ (.Y(_0613_),
    .A(_0612_));
 sg13g2_xnor2_1 _1451_ (.Y(_0614_),
    .A(_0604_),
    .B(_0613_));
 sg13g2_a21oi_1 _1452_ (.A1(net182),
    .A2(net85),
    .Y(_0615_),
    .B1(net102));
 sg13g2_o21ai_1 _1453_ (.B1(_0615_),
    .Y(_0073_),
    .A1(net84),
    .A2(_0614_));
 sg13g2_a21oi_1 _1454_ (.A1(_0604_),
    .A2(_0613_),
    .Y(_0616_),
    .B1(_0611_));
 sg13g2_nand2_1 _1455_ (.Y(_0617_),
    .A(_0121_),
    .B(_0607_));
 sg13g2_xnor2_1 _1456_ (.Y(_0618_),
    .A(_0121_),
    .B(_0607_));
 sg13g2_xor2_1 _1457_ (.B(_0605_),
    .A(_0007_),
    .X(_0619_));
 sg13g2_nor2_1 _1458_ (.A(net88),
    .B(_0619_),
    .Y(_0620_));
 sg13g2_a21oi_1 _1459_ (.A1(net88),
    .A2(_0618_),
    .Y(_0621_),
    .B1(_0620_));
 sg13g2_xnor2_1 _1460_ (.Y(_0622_),
    .A(_0012_),
    .B(_0621_));
 sg13g2_xnor2_1 _1461_ (.Y(_0623_),
    .A(_0616_),
    .B(_0622_));
 sg13g2_a21oi_1 _1462_ (.A1(net167),
    .A2(net84),
    .Y(_0624_),
    .B1(net102));
 sg13g2_o21ai_1 _1463_ (.B1(_0624_),
    .Y(_0074_),
    .A1(net85),
    .A2(_0623_));
 sg13g2_nor3_1 _1464_ (.A(_0007_),
    .B(net88),
    .C(_0605_),
    .Y(_0625_));
 sg13g2_o21ai_1 _1465_ (.B1(net88),
    .Y(_0626_),
    .A1(\lif2.state[7] ),
    .A2(_0617_));
 sg13g2_a21oi_1 _1466_ (.A1(\lif2.state[7] ),
    .A2(_0617_),
    .Y(_0627_),
    .B1(_0626_));
 sg13g2_or2_1 _1467_ (.X(_0628_),
    .B(_0627_),
    .A(_0625_));
 sg13g2_nor2_1 _1468_ (.A(_0096_),
    .B(_0628_),
    .Y(_0629_));
 sg13g2_and2_1 _1469_ (.A(_0096_),
    .B(_0628_),
    .X(_0630_));
 sg13g2_inv_1 _1470_ (.Y(_0631_),
    .A(_0630_));
 sg13g2_nor2_1 _1471_ (.A(_0629_),
    .B(_0630_),
    .Y(_0632_));
 sg13g2_or2_1 _1472_ (.X(_0633_),
    .B(_0621_),
    .A(_0097_));
 sg13g2_o21ai_1 _1473_ (.B1(_0633_),
    .Y(_0634_),
    .A1(_0616_),
    .A2(_0622_));
 sg13g2_xnor2_1 _1474_ (.Y(_0635_),
    .A(_0632_),
    .B(_0634_));
 sg13g2_a21oi_1 _1475_ (.A1(net169),
    .A2(net84),
    .Y(_0636_),
    .B1(net102));
 sg13g2_o21ai_1 _1476_ (.B1(_0636_),
    .Y(_0075_),
    .A1(net84),
    .A2(_0635_));
 sg13g2_xnor2_1 _1477_ (.Y(_0637_),
    .A(\lif2.adapt_threshold[6] ),
    .B(_0626_));
 sg13g2_a21oi_1 _1478_ (.A1(_0631_),
    .A2(_0634_),
    .Y(_0638_),
    .B1(_0629_));
 sg13g2_nor2_1 _1479_ (.A(_0637_),
    .B(_0638_),
    .Y(_0639_));
 sg13g2_a21o_1 _1480_ (.A2(_0638_),
    .A1(_0637_),
    .B1(net84),
    .X(_0640_));
 sg13g2_a21oi_1 _1481_ (.A1(net201),
    .A2(net84),
    .Y(_0641_),
    .B1(net102));
 sg13g2_o21ai_1 _1482_ (.B1(_0641_),
    .Y(_0076_),
    .A1(_0639_),
    .A2(_0640_));
 sg13g2_a21oi_1 _1483_ (.A1(\lif2.adapt_threshold[6] ),
    .A2(_0626_),
    .Y(_0642_),
    .B1(_0639_));
 sg13g2_xnor2_1 _1484_ (.Y(_0643_),
    .A(net186),
    .B(_0626_));
 sg13g2_xnor2_1 _1485_ (.Y(_0644_),
    .A(_0642_),
    .B(_0643_));
 sg13g2_a21oi_1 _1486_ (.A1(net186),
    .A2(net84),
    .Y(_0645_),
    .B1(net102));
 sg13g2_o21ai_1 _1487_ (.B1(_0645_),
    .Y(_0077_),
    .A1(net84),
    .A2(_0644_));
 sg13g2_o21ai_1 _1488_ (.B1(net91),
    .Y(_0646_),
    .A1(_0120_),
    .A2(_0121_));
 sg13g2_inv_1 _1489_ (.Y(_0647_),
    .A(_0646_));
 sg13g2_and2_1 _1490_ (.A(net91),
    .B(\lif2.state[4] ),
    .X(_0648_));
 sg13g2_xor2_1 _1491_ (.B(\lif2.state[4] ),
    .A(net91),
    .X(_0649_));
 sg13g2_a21oi_2 _1492_ (.B1(_0648_),
    .Y(_0650_),
    .A2(_0649_),
    .A1(\lif2.state[6] ));
 sg13g2_xor2_1 _1493_ (.B(net91),
    .A(\lif2.state[6] ),
    .X(_0651_));
 sg13g2_xnor2_1 _1494_ (.Y(_0652_),
    .A(\lif2.state[7] ),
    .B(_0651_));
 sg13g2_nand2_1 _1495_ (.Y(_0653_),
    .A(_0650_),
    .B(_0652_));
 sg13g2_or2_1 _1496_ (.X(_0654_),
    .B(_0652_),
    .A(_0650_));
 sg13g2_xnor2_1 _1497_ (.Y(_0655_),
    .A(\lif2.state[6] ),
    .B(_0649_));
 sg13g2_nor2_1 _1498_ (.A(_0118_),
    .B(_0123_),
    .Y(_0656_));
 sg13g2_xor2_1 _1499_ (.B(\lif2.state[4] ),
    .A(\lif2.state[3] ),
    .X(_0657_));
 sg13g2_a21oi_1 _1500_ (.A1(\lif2.state[5] ),
    .A2(_0657_),
    .Y(_0658_),
    .B1(_0656_));
 sg13g2_nor2_1 _1501_ (.A(_0655_),
    .B(_0658_),
    .Y(_0659_));
 sg13g2_xnor2_1 _1502_ (.Y(_0660_),
    .A(net91),
    .B(_0657_));
 sg13g2_inv_1 _1503_ (.Y(_0661_),
    .A(_0660_));
 sg13g2_nand2_1 _1504_ (.Y(_0662_),
    .A(_0586_),
    .B(_0597_));
 sg13g2_nor2_1 _1505_ (.A(_0661_),
    .B(_0662_),
    .Y(_0663_));
 sg13g2_a21oi_1 _1506_ (.A1(\lif2.state[3] ),
    .A2(\lif2.state[2] ),
    .Y(_0664_),
    .B1(\lif2.state[1] ));
 sg13g2_nor2_1 _1507_ (.A(_0585_),
    .B(_0664_),
    .Y(_0665_));
 sg13g2_xnor2_1 _1508_ (.Y(_0666_),
    .A(net92),
    .B(_0657_));
 sg13g2_nor3_1 _1509_ (.A(_0585_),
    .B(_0664_),
    .C(_0666_),
    .Y(_0667_));
 sg13g2_nand3_1 _1510_ (.B(\lif2.state[3] ),
    .C(net92),
    .A(\lif2.state[1] ),
    .Y(_0668_));
 sg13g2_nor2_1 _1511_ (.A(\lif2.state[1] ),
    .B(net92),
    .Y(_0669_));
 sg13g2_nand2_1 _1512_ (.Y(_0670_),
    .A(\lif2.state[0] ),
    .B(_0118_));
 sg13g2_o21ai_1 _1513_ (.B1(_0668_),
    .Y(_0671_),
    .A1(_0669_),
    .A2(_0670_));
 sg13g2_nand2b_1 _1514_ (.Y(_0672_),
    .B(_0666_),
    .A_N(_0665_));
 sg13g2_xnor2_1 _1515_ (.Y(_0673_),
    .A(_0665_),
    .B(_0666_));
 sg13g2_a21oi_1 _1516_ (.A1(_0671_),
    .A2(_0672_),
    .Y(_0674_),
    .B1(_0667_));
 sg13g2_a221oi_1 _1517_ (.B2(_0672_),
    .C1(_0667_),
    .B1(_0671_),
    .A1(_0661_),
    .Y(_0675_),
    .A2(_0662_));
 sg13g2_xnor2_1 _1518_ (.Y(_0676_),
    .A(_0655_),
    .B(_0658_));
 sg13g2_nor3_1 _1519_ (.A(_0663_),
    .B(_0675_),
    .C(_0676_),
    .Y(_0677_));
 sg13g2_nor2_1 _1520_ (.A(_0659_),
    .B(_0677_),
    .Y(_0678_));
 sg13g2_nand2_1 _1521_ (.Y(_0679_),
    .A(_0653_),
    .B(_0659_));
 sg13g2_xor2_1 _1522_ (.B(_0652_),
    .A(_0650_),
    .X(_0680_));
 sg13g2_inv_1 _1523_ (.Y(_0681_),
    .A(_0680_));
 sg13g2_or4_1 _1524_ (.A(_0663_),
    .B(_0675_),
    .C(_0676_),
    .D(_0681_),
    .X(_0682_));
 sg13g2_nand3_1 _1525_ (.B(_0679_),
    .C(_0682_),
    .A(_0654_),
    .Y(_0683_));
 sg13g2_o21ai_1 _1526_ (.B1(\lif2.state[6] ),
    .Y(_0684_),
    .A1(_0647_),
    .A2(_0683_));
 sg13g2_nand4_1 _1527_ (.B(_0121_),
    .C(_0122_),
    .A(\lif2.state[7] ),
    .Y(_0685_),
    .D(_0678_));
 sg13g2_a21oi_2 _1528_ (.B1(_0134_),
    .Y(_0686_),
    .A2(_0685_),
    .A1(_0684_));
 sg13g2_nor2_1 _1529_ (.A(_0651_),
    .B(_0683_),
    .Y(_0687_));
 sg13g2_nor2_1 _1530_ (.A(_0120_),
    .B(_0687_),
    .Y(_0688_));
 sg13g2_nor2_1 _1531_ (.A(net9),
    .B(_0688_),
    .Y(_0689_));
 sg13g2_nor3_1 _1532_ (.A(net9),
    .B(_0686_),
    .C(_0688_),
    .Y(_0690_));
 sg13g2_o21ai_1 _1533_ (.B1(_0646_),
    .Y(_0691_),
    .A1(\lif2.state[7] ),
    .A2(\lif2.state[6] ));
 sg13g2_xor2_1 _1534_ (.B(_0691_),
    .A(_0683_),
    .X(_0692_));
 sg13g2_nand2b_1 _1535_ (.Y(_0693_),
    .B(net7),
    .A_N(_0692_));
 sg13g2_and3_1 _1536_ (.X(_0694_),
    .A(_0134_),
    .B(_0684_),
    .C(_0685_));
 sg13g2_nor3_1 _1537_ (.A(_0686_),
    .B(_0693_),
    .C(_0694_),
    .Y(_0695_));
 sg13g2_o21ai_1 _1538_ (.B1(_0693_),
    .Y(_0696_),
    .A1(_0686_),
    .A2(_0694_));
 sg13g2_nor2b_1 _1539_ (.A(_0695_),
    .B_N(_0696_),
    .Y(_0697_));
 sg13g2_xnor2_1 _1540_ (.Y(_0698_),
    .A(net7),
    .B(_0692_));
 sg13g2_xnor2_1 _1541_ (.Y(_0699_),
    .A(_0678_),
    .B(_0680_));
 sg13g2_or2_1 _1542_ (.X(_0700_),
    .B(_0699_),
    .A(net6));
 sg13g2_or2_1 _1543_ (.X(_0701_),
    .B(_0700_),
    .A(_0698_));
 sg13g2_inv_1 _1544_ (.Y(_0702_),
    .A(_0701_));
 sg13g2_nand2_1 _1545_ (.Y(_0703_),
    .A(_0698_),
    .B(_0700_));
 sg13g2_o21ai_1 _1546_ (.B1(_0676_),
    .Y(_0704_),
    .A1(_0663_),
    .A2(_0675_));
 sg13g2_nor2b_1 _1547_ (.A(_0677_),
    .B_N(_0704_),
    .Y(_0705_));
 sg13g2_nand2_1 _1548_ (.Y(_0706_),
    .A(net5),
    .B(_0705_));
 sg13g2_xnor2_1 _1549_ (.Y(_0707_),
    .A(net6),
    .B(_0699_));
 sg13g2_nor2b_1 _1550_ (.A(_0706_),
    .B_N(_0707_),
    .Y(_0708_));
 sg13g2_xnor2_1 _1551_ (.Y(_0709_),
    .A(_0660_),
    .B(_0662_));
 sg13g2_xnor2_1 _1552_ (.Y(_0710_),
    .A(_0674_),
    .B(_0709_));
 sg13g2_nor2_1 _1553_ (.A(net4),
    .B(_0710_),
    .Y(_0711_));
 sg13g2_xnor2_1 _1554_ (.Y(_0712_),
    .A(net5),
    .B(_0705_));
 sg13g2_nor2_1 _1555_ (.A(_0711_),
    .B(_0712_),
    .Y(_0713_));
 sg13g2_xnor2_1 _1556_ (.Y(_0714_),
    .A(_0671_),
    .B(_0673_));
 sg13g2_inv_1 _1557_ (.Y(_0715_),
    .A(_0714_));
 sg13g2_nand2_1 _1558_ (.Y(_0716_),
    .A(net3),
    .B(_0715_));
 sg13g2_xnor2_1 _1559_ (.Y(_0717_),
    .A(net4),
    .B(_0710_));
 sg13g2_nand2b_1 _1560_ (.Y(_0718_),
    .B(_0717_),
    .A_N(_0716_));
 sg13g2_nor2_1 _1561_ (.A(\lif2.state[0] ),
    .B(_0669_),
    .Y(_0719_));
 sg13g2_xnor2_1 _1562_ (.Y(_0720_),
    .A(\lif2.state[3] ),
    .B(_0719_));
 sg13g2_nand2b_1 _1563_ (.Y(_0721_),
    .B(net2),
    .A_N(_0720_));
 sg13g2_xor2_1 _1564_ (.B(_0714_),
    .A(net3),
    .X(_0722_));
 sg13g2_or2_1 _1565_ (.X(_0723_),
    .B(_0722_),
    .A(_0721_));
 sg13g2_xor2_1 _1566_ (.B(_0717_),
    .A(_0716_),
    .X(_0724_));
 sg13g2_o21ai_1 _1567_ (.B1(_0718_),
    .Y(_0725_),
    .A1(_0723_),
    .A2(_0724_));
 sg13g2_xor2_1 _1568_ (.B(_0712_),
    .A(_0711_),
    .X(_0726_));
 sg13g2_a21o_1 _1569_ (.A2(_0726_),
    .A1(_0725_),
    .B1(_0713_),
    .X(_0727_));
 sg13g2_xnor2_1 _1570_ (.Y(_0728_),
    .A(_0706_),
    .B(_0707_));
 sg13g2_a21oi_1 _1571_ (.A1(_0727_),
    .A2(_0728_),
    .Y(_0729_),
    .B1(_0708_));
 sg13g2_nand2_1 _1572_ (.Y(_0730_),
    .A(_0701_),
    .B(_0703_));
 sg13g2_a21oi_1 _1573_ (.A1(_0703_),
    .A2(_0729_),
    .Y(_0731_),
    .B1(_0702_));
 sg13g2_a21oi_1 _1574_ (.A1(_0697_),
    .A2(_0731_),
    .Y(_0732_),
    .B1(_0695_));
 sg13g2_nor2b_1 _1575_ (.A(_0689_),
    .B_N(_0686_),
    .Y(_0733_));
 sg13g2_a21oi_1 _1576_ (.A1(net9),
    .A2(_0688_),
    .Y(_0734_),
    .B1(_0733_));
 sg13g2_a21o_2 _1577_ (.A2(_0734_),
    .A1(_0732_),
    .B1(_0690_),
    .X(_0735_));
 sg13g2_xor2_1 _1578_ (.B(_0720_),
    .A(net2),
    .X(_0736_));
 sg13g2_a21oi_1 _1579_ (.A1(_0735_),
    .A2(_0736_),
    .Y(_0078_),
    .B1(net105));
 sg13g2_xnor2_1 _1580_ (.Y(_0737_),
    .A(_0721_),
    .B(_0722_));
 sg13g2_a21oi_1 _1581_ (.A1(_0735_),
    .A2(_0737_),
    .Y(_0079_),
    .B1(net105));
 sg13g2_xnor2_1 _1582_ (.Y(_0738_),
    .A(_0723_),
    .B(_0724_));
 sg13g2_a21oi_1 _1583_ (.A1(_0735_),
    .A2(_0738_),
    .Y(_0080_),
    .B1(net105));
 sg13g2_xnor2_1 _1584_ (.Y(_0739_),
    .A(_0725_),
    .B(_0726_));
 sg13g2_a21oi_1 _1585_ (.A1(_0735_),
    .A2(_0739_),
    .Y(_0081_),
    .B1(net105));
 sg13g2_xnor2_1 _1586_ (.Y(_0740_),
    .A(_0727_),
    .B(_0728_));
 sg13g2_a21oi_1 _1587_ (.A1(_0735_),
    .A2(_0740_),
    .Y(_0082_),
    .B1(net105));
 sg13g2_xnor2_1 _1588_ (.Y(_0741_),
    .A(_0729_),
    .B(_0730_));
 sg13g2_a21oi_1 _1589_ (.A1(_0735_),
    .A2(_0741_),
    .Y(_0083_),
    .B1(_0133_));
 sg13g2_xnor2_1 _1590_ (.Y(_0742_),
    .A(_0697_),
    .B(_0731_));
 sg13g2_a21oi_1 _1591_ (.A1(_0735_),
    .A2(_0742_),
    .Y(_0084_),
    .B1(net102));
 sg13g2_a21oi_1 _1592_ (.A1(_0690_),
    .A2(_0732_),
    .Y(_0085_),
    .B1(net101));
 sg13g2_nand2b_2 _1593_ (.Y(_0743_),
    .B(net106),
    .A_N(\lif2.spike ));
 sg13g2_nor2_1 _1594_ (.A(_0136_),
    .B(_0743_),
    .Y(_0086_));
 sg13g2_xnor2_1 _1595_ (.Y(_0744_),
    .A(\lif2.spike_counter[1] ),
    .B(net157));
 sg13g2_nor2_1 _1596_ (.A(_0743_),
    .B(net158),
    .Y(_0087_));
 sg13g2_and3_1 _1597_ (.X(_0745_),
    .A(net140),
    .B(\lif2.spike_counter[1] ),
    .C(net157));
 sg13g2_nand3_1 _1598_ (.B(\lif2.spike_counter[1] ),
    .C(net157),
    .A(net140),
    .Y(_0746_));
 sg13g2_a21oi_1 _1599_ (.A1(\lif2.spike_counter[1] ),
    .A2(\lif2.spike_counter[0] ),
    .Y(_0747_),
    .B1(net140));
 sg13g2_nor3_1 _1600_ (.A(_0743_),
    .B(_0745_),
    .C(net141),
    .Y(_0088_));
 sg13g2_xnor2_1 _1601_ (.Y(_0748_),
    .A(net180),
    .B(_0745_));
 sg13g2_nor2_1 _1602_ (.A(_0743_),
    .B(net181),
    .Y(_0089_));
 sg13g2_a21oi_1 _1603_ (.A1(\lif2.spike_counter[3] ),
    .A2(_0745_),
    .Y(_0749_),
    .B1(net143));
 sg13g2_nor2_1 _1604_ (.A(_0583_),
    .B(_0746_),
    .Y(_0750_));
 sg13g2_nor3_1 _1605_ (.A(_0743_),
    .B(net144),
    .C(_0750_),
    .Y(_0090_));
 sg13g2_xnor2_1 _1606_ (.Y(_0751_),
    .A(net179),
    .B(_0750_));
 sg13g2_nor2_1 _1607_ (.A(_0743_),
    .B(_0751_),
    .Y(_0091_));
 sg13g2_nor2_1 _1608_ (.A(_0605_),
    .B(_0746_),
    .Y(_0752_));
 sg13g2_a21oi_1 _1609_ (.A1(\lif2.spike_counter[5] ),
    .A2(_0750_),
    .Y(_0753_),
    .B1(net123));
 sg13g2_nor3_1 _1610_ (.A(_0743_),
    .B(_0752_),
    .C(net124),
    .Y(_0092_));
 sg13g2_xnor2_1 _1611_ (.Y(_0754_),
    .A(net135),
    .B(_0752_));
 sg13g2_nor2_1 _1612_ (.A(_0743_),
    .B(net136),
    .Y(_0093_));
 sg13g2_dfrbp_1 _1613_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net111),
    .D(net152),
    .Q_N(_0002_),
    .Q(\lif3.adapt_threshold[0] ));
 sg13g2_dfrbp_1 _1614_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net25),
    .D(_0023_),
    .Q_N(_0804_),
    .Q(\lif3.adapt_threshold[1] ));
 sg13g2_dfrbp_1 _1615_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net23),
    .D(net190),
    .Q_N(_0015_),
    .Q(\lif3.adapt_threshold[2] ));
 sg13g2_dfrbp_1 _1616_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net118),
    .D(net177),
    .Q_N(_0016_),
    .Q(\lif3.adapt_threshold[3] ));
 sg13g2_dfrbp_1 _1617_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net116),
    .D(net174),
    .Q_N(_0013_),
    .Q(\lif3.adapt_threshold[4] ));
 sg13g2_dfrbp_1 _1618_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net114),
    .D(_0027_),
    .Q_N(_0803_),
    .Q(\lif3.adapt_threshold[5] ));
 sg13g2_dfrbp_1 _1619_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net112),
    .D(_0028_),
    .Q_N(_0802_),
    .Q(\lif3.adapt_threshold[6] ));
 sg13g2_dfrbp_1 _1620_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net110),
    .D(_0029_),
    .Q_N(_0801_),
    .Q(\lif3.adapt_threshold[7] ));
 sg13g2_dfrbp_1 _1621_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net108),
    .D(_0030_),
    .Q_N(_0800_),
    .Q(\lif3.state[0] ));
 sg13g2_dfrbp_1 _1622_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net82),
    .D(_0031_),
    .Q_N(_0799_),
    .Q(\lif3.state[1] ));
 sg13g2_dfrbp_1 _1623_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net81),
    .D(_0032_),
    .Q_N(_0003_),
    .Q(\lif3.state[2] ));
 sg13g2_dfrbp_1 _1624_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net80),
    .D(_0033_),
    .Q_N(_0798_),
    .Q(\lif3.state[3] ));
 sg13g2_dfrbp_1 _1625_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net79),
    .D(_0034_),
    .Q_N(_0797_),
    .Q(\lif3.state[4] ));
 sg13g2_dfrbp_1 _1626_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net78),
    .D(_0035_),
    .Q_N(_0796_),
    .Q(\lif3.state[5] ));
 sg13g2_dfrbp_1 _1627_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net77),
    .D(_0036_),
    .Q_N(_0795_),
    .Q(\lif3.state[6] ));
 sg13g2_dfrbp_1 _1628_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net76),
    .D(_0037_),
    .Q_N(_0794_),
    .Q(\lif3.state[7] ));
 sg13g2_dfrbp_1 _1629_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net75),
    .D(_0038_),
    .Q_N(_0021_),
    .Q(\lif3.spike_counter[0] ));
 sg13g2_dfrbp_1 _1630_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net74),
    .D(_0039_),
    .Q_N(_0793_),
    .Q(\lif3.spike_counter[1] ));
 sg13g2_dfrbp_1 _1631_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net73),
    .D(net128),
    .Q_N(_0792_),
    .Q(\lif3.spike_counter[2] ));
 sg13g2_dfrbp_1 _1632_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net72),
    .D(_0041_),
    .Q_N(_0791_),
    .Q(\lif3.spike_counter[3] ));
 sg13g2_dfrbp_1 _1633_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net71),
    .D(net149),
    .Q_N(_0790_),
    .Q(\lif3.spike_counter[4] ));
 sg13g2_dfrbp_1 _1634_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net70),
    .D(_0043_),
    .Q_N(_0789_),
    .Q(\lif3.spike_counter[5] ));
 sg13g2_dfrbp_1 _1635_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net69),
    .D(_0044_),
    .Q_N(_0014_),
    .Q(\lif3.spike_counter[6] ));
 sg13g2_dfrbp_1 _1636_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net68),
    .D(_0045_),
    .Q_N(_0004_),
    .Q(\lif3.spike_counter[7] ));
 sg13g2_dfrbp_1 _1637_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net67),
    .D(_0046_),
    .Q_N(_0008_),
    .Q(\lif1.adapt_threshold[0] ));
 sg13g2_dfrbp_1 _1638_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net65),
    .D(net200),
    .Q_N(_0788_),
    .Q(\lif1.adapt_threshold[1] ));
 sg13g2_dfrbp_1 _1639_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net63),
    .D(_0048_),
    .Q_N(_0017_),
    .Q(\lif1.adapt_threshold[2] ));
 sg13g2_dfrbp_1 _1640_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net61),
    .D(net185),
    .Q_N(_0018_),
    .Q(\lif1.adapt_threshold[3] ));
 sg13g2_dfrbp_1 _1641_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net59),
    .D(net164),
    .Q_N(_0011_),
    .Q(\lif1.adapt_threshold[4] ));
 sg13g2_dfrbp_1 _1642_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net57),
    .D(_0051_),
    .Q_N(_0787_),
    .Q(\lif1.adapt_threshold[5] ));
 sg13g2_dfrbp_1 _1643_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net55),
    .D(_0052_),
    .Q_N(_0786_),
    .Q(\lif1.adapt_threshold[6] ));
 sg13g2_dfrbp_1 _1644_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net53),
    .D(net196),
    .Q_N(_0785_),
    .Q(\lif1.adapt_threshold[7] ));
 sg13g2_dfrbp_1 _1645_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net51),
    .D(_0054_),
    .Q_N(_0784_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1646_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net50),
    .D(_0055_),
    .Q_N(_0783_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1647_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net49),
    .D(_0056_),
    .Q_N(_0009_),
    .Q(net98));
 sg13g2_dfrbp_1 _1648_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net48),
    .D(_0057_),
    .Q_N(_0782_),
    .Q(net96));
 sg13g2_dfrbp_1 _1649_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net47),
    .D(_0058_),
    .Q_N(_0781_),
    .Q(net95));
 sg13g2_dfrbp_1 _1650_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net46),
    .D(_0059_),
    .Q_N(_0780_),
    .Q(net93));
 sg13g2_dfrbp_1 _1651_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net45),
    .D(_0060_),
    .Q_N(_0779_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1652_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net44),
    .D(_0061_),
    .Q_N(_0778_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _1653_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net43),
    .D(_0062_),
    .Q_N(_0020_),
    .Q(\lif1.spike_counter[0] ));
 sg13g2_dfrbp_1 _1654_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net42),
    .D(_0063_),
    .Q_N(_0777_),
    .Q(\lif1.spike_counter[1] ));
 sg13g2_dfrbp_1 _1655_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net41),
    .D(net139),
    .Q_N(_0776_),
    .Q(\lif1.spike_counter[2] ));
 sg13g2_dfrbp_1 _1656_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net40),
    .D(_0065_),
    .Q_N(_0775_),
    .Q(\lif1.spike_counter[3] ));
 sg13g2_dfrbp_1 _1657_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net39),
    .D(_0066_),
    .Q_N(_0774_),
    .Q(\lif1.spike_counter[4] ));
 sg13g2_dfrbp_1 _1658_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net38),
    .D(_0067_),
    .Q_N(_0773_),
    .Q(\lif1.spike_counter[5] ));
 sg13g2_dfrbp_1 _1659_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net37),
    .D(_0068_),
    .Q_N(_0772_),
    .Q(\lif1.spike_counter[6] ));
 sg13g2_dfrbp_1 _1660_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net36),
    .D(_0069_),
    .Q_N(_0010_),
    .Q(\lif1.spike_counter[7] ));
 sg13g2_dfrbp_1 _1661_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net35),
    .D(net134),
    .Q_N(_0005_),
    .Q(\lif2.adapt_threshold[0] ));
 sg13g2_dfrbp_1 _1662_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net33),
    .D(net198),
    .Q_N(_0771_),
    .Q(\lif2.adapt_threshold[1] ));
 sg13g2_dfrbp_1 _1663_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net31),
    .D(_0072_),
    .Q_N(_0000_),
    .Q(\lif2.adapt_threshold[2] ));
 sg13g2_dfrbp_1 _1664_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net29),
    .D(net183),
    .Q_N(_0001_),
    .Q(\lif2.adapt_threshold[3] ));
 sg13g2_dfrbp_1 _1665_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net27),
    .D(net168),
    .Q_N(_0012_),
    .Q(\lif2.adapt_threshold[4] ));
 sg13g2_dfrbp_1 _1666_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net24),
    .D(_0075_),
    .Q_N(_0770_),
    .Q(\lif2.adapt_threshold[5] ));
 sg13g2_dfrbp_1 _1667_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net117),
    .D(_0076_),
    .Q_N(_0769_),
    .Q(\lif2.adapt_threshold[6] ));
 sg13g2_dfrbp_1 _1668_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net113),
    .D(_0077_),
    .Q_N(_0768_),
    .Q(\lif2.adapt_threshold[7] ));
 sg13g2_dfrbp_1 _1669_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net109),
    .D(_0078_),
    .Q_N(_0767_),
    .Q(\lif2.state[0] ));
 sg13g2_dfrbp_1 _1670_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net66),
    .D(_0079_),
    .Q_N(_0766_),
    .Q(\lif2.state[1] ));
 sg13g2_dfrbp_1 _1671_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net64),
    .D(_0080_),
    .Q_N(_0006_),
    .Q(\lif2.state[2] ));
 sg13g2_dfrbp_1 _1672_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net62),
    .D(_0081_),
    .Q_N(_0765_),
    .Q(\lif2.state[3] ));
 sg13g2_dfrbp_1 _1673_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net60),
    .D(_0082_),
    .Q_N(_0764_),
    .Q(\lif2.state[4] ));
 sg13g2_dfrbp_1 _1674_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net58),
    .D(_0083_),
    .Q_N(_0763_),
    .Q(\lif2.state[5] ));
 sg13g2_dfrbp_1 _1675_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net56),
    .D(_0084_),
    .Q_N(_0762_),
    .Q(\lif2.state[6] ));
 sg13g2_dfrbp_1 _1676_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net54),
    .D(_0085_),
    .Q_N(_0761_),
    .Q(\lif2.state[7] ));
 sg13g2_dfrbp_1 _1677_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net52),
    .D(_0086_),
    .Q_N(_0019_),
    .Q(\lif2.spike_counter[0] ));
 sg13g2_dfrbp_1 _1678_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net34),
    .D(_0087_),
    .Q_N(_0760_),
    .Q(\lif2.spike_counter[1] ));
 sg13g2_dfrbp_1 _1679_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net32),
    .D(net142),
    .Q_N(_0759_),
    .Q(\lif2.spike_counter[2] ));
 sg13g2_dfrbp_1 _1680_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net30),
    .D(_0089_),
    .Q_N(_0758_),
    .Q(\lif2.spike_counter[3] ));
 sg13g2_dfrbp_1 _1681_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net28),
    .D(_0090_),
    .Q_N(_0757_),
    .Q(\lif2.spike_counter[4] ));
 sg13g2_dfrbp_1 _1682_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net26),
    .D(_0091_),
    .Q_N(_0756_),
    .Q(\lif2.spike_counter[5] ));
 sg13g2_dfrbp_1 _1683_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net22),
    .D(net125),
    .Q_N(_0755_),
    .Q(\lif2.spike_counter[6] ));
 sg13g2_dfrbp_1 _1684_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net115),
    .D(_0093_),
    .Q_N(_0007_),
    .Q(\lif2.spike_counter[7] ));
 sg13g2_tiehi _1615__23 (.L_HI(net23));
 sg13g2_tiehi _1666__24 (.L_HI(net24));
 sg13g2_tiehi _1614__25 (.L_HI(net25));
 sg13g2_tiehi _1682__26 (.L_HI(net26));
 sg13g2_tiehi _1665__27 (.L_HI(net27));
 sg13g2_tiehi _1681__28 (.L_HI(net28));
 sg13g2_tiehi _1664__29 (.L_HI(net29));
 sg13g2_tiehi _1680__30 (.L_HI(net30));
 sg13g2_tiehi _1663__31 (.L_HI(net31));
 sg13g2_tiehi _1679__32 (.L_HI(net32));
 sg13g2_tiehi _1662__33 (.L_HI(net33));
 sg13g2_tiehi _1678__34 (.L_HI(net34));
 sg13g2_tiehi _1661__35 (.L_HI(net35));
 sg13g2_tiehi _1660__36 (.L_HI(net36));
 sg13g2_tiehi _1659__37 (.L_HI(net37));
 sg13g2_tiehi _1658__38 (.L_HI(net38));
 sg13g2_tiehi _1657__39 (.L_HI(net39));
 sg13g2_tiehi _1656__40 (.L_HI(net40));
 sg13g2_tiehi _1655__41 (.L_HI(net41));
 sg13g2_tiehi _1654__42 (.L_HI(net42));
 sg13g2_tiehi _1653__43 (.L_HI(net43));
 sg13g2_tiehi _1652__44 (.L_HI(net44));
 sg13g2_tiehi _1651__45 (.L_HI(net45));
 sg13g2_tiehi _1650__46 (.L_HI(net46));
 sg13g2_tiehi _1649__47 (.L_HI(net47));
 sg13g2_tiehi _1648__48 (.L_HI(net48));
 sg13g2_tiehi _1647__49 (.L_HI(net49));
 sg13g2_tiehi _1646__50 (.L_HI(net50));
 sg13g2_tiehi _1645__51 (.L_HI(net51));
 sg13g2_tiehi _1677__52 (.L_HI(net52));
 sg13g2_tiehi _1644__53 (.L_HI(net53));
 sg13g2_tiehi _1676__54 (.L_HI(net54));
 sg13g2_tiehi _1643__55 (.L_HI(net55));
 sg13g2_tiehi _1675__56 (.L_HI(net56));
 sg13g2_tiehi _1642__57 (.L_HI(net57));
 sg13g2_tiehi _1674__58 (.L_HI(net58));
 sg13g2_tiehi _1641__59 (.L_HI(net59));
 sg13g2_tiehi _1673__60 (.L_HI(net60));
 sg13g2_tiehi _1640__61 (.L_HI(net61));
 sg13g2_tiehi _1672__62 (.L_HI(net62));
 sg13g2_tiehi _1639__63 (.L_HI(net63));
 sg13g2_tiehi _1671__64 (.L_HI(net64));
 sg13g2_tiehi _1638__65 (.L_HI(net65));
 sg13g2_tiehi _1670__66 (.L_HI(net66));
 sg13g2_tiehi _1637__67 (.L_HI(net67));
 sg13g2_tiehi _1636__68 (.L_HI(net68));
 sg13g2_tiehi _1635__69 (.L_HI(net69));
 sg13g2_tiehi _1634__70 (.L_HI(net70));
 sg13g2_tiehi _1633__71 (.L_HI(net71));
 sg13g2_tiehi _1632__72 (.L_HI(net72));
 sg13g2_tiehi _1631__73 (.L_HI(net73));
 sg13g2_tiehi _1630__74 (.L_HI(net74));
 sg13g2_tiehi _1629__75 (.L_HI(net75));
 sg13g2_tiehi _1628__76 (.L_HI(net76));
 sg13g2_tiehi _1627__77 (.L_HI(net77));
 sg13g2_tiehi _1626__78 (.L_HI(net78));
 sg13g2_tiehi _1625__79 (.L_HI(net79));
 sg13g2_tiehi _1624__80 (.L_HI(net80));
 sg13g2_tiehi _1623__81 (.L_HI(net81));
 sg13g2_tiehi _1622__82 (.L_HI(net82));
 sg13g2_tiehi _1621__83 (.L_HI(net108));
 sg13g2_tiehi _1669__84 (.L_HI(net109));
 sg13g2_tiehi _1620__85 (.L_HI(net110));
 sg13g2_tiehi _1613__86 (.L_HI(net111));
 sg13g2_tiehi _1619__87 (.L_HI(net112));
 sg13g2_tiehi _1668__88 (.L_HI(net113));
 sg13g2_tiehi _1618__89 (.L_HI(net114));
 sg13g2_tiehi _1684__90 (.L_HI(net115));
 sg13g2_tiehi _1617__91 (.L_HI(net116));
 sg13g2_tiehi _1667__92 (.L_HI(net117));
 sg13g2_tiehi _1616__93 (.L_HI(net118));
 sg13g2_tiehi tt_um_alif_94 (.L_HI(net119));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_alif_11 (.L_LO(net11));
 sg13g2_tielo tt_um_alif_12 (.L_LO(net12));
 sg13g2_tielo tt_um_alif_13 (.L_LO(net13));
 sg13g2_tielo tt_um_alif_14 (.L_LO(net14));
 sg13g2_tielo tt_um_alif_15 (.L_LO(net15));
 sg13g2_tielo tt_um_alif_16 (.L_LO(net16));
 sg13g2_tielo tt_um_alif_17 (.L_LO(net17));
 sg13g2_tielo tt_um_alif_18 (.L_LO(net18));
 sg13g2_tielo tt_um_alif_19 (.L_LO(net19));
 sg13g2_tielo tt_um_alif_20 (.L_LO(net20));
 sg13g2_tielo tt_um_alif_21 (.L_LO(net21));
 sg13g2_tiehi _1683__22 (.L_HI(net22));
 sg13g2_buf_2 _1770_ (.A(\lif3.spike ),
    .X(uio_out[5]));
 sg13g2_buf_1 _1771_ (.A(\lif2.spike ),
    .X(uio_out[6]));
 sg13g2_buf_1 _1772_ (.A(\lif1.spike ),
    .X(uio_out[7]));
 sg13g2_buf_2 fanout83 (.A(_0182_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(net85),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0577_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(net87),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0367_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0571_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0361_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0175_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(\lif2.state[5] ),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(\lif2.state[2] ),
    .X(net92));
 sg13g2_buf_4 fanout93 (.X(uo_out[5]),
    .A(net93));
 sg13g2_buf_1 fanout94 (.A(net93),
    .X(net94));
 sg13g2_buf_4 fanout95 (.X(uo_out[4]),
    .A(net95));
 sg13g2_buf_2 fanout96 (.A(net97),
    .X(uo_out[3]));
 sg13g2_buf_2 fanout97 (.A(net96),
    .X(net97));
 sg13g2_buf_4 fanout98 (.X(uo_out[2]),
    .A(net98));
 sg13g2_buf_2 fanout99 (.A(\lif3.state[6] ),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(\lif3.state[5] ),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(net102),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_0133_),
    .X(net102));
 sg13g2_buf_4 fanout103 (.X(net103),
    .A(net104));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(net105));
 sg13g2_buf_2 fanout105 (.A(_0133_),
    .X(net105));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(net107));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(net1));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[0]));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[1]));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[2]));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[3]));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[4]));
 sg13g2_buf_2 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_4 input9 (.X(net9),
    .A(ui_in[7]));
 sg13g2_tielo tt_um_alif_10 (.L_LO(net10));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0019_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0021_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0020_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold4 (.A(\lif2.spike_counter[6] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0753_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0092_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold7 (.A(\lif3.spike_counter[2] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0344_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0040_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold10 (.A(\lif3.spike_counter[7] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0352_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold12 (.A(\lif1.spike_counter[7] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0562_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold14 (.A(\lif2.adapt_threshold[0] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0070_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold16 (.A(\lif2.spike_counter[7] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0754_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold18 (.A(\lif1.spike_counter[2] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0555_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0064_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold21 (.A(\lif2.spike_counter[2] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0747_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0088_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold24 (.A(\lif2.spike_counter[4] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0749_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold26 (.A(\lif1.spike_counter[6] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0561_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold28 (.A(\lif3.spike_counter[4] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0346_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0042_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0002_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0185_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0022_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold34 (.A(\lif3.spike_counter[5] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0349_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold36 (.A(\lif3.spike_counter[6] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0350_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold38 (.A(\lif2.spike_counter[0] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0744_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold40 (.A(\lif1.spike_counter[4] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0557_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold42 (.A(\lif3.spike_counter[0] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0341_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold44 (.A(\lif1.adapt_threshold[4] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0050_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold46 (.A(\lif1.spike_counter[0] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0552_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold48 (.A(\lif2.adapt_threshold[4] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0074_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold50 (.A(\lif2.adapt_threshold[5] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold51 (.A(\lif1.adapt_threshold[5] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold52 (.A(\lif1.spike_counter[5] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0559_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold54 (.A(\lif3.adapt_threshold[4] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0026_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold56 (.A(\lif3.adapt_threshold[1] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold57 (.A(\lif3.adapt_threshold[3] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0025_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold59 (.A(\lif3.adapt_threshold[7] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold60 (.A(\lif2.spike_counter[5] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold61 (.A(\lif2.spike_counter[3] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0748_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold63 (.A(\lif2.adapt_threshold[3] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0073_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold65 (.A(\lif1.adapt_threshold[3] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0049_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold67 (.A(\lif2.adapt_threshold[7] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold68 (.A(\lif3.spike_counter[3] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0345_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold70 (.A(\lif3.adapt_threshold[2] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0024_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold72 (.A(\lif3.adapt_threshold[5] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold73 (.A(\lif1.spike_counter[3] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0556_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold75 (.A(\lif3.adapt_threshold[6] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold76 (.A(\lif1.adapt_threshold[7] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0053_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold78 (.A(\lif2.adapt_threshold[1] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0071_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold80 (.A(\lif1.adapt_threshold[1] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0047_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold82 (.A(\lif2.adapt_threshold[6] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold83 (.A(\lif2.adapt_threshold[2] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0602_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold85 (.A(\lif1.adapt_threshold[6] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold86 (.A(\lif1.adapt_threshold[0] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0371_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold88 (.A(\lif1.adapt_threshold[2] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold89 (.A(\lif3.adapt_threshold[7] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold90 (.A(\lif3.spike_counter[0] ),
    .X(net209));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_4 FILLER_8_168 ();
 sg13g2_fill_1 FILLER_8_172 ();
 sg13g2_decap_8 FILLER_8_181 ();
 sg13g2_decap_8 FILLER_8_188 ();
 sg13g2_decap_8 FILLER_8_195 ();
 sg13g2_decap_8 FILLER_8_202 ();
 sg13g2_decap_8 FILLER_8_209 ();
 sg13g2_decap_8 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_223 ();
 sg13g2_decap_8 FILLER_8_230 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_decap_8 FILLER_8_251 ();
 sg13g2_decap_8 FILLER_8_258 ();
 sg13g2_decap_8 FILLER_8_265 ();
 sg13g2_decap_8 FILLER_8_272 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_decap_8 FILLER_8_286 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_321 ();
 sg13g2_decap_8 FILLER_8_328 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_4 FILLER_9_157 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_decap_4 FILLER_9_171 ();
 sg13g2_fill_2 FILLER_9_184 ();
 sg13g2_decap_8 FILLER_9_191 ();
 sg13g2_decap_8 FILLER_9_198 ();
 sg13g2_decap_8 FILLER_9_205 ();
 sg13g2_decap_8 FILLER_9_212 ();
 sg13g2_decap_8 FILLER_9_219 ();
 sg13g2_decap_8 FILLER_9_226 ();
 sg13g2_decap_8 FILLER_9_233 ();
 sg13g2_decap_8 FILLER_9_240 ();
 sg13g2_decap_8 FILLER_9_247 ();
 sg13g2_decap_8 FILLER_9_254 ();
 sg13g2_decap_8 FILLER_9_261 ();
 sg13g2_decap_8 FILLER_9_268 ();
 sg13g2_decap_8 FILLER_9_275 ();
 sg13g2_decap_8 FILLER_9_282 ();
 sg13g2_decap_8 FILLER_9_289 ();
 sg13g2_decap_8 FILLER_9_296 ();
 sg13g2_decap_8 FILLER_9_303 ();
 sg13g2_decap_8 FILLER_9_310 ();
 sg13g2_decap_8 FILLER_9_317 ();
 sg13g2_decap_8 FILLER_9_324 ();
 sg13g2_decap_8 FILLER_9_331 ();
 sg13g2_decap_8 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_345 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_decap_8 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_fill_2 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_220 ();
 sg13g2_decap_8 FILLER_10_227 ();
 sg13g2_decap_8 FILLER_10_234 ();
 sg13g2_decap_8 FILLER_10_241 ();
 sg13g2_decap_8 FILLER_10_248 ();
 sg13g2_decap_8 FILLER_10_255 ();
 sg13g2_decap_8 FILLER_10_262 ();
 sg13g2_decap_8 FILLER_10_269 ();
 sg13g2_decap_8 FILLER_10_276 ();
 sg13g2_decap_8 FILLER_10_283 ();
 sg13g2_decap_8 FILLER_10_290 ();
 sg13g2_decap_8 FILLER_10_297 ();
 sg13g2_decap_8 FILLER_10_304 ();
 sg13g2_decap_8 FILLER_10_311 ();
 sg13g2_decap_8 FILLER_10_318 ();
 sg13g2_decap_8 FILLER_10_325 ();
 sg13g2_decap_8 FILLER_10_332 ();
 sg13g2_decap_8 FILLER_10_339 ();
 sg13g2_decap_8 FILLER_10_346 ();
 sg13g2_decap_8 FILLER_10_353 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_4 FILLER_11_119 ();
 sg13g2_fill_1 FILLER_11_128 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_fill_2 FILLER_11_140 ();
 sg13g2_fill_2 FILLER_11_154 ();
 sg13g2_fill_1 FILLER_11_156 ();
 sg13g2_fill_1 FILLER_11_183 ();
 sg13g2_decap_8 FILLER_11_226 ();
 sg13g2_decap_8 FILLER_11_233 ();
 sg13g2_decap_8 FILLER_11_240 ();
 sg13g2_decap_8 FILLER_11_247 ();
 sg13g2_decap_8 FILLER_11_254 ();
 sg13g2_decap_8 FILLER_11_261 ();
 sg13g2_decap_8 FILLER_11_268 ();
 sg13g2_decap_8 FILLER_11_275 ();
 sg13g2_decap_8 FILLER_11_282 ();
 sg13g2_decap_8 FILLER_11_289 ();
 sg13g2_decap_8 FILLER_11_296 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_decap_8 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_317 ();
 sg13g2_decap_8 FILLER_11_324 ();
 sg13g2_decap_8 FILLER_11_331 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_decap_8 FILLER_11_345 ();
 sg13g2_decap_8 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_fill_2 FILLER_12_116 ();
 sg13g2_fill_2 FILLER_12_201 ();
 sg13g2_fill_1 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_4 FILLER_13_84 ();
 sg13g2_fill_1 FILLER_13_88 ();
 sg13g2_fill_2 FILLER_13_141 ();
 sg13g2_fill_1 FILLER_13_162 ();
 sg13g2_fill_1 FILLER_13_187 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_4 FILLER_14_95 ();
 sg13g2_fill_1 FILLER_14_99 ();
 sg13g2_fill_2 FILLER_14_104 ();
 sg13g2_fill_1 FILLER_14_106 ();
 sg13g2_fill_1 FILLER_14_133 ();
 sg13g2_fill_2 FILLER_14_138 ();
 sg13g2_decap_4 FILLER_14_152 ();
 sg13g2_fill_1 FILLER_14_172 ();
 sg13g2_fill_2 FILLER_14_190 ();
 sg13g2_fill_1 FILLER_14_192 ();
 sg13g2_fill_1 FILLER_14_206 ();
 sg13g2_fill_2 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_251 ();
 sg13g2_decap_8 FILLER_14_258 ();
 sg13g2_decap_8 FILLER_14_265 ();
 sg13g2_decap_8 FILLER_14_272 ();
 sg13g2_decap_8 FILLER_14_279 ();
 sg13g2_decap_8 FILLER_14_286 ();
 sg13g2_decap_8 FILLER_14_293 ();
 sg13g2_decap_8 FILLER_14_300 ();
 sg13g2_decap_8 FILLER_14_307 ();
 sg13g2_decap_8 FILLER_14_314 ();
 sg13g2_decap_8 FILLER_14_321 ();
 sg13g2_decap_8 FILLER_14_328 ();
 sg13g2_decap_8 FILLER_14_335 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_356 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_fill_2 FILLER_15_63 ();
 sg13g2_fill_1 FILLER_15_74 ();
 sg13g2_fill_2 FILLER_15_106 ();
 sg13g2_fill_1 FILLER_15_108 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_196 ();
 sg13g2_fill_1 FILLER_15_207 ();
 sg13g2_fill_1 FILLER_15_221 ();
 sg13g2_fill_2 FILLER_15_231 ();
 sg13g2_fill_1 FILLER_15_233 ();
 sg13g2_decap_8 FILLER_15_258 ();
 sg13g2_decap_8 FILLER_15_265 ();
 sg13g2_decap_8 FILLER_15_272 ();
 sg13g2_decap_8 FILLER_15_279 ();
 sg13g2_decap_8 FILLER_15_286 ();
 sg13g2_decap_8 FILLER_15_293 ();
 sg13g2_decap_8 FILLER_15_300 ();
 sg13g2_decap_8 FILLER_15_307 ();
 sg13g2_decap_8 FILLER_15_314 ();
 sg13g2_decap_8 FILLER_15_321 ();
 sg13g2_decap_8 FILLER_15_328 ();
 sg13g2_decap_8 FILLER_15_335 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_decap_8 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_49 ();
 sg13g2_fill_1 FILLER_16_79 ();
 sg13g2_fill_1 FILLER_16_99 ();
 sg13g2_decap_4 FILLER_16_117 ();
 sg13g2_fill_1 FILLER_16_130 ();
 sg13g2_fill_1 FILLER_16_150 ();
 sg13g2_fill_2 FILLER_16_160 ();
 sg13g2_fill_1 FILLER_16_162 ();
 sg13g2_decap_4 FILLER_16_204 ();
 sg13g2_decap_4 FILLER_16_213 ();
 sg13g2_fill_1 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_262 ();
 sg13g2_decap_8 FILLER_16_269 ();
 sg13g2_decap_8 FILLER_16_276 ();
 sg13g2_decap_8 FILLER_16_283 ();
 sg13g2_decap_8 FILLER_16_290 ();
 sg13g2_decap_8 FILLER_16_297 ();
 sg13g2_decap_8 FILLER_16_304 ();
 sg13g2_decap_8 FILLER_16_311 ();
 sg13g2_decap_8 FILLER_16_318 ();
 sg13g2_decap_8 FILLER_16_325 ();
 sg13g2_decap_8 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_4 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_60 ();
 sg13g2_fill_1 FILLER_17_92 ();
 sg13g2_fill_1 FILLER_17_106 ();
 sg13g2_fill_2 FILLER_17_117 ();
 sg13g2_fill_2 FILLER_17_124 ();
 sg13g2_fill_1 FILLER_17_134 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_fill_2 FILLER_17_150 ();
 sg13g2_fill_1 FILLER_17_152 ();
 sg13g2_fill_2 FILLER_17_183 ();
 sg13g2_fill_1 FILLER_17_185 ();
 sg13g2_fill_2 FILLER_17_190 ();
 sg13g2_fill_1 FILLER_17_192 ();
 sg13g2_decap_4 FILLER_17_214 ();
 sg13g2_decap_4 FILLER_17_223 ();
 sg13g2_fill_2 FILLER_17_227 ();
 sg13g2_fill_2 FILLER_17_239 ();
 sg13g2_fill_1 FILLER_17_241 ();
 sg13g2_fill_1 FILLER_17_251 ();
 sg13g2_decap_8 FILLER_17_269 ();
 sg13g2_decap_8 FILLER_17_276 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_decap_8 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_297 ();
 sg13g2_decap_8 FILLER_17_304 ();
 sg13g2_decap_8 FILLER_17_311 ();
 sg13g2_decap_8 FILLER_17_318 ();
 sg13g2_decap_8 FILLER_17_325 ();
 sg13g2_decap_8 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_fill_2 FILLER_18_61 ();
 sg13g2_fill_1 FILLER_18_97 ();
 sg13g2_fill_2 FILLER_18_118 ();
 sg13g2_fill_1 FILLER_18_135 ();
 sg13g2_decap_8 FILLER_18_156 ();
 sg13g2_decap_4 FILLER_18_163 ();
 sg13g2_fill_1 FILLER_18_167 ();
 sg13g2_fill_2 FILLER_18_172 ();
 sg13g2_fill_1 FILLER_18_174 ();
 sg13g2_fill_2 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_decap_8 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_229 ();
 sg13g2_decap_8 FILLER_18_265 ();
 sg13g2_decap_8 FILLER_18_272 ();
 sg13g2_decap_8 FILLER_18_279 ();
 sg13g2_decap_8 FILLER_18_286 ();
 sg13g2_decap_8 FILLER_18_293 ();
 sg13g2_decap_8 FILLER_18_300 ();
 sg13g2_decap_8 FILLER_18_307 ();
 sg13g2_decap_8 FILLER_18_314 ();
 sg13g2_decap_8 FILLER_18_321 ();
 sg13g2_decap_8 FILLER_18_328 ();
 sg13g2_decap_8 FILLER_18_335 ();
 sg13g2_decap_8 FILLER_18_342 ();
 sg13g2_decap_8 FILLER_18_349 ();
 sg13g2_decap_8 FILLER_18_356 ();
 sg13g2_decap_8 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_18_370 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_4 FILLER_19_42 ();
 sg13g2_decap_4 FILLER_19_50 ();
 sg13g2_fill_1 FILLER_19_54 ();
 sg13g2_decap_4 FILLER_19_77 ();
 sg13g2_fill_2 FILLER_19_89 ();
 sg13g2_fill_2 FILLER_19_104 ();
 sg13g2_decap_4 FILLER_19_115 ();
 sg13g2_fill_2 FILLER_19_137 ();
 sg13g2_fill_1 FILLER_19_139 ();
 sg13g2_fill_2 FILLER_19_143 ();
 sg13g2_decap_8 FILLER_19_166 ();
 sg13g2_decap_4 FILLER_19_173 ();
 sg13g2_fill_1 FILLER_19_193 ();
 sg13g2_fill_2 FILLER_19_212 ();
 sg13g2_fill_2 FILLER_19_223 ();
 sg13g2_fill_1 FILLER_19_225 ();
 sg13g2_decap_8 FILLER_19_233 ();
 sg13g2_fill_2 FILLER_19_258 ();
 sg13g2_fill_1 FILLER_19_260 ();
 sg13g2_decap_8 FILLER_19_265 ();
 sg13g2_decap_8 FILLER_19_272 ();
 sg13g2_decap_8 FILLER_19_279 ();
 sg13g2_decap_8 FILLER_19_286 ();
 sg13g2_decap_8 FILLER_19_293 ();
 sg13g2_decap_8 FILLER_19_300 ();
 sg13g2_decap_8 FILLER_19_307 ();
 sg13g2_decap_8 FILLER_19_314 ();
 sg13g2_decap_8 FILLER_19_321 ();
 sg13g2_decap_8 FILLER_19_328 ();
 sg13g2_decap_8 FILLER_19_335 ();
 sg13g2_decap_8 FILLER_19_342 ();
 sg13g2_decap_8 FILLER_19_349 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_19_370 ();
 sg13g2_decap_8 FILLER_19_377 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_fill_1 FILLER_20_21 ();
 sg13g2_fill_1 FILLER_20_26 ();
 sg13g2_fill_2 FILLER_20_55 ();
 sg13g2_fill_1 FILLER_20_61 ();
 sg13g2_fill_1 FILLER_20_78 ();
 sg13g2_fill_2 FILLER_20_105 ();
 sg13g2_fill_2 FILLER_20_124 ();
 sg13g2_fill_1 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_136 ();
 sg13g2_decap_4 FILLER_20_143 ();
 sg13g2_fill_1 FILLER_20_147 ();
 sg13g2_decap_4 FILLER_20_176 ();
 sg13g2_decap_4 FILLER_20_193 ();
 sg13g2_fill_1 FILLER_20_201 ();
 sg13g2_decap_4 FILLER_20_227 ();
 sg13g2_fill_2 FILLER_20_231 ();
 sg13g2_fill_2 FILLER_20_247 ();
 sg13g2_fill_1 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_276 ();
 sg13g2_decap_8 FILLER_20_283 ();
 sg13g2_decap_8 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_297 ();
 sg13g2_decap_8 FILLER_20_304 ();
 sg13g2_decap_8 FILLER_20_311 ();
 sg13g2_decap_4 FILLER_20_318 ();
 sg13g2_fill_1 FILLER_20_327 ();
 sg13g2_decap_8 FILLER_20_332 ();
 sg13g2_decap_8 FILLER_20_339 ();
 sg13g2_decap_4 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_15 ();
 sg13g2_fill_1 FILLER_21_17 ();
 sg13g2_fill_2 FILLER_21_44 ();
 sg13g2_fill_1 FILLER_21_46 ();
 sg13g2_fill_1 FILLER_21_73 ();
 sg13g2_decap_8 FILLER_21_79 ();
 sg13g2_fill_2 FILLER_21_86 ();
 sg13g2_fill_1 FILLER_21_88 ();
 sg13g2_decap_8 FILLER_21_93 ();
 sg13g2_decap_8 FILLER_21_100 ();
 sg13g2_decap_8 FILLER_21_107 ();
 sg13g2_fill_2 FILLER_21_114 ();
 sg13g2_fill_1 FILLER_21_116 ();
 sg13g2_fill_2 FILLER_21_120 ();
 sg13g2_fill_1 FILLER_21_122 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_fill_1 FILLER_21_189 ();
 sg13g2_fill_2 FILLER_21_214 ();
 sg13g2_fill_1 FILLER_21_216 ();
 sg13g2_fill_2 FILLER_21_238 ();
 sg13g2_fill_1 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_272 ();
 sg13g2_decap_8 FILLER_21_279 ();
 sg13g2_decap_8 FILLER_21_286 ();
 sg13g2_decap_4 FILLER_21_314 ();
 sg13g2_decap_8 FILLER_21_374 ();
 sg13g2_decap_8 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_4 ();
 sg13g2_fill_1 FILLER_22_36 ();
 sg13g2_fill_2 FILLER_22_60 ();
 sg13g2_fill_1 FILLER_22_62 ();
 sg13g2_decap_4 FILLER_22_115 ();
 sg13g2_decap_4 FILLER_22_123 ();
 sg13g2_fill_1 FILLER_22_127 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_fill_2 FILLER_22_147 ();
 sg13g2_fill_1 FILLER_22_157 ();
 sg13g2_decap_8 FILLER_22_166 ();
 sg13g2_decap_4 FILLER_22_173 ();
 sg13g2_fill_2 FILLER_22_177 ();
 sg13g2_decap_8 FILLER_22_184 ();
 sg13g2_decap_8 FILLER_22_191 ();
 sg13g2_decap_4 FILLER_22_198 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_decap_8 FILLER_22_211 ();
 sg13g2_decap_4 FILLER_22_218 ();
 sg13g2_fill_2 FILLER_22_222 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_fill_2 FILLER_22_235 ();
 sg13g2_fill_1 FILLER_22_237 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_260 ();
 sg13g2_decap_8 FILLER_22_267 ();
 sg13g2_decap_4 FILLER_22_274 ();
 sg13g2_fill_1 FILLER_22_278 ();
 sg13g2_decap_4 FILLER_22_284 ();
 sg13g2_fill_1 FILLER_22_288 ();
 sg13g2_fill_2 FILLER_22_319 ();
 sg13g2_fill_1 FILLER_22_321 ();
 sg13g2_fill_1 FILLER_22_331 ();
 sg13g2_fill_2 FILLER_22_359 ();
 sg13g2_fill_1 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_4 FILLER_23_90 ();
 sg13g2_decap_4 FILLER_23_124 ();
 sg13g2_decap_8 FILLER_23_141 ();
 sg13g2_decap_8 FILLER_23_148 ();
 sg13g2_fill_2 FILLER_23_155 ();
 sg13g2_fill_1 FILLER_23_157 ();
 sg13g2_fill_2 FILLER_23_210 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_fill_1 FILLER_23_239 ();
 sg13g2_decap_4 FILLER_23_258 ();
 sg13g2_fill_1 FILLER_23_262 ();
 sg13g2_fill_1 FILLER_23_301 ();
 sg13g2_fill_2 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_51 ();
 sg13g2_fill_1 FILLER_24_62 ();
 sg13g2_fill_2 FILLER_24_72 ();
 sg13g2_decap_4 FILLER_24_95 ();
 sg13g2_fill_1 FILLER_24_109 ();
 sg13g2_decap_8 FILLER_24_115 ();
 sg13g2_decap_8 FILLER_24_122 ();
 sg13g2_decap_4 FILLER_24_144 ();
 sg13g2_fill_1 FILLER_24_148 ();
 sg13g2_fill_2 FILLER_24_167 ();
 sg13g2_decap_8 FILLER_24_173 ();
 sg13g2_fill_2 FILLER_24_180 ();
 sg13g2_fill_1 FILLER_24_182 ();
 sg13g2_fill_1 FILLER_24_188 ();
 sg13g2_fill_2 FILLER_24_209 ();
 sg13g2_decap_8 FILLER_24_216 ();
 sg13g2_fill_2 FILLER_24_223 ();
 sg13g2_fill_2 FILLER_24_238 ();
 sg13g2_fill_1 FILLER_24_240 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_fill_2 FILLER_24_266 ();
 sg13g2_fill_1 FILLER_24_314 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_4 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_102 ();
 sg13g2_fill_1 FILLER_25_122 ();
 sg13g2_fill_1 FILLER_25_146 ();
 sg13g2_decap_4 FILLER_25_167 ();
 sg13g2_fill_1 FILLER_25_171 ();
 sg13g2_fill_2 FILLER_25_189 ();
 sg13g2_fill_2 FILLER_25_236 ();
 sg13g2_decap_8 FILLER_25_246 ();
 sg13g2_decap_8 FILLER_25_253 ();
 sg13g2_fill_2 FILLER_25_260 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_fill_2 FILLER_25_273 ();
 sg13g2_fill_2 FILLER_25_280 ();
 sg13g2_fill_2 FILLER_25_291 ();
 sg13g2_fill_2 FILLER_25_297 ();
 sg13g2_fill_1 FILLER_25_303 ();
 sg13g2_fill_2 FILLER_25_321 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_328 ();
 sg13g2_fill_2 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_68 ();
 sg13g2_fill_2 FILLER_26_85 ();
 sg13g2_fill_1 FILLER_26_95 ();
 sg13g2_fill_2 FILLER_26_110 ();
 sg13g2_decap_8 FILLER_26_120 ();
 sg13g2_fill_2 FILLER_26_127 ();
 sg13g2_fill_1 FILLER_26_129 ();
 sg13g2_fill_1 FILLER_26_148 ();
 sg13g2_fill_2 FILLER_26_158 ();
 sg13g2_fill_1 FILLER_26_160 ();
 sg13g2_fill_2 FILLER_26_166 ();
 sg13g2_fill_1 FILLER_26_176 ();
 sg13g2_decap_8 FILLER_26_190 ();
 sg13g2_decap_4 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_decap_4 FILLER_26_223 ();
 sg13g2_fill_2 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_249 ();
 sg13g2_fill_1 FILLER_26_251 ();
 sg13g2_fill_1 FILLER_26_278 ();
 sg13g2_fill_2 FILLER_26_284 ();
 sg13g2_fill_1 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_292 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_fill_2 FILLER_26_316 ();
 sg13g2_fill_1 FILLER_26_318 ();
 sg13g2_fill_1 FILLER_26_345 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_fill_2 FILLER_26_384 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_fill_2 FILLER_27_47 ();
 sg13g2_fill_1 FILLER_27_70 ();
 sg13g2_fill_2 FILLER_27_89 ();
 sg13g2_fill_1 FILLER_27_101 ();
 sg13g2_fill_2 FILLER_27_128 ();
 sg13g2_fill_2 FILLER_27_133 ();
 sg13g2_fill_1 FILLER_27_135 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_fill_1 FILLER_27_147 ();
 sg13g2_fill_2 FILLER_27_156 ();
 sg13g2_decap_8 FILLER_27_184 ();
 sg13g2_fill_2 FILLER_27_191 ();
 sg13g2_fill_1 FILLER_27_193 ();
 sg13g2_fill_1 FILLER_27_215 ();
 sg13g2_decap_4 FILLER_27_234 ();
 sg13g2_fill_2 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_280 ();
 sg13g2_fill_1 FILLER_27_314 ();
 sg13g2_decap_4 FILLER_27_329 ();
 sg13g2_fill_1 FILLER_27_351 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_49 ();
 sg13g2_fill_2 FILLER_28_60 ();
 sg13g2_fill_1 FILLER_28_62 ();
 sg13g2_fill_2 FILLER_28_81 ();
 sg13g2_fill_2 FILLER_28_108 ();
 sg13g2_fill_1 FILLER_28_110 ();
 sg13g2_decap_8 FILLER_28_117 ();
 sg13g2_fill_1 FILLER_28_124 ();
 sg13g2_decap_4 FILLER_28_151 ();
 sg13g2_decap_4 FILLER_28_163 ();
 sg13g2_fill_2 FILLER_28_167 ();
 sg13g2_decap_8 FILLER_28_173 ();
 sg13g2_decap_4 FILLER_28_180 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_decap_4 FILLER_28_194 ();
 sg13g2_fill_2 FILLER_28_198 ();
 sg13g2_decap_8 FILLER_28_208 ();
 sg13g2_decap_8 FILLER_28_215 ();
 sg13g2_fill_2 FILLER_28_222 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_fill_2 FILLER_28_249 ();
 sg13g2_fill_1 FILLER_28_290 ();
 sg13g2_decap_4 FILLER_28_296 ();
 sg13g2_fill_2 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_311 ();
 sg13g2_decap_4 FILLER_28_318 ();
 sg13g2_fill_2 FILLER_28_322 ();
 sg13g2_fill_1 FILLER_28_342 ();
 sg13g2_fill_1 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_4 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_25 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_fill_2 FILLER_29_84 ();
 sg13g2_fill_1 FILLER_29_96 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_fill_2 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_152 ();
 sg13g2_fill_2 FILLER_29_159 ();
 sg13g2_fill_1 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_166 ();
 sg13g2_fill_2 FILLER_29_173 ();
 sg13g2_decap_8 FILLER_29_207 ();
 sg13g2_fill_2 FILLER_29_214 ();
 sg13g2_fill_2 FILLER_29_266 ();
 sg13g2_fill_1 FILLER_29_280 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_fill_2 FILLER_29_302 ();
 sg13g2_fill_2 FILLER_29_329 ();
 sg13g2_fill_1 FILLER_29_331 ();
 sg13g2_fill_2 FILLER_29_372 ();
 sg13g2_fill_2 FILLER_30_46 ();
 sg13g2_fill_1 FILLER_30_48 ();
 sg13g2_fill_2 FILLER_30_53 ();
 sg13g2_fill_1 FILLER_30_78 ();
 sg13g2_fill_1 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_97 ();
 sg13g2_fill_1 FILLER_30_185 ();
 sg13g2_decap_4 FILLER_30_199 ();
 sg13g2_fill_1 FILLER_30_224 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_fill_1 FILLER_30_269 ();
 sg13g2_decap_4 FILLER_30_298 ();
 sg13g2_fill_1 FILLER_30_302 ();
 sg13g2_fill_1 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_67 ();
 sg13g2_fill_2 FILLER_31_79 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_fill_1 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_172 ();
 sg13g2_fill_1 FILLER_31_174 ();
 sg13g2_fill_2 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_209 ();
 sg13g2_decap_8 FILLER_31_220 ();
 sg13g2_decap_8 FILLER_31_227 ();
 sg13g2_decap_4 FILLER_31_234 ();
 sg13g2_fill_1 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_243 ();
 sg13g2_fill_1 FILLER_31_250 ();
 sg13g2_decap_8 FILLER_31_265 ();
 sg13g2_decap_4 FILLER_31_272 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_decap_4 FILLER_31_291 ();
 sg13g2_fill_2 FILLER_31_330 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_fill_2 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_27 ();
 sg13g2_fill_1 FILLER_32_48 ();
 sg13g2_fill_1 FILLER_32_54 ();
 sg13g2_decap_8 FILLER_32_58 ();
 sg13g2_fill_2 FILLER_32_65 ();
 sg13g2_fill_1 FILLER_32_67 ();
 sg13g2_fill_2 FILLER_32_72 ();
 sg13g2_fill_1 FILLER_32_74 ();
 sg13g2_fill_1 FILLER_32_79 ();
 sg13g2_fill_2 FILLER_32_96 ();
 sg13g2_decap_4 FILLER_32_110 ();
 sg13g2_fill_1 FILLER_32_114 ();
 sg13g2_decap_4 FILLER_32_128 ();
 sg13g2_fill_2 FILLER_32_132 ();
 sg13g2_decap_4 FILLER_32_151 ();
 sg13g2_fill_2 FILLER_32_155 ();
 sg13g2_decap_8 FILLER_32_174 ();
 sg13g2_decap_8 FILLER_32_181 ();
 sg13g2_decap_4 FILLER_32_200 ();
 sg13g2_fill_2 FILLER_32_204 ();
 sg13g2_decap_4 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_249 ();
 sg13g2_fill_2 FILLER_32_261 ();
 sg13g2_decap_4 FILLER_32_279 ();
 sg13g2_fill_2 FILLER_32_283 ();
 sg13g2_fill_1 FILLER_32_290 ();
 sg13g2_decap_4 FILLER_32_301 ();
 sg13g2_fill_1 FILLER_32_305 ();
 sg13g2_decap_8 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_345 ();
 sg13g2_fill_1 FILLER_32_358 ();
 sg13g2_fill_2 FILLER_33_73 ();
 sg13g2_fill_2 FILLER_33_83 ();
 sg13g2_fill_1 FILLER_33_85 ();
 sg13g2_decap_4 FILLER_33_104 ();
 sg13g2_decap_8 FILLER_33_129 ();
 sg13g2_fill_2 FILLER_33_136 ();
 sg13g2_fill_1 FILLER_33_138 ();
 sg13g2_fill_2 FILLER_33_157 ();
 sg13g2_fill_1 FILLER_33_159 ();
 sg13g2_fill_1 FILLER_33_172 ();
 sg13g2_decap_4 FILLER_33_185 ();
 sg13g2_fill_2 FILLER_33_189 ();
 sg13g2_decap_4 FILLER_33_212 ();
 sg13g2_fill_2 FILLER_33_216 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_233 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_fill_1 FILLER_33_245 ();
 sg13g2_fill_2 FILLER_33_268 ();
 sg13g2_fill_2 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_286 ();
 sg13g2_decap_4 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_decap_4 FILLER_33_311 ();
 sg13g2_fill_1 FILLER_33_315 ();
 sg13g2_fill_1 FILLER_33_329 ();
 sg13g2_decap_4 FILLER_33_333 ();
 sg13g2_fill_1 FILLER_33_337 ();
 sg13g2_fill_2 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_fill_2 FILLER_33_370 ();
 sg13g2_fill_2 FILLER_33_392 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_16 ();
 sg13g2_fill_1 FILLER_34_40 ();
 sg13g2_fill_2 FILLER_34_55 ();
 sg13g2_decap_8 FILLER_34_62 ();
 sg13g2_fill_2 FILLER_34_72 ();
 sg13g2_fill_1 FILLER_34_74 ();
 sg13g2_decap_8 FILLER_34_104 ();
 sg13g2_decap_4 FILLER_34_111 ();
 sg13g2_fill_1 FILLER_34_115 ();
 sg13g2_fill_2 FILLER_34_125 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_decap_8 FILLER_34_137 ();
 sg13g2_fill_1 FILLER_34_144 ();
 sg13g2_decap_4 FILLER_34_157 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_decap_4 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_decap_4 FILLER_34_210 ();
 sg13g2_fill_1 FILLER_34_222 ();
 sg13g2_decap_8 FILLER_34_239 ();
 sg13g2_decap_8 FILLER_34_254 ();
 sg13g2_fill_2 FILLER_34_261 ();
 sg13g2_decap_8 FILLER_34_281 ();
 sg13g2_fill_2 FILLER_34_308 ();
 sg13g2_fill_1 FILLER_34_310 ();
 sg13g2_decap_4 FILLER_34_335 ();
 sg13g2_fill_1 FILLER_34_339 ();
 sg13g2_decap_8 FILLER_34_351 ();
 sg13g2_decap_4 FILLER_34_358 ();
 sg13g2_fill_2 FILLER_34_373 ();
 sg13g2_decap_4 FILLER_34_391 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_fill_2 FILLER_35_48 ();
 sg13g2_fill_1 FILLER_35_50 ();
 sg13g2_fill_1 FILLER_35_64 ();
 sg13g2_fill_1 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_83 ();
 sg13g2_fill_2 FILLER_35_93 ();
 sg13g2_fill_1 FILLER_35_95 ();
 sg13g2_fill_2 FILLER_35_122 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_4 FILLER_35_171 ();
 sg13g2_fill_1 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_185 ();
 sg13g2_fill_1 FILLER_35_192 ();
 sg13g2_decap_8 FILLER_35_201 ();
 sg13g2_decap_8 FILLER_35_208 ();
 sg13g2_decap_8 FILLER_35_215 ();
 sg13g2_fill_1 FILLER_35_222 ();
 sg13g2_fill_2 FILLER_35_232 ();
 sg13g2_fill_1 FILLER_35_234 ();
 sg13g2_fill_2 FILLER_35_243 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_261 ();
 sg13g2_decap_8 FILLER_35_274 ();
 sg13g2_decap_8 FILLER_35_281 ();
 sg13g2_decap_4 FILLER_35_288 ();
 sg13g2_fill_1 FILLER_35_292 ();
 sg13g2_fill_1 FILLER_35_301 ();
 sg13g2_fill_2 FILLER_35_307 ();
 sg13g2_fill_1 FILLER_35_309 ();
 sg13g2_decap_4 FILLER_35_326 ();
 sg13g2_fill_2 FILLER_35_342 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_fill_2 FILLER_35_371 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_22 ();
 sg13g2_fill_2 FILLER_36_33 ();
 sg13g2_decap_8 FILLER_36_88 ();
 sg13g2_decap_8 FILLER_36_95 ();
 sg13g2_decap_4 FILLER_36_102 ();
 sg13g2_fill_2 FILLER_36_110 ();
 sg13g2_fill_1 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_122 ();
 sg13g2_fill_1 FILLER_36_129 ();
 sg13g2_decap_8 FILLER_36_134 ();
 sg13g2_decap_4 FILLER_36_141 ();
 sg13g2_fill_1 FILLER_36_145 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_decap_4 FILLER_36_194 ();
 sg13g2_fill_2 FILLER_36_198 ();
 sg13g2_decap_8 FILLER_36_205 ();
 sg13g2_decap_4 FILLER_36_212 ();
 sg13g2_decap_4 FILLER_36_234 ();
 sg13g2_fill_2 FILLER_36_238 ();
 sg13g2_fill_2 FILLER_36_253 ();
 sg13g2_fill_2 FILLER_36_267 ();
 sg13g2_fill_1 FILLER_36_269 ();
 sg13g2_fill_2 FILLER_36_278 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_fill_2 FILLER_36_298 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_fill_2 FILLER_36_309 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_fill_2 FILLER_36_320 ();
 sg13g2_fill_2 FILLER_36_327 ();
 sg13g2_fill_1 FILLER_36_337 ();
 sg13g2_decap_4 FILLER_36_351 ();
 sg13g2_fill_1 FILLER_36_363 ();
 sg13g2_fill_2 FILLER_36_390 ();
 sg13g2_fill_1 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_fill_1 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_39 ();
 sg13g2_decap_8 FILLER_37_46 ();
 sg13g2_fill_1 FILLER_37_53 ();
 sg13g2_fill_2 FILLER_37_92 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_fill_2 FILLER_37_121 ();
 sg13g2_decap_4 FILLER_37_130 ();
 sg13g2_fill_1 FILLER_37_168 ();
 sg13g2_fill_1 FILLER_37_219 ();
 sg13g2_fill_2 FILLER_37_233 ();
 sg13g2_fill_2 FILLER_37_247 ();
 sg13g2_fill_2 FILLER_37_257 ();
 sg13g2_decap_4 FILLER_37_272 ();
 sg13g2_decap_4 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_297 ();
 sg13g2_fill_2 FILLER_37_304 ();
 sg13g2_fill_2 FILLER_37_326 ();
 sg13g2_fill_1 FILLER_37_347 ();
 sg13g2_decap_4 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_4 FILLER_38_42 ();
 sg13g2_fill_2 FILLER_38_85 ();
 sg13g2_fill_1 FILLER_38_87 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_108 ();
 sg13g2_fill_2 FILLER_38_139 ();
 sg13g2_fill_1 FILLER_38_141 ();
 sg13g2_fill_1 FILLER_38_155 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_4 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_202 ();
 sg13g2_decap_8 FILLER_38_209 ();
 sg13g2_decap_4 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_fill_2 FILLER_38_262 ();
 sg13g2_fill_1 FILLER_38_264 ();
 sg13g2_decap_4 FILLER_38_291 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_309 ();
 sg13g2_fill_1 FILLER_38_382 ();
 assign uio_oe[0] = net119;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
endmodule

module tt_um_wokwi_group_5 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire clk_regs;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire net109;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire \proj_10.net10 ;
 wire \proj_10.net17 ;
 wire \proj_10.net18 ;
 wire \proj_10.net19 ;
 wire \proj_10.net20 ;
 wire \proj_10.net9 ;
 wire \proj_11.net3 ;
 wire \proj_11.net4 ;
 wire \proj_12.net10 ;
 wire \proj_12.net11 ;
 wire \proj_12.net12 ;
 wire \proj_12.net13 ;
 wire \proj_13.net14 ;
 wire \proj_13.net15 ;
 wire \proj_13.net16 ;
 wire \proj_13.net17 ;
 wire \proj_13.net18 ;
 wire \proj_13.net4 ;
 wire \proj_13.net5 ;
 wire \proj_13.net6 ;
 wire \proj_13.net7 ;
 wire \proj_13.net8 ;
 wire \proj_14.net11 ;
 wire \proj_14.net12 ;
 wire \proj_14.net13 ;
 wire \proj_14.net4 ;
 wire \proj_14.net5 ;
 wire \proj__0.net14 ;
 wire \proj__0.net3 ;
 wire \proj__0.net4 ;
 wire \proj__0.net5 ;
 wire \proj__0.net6 ;
 wire \proj__0.net7 ;
 wire \proj__0.net8 ;
 wire \proj__1.net10 ;
 wire \proj__1.net11 ;
 wire \proj__1.net12 ;
 wire \proj__1.net9 ;
 wire \proj__2.net12 ;
 wire \proj__2.net13 ;
 wire \proj__2.net14 ;
 wire \proj__2.net15 ;
 wire \proj__2.net16 ;
 wire \proj__2.net17 ;
 wire \proj__2.net18 ;
 wire \proj__2.net19 ;
 wire \proj__2.net2 ;
 wire \proj__2.net20 ;
 wire \proj__2.net21 ;
 wire \proj__2.net22 ;
 wire \proj__2.net23 ;
 wire \proj__2.net24 ;
 wire \proj__2.net25 ;
 wire \proj__2.net26 ;
 wire \proj__2.net27 ;
 wire \proj__2.net28 ;
 wire \proj__2.net29 ;
 wire \proj__2.net3 ;
 wire \proj__2.net30 ;
 wire \proj__2.net31 ;
 wire \proj__2.net32 ;
 wire \proj__2.net33 ;
 wire \proj__2.net34 ;
 wire \proj__2.net4 ;
 wire \proj__2.net5 ;
 wire \proj__2.net6 ;
 wire \proj__3.net9 ;
 wire \proj__4.net10 ;
 wire \proj__4.net11 ;
 wire \proj__4.net12 ;
 wire \proj__4.net9 ;
 wire \proj__5.net10 ;
 wire \proj__5.net9 ;
 wire \proj__6.net11 ;
 wire \proj__6.net12 ;
 wire \proj__6.net5 ;
 wire \proj__7.net10 ;
 wire \proj__7.net100 ;
 wire \proj__7.net101 ;
 wire \proj__7.net102 ;
 wire \proj__7.net103 ;
 wire \proj__7.net104 ;
 wire \proj__7.net105 ;
 wire \proj__7.net106 ;
 wire \proj__7.net107 ;
 wire \proj__7.net108 ;
 wire \proj__7.net109 ;
 wire \proj__7.net11 ;
 wire \proj__7.net110 ;
 wire \proj__7.net112 ;
 wire \proj__7.net113 ;
 wire \proj__7.net114 ;
 wire \proj__7.net115 ;
 wire \proj__7.net116 ;
 wire \proj__7.net117 ;
 wire \proj__7.net118 ;
 wire \proj__7.net119 ;
 wire \proj__7.net12 ;
 wire \proj__7.net120 ;
 wire \proj__7.net121 ;
 wire \proj__7.net122 ;
 wire \proj__7.net123 ;
 wire \proj__7.net124 ;
 wire \proj__7.net125 ;
 wire \proj__7.net126 ;
 wire \proj__7.net127 ;
 wire \proj__7.net128 ;
 wire \proj__7.net129 ;
 wire \proj__7.net13 ;
 wire \proj__7.net130 ;
 wire \proj__7.net131 ;
 wire \proj__7.net132 ;
 wire \proj__7.net133 ;
 wire \proj__7.net134 ;
 wire \proj__7.net135 ;
 wire \proj__7.net136 ;
 wire \proj__7.net137 ;
 wire \proj__7.net138 ;
 wire \proj__7.net139 ;
 wire \proj__7.net14 ;
 wire \proj__7.net140 ;
 wire \proj__7.net141 ;
 wire \proj__7.net142 ;
 wire \proj__7.net143 ;
 wire \proj__7.net145 ;
 wire \proj__7.net146 ;
 wire \proj__7.net147 ;
 wire \proj__7.net148 ;
 wire \proj__7.net149 ;
 wire \proj__7.net15 ;
 wire \proj__7.net150 ;
 wire \proj__7.net151 ;
 wire \proj__7.net152 ;
 wire \proj__7.net153 ;
 wire \proj__7.net154 ;
 wire \proj__7.net155 ;
 wire \proj__7.net156 ;
 wire \proj__7.net157 ;
 wire \proj__7.net158 ;
 wire \proj__7.net159 ;
 wire \proj__7.net160 ;
 wire \proj__7.net161 ;
 wire \proj__7.net162 ;
 wire \proj__7.net163 ;
 wire \proj__7.net164 ;
 wire \proj__7.net165 ;
 wire \proj__7.net166 ;
 wire \proj__7.net167 ;
 wire \proj__7.net168 ;
 wire \proj__7.net170 ;
 wire \proj__7.net171 ;
 wire \proj__7.net172 ;
 wire \proj__7.net173 ;
 wire \proj__7.net174 ;
 wire \proj__7.net21 ;
 wire \proj__7.net22 ;
 wire \proj__7.net23 ;
 wire \proj__7.net24 ;
 wire \proj__7.net25 ;
 wire \proj__7.net26 ;
 wire \proj__7.net27 ;
 wire \proj__7.net28 ;
 wire \proj__7.net29 ;
 wire \proj__7.net30 ;
 wire \proj__7.net31 ;
 wire \proj__7.net32 ;
 wire \proj__7.net33 ;
 wire \proj__7.net34 ;
 wire \proj__7.net35 ;
 wire \proj__7.net36 ;
 wire \proj__7.net37 ;
 wire \proj__7.net38 ;
 wire \proj__7.net39 ;
 wire \proj__7.net40 ;
 wire \proj__7.net42 ;
 wire \proj__7.net43 ;
 wire \proj__7.net44 ;
 wire \proj__7.net45 ;
 wire \proj__7.net46 ;
 wire \proj__7.net47 ;
 wire \proj__7.net48 ;
 wire \proj__7.net49 ;
 wire \proj__7.net50 ;
 wire \proj__7.net51 ;
 wire \proj__7.net52 ;
 wire \proj__7.net53 ;
 wire \proj__7.net54 ;
 wire \proj__7.net55 ;
 wire \proj__7.net56 ;
 wire \proj__7.net58 ;
 wire \proj__7.net59 ;
 wire \proj__7.net60 ;
 wire \proj__7.net61 ;
 wire \proj__7.net62 ;
 wire \proj__7.net63 ;
 wire \proj__7.net64 ;
 wire \proj__7.net65 ;
 wire \proj__7.net66 ;
 wire \proj__7.net67 ;
 wire \proj__7.net68 ;
 wire \proj__7.net69 ;
 wire \proj__7.net70 ;
 wire \proj__7.net71 ;
 wire \proj__7.net72 ;
 wire \proj__7.net73 ;
 wire \proj__7.net74 ;
 wire \proj__7.net75 ;
 wire \proj__7.net76 ;
 wire \proj__7.net77 ;
 wire \proj__7.net78 ;
 wire \proj__7.net79 ;
 wire \proj__7.net80 ;
 wire \proj__7.net81 ;
 wire \proj__7.net82 ;
 wire \proj__7.net83 ;
 wire \proj__7.net84 ;
 wire \proj__7.net85 ;
 wire \proj__7.net86 ;
 wire \proj__7.net87 ;
 wire \proj__7.net88 ;
 wire \proj__7.net89 ;
 wire \proj__7.net9 ;
 wire \proj__7.net90 ;
 wire \proj__7.net91 ;
 wire \proj__7.net93 ;
 wire \proj__7.net94 ;
 wire \proj__7.net95 ;
 wire \proj__7.net96 ;
 wire \proj__7.net97 ;
 wire \proj__7.net98 ;
 wire \proj__7.net99 ;
 wire \proj__9.net10 ;
 wire \proj__9.net11 ;
 wire \proj__9.net12 ;
 wire \proj__9.net13 ;
 wire \proj__9.net14 ;
 wire \proj__9.net20 ;
 wire \proj__9.net21 ;
 wire \proj__9.net22 ;
 wire \proj__9.net23 ;
 wire \proj__9.net24 ;
 wire \proj__9.net25 ;
 wire \proj__9.net26 ;
 wire \proj__9.net27 ;
 wire \proj__9.net7 ;
 wire \proj__9.net8 ;
 wire \proj__9.net9 ;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire \proj__0.flop1/_0_ ;
 wire \proj__0.flop1/_1_ ;
 wire net97;
 wire net98;
 wire \proj__0.flop1/notq ;
 wire \proj__0.flop2/_0_ ;
 wire \proj__0.flop2/_1_ ;
 wire net99;
 wire net100;
 wire \proj__0.flop2/notq ;
 wire \proj__0.flop3/_0_ ;
 wire \proj__0.flop3/_1_ ;
 wire net101;
 wire net102;
 wire \proj__0.flop3/notq ;
 wire \proj__0.flop4/_0_ ;
 wire \proj__0.flop4/_1_ ;
 wire net103;
 wire net104;
 wire \proj__0.flop4/notq ;
 wire \proj__0.flop5/_0_ ;
 wire \proj__0.flop5/_1_ ;
 wire net105;
 wire net106;
 wire \proj__0.flop5/notq ;
 wire \proj__0.flop6/_0_ ;
 wire \proj__0.flop6/_1_ ;
 wire net107;
 wire net108;
 wire \proj__0.flop6/notq ;
 wire net110;
 wire net111;
 wire net112;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_1_0__leaf_clk_regs;
 wire clknet_1_1__leaf_clk_regs;
 wire clknet_0__005_;
 wire clknet_1_0__leaf__005_;
 wire clknet_1_1__leaf__005_;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;

 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_nor2_2 _142_ (.A(net9),
    .B(net10),
    .Y(_064_));
 sg13g2_nor2_2 _143_ (.A(net7),
    .B(net8),
    .Y(_065_));
 sg13g2_and2_1 _144_ (.A(_064_),
    .B(_065_),
    .X(_066_));
 sg13g2_nand2_1 _145_ (.Y(_067_),
    .A(_064_),
    .B(_065_));
 sg13g2_nor2b_2 _146_ (.A(net7),
    .B_N(net8),
    .Y(_068_));
 sg13g2_and2_2 _147_ (.A(_064_),
    .B(_068_),
    .X(_069_));
 sg13g2_a21oi_2 _148_ (.B1(net35),
    .Y(_070_),
    .A2(_069_),
    .A1(\proj__2.net2 ));
 sg13g2_nor2b_2 _149_ (.A(net10),
    .B_N(net9),
    .Y(_071_));
 sg13g2_and2_1 _150_ (.A(_068_),
    .B(_071_),
    .X(_072_));
 sg13g2_and2_2 _151_ (.A(net7),
    .B(net8),
    .X(_073_));
 sg13g2_and2_2 _152_ (.A(_071_),
    .B(_073_),
    .X(_074_));
 sg13g2_a22oi_1 _153_ (.Y(_075_),
    .B1(_074_),
    .B2(\proj__7.net9 ),
    .A2(_072_),
    .A1(\proj__6.net5 ));
 sg13g2_nor2b_2 _154_ (.A(net8),
    .B_N(net7),
    .Y(_076_));
 sg13g2_nand3_1 _155_ (.B(_071_),
    .C(_076_),
    .A(\proj__5.net9 ),
    .Y(_077_));
 sg13g2_nor2b_2 _156_ (.A(net9),
    .B_N(net10),
    .Y(_078_));
 sg13g2_nand3_1 _157_ (.B(_073_),
    .C(_078_),
    .A(\proj_11.net3 ),
    .Y(_079_));
 sg13g2_and4_1 _158_ (.A(_070_),
    .B(_075_),
    .C(_077_),
    .D(_079_),
    .X(_080_));
 sg13g2_and2_1 _159_ (.A(_064_),
    .B(_076_),
    .X(_081_));
 sg13g2_and2_1 _160_ (.A(_065_),
    .B(_071_),
    .X(_000_));
 sg13g2_a22oi_1 _161_ (.Y(_001_),
    .B1(_000_),
    .B2(\proj__4.net9 ),
    .A2(_081_),
    .A1(\proj__1.net9 ));
 sg13g2_and2_1 _162_ (.A(_064_),
    .B(_073_),
    .X(_002_));
 sg13g2_nand3_1 _163_ (.B(_064_),
    .C(_073_),
    .A(net43),
    .Y(_003_));
 sg13g2_and2_2 _164_ (.A(net9),
    .B(net10),
    .X(_004_));
 sg13g2_nand3_1 _165_ (.B(_065_),
    .C(_004_),
    .A(\proj_12.net10 ),
    .Y(_005_));
 sg13g2_and2_1 _166_ (.A(_003_),
    .B(clknet_1_0__leaf__005_),
    .X(_006_));
 sg13g2_and2_1 _167_ (.A(_068_),
    .B(_078_),
    .X(_007_));
 sg13g2_and2_2 _168_ (.A(_076_),
    .B(_078_),
    .X(_008_));
 sg13g2_a22oi_1 _169_ (.Y(_009_),
    .B1(_008_),
    .B2(\proj__9.net7 ),
    .A2(_007_),
    .A1(\proj_10.net9 ));
 sg13g2_and2_2 _170_ (.A(_076_),
    .B(_004_),
    .X(_010_));
 sg13g2_nand2_1 _171_ (.Y(_011_),
    .A(\proj_13.net4 ),
    .B(_010_));
 sg13g2_and2_1 _172_ (.A(_068_),
    .B(_004_),
    .X(_012_));
 sg13g2_a22oi_1 _173_ (.Y(_013_),
    .B1(_012_),
    .B2(\proj_14.net4 ),
    .A2(_010_),
    .A1(\proj_13.net4 ));
 sg13g2_and4_1 _174_ (.A(_001_),
    .B(_006_),
    .C(_009_),
    .D(_013_),
    .X(_014_));
 sg13g2_a22oi_1 _175_ (.Y(uo_out[0]),
    .B1(_080_),
    .B2(_014_),
    .A2(_066_),
    .A1(_057_));
 sg13g2_nand3_1 _176_ (.B(_071_),
    .C(_076_),
    .A(\proj__5.net10 ),
    .Y(_015_));
 sg13g2_nand3_1 _177_ (.B(_073_),
    .C(_078_),
    .A(\proj_11.net4 ),
    .Y(_016_));
 sg13g2_nand2_1 _178_ (.Y(_017_),
    .A(\proj__7.net10 ),
    .B(_074_));
 sg13g2_nand3_1 _179_ (.B(_065_),
    .C(_004_),
    .A(\proj_12.net11 ),
    .Y(_018_));
 sg13g2_and4_1 _180_ (.A(_015_),
    .B(_016_),
    .C(_017_),
    .D(_018_),
    .X(_019_));
 sg13g2_a22oi_1 _181_ (.Y(_020_),
    .B1(_000_),
    .B2(\proj__4.net10 ),
    .A2(_081_),
    .A1(\proj__1.net10 ));
 sg13g2_a22oi_1 _182_ (.Y(_021_),
    .B1(_012_),
    .B2(\proj_14.net5 ),
    .A2(_008_),
    .A1(\proj__9.net8 ));
 sg13g2_a22oi_1 _183_ (.Y(_022_),
    .B1(_010_),
    .B2(\proj_13.net5 ),
    .A2(_002_),
    .A1(\proj__3.net9 ));
 sg13g2_and4_1 _184_ (.A(_070_),
    .B(_020_),
    .C(_021_),
    .D(_022_),
    .X(_023_));
 sg13g2_a22oi_1 _185_ (.Y(uo_out[1]),
    .B1(_019_),
    .B2(_023_),
    .A2(net35),
    .A1(_058_));
 sg13g2_nand2_1 _186_ (.Y(_024_),
    .A(\proj__4.net11 ),
    .B(_000_));
 sg13g2_a22oi_1 _187_ (.Y(_025_),
    .B1(_076_),
    .B2(_071_),
    .A2(_073_),
    .A1(_064_));
 sg13g2_nand2b_1 _188_ (.Y(_026_),
    .B(net37),
    .A_N(_025_));
 sg13g2_a22oi_1 _189_ (.Y(_027_),
    .B1(_010_),
    .B2(\proj_13.net6 ),
    .A2(_074_),
    .A1(\proj__7.net11 ));
 sg13g2_and3_1 _190_ (.X(_028_),
    .A(\proj_12.net12 ),
    .B(_065_),
    .C(_004_));
 sg13g2_a21oi_1 _191_ (.A1(\proj__9.net9 ),
    .A2(_008_),
    .Y(_029_),
    .B1(net35));
 sg13g2_a221oi_1 _192_ (.B2(\proj__1.net11 ),
    .C1(_028_),
    .B1(_081_),
    .A1(\proj__2.net3 ),
    .Y(_030_),
    .A2(_069_));
 sg13g2_and4_1 _193_ (.A(_024_),
    .B(_026_),
    .C(_027_),
    .D(_030_),
    .X(_031_));
 sg13g2_a22oi_1 _194_ (.Y(uo_out[2]),
    .B1(_029_),
    .B2(_031_),
    .A2(net35),
    .A1(_059_));
 sg13g2_nand3_1 _195_ (.B(_065_),
    .C(_004_),
    .A(\proj_12.net13 ),
    .Y(_032_));
 sg13g2_nand2_1 _196_ (.Y(_033_),
    .A(\proj__9.net10 ),
    .B(_008_));
 sg13g2_a22oi_1 _197_ (.Y(_034_),
    .B1(_074_),
    .B2(\proj__7.net12 ),
    .A2(_069_),
    .A1(\proj__2.net4 ));
 sg13g2_and3_1 _198_ (.X(_035_),
    .A(_032_),
    .B(_033_),
    .C(_034_));
 sg13g2_nand2b_1 _199_ (.Y(_036_),
    .B(net36),
    .A_N(_025_));
 sg13g2_a22oi_1 _200_ (.Y(_037_),
    .B1(_000_),
    .B2(\proj__4.net12 ),
    .A2(_081_),
    .A1(\proj__1.net12 ));
 sg13g2_and4_1 _201_ (.A(_067_),
    .B(_011_),
    .C(_036_),
    .D(_037_),
    .X(_038_));
 sg13g2_a22oi_1 _202_ (.Y(uo_out[3]),
    .B1(_035_),
    .B2(_038_),
    .A2(net35),
    .A1(_060_));
 sg13g2_a22oi_1 _203_ (.Y(_039_),
    .B1(_071_),
    .B2(_056_),
    .A2(_064_),
    .A1(net7));
 sg13g2_nand2b_1 _204_ (.Y(_040_),
    .B(net3),
    .A_N(_039_));
 sg13g2_a22oi_1 _205_ (.Y(_041_),
    .B1(_008_),
    .B2(\proj__9.net11 ),
    .A2(_069_),
    .A1(\proj__2.net5 ));
 sg13g2_a22oi_1 _206_ (.Y(_042_),
    .B1(_010_),
    .B2(\proj_13.net7 ),
    .A2(_074_),
    .A1(\proj__7.net13 ));
 sg13g2_and4_1 _207_ (.A(_067_),
    .B(_018_),
    .C(_041_),
    .D(_042_),
    .X(_043_));
 sg13g2_a22oi_1 _208_ (.Y(uo_out[4]),
    .B1(_040_),
    .B2(_043_),
    .A2(net35),
    .A1(_061_));
 sg13g2_nand2b_1 _209_ (.Y(_044_),
    .B(net4),
    .A_N(_039_));
 sg13g2_nand2_1 _210_ (.Y(_045_),
    .A(\proj__7.net14 ),
    .B(_074_));
 sg13g2_a22oi_1 _211_ (.Y(_046_),
    .B1(_010_),
    .B2(\proj_13.net8 ),
    .A2(_008_),
    .A1(\proj__9.net12 ));
 sg13g2_and4_1 _212_ (.A(_070_),
    .B(_032_),
    .C(_045_),
    .D(_046_),
    .X(_047_));
 sg13g2_a22oi_1 _213_ (.Y(uo_out[5]),
    .B1(_044_),
    .B2(_047_),
    .A2(net35),
    .A1(_062_));
 sg13g2_nand2b_1 _214_ (.Y(_048_),
    .B(net5),
    .A_N(_039_));
 sg13g2_a22oi_1 _215_ (.Y(_049_),
    .B1(_008_),
    .B2(\proj__9.net13 ),
    .A2(_069_),
    .A1(\proj__2.net6 ));
 sg13g2_a22oi_1 _216_ (.Y(_050_),
    .B1(_010_),
    .B2(net43),
    .A2(_074_),
    .A1(\proj__7.net15 ));
 sg13g2_nand4_1 _217_ (.B(_048_),
    .C(_049_),
    .A(clknet_1_1__leaf__005_),
    .Y(uo_out[6]),
    .D(_050_));
 sg13g2_a22oi_1 _218_ (.Y(_051_),
    .B1(_004_),
    .B2(_065_),
    .A2(_073_),
    .A1(_071_));
 sg13g2_nand2_1 _219_ (.Y(_052_),
    .A(_039_),
    .B(_051_));
 sg13g2_nand3_1 _220_ (.B(_068_),
    .C(_078_),
    .A(\proj_10.net10 ),
    .Y(_053_));
 sg13g2_nand2_1 _221_ (.Y(_054_),
    .A(_067_),
    .B(_053_));
 sg13g2_a221oi_1 _222_ (.B2(net6),
    .C1(_054_),
    .B1(_052_),
    .A1(\proj__9.net14 ),
    .Y(_055_),
    .A2(_008_));
 sg13g2_a21oi_1 _223_ (.A1(net112),
    .A2(net35),
    .Y(uo_out[7]),
    .B1(_055_));
 sg13g2_inv_1 _224_ (.Y(_056_),
    .A(net8));
 sg13g2_inv_1 _225_ (.Y(_057_),
    .A(\proj__0.net3 ));
 sg13g2_inv_1 _226_ (.Y(_058_),
    .A(\proj__0.net4 ));
 sg13g2_inv_1 _227_ (.Y(_059_),
    .A(\proj__0.net5 ));
 sg13g2_inv_1 _228_ (.Y(_060_),
    .A(\proj__0.net6 ));
 sg13g2_inv_1 _229_ (.Y(_061_),
    .A(\proj__0.net7 ));
 sg13g2_inv_1 _230_ (.Y(_062_),
    .A(\proj__0.net8 ));
 sg13g2_tiehi \proj__2.flop1/_1__98  (.L_HI(net109));
 sg13g2_tielo \proj__0.flop2/_4__12  (.L_LO(net12));
 sg13g2_tielo \proj__0.flop3/_4__13  (.L_LO(net13));
 sg13g2_tielo \proj__0.flop4/_5__14  (.L_LO(net14));
 sg13g2_tielo \proj__0.flop5/_4__15  (.L_LO(net15));
 sg13g2_tielo \proj__0.flop6/_4__16  (.L_LO(net16));
 sg13g2_tielo \proj__7.or10/_0__17  (.L_LO(net17));
 sg13g2_tielo \proj__7.or11/_0__18  (.L_LO(net18));
 sg13g2_tielo \proj__7.or12/_0__19  (.L_LO(net19));
 sg13g2_tielo \proj__7.or13/_0__20  (.L_LO(net20));
 sg13g2_tielo \proj__7.or16/_0__21  (.L_LO(net21));
 sg13g2_tielo \proj__7.or17/_0__22  (.L_LO(net22));
 sg13g2_tielo \proj__7.or17/_0__23  (.L_LO(net23));
 sg13g2_tielo \proj__7.or18/_0__24  (.L_LO(net24));
 sg13g2_tielo \proj__7.or19/_0__25  (.L_LO(net25));
 sg13g2_tielo \proj__7.or2/_0__26  (.L_LO(net26));
 sg13g2_tielo \proj__7.or20/_0__27  (.L_LO(net27));
 sg13g2_tielo \proj__7.or21/_0__28  (.L_LO(net28));
 sg13g2_tielo \proj__7.or22/_0__29  (.L_LO(net29));
 sg13g2_tielo \proj__7.or23/_0__30  (.L_LO(net30));
 sg13g2_tielo \proj__7.or24/_0__31  (.L_LO(net31));
 sg13g2_tielo \proj__7.or25/_0__32  (.L_LO(net32));
 sg13g2_tielo \proj__7.or26/_0__33  (.L_LO(net33));
 sg13g2_tielo \proj__7.or27/_0__34  (.L_LO(net34));
 sg13g2_tielo \proj__7.or28/_0__35  (.L_LO(net46));
 sg13g2_tielo \proj__7.or29/_0__36  (.L_LO(net47));
 sg13g2_tielo \proj__7.or3/_0__37  (.L_LO(net48));
 sg13g2_tielo \proj__7.or3/_0__38  (.L_LO(net49));
 sg13g2_tielo \proj__7.or30/_0__39  (.L_LO(net50));
 sg13g2_tielo \proj__7.or32/_0__40  (.L_LO(net51));
 sg13g2_tielo \proj__7.or33/_0__41  (.L_LO(net52));
 sg13g2_tielo \proj__7.or34/_0__42  (.L_LO(net53));
 sg13g2_tielo \proj__7.or35/_0__43  (.L_LO(net54));
 sg13g2_tielo \proj__7.or36/_0__44  (.L_LO(net55));
 sg13g2_tielo \proj__7.or37/_0__45  (.L_LO(net56));
 sg13g2_tielo \proj__7.or39/_0__46  (.L_LO(net57));
 sg13g2_tielo \proj__7.or4/_0__47  (.L_LO(net58));
 sg13g2_tielo \proj__7.or40/_0__48  (.L_LO(net59));
 sg13g2_tielo \proj__7.or41/_0__49  (.L_LO(net60));
 sg13g2_tielo \proj__7.or42/_0__50  (.L_LO(net61));
 sg13g2_tielo \proj__7.or43/_0__51  (.L_LO(net62));
 sg13g2_tielo \proj__7.or44/_0__52  (.L_LO(net63));
 sg13g2_tielo \proj__7.or45/_0__53  (.L_LO(net64));
 sg13g2_tielo \proj__7.or46/_0__54  (.L_LO(net65));
 sg13g2_tielo \proj__7.or47/_0__55  (.L_LO(net66));
 sg13g2_tielo \proj__7.or48/_0__56  (.L_LO(net67));
 sg13g2_tielo \proj__7.or49/_0__57  (.L_LO(net68));
 sg13g2_tielo \proj__7.or5/_0__58  (.L_LO(net69));
 sg13g2_tielo \proj__7.or50/_0__59  (.L_LO(net70));
 sg13g2_tielo \proj__7.or51/_0__60  (.L_LO(net71));
 sg13g2_tielo \proj__7.or52/_0__61  (.L_LO(net72));
 sg13g2_tielo \proj__7.or6/_0__62  (.L_LO(net73));
 sg13g2_tielo \proj__7.or61/_0__63  (.L_LO(net74));
 sg13g2_tielo \proj__7.or79/_0__64  (.L_LO(net75));
 sg13g2_tielo \proj__7.or8/_0__65  (.L_LO(net76));
 sg13g2_tielo \proj__7.or8/_0__66  (.L_LO(net77));
 sg13g2_tielo \proj__7.or87/_0__67  (.L_LO(net78));
 sg13g2_tielo \proj__7.or9/_0__68  (.L_LO(net79));
 sg13g2_tielo tt_um_wokwi_group_5_69 (.L_LO(net80));
 sg13g2_tielo tt_um_wokwi_group_5_70 (.L_LO(net81));
 sg13g2_tielo tt_um_wokwi_group_5_71 (.L_LO(net82));
 sg13g2_tielo tt_um_wokwi_group_5_72 (.L_LO(net83));
 sg13g2_tielo tt_um_wokwi_group_5_73 (.L_LO(net84));
 sg13g2_tielo tt_um_wokwi_group_5_74 (.L_LO(net85));
 sg13g2_tielo tt_um_wokwi_group_5_75 (.L_LO(net86));
 sg13g2_tielo tt_um_wokwi_group_5_76 (.L_LO(net87));
 sg13g2_tielo tt_um_wokwi_group_5_77 (.L_LO(net88));
 sg13g2_tielo tt_um_wokwi_group_5_78 (.L_LO(net89));
 sg13g2_tielo tt_um_wokwi_group_5_79 (.L_LO(net90));
 sg13g2_tielo tt_um_wokwi_group_5_80 (.L_LO(net91));
 sg13g2_tielo tt_um_wokwi_group_5_81 (.L_LO(net92));
 sg13g2_tielo tt_um_wokwi_group_5_82 (.L_LO(net93));
 sg13g2_tielo tt_um_wokwi_group_5_83 (.L_LO(net94));
 sg13g2_tielo tt_um_wokwi_group_5_84 (.L_LO(net95));
 sg13g2_tielo \proj__0.flop1/dffsr_85  (.L_LO(net96));
 sg13g2_or2_1 \proj_10.or2/_0_  (.X(\proj_10.net10 ),
    .B(\proj_10.net17 ),
    .A(\proj_10.net18 ));
 sg13g2_or2_1 \proj_10.or4/_0_  (.X(\proj_10.net19 ),
    .B(net3),
    .A(net5));
 sg13g2_or2_1 \proj_10.or5/_0_  (.X(\proj_10.net20 ),
    .B(net43),
    .A(net37));
 sg13g2_or2_1 \proj_10.or6/_0_  (.X(\proj_10.net9 ),
    .B(\proj_10.net20 ),
    .A(\proj_10.net19 ));
 sg13g2_or2_1 \proj_10.or7/_0_  (.X(\proj_10.net18 ),
    .B(net4),
    .A(net6));
 sg13g2_or2_1 \proj_10.or8/_0_  (.X(\proj_10.net17 ),
    .B(net41),
    .A(net36));
 sg13g2_and2_1 \proj_11.and1/_0_  (.A(net44),
    .B(net41),
    .X(\proj_11.net4 ));
 sg13g2_xor2_1 \proj_11.xor1/_0_  (.B(net44),
    .A(net40),
    .X(\proj_11.net3 ));
 sg13g2_and2_1 \proj_12.and1/_0_  (.A(net42),
    .B(clknet_1_0__leaf_clk),
    .X(\proj_12.net10 ));
 sg13g2_and2_1 \proj_12.and2/_0_  (.A(net36),
    .B(net37),
    .X(\proj_12.net11 ));
 sg13g2_mux2_1 \proj_12.mux1/_0_  (.A0(net4),
    .A1(net5),
    .S(net6),
    .X(\proj_12.net13 ));
 sg13g2_or2_1 \proj_12.or1/_0_  (.X(\proj_12.net12 ),
    .B(net1),
    .A(net41));
 sg13g2_and2_1 \proj_13.and1/_0_  (.A(\proj_13.net14 ),
    .B(\proj_13.net17 ),
    .X(\proj_13.net8 ));
 sg13g2_inv_1 \proj_13.not1/_0_  (.Y(\proj_13.net14 ),
    .A(net39));
 sg13g2_inv_1 \proj_13.not2/_0_  (.Y(\proj_13.net15 ),
    .A(net39));
 sg13g2_inv_1 \proj_13.not3/_0_  (.Y(\proj_13.net16 ),
    .A(net43));
 sg13g2_inv_1 \proj_13.not4/_0_  (.Y(\proj_13.net7 ),
    .A(net39));
 sg13g2_inv_1 \proj_13.not5/_0_  (.Y(\proj_13.net17 ),
    .A(net42));
 sg13g2_inv_1 \proj_13.not6/_0_  (.Y(\proj_13.net18 ),
    .A(net6));
 sg13g2_or2_1 \proj_13.or1/_0_  (.X(\proj_13.net4 ),
    .B(net42),
    .A(\proj_13.net15 ));
 sg13g2_or2_1 \proj_13.or2/_0_  (.X(\proj_13.net6 ),
    .B(\proj_13.net16 ),
    .A(net39));
 sg13g2_or2_1 \proj_13.or3/_0_  (.X(\proj_13.net5 ),
    .B(\proj_13.net18 ),
    .A(net6));
 sg13g2_and2_1 \proj_14.and1/_0_  (.A(net37),
    .B(\proj_14.net11 ),
    .X(\proj_14.net12 ));
 sg13g2_and2_1 \proj_14.and2/_0_  (.A(net42),
    .B(net39),
    .X(\proj_14.net13 ));
 sg13g2_or2_1 \proj_14.or1/_0_  (.X(\proj_14.net5 ),
    .B(\proj_14.net12 ),
    .A(\proj_14.net13 ));
 sg13g2_xor2_1 \proj_14.xor1/_0_  (.B(net42),
    .A(net39),
    .X(\proj_14.net11 ));
 sg13g2_xor2_1 \proj_14.xor2/_0_  (.B(\proj_14.net11 ),
    .A(net37),
    .X(\proj_14.net4 ));
 sg13g2_inv_1 \proj__0.flop1/_4_  (.Y(\proj__0.flop1/_1_ ),
    .A(net11));
 sg13g2_inv_1 \proj__0.flop1/_5_  (.Y(\proj__0.flop1/_0_ ),
    .A(\proj__0.net14 ));
 sg13g2_tielo \proj__0.flop1/dffsr_86  (.L_LO(net97));
 sg13g2_tielo \proj__0.flop2/dffsr_87  (.L_LO(net98));
 sg13g2_sdfbbp_1 \proj__0.flop1/dffsr  (.Q(\proj__0.net7 ),
    .Q_N(\proj__0.flop1/notq ),
    .RESET_B(\proj__0.flop1/_0_ ),
    .SET_B(\proj__0.flop1/_1_ ),
    .D(net118),
    .SCE(net97),
    .SCD(net96),
    .CLK(clknet_1_0__leaf_clk_regs));
 sg13g2_inv_1 \proj__0.flop2/_4_  (.Y(\proj__0.flop2/_1_ ),
    .A(net12));
 sg13g2_inv_1 \proj__0.flop2/_5_  (.Y(\proj__0.flop2/_0_ ),
    .A(\proj__0.net14 ));
 sg13g2_tielo \proj__0.flop2/dffsr_88  (.L_LO(net99));
 sg13g2_tielo \proj__0.flop3/dffsr_89  (.L_LO(net100));
 sg13g2_sdfbbp_1 \proj__0.flop2/dffsr  (.Q(\proj__0.net8 ),
    .Q_N(\proj__0.flop2/notq ),
    .RESET_B(\proj__0.flop2/_0_ ),
    .SET_B(\proj__0.flop2/_1_ ),
    .D(net116),
    .SCE(net99),
    .SCD(net98),
    .CLK(clknet_1_0__leaf_clk_regs));
 sg13g2_inv_1 \proj__0.flop3/_4_  (.Y(\proj__0.flop3/_1_ ),
    .A(net13));
 sg13g2_inv_1 \proj__0.flop3/_5_  (.Y(\proj__0.flop3/_0_ ),
    .A(\proj__0.net14 ));
 sg13g2_tielo \proj__0.flop3/dffsr_90  (.L_LO(net101));
 sg13g2_tielo \proj__0.flop4/dffsr_91  (.L_LO(net102));
 sg13g2_sdfbbp_1 \proj__0.flop3/dffsr  (.Q(\proj__0.net3 ),
    .Q_N(\proj__0.flop3/notq ),
    .RESET_B(\proj__0.flop3/_0_ ),
    .SET_B(\proj__0.flop3/_1_ ),
    .D(net114),
    .SCE(net101),
    .SCD(net100),
    .CLK(clknet_1_0__leaf_clk_regs));
 sg13g2_inv_1 \proj__0.flop4/_4_  (.Y(\proj__0.flop4/_1_ ),
    .A(\proj__0.net14 ));
 sg13g2_inv_1 \proj__0.flop4/_5_  (.Y(\proj__0.flop4/_0_ ),
    .A(net14));
 sg13g2_tielo \proj__0.flop4/dffsr_92  (.L_LO(net103));
 sg13g2_tielo \proj__0.flop5/dffsr_93  (.L_LO(net104));
 sg13g2_sdfbbp_1 \proj__0.flop4/dffsr  (.Q(\proj__0.net6 ),
    .Q_N(\proj__0.flop4/notq ),
    .RESET_B(\proj__0.flop4/_0_ ),
    .SET_B(\proj__0.flop4/_1_ ),
    .D(net115),
    .SCE(net103),
    .SCD(net102),
    .CLK(clknet_1_1__leaf_clk_regs));
 sg13g2_inv_1 \proj__0.flop5/_4_  (.Y(\proj__0.flop5/_1_ ),
    .A(net15));
 sg13g2_inv_1 \proj__0.flop5/_5_  (.Y(\proj__0.flop5/_0_ ),
    .A(\proj__0.net14 ));
 sg13g2_tielo \proj__0.flop5/dffsr_94  (.L_LO(net105));
 sg13g2_tielo \proj__0.flop6/dffsr_95  (.L_LO(net106));
 sg13g2_sdfbbp_1 \proj__0.flop5/dffsr  (.Q(\proj__0.net4 ),
    .Q_N(\proj__0.flop5/notq ),
    .RESET_B(\proj__0.flop5/_0_ ),
    .SET_B(\proj__0.flop5/_1_ ),
    .D(net117),
    .SCE(net105),
    .SCD(net104),
    .CLK(clknet_1_0__leaf_clk_regs));
 sg13g2_inv_1 \proj__0.flop6/_4_  (.Y(\proj__0.flop6/_1_ ),
    .A(net16));
 sg13g2_inv_1 \proj__0.flop6/_5_  (.Y(\proj__0.flop6/_0_ ),
    .A(\proj__0.net14 ));
 sg13g2_tielo \proj__0.flop6/dffsr_96  (.L_LO(net107));
 sg13g2_tiehi \proj__7.and22/_0__97  (.L_HI(net108));
 sg13g2_sdfbbp_1 \proj__0.flop6/dffsr  (.Q(\proj__0.net5 ),
    .Q_N(\proj__0.flop6/notq ),
    .RESET_B(\proj__0.flop6/_0_ ),
    .SET_B(\proj__0.flop6/_1_ ),
    .D(net119),
    .SCE(net107),
    .SCD(net106),
    .CLK(clknet_1_1__leaf_clk_regs));
 sg13g2_inv_2 \proj__0.not4/_0_  (.Y(\proj__0.net14 ),
    .A(net1));
 sg13g2_inv_1 \proj__1.not1/_0_  (.Y(\proj__1.net9 ),
    .A(net43));
 sg13g2_inv_1 \proj__1.not2/_0_  (.Y(\proj__1.net10 ),
    .A(net39));
 sg13g2_inv_1 \proj__1.not3/_0_  (.Y(\proj__1.net11 ),
    .A(net37));
 sg13g2_inv_1 \proj__1.not4/_0_  (.Y(\proj__1.net12 ),
    .A(net36));
 sg13g2_and2_1 \proj__2.and1/_0_  (.A(\proj__2.net18 ),
    .B(\proj__2.net19 ),
    .X(\proj__2.net2 ));
 sg13g2_and2_1 \proj__2.and2/_0_  (.A(\proj__2.net20 ),
    .B(\proj__2.net21 ),
    .X(\proj__2.net22 ));
 sg13g2_and2_1 \proj__2.and3/_0_  (.A(\proj__2.net15 ),
    .B(\proj__2.net22 ),
    .X(\proj__2.net23 ));
 sg13g2_and2_1 \proj__2.and4/_0_  (.A(\proj__2.net13 ),
    .B(\proj__2.net15 ),
    .X(\proj__2.net25 ));
 sg13g2_and2_1 \proj__2.and5/_0_  (.A(\proj__2.net25 ),
    .B(\proj__2.net24 ),
    .X(\proj__2.net4 ));
 sg13g2_and2_1 \proj__2.and6/_0_  (.A(\proj__2.net26 ),
    .B(\proj__2.net27 ),
    .X(\proj__2.net28 ));
 sg13g2_and2_1 \proj__2.and7/_0_  (.A(\proj__2.net28 ),
    .B(\proj__2.net17 ),
    .X(\proj__2.net29 ));
 sg13g2_dfrbp_1 \proj__2.flop1/_1_  (.CLK(clknet_1_1__leaf_clk_regs),
    .RESET_B(net109),
    .D(net113),
    .Q_N(\proj__2.net12 ),
    .Q(\proj__2.net13 ));
 sg13g2_tiehi \proj__2.flop2/_1__99  (.L_HI(net110));
 sg13g2_dfrbp_1 \proj__2.flop2/_1_  (.CLK(\proj__2.net12 ),
    .RESET_B(net110),
    .D(\proj__2.net14 ),
    .Q_N(\proj__2.net14 ),
    .Q(\proj__2.net15 ));
 sg13g2_tiehi \proj__2.flop3/_1__100  (.L_HI(net111));
 sg13g2_dfrbp_1 \proj__2.flop3/_1_  (.CLK(\proj__2.net14 ),
    .RESET_B(net111),
    .D(\proj__2.net16 ),
    .Q_N(\proj__2.net16 ),
    .Q(\proj__2.net17 ));
 sg13g2_inv_1 _141__1 (.Y(net112),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 \proj__2.not1/_0_  (.Y(\proj__2.net18 ),
    .A(\proj__2.net15 ));
 sg13g2_inv_1 \proj__2.not2/_0_  (.Y(\proj__2.net19 ),
    .A(\proj__2.net17 ));
 sg13g2_inv_1 \proj__2.not3/_0_  (.Y(\proj__2.net20 ),
    .A(\proj__2.net13 ));
 sg13g2_inv_1 \proj__2.not4/_0_  (.Y(\proj__2.net21 ),
    .A(\proj__2.net17 ));
 sg13g2_inv_1 \proj__2.not5/_0_  (.Y(\proj__2.net24 ),
    .A(\proj__2.net17 ));
 sg13g2_inv_1 \proj__2.not6/_0_  (.Y(\proj__2.net26 ),
    .A(\proj__2.net13 ));
 sg13g2_inv_1 \proj__2.not7/_0_  (.Y(\proj__2.net27 ),
    .A(\proj__2.net15 ));
 sg13g2_or2_1 \proj__2.or1/_0_  (.X(\proj__2.net6 ),
    .B(\proj__2.net30 ),
    .A(\proj__2.net2 ));
 sg13g2_or2_1 \proj__2.or2/_0_  (.X(\proj__2.net5 ),
    .B(\proj__2.net31 ),
    .A(\proj__2.net2 ));
 sg13g2_or2_1 \proj__2.or3/_0_  (.X(\proj__2.net3 ),
    .B(\proj__2.net32 ),
    .A(\proj__2.net2 ));
 sg13g2_or2_1 \proj__2.or4/_0_  (.X(\proj__2.net31 ),
    .B(\proj__2.net33 ),
    .A(\proj__2.net23 ));
 sg13g2_or2_1 \proj__2.or5/_0_  (.X(\proj__2.net30 ),
    .B(\proj__2.net34 ),
    .A(\proj__2.net23 ));
 sg13g2_or2_1 \proj__2.or6/_0_  (.X(\proj__2.net34 ),
    .B(\proj__2.net29 ),
    .A(\proj__2.net4 ));
 sg13g2_or2_1 \proj__2.or7/_0_  (.X(\proj__2.net32 ),
    .B(\proj__2.net29 ),
    .A(\proj__2.net4 ));
 sg13g2_or2_1 \proj__2.or8/_0_  (.X(\proj__2.net33 ),
    .B(\proj__2.net29 ),
    .A(\proj__2.net4 ));
 sg13g2_or2_1 \proj__3.or1/_0_  (.X(\proj__3.net9 ),
    .B(net42),
    .A(net41));
 sg13g2_inv_1 \proj__4.not1/_0_  (.Y(\proj__4.net9 ),
    .A(net43));
 sg13g2_inv_1 \proj__4.not2/_0_  (.Y(\proj__4.net10 ),
    .A(net39));
 sg13g2_inv_1 \proj__4.not3/_0_  (.Y(\proj__4.net11 ),
    .A(net37));
 sg13g2_inv_1 \proj__4.not4/_0_  (.Y(\proj__4.net12 ),
    .A(net36));
 sg13g2_and2_1 \proj__5.and1/_0_  (.A(net41),
    .B(net44),
    .X(\proj__5.net9 ));
 sg13g2_xor2_1 \proj__5.xor1/_0_  (.B(net44),
    .A(net40),
    .X(\proj__5.net10 ));
 sg13g2_and2_1 \proj__6.and1/_0_  (.A(net38),
    .B(net44),
    .X(\proj__6.net11 ));
 sg13g2_and2_1 \proj__6.and2/_0_  (.A(net2),
    .B(\proj__6.net11 ),
    .X(\proj__6.net12 ));
 sg13g2_and2_1 \proj__6.and3/_0_  (.A(net3),
    .B(\proj__6.net12 ),
    .X(\proj__6.net5 ));
 sg13g2_and2_2 \proj__7.and1/_0_  (.A(\proj__7.net36 ),
    .B(net40),
    .X(\proj__7.net37 ));
 sg13g2_and2_1 \proj__7.and10/_0_  (.A(\proj__7.net38 ),
    .B(\proj__7.net21 ),
    .X(\proj__7.net36 ));
 sg13g2_and2_1 \proj__7.and11/_0_  (.A(\proj__7.net29 ),
    .B(\proj__7.net32 ),
    .X(\proj__7.net38 ));
 sg13g2_and2_1 \proj__7.and12/_0_  (.A(\proj__7.net38 ),
    .B(\proj__7.net39 ),
    .X(\proj__7.net40 ));
 sg13g2_and2_1 \proj__7.and13/_0_  (.A(\proj__7.net83 ),
    .B(\proj__7.net32 ),
    .X(\proj__7.net84 ));
 sg13g2_and2_1 \proj__7.and14/_0_  (.A(\proj__7.net22 ),
    .B(\proj__7.net21 ),
    .X(\proj__7.net83 ));
 sg13g2_and2_1 \proj__7.and15/_0_  (.A(\proj__7.net24 ),
    .B(\proj__7.net84 ),
    .X(\proj__7.net85 ));
 sg13g2_and2_1 \proj__7.and16/_0_  (.A(net38),
    .B(\proj__7.net85 ),
    .X(\proj__7.net82 ));
 sg13g2_and2_1 \proj__7.and17/_0_  (.A(\proj__7.net83 ),
    .B(\proj__7.net32 ),
    .X(\proj__7.net86 ));
 sg13g2_and2_1 \proj__7.and18/_0_  (.A(net36),
    .B(\proj__7.net23 ),
    .X(\proj__7.net87 ));
 sg13g2_and2_1 \proj__7.and19/_0_  (.A(\proj__7.net86 ),
    .B(\proj__7.net87 ),
    .X(\proj__7.net88 ));
 sg13g2_and2_1 \proj__7.and2/_0_  (.A(\proj__7.net24 ),
    .B(\proj__7.net23 ),
    .X(\proj__7.net29 ));
 sg13g2_and2_1 \proj__7.and20/_0_  (.A(net38),
    .B(net45),
    .X(\proj__7.net90 ));
 sg13g2_and2_1 \proj__7.and21/_0_  (.A(\proj__7.net22 ),
    .B(\proj__7.net24 ),
    .X(\proj__7.net91 ));
 sg13g2_and2_1 \proj__7.and22/_0_  (.A(\proj__7.net32 ),
    .B(net108),
    .X(\proj__7.net93 ));
 sg13g2_and2_1 \proj__7.and23/_0_  (.A(\proj__7.net90 ),
    .B(\proj__7.net91 ),
    .X(\proj__7.net94 ));
 sg13g2_and2_1 \proj__7.and24/_0_  (.A(\proj__7.net94 ),
    .B(\proj__7.net93 ),
    .X(\proj__7.net89 ));
 sg13g2_and2_1 \proj__7.and25/_0_  (.A(\proj__7.net31 ),
    .B(\proj__7.net102 ),
    .X(\proj__7.net103 ));
 sg13g2_and2_1 \proj__7.and26/_0_  (.A(\proj__7.net29 ),
    .B(\proj__7.net83 ),
    .X(\proj__7.net102 ));
 sg13g2_and2_1 \proj__7.and27/_0_  (.A(\proj__7.net26 ),
    .B(net3),
    .X(\proj__7.net104 ));
 sg13g2_and2_1 \proj__7.and28/_0_  (.A(\proj__7.net104 ),
    .B(\proj__7.net103 ),
    .X(\proj__7.net105 ));
 sg13g2_and2_1 \proj__7.and29/_0_  (.A(\proj__7.net31 ),
    .B(\proj__7.net102 ),
    .X(\proj__7.net106 ));
 sg13g2_and2_1 \proj__7.and3/_0_  (.A(\proj__7.net26 ),
    .B(\proj__7.net25 ),
    .X(\proj__7.net30 ));
 sg13g2_and2_1 \proj__7.and30/_0_  (.A(\proj__7.net25 ),
    .B(net4),
    .X(\proj__7.net107 ));
 sg13g2_and2_1 \proj__7.and31/_0_  (.A(\proj__7.net107 ),
    .B(\proj__7.net106 ),
    .X(\proj__7.net56 ));
 sg13g2_and2_1 \proj__7.and32/_0_  (.A(\proj__7.net30 ),
    .B(\proj__7.net102 ),
    .X(\proj__7.net108 ));
 sg13g2_and2_1 \proj__7.and33/_0_  (.A(net5),
    .B(\proj__7.net28 ),
    .X(\proj__7.net109 ));
 sg13g2_and2_2 \proj__7.and34/_0_  (.A(\proj__7.net109 ),
    .B(\proj__7.net108 ),
    .X(\proj__7.net95 ));
 sg13g2_and2_1 \proj__7.and35/_0_  (.A(\proj__7.net22 ),
    .B(\proj__7.net29 ),
    .X(\proj__7.net117 ));
 sg13g2_and2_1 \proj__7.and36/_0_  (.A(\proj__7.net30 ),
    .B(\proj__7.net28 ),
    .X(\proj__7.net118 ));
 sg13g2_and2_1 \proj__7.and37/_0_  (.A(\proj__7.net118 ),
    .B(\proj__7.net117 ),
    .X(\proj__7.net119 ));
 sg13g2_and2_1 \proj__7.and38/_0_  (.A(net5),
    .B(\proj__7.net119 ),
    .X(\proj__7.net120 ));
 sg13g2_and2_1 \proj__7.and39/_0_  (.A(net44),
    .B(\proj__7.net120 ),
    .X(\proj__7.net121 ));
 sg13g2_and2_1 \proj__7.and4/_0_  (.A(net40),
    .B(net45),
    .X(\proj__7.net39 ));
 sg13g2_and2_1 \proj__7.and40/_0_  (.A(\proj__7.net24 ),
    .B(\proj__7.net83 ),
    .X(\proj__7.net122 ));
 sg13g2_and2_1 \proj__7.and41/_0_  (.A(\proj__7.net28 ),
    .B(\proj__7.net31 ),
    .X(\proj__7.net123 ));
 sg13g2_and2_1 \proj__7.and42/_0_  (.A(\proj__7.net123 ),
    .B(\proj__7.net122 ),
    .X(\proj__7.net124 ));
 sg13g2_and2_1 \proj__7.and43/_0_  (.A(net3),
    .B(net38),
    .X(\proj__7.net125 ));
 sg13g2_and2_1 \proj__7.and44/_0_  (.A(\proj__7.net124 ),
    .B(\proj__7.net125 ),
    .X(\proj__7.net126 ));
 sg13g2_and2_1 \proj__7.and45/_0_  (.A(net4),
    .B(net40),
    .X(\proj__7.net129 ));
 sg13g2_and2_1 \proj__7.and46/_0_  (.A(\proj__7.net130 ),
    .B(\proj__7.net29 ),
    .X(\proj__7.net131 ));
 sg13g2_and2_1 \proj__7.and47/_0_  (.A(\proj__7.net132 ),
    .B(\proj__7.net21 ),
    .X(\proj__7.net133 ));
 sg13g2_and2_1 \proj__7.and48/_0_  (.A(\proj__7.net131 ),
    .B(\proj__7.net129 ),
    .X(\proj__7.net132 ));
 sg13g2_and2_1 \proj__7.and49/_0_  (.A(\proj__7.net133 ),
    .B(\proj__7.net25 ),
    .X(\proj__7.net128 ));
 sg13g2_and2_1 \proj__7.and5/_0_  (.A(\proj__7.net28 ),
    .B(\proj__7.net27 ),
    .X(\proj__7.net31 ));
 sg13g2_and2_1 \proj__7.and50/_0_  (.A(\proj__7.net32 ),
    .B(\proj__7.net24 ),
    .X(\proj__7.net171 ));
 sg13g2_and2_1 \proj__7.and51/_0_  (.A(\proj__7.net28 ),
    .B(\proj__7.net27 ),
    .X(\proj__7.net130 ));
 sg13g2_and2_1 \proj__7.and52/_0_  (.A(net40),
    .B(\proj__7.net21 ),
    .X(\proj__7.net172 ));
 sg13g2_and2_1 \proj__7.and54/_0_  (.A(\proj__7.net172 ),
    .B(\proj__7.net171 ),
    .X(\proj__7.net173 ));
 sg13g2_and2_1 \proj__7.and55/_0_  (.A(\proj__7.net173 ),
    .B(net38),
    .X(\proj__7.net174 ));
 sg13g2_and2_2 \proj__7.and6/_0_  (.A(\proj__7.net31 ),
    .B(\proj__7.net30 ),
    .X(\proj__7.net32 ));
 sg13g2_and2_1 \proj__7.and7/_0_  (.A(\proj__7.net29 ),
    .B(\proj__7.net22 ),
    .X(\proj__7.net33 ));
 sg13g2_and2_1 \proj__7.and8/_0_  (.A(\proj__7.net32 ),
    .B(\proj__7.net33 ),
    .X(\proj__7.net34 ));
 sg13g2_and2_2 \proj__7.and9/_0_  (.A(\proj__7.net34 ),
    .B(net45),
    .X(\proj__7.net35 ));
 sg13g2_inv_1 \proj__7.not1/_0_  (.Y(\proj__7.net21 ),
    .A(net44));
 sg13g2_inv_1 \proj__7.not2/_0_  (.Y(\proj__7.net22 ),
    .A(net40));
 sg13g2_inv_1 \proj__7.not3/_0_  (.Y(\proj__7.net23 ),
    .A(net38));
 sg13g2_inv_1 \proj__7.not4/_0_  (.Y(\proj__7.net24 ),
    .A(net36));
 sg13g2_inv_1 \proj__7.not5/_0_  (.Y(\proj__7.net25 ),
    .A(net3));
 sg13g2_inv_1 \proj__7.not6/_0_  (.Y(\proj__7.net26 ),
    .A(net4));
 sg13g2_inv_1 \proj__7.not7/_0_  (.Y(\proj__7.net27 ),
    .A(net5));
 sg13g2_inv_1 \proj__7.not8/_0_  (.Y(\proj__7.net28 ),
    .A(net6));
 sg13g2_or2_1 \proj__7.or1/_0_  (.X(\proj__7.net50 ),
    .B(\proj__7.net40 ),
    .A(\proj__7.net82 ));
 sg13g2_or2_1 \proj__7.or10/_0_  (.X(\proj__7.net48 ),
    .B(\proj__7.net35 ),
    .A(net17));
 sg13g2_or2_1 \proj__7.or11/_0_  (.X(\proj__7.net51 ),
    .B(\proj__7.net50 ),
    .A(net18));
 sg13g2_or2_1 \proj__7.or12/_0_  (.X(\proj__7.net52 ),
    .B(\proj__7.net50 ),
    .A(net19));
 sg13g2_or2_1 \proj__7.or13/_0_  (.X(\proj__7.net53 ),
    .B(\proj__7.net50 ),
    .A(net20));
 sg13g2_or2_1 \proj__7.or14/_0_  (.X(\proj__7.net135 ),
    .B(\proj__7.net134 ),
    .A(\proj__7.net80 ));
 sg13g2_or2_1 \proj__7.or15/_0_  (.X(\proj__7.net136 ),
    .B(\proj__7.net97 ),
    .A(\proj__7.net59 ));
 sg13g2_or2_1 \proj__7.or16/_0_  (.X(\proj__7.net54 ),
    .B(\proj__7.net50 ),
    .A(net21));
 sg13g2_or2_1 \proj__7.or17/_0_  (.X(\proj__7.net55 ),
    .B(net22),
    .A(net23));
 sg13g2_or2_1 \proj__7.or18/_0_  (.X(\proj__7.net112 ),
    .B(\proj__7.net110 ),
    .A(net24));
 sg13g2_or2_1 \proj__7.or19/_0_  (.X(\proj__7.net96 ),
    .B(\proj__7.net95 ),
    .A(net25));
 sg13g2_or2_1 \proj__7.or2/_0_  (.X(\proj__7.net42 ),
    .B(\proj__7.net35 ),
    .A(net26));
 sg13g2_or2_1 \proj__7.or20/_0_  (.X(\proj__7.net58 ),
    .B(\proj__7.net56 ),
    .A(net27));
 sg13g2_or2_1 \proj__7.or21/_0_  (.X(\proj__7.net59 ),
    .B(\proj__7.net56 ),
    .A(net28));
 sg13g2_or2_1 \proj__7.or22/_0_  (.X(\proj__7.net60 ),
    .B(\proj__7.net56 ),
    .A(net29));
 sg13g2_or2_1 \proj__7.or23/_0_  (.X(\proj__7.net97 ),
    .B(\proj__7.net95 ),
    .A(net30));
 sg13g2_or2_1 \proj__7.or24/_0_  (.X(\proj__7.net61 ),
    .B(\proj__7.net56 ),
    .A(net31));
 sg13g2_or2_1 \proj__7.or25/_0_  (.X(\proj__7.net113 ),
    .B(\proj__7.net110 ),
    .A(net32));
 sg13g2_or2_1 \proj__7.or26/_0_  (.X(\proj__7.net62 ),
    .B(\proj__7.net37 ),
    .A(net33));
 sg13g2_or2_1 \proj__7.or27/_0_  (.X(\proj__7.net63 ),
    .B(\proj__7.net37 ),
    .A(net34));
 sg13g2_or2_1 \proj__7.or28/_0_  (.X(\proj__7.net64 ),
    .B(\proj__7.net37 ),
    .A(net46));
 sg13g2_or2_1 \proj__7.or29/_0_  (.X(\proj__7.net65 ),
    .B(\proj__7.net37 ),
    .A(net47));
 sg13g2_or2_1 \proj__7.or3/_0_  (.X(\proj__7.net43 ),
    .B(net48),
    .A(net49));
 sg13g2_or2_1 \proj__7.or30/_0_  (.X(\proj__7.net66 ),
    .B(\proj__7.net37 ),
    .A(net50));
 sg13g2_or2_1 \proj__7.or31/_0_  (.X(\proj__7.net137 ),
    .B(\proj__7.net79 ),
    .A(\proj__7.net136 ));
 sg13g2_or2_1 \proj__7.or32/_0_  (.X(\proj__7.net67 ),
    .B(\proj__7.net37 ),
    .A(net51));
 sg13g2_or2_1 \proj__7.or33/_0_  (.X(\proj__7.net68 ),
    .B(\proj__7.net37 ),
    .A(net52));
 sg13g2_or2_1 \proj__7.or34/_0_  (.X(\proj__7.net70 ),
    .B(net53),
    .A(\proj__7.net69 ));
 sg13g2_or2_1 \proj__7.or35/_0_  (.X(\proj__7.net71 ),
    .B(net54),
    .A(\proj__7.net69 ));
 sg13g2_or2_1 \proj__7.or36/_0_  (.X(\proj__7.net72 ),
    .B(net55),
    .A(\proj__7.net69 ));
 sg13g2_or2_1 \proj__7.or37/_0_  (.X(\proj__7.net73 ),
    .B(net56),
    .A(\proj__7.net69 ));
 sg13g2_or2_2 \proj__7.or38/_0_  (.X(\proj__7.net69 ),
    .B(\proj__7.net89 ),
    .A(\proj__7.net88 ));
 sg13g2_or2_1 \proj__7.or39/_0_  (.X(\proj__7.net114 ),
    .B(\proj__7.net110 ),
    .A(net57));
 sg13g2_or2_1 \proj__7.or4/_0_  (.X(\proj__7.net44 ),
    .B(\proj__7.net35 ),
    .A(net58));
 sg13g2_or2_1 \proj__7.or40/_0_  (.X(\proj__7.net74 ),
    .B(net59),
    .A(\proj__7.net69 ));
 sg13g2_or2_1 \proj__7.or41/_0_  (.X(\proj__7.net75 ),
    .B(net60),
    .A(\proj__7.net69 ));
 sg13g2_or2_1 \proj__7.or42/_0_  (.X(\proj__7.net98 ),
    .B(\proj__7.net95 ),
    .A(net61));
 sg13g2_or2_1 \proj__7.or43/_0_  (.X(\proj__7.net77 ),
    .B(\proj__7.net76 ),
    .A(net62));
 sg13g2_or2_1 \proj__7.or44/_0_  (.X(\proj__7.net78 ),
    .B(\proj__7.net76 ),
    .A(net63));
 sg13g2_or2_1 \proj__7.or45/_0_  (.X(\proj__7.net79 ),
    .B(\proj__7.net76 ),
    .A(net64));
 sg13g2_or2_1 \proj__7.or46/_0_  (.X(\proj__7.net80 ),
    .B(\proj__7.net76 ),
    .A(net65));
 sg13g2_or2_1 \proj__7.or47/_0_  (.X(\proj__7.net99 ),
    .B(\proj__7.net95 ),
    .A(net66));
 sg13g2_or2_1 \proj__7.or48/_0_  (.X(\proj__7.net81 ),
    .B(\proj__7.net76 ),
    .A(net67));
 sg13g2_or2_1 \proj__7.or49/_0_  (.X(\proj__7.net100 ),
    .B(\proj__7.net95 ),
    .A(net68));
 sg13g2_or2_1 \proj__7.or5/_0_  (.X(\proj__7.net45 ),
    .B(\proj__7.net35 ),
    .A(net69));
 sg13g2_or2_1 \proj__7.or50/_0_  (.X(\proj__7.net101 ),
    .B(\proj__7.net95 ),
    .A(net70));
 sg13g2_or2_1 \proj__7.or51/_0_  (.X(\proj__7.net115 ),
    .B(\proj__7.net110 ),
    .A(net71));
 sg13g2_or2_1 \proj__7.or52/_0_  (.X(\proj__7.net116 ),
    .B(\proj__7.net110 ),
    .A(net72));
 sg13g2_or2_1 \proj__7.or53/_0_  (.X(\proj__7.net127 ),
    .B(\proj__7.net121 ),
    .A(\proj__7.net126 ));
 sg13g2_or2_2 \proj__7.or54/_0_  (.X(\proj__7.net110 ),
    .B(\proj__7.net127 ),
    .A(\proj__7.net128 ));
 sg13g2_or2_1 \proj__7.or55/_0_  (.X(\proj__7.net138 ),
    .B(\proj__7.net61 ),
    .A(\proj__7.net101 ));
 sg13g2_or2_1 \proj__7.or56/_0_  (.X(\proj__7.net139 ),
    .B(\proj__7.net138 ),
    .A(\proj__7.net81 ));
 sg13g2_or2_1 \proj__7.or57/_0_  (.X(\proj__7.net140 ),
    .B(\proj__7.net98 ),
    .A(\proj__7.net77 ));
 sg13g2_or2_1 \proj__7.or58/_0_  (.X(\proj__7.net141 ),
    .B(\proj__7.net78 ),
    .A(\proj__7.net58 ));
 sg13g2_or2_1 \proj__7.or59/_0_  (.X(\proj__7.net142 ),
    .B(\proj__7.net112 ),
    .A(\proj__7.net100 ));
 sg13g2_or2_1 \proj__7.or6/_0_  (.X(\proj__7.net46 ),
    .B(\proj__7.net35 ),
    .A(net73));
 sg13g2_or2_1 \proj__7.or60/_0_  (.X(\proj__7.net143 ),
    .B(\proj__7.net113 ),
    .A(\proj__7.net99 ));
 sg13g2_or2_1 \proj__7.or61/_0_  (.X(\proj__7.net145 ),
    .B(\proj__7.net140 ),
    .A(net74));
 sg13g2_or2_1 \proj__7.or62/_0_  (.X(\proj__7.net146 ),
    .B(\proj__7.net114 ),
    .A(\proj__7.net141 ));
 sg13g2_or2_1 \proj__7.or63/_0_  (.X(\proj__7.net147 ),
    .B(\proj__7.net70 ),
    .A(\proj__7.net49 ));
 sg13g2_or2_1 \proj__7.or64/_0_  (.X(\proj__7.net148 ),
    .B(\proj__7.net51 ),
    .A(\proj__7.net71 ));
 sg13g2_or2_1 \proj__7.or65/_0_  (.X(\proj__7.net149 ),
    .B(\proj__7.net52 ),
    .A(\proj__7.net72 ));
 sg13g2_or2_1 \proj__7.or66/_0_  (.X(\proj__7.net150 ),
    .B(\proj__7.net73 ),
    .A(\proj__7.net53 ));
 sg13g2_or2_1 \proj__7.or67/_0_  (.X(\proj__7.net151 ),
    .B(\proj__7.net54 ),
    .A(\proj__7.net74 ));
 sg13g2_or2_1 \proj__7.or68/_0_  (.X(\proj__7.net152 ),
    .B(\proj__7.net75 ),
    .A(\proj__7.net55 ));
 sg13g2_or2_1 \proj__7.or69/_0_  (.X(\proj__7.net10 ),
    .B(\proj__7.net142 ),
    .A(\proj__7.net168 ));
 sg13g2_or2_1 \proj__7.or7/_0_  (.X(\proj__7.net134 ),
    .B(\proj__7.net96 ),
    .A(\proj__7.net60 ));
 sg13g2_or2_1 \proj__7.or70/_0_  (.X(\proj__7.net153 ),
    .B(\proj__7.net42 ),
    .A(\proj__7.net62 ));
 sg13g2_or2_1 \proj__7.or71/_0_  (.X(\proj__7.net154 ),
    .B(\proj__7.net43 ),
    .A(\proj__7.net63 ));
 sg13g2_or2_1 \proj__7.or72/_0_  (.X(\proj__7.net155 ),
    .B(\proj__7.net44 ),
    .A(\proj__7.net64 ));
 sg13g2_or2_1 \proj__7.or73/_0_  (.X(\proj__7.net156 ),
    .B(\proj__7.net45 ),
    .A(\proj__7.net65 ));
 sg13g2_or2_1 \proj__7.or74/_0_  (.X(\proj__7.net157 ),
    .B(\proj__7.net67 ),
    .A(\proj__7.net47 ));
 sg13g2_or2_1 \proj__7.or75/_0_  (.X(\proj__7.net158 ),
    .B(\proj__7.net68 ),
    .A(\proj__7.net48 ));
 sg13g2_or2_1 \proj__7.or76/_0_  (.X(\proj__7.net159 ),
    .B(\proj__7.net46 ),
    .A(\proj__7.net66 ));
 sg13g2_or2_1 \proj__7.or77/_0_  (.X(\proj__7.net160 ),
    .B(\proj__7.net115 ),
    .A(\proj__7.net137 ));
 sg13g2_or2_1 \proj__7.or78/_0_  (.X(\proj__7.net161 ),
    .B(\proj__7.net116 ),
    .A(\proj__7.net135 ));
 sg13g2_or2_1 \proj__7.or79/_0_  (.X(\proj__7.net162 ),
    .B(\proj__7.net139 ),
    .A(net75));
 sg13g2_or2_1 \proj__7.or8/_0_  (.X(\proj__7.net49 ),
    .B(net76),
    .A(net77));
 sg13g2_or2_1 \proj__7.or81/_0_  (.X(\proj__7.net163 ),
    .B(\proj__7.net147 ),
    .A(\proj__7.net153 ));
 sg13g2_or2_1 \proj__7.or82/_0_  (.X(\proj__7.net164 ),
    .B(\proj__7.net148 ),
    .A(\proj__7.net154 ));
 sg13g2_or2_1 \proj__7.or83/_0_  (.X(\proj__7.net165 ),
    .B(\proj__7.net149 ),
    .A(\proj__7.net155 ));
 sg13g2_or2_1 \proj__7.or84/_0_  (.X(\proj__7.net166 ),
    .B(\proj__7.net150 ),
    .A(\proj__7.net156 ));
 sg13g2_or2_1 \proj__7.or85/_0_  (.X(\proj__7.net167 ),
    .B(\proj__7.net151 ),
    .A(\proj__7.net157 ));
 sg13g2_or2_1 \proj__7.or86/_0_  (.X(\proj__7.net168 ),
    .B(\proj__7.net152 ),
    .A(\proj__7.net158 ));
 sg13g2_or2_1 \proj__7.or87/_0_  (.X(\proj__7.net170 ),
    .B(net78),
    .A(\proj__7.net159 ));
 sg13g2_or2_1 \proj__7.or88/_0_  (.X(\proj__7.net11 ),
    .B(\proj__7.net143 ),
    .A(\proj__7.net163 ));
 sg13g2_or2_1 \proj__7.or89/_0_  (.X(\proj__7.net12 ),
    .B(\proj__7.net145 ),
    .A(\proj__7.net164 ));
 sg13g2_or2_1 \proj__7.or9/_0_  (.X(\proj__7.net47 ),
    .B(\proj__7.net35 ),
    .A(net79));
 sg13g2_or2_1 \proj__7.or90/_0_  (.X(\proj__7.net13 ),
    .B(\proj__7.net146 ),
    .A(\proj__7.net165 ));
 sg13g2_or2_1 \proj__7.or91/_0_  (.X(\proj__7.net14 ),
    .B(\proj__7.net160 ),
    .A(\proj__7.net166 ));
 sg13g2_or2_1 \proj__7.or92/_0_  (.X(\proj__7.net9 ),
    .B(\proj__7.net162 ),
    .A(\proj__7.net167 ));
 sg13g2_or2_1 \proj__7.or93/_0_  (.X(\proj__7.net15 ),
    .B(\proj__7.net161 ),
    .A(\proj__7.net170 ));
 sg13g2_or2_1 \proj__7.or94/_0_  (.X(\proj__7.net76 ),
    .B(\proj__7.net105 ),
    .A(\proj__7.net174 ));
 sg13g2_and2_1 \proj__9.and1/_0_  (.A(\proj__9.net21 ),
    .B(\proj__9.net20 ),
    .X(\proj__9.net7 ));
 sg13g2_and2_1 \proj__9.and2/_0_  (.A(\proj__9.net26 ),
    .B(\proj__9.net20 ),
    .X(\proj__9.net8 ));
 sg13g2_and2_1 \proj__9.and3/_0_  (.A(\proj__9.net26 ),
    .B(\proj__9.net20 ),
    .X(\proj__9.net9 ));
 sg13g2_and2_1 \proj__9.and4/_0_  (.A(\proj__9.net21 ),
    .B(\proj__9.net20 ),
    .X(\proj__9.net10 ));
 sg13g2_and2_1 \proj__9.and5/_0_  (.A(\proj__9.net21 ),
    .B(\proj__9.net20 ),
    .X(\proj__9.net11 ));
 sg13g2_and2_1 \proj__9.and6/_0_  (.A(\proj__9.net21 ),
    .B(\proj__9.net20 ),
    .X(\proj__9.net12 ));
 sg13g2_and2_1 \proj__9.and7/_0_  (.A(\proj__9.net21 ),
    .B(\proj__9.net20 ),
    .X(\proj__9.net13 ));
 sg13g2_and2_1 \proj__9.and8/_0_  (.A(\proj__9.net21 ),
    .B(\proj__9.net20 ),
    .X(\proj__9.net14 ));
 sg13g2_inv_2 \proj__9.not1/_0_  (.Y(\proj__9.net21 ),
    .A(net42));
 sg13g2_inv_1 \proj__9.not2/_0_  (.Y(\proj__9.net27 ),
    .A(net42));
 sg13g2_inv_1 \proj__9.not3/_0_  (.Y(\proj__9.net26 ),
    .A(\proj__9.net27 ));
 sg13g2_or2_1 \proj__9.or1/_0_  (.X(\proj__9.net22 ),
    .B(net40),
    .A(net44));
 sg13g2_or2_1 \proj__9.or2/_0_  (.X(\proj__9.net23 ),
    .B(\proj__9.net22 ),
    .A(net37));
 sg13g2_or2_1 \proj__9.or3/_0_  (.X(\proj__9.net24 ),
    .B(\proj__9.net23 ),
    .A(net36));
 sg13g2_or2_1 \proj__9.or4/_0_  (.X(\proj__9.net25 ),
    .B(\proj__9.net24 ),
    .A(net3));
 sg13g2_or2_2 \proj__9.or5/_0_  (.X(\proj__9.net20 ),
    .B(\proj__9.net25 ),
    .A(net4));
 sg13g2_buf_2 fanout35 (.A(_066_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(net2),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(ui_in[2]),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(ui_in[2]),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(net41),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(net41),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(ui_in[1]),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(net43),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(net45),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(net45),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(ui_in[0]),
    .X(net45));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[0]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_tielo \proj__0.flop1/_4__11  (.L_LO(net11));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_1_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_1_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_1_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_1_1__leaf_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_1_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_0__005_ (.A(_005_),
    .X(clknet_0__005_));
 sg13g2_buf_2 clkbuf_1_0__f__005_ (.A(clknet_0__005_),
    .X(clknet_1_0__leaf__005_));
 sg13g2_buf_2 clkbuf_1_1__f__005_ (.A(clknet_0__005_),
    .X(clknet_1_1__leaf__005_));
 sg13g2_buf_1 clkload2 (.A(clknet_1_0__leaf__005_));
 sg13g2_dlygate4sd3_1 hold1 (.A(\proj__2.net12 ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold2 (.A(\proj__0.net8 ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold3 (.A(\proj__0.net5 ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold4 (.A(\proj__0.net7 ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold5 (.A(\proj__0.net3 ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold6 (.A(\proj__0.net6 ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold7 (.A(\proj__0.net4 ),
    .X(net119));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_fill_2 FILLER_17_98 ();
 sg13g2_fill_1 FILLER_17_100 ();
 sg13g2_decap_8 FILLER_17_106 ();
 sg13g2_decap_8 FILLER_17_113 ();
 sg13g2_decap_8 FILLER_17_120 ();
 sg13g2_decap_8 FILLER_17_127 ();
 sg13g2_decap_8 FILLER_17_134 ();
 sg13g2_decap_8 FILLER_17_141 ();
 sg13g2_decap_8 FILLER_17_148 ();
 sg13g2_decap_8 FILLER_17_155 ();
 sg13g2_decap_8 FILLER_17_162 ();
 sg13g2_decap_8 FILLER_17_169 ();
 sg13g2_decap_8 FILLER_17_176 ();
 sg13g2_decap_8 FILLER_17_183 ();
 sg13g2_decap_8 FILLER_17_190 ();
 sg13g2_decap_8 FILLER_17_197 ();
 sg13g2_decap_8 FILLER_17_204 ();
 sg13g2_decap_8 FILLER_17_211 ();
 sg13g2_decap_8 FILLER_17_218 ();
 sg13g2_decap_8 FILLER_17_225 ();
 sg13g2_decap_8 FILLER_17_232 ();
 sg13g2_decap_8 FILLER_17_239 ();
 sg13g2_decap_8 FILLER_17_246 ();
 sg13g2_decap_8 FILLER_17_253 ();
 sg13g2_decap_8 FILLER_17_260 ();
 sg13g2_decap_8 FILLER_17_267 ();
 sg13g2_decap_8 FILLER_17_274 ();
 sg13g2_decap_8 FILLER_17_281 ();
 sg13g2_decap_8 FILLER_17_288 ();
 sg13g2_decap_8 FILLER_17_295 ();
 sg13g2_decap_8 FILLER_17_302 ();
 sg13g2_decap_8 FILLER_17_309 ();
 sg13g2_decap_8 FILLER_17_316 ();
 sg13g2_decap_8 FILLER_17_323 ();
 sg13g2_decap_8 FILLER_17_330 ();
 sg13g2_decap_8 FILLER_17_337 ();
 sg13g2_decap_8 FILLER_17_344 ();
 sg13g2_decap_8 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_358 ();
 sg13g2_decap_8 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_fill_2 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_244 ();
 sg13g2_decap_8 FILLER_23_251 ();
 sg13g2_decap_8 FILLER_23_258 ();
 sg13g2_decap_8 FILLER_23_265 ();
 sg13g2_decap_8 FILLER_23_272 ();
 sg13g2_decap_8 FILLER_23_279 ();
 sg13g2_decap_8 FILLER_23_286 ();
 sg13g2_decap_8 FILLER_23_293 ();
 sg13g2_decap_8 FILLER_23_300 ();
 sg13g2_decap_8 FILLER_23_307 ();
 sg13g2_decap_8 FILLER_23_314 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_decap_8 FILLER_23_335 ();
 sg13g2_decap_8 FILLER_23_342 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_262 ();
 sg13g2_decap_8 FILLER_24_269 ();
 sg13g2_decap_8 FILLER_24_276 ();
 sg13g2_decap_8 FILLER_24_283 ();
 sg13g2_decap_8 FILLER_24_290 ();
 sg13g2_decap_8 FILLER_24_297 ();
 sg13g2_decap_8 FILLER_24_304 ();
 sg13g2_decap_8 FILLER_24_311 ();
 sg13g2_decap_8 FILLER_24_318 ();
 sg13g2_decap_8 FILLER_24_325 ();
 sg13g2_decap_8 FILLER_24_332 ();
 sg13g2_decap_8 FILLER_24_339 ();
 sg13g2_decap_8 FILLER_24_346 ();
 sg13g2_decap_8 FILLER_24_353 ();
 sg13g2_decap_8 FILLER_24_360 ();
 sg13g2_decap_8 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_decap_4 FILLER_25_215 ();
 sg13g2_fill_1 FILLER_25_219 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_fill_2 FILLER_25_231 ();
 sg13g2_fill_2 FILLER_25_236 ();
 sg13g2_fill_1 FILLER_25_238 ();
 sg13g2_fill_1 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_260 ();
 sg13g2_decap_8 FILLER_25_267 ();
 sg13g2_decap_8 FILLER_25_274 ();
 sg13g2_decap_8 FILLER_25_281 ();
 sg13g2_decap_8 FILLER_25_288 ();
 sg13g2_decap_8 FILLER_25_295 ();
 sg13g2_decap_8 FILLER_25_302 ();
 sg13g2_decap_8 FILLER_25_309 ();
 sg13g2_decap_8 FILLER_25_316 ();
 sg13g2_decap_8 FILLER_25_323 ();
 sg13g2_decap_8 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_25_337 ();
 sg13g2_decap_8 FILLER_25_344 ();
 sg13g2_decap_8 FILLER_25_351 ();
 sg13g2_decap_8 FILLER_25_358 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_fill_2 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_174 ();
 sg13g2_decap_8 FILLER_26_181 ();
 sg13g2_decap_8 FILLER_26_188 ();
 sg13g2_decap_4 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_199 ();
 sg13g2_decap_8 FILLER_26_226 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_fill_1 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_269 ();
 sg13g2_decap_8 FILLER_26_276 ();
 sg13g2_decap_8 FILLER_26_283 ();
 sg13g2_decap_8 FILLER_26_290 ();
 sg13g2_decap_8 FILLER_26_297 ();
 sg13g2_decap_8 FILLER_26_304 ();
 sg13g2_decap_8 FILLER_26_311 ();
 sg13g2_decap_8 FILLER_26_318 ();
 sg13g2_decap_8 FILLER_26_325 ();
 sg13g2_decap_8 FILLER_26_332 ();
 sg13g2_decap_8 FILLER_26_339 ();
 sg13g2_decap_8 FILLER_26_346 ();
 sg13g2_decap_8 FILLER_26_353 ();
 sg13g2_decap_8 FILLER_26_360 ();
 sg13g2_decap_8 FILLER_26_367 ();
 sg13g2_decap_8 FILLER_26_374 ();
 sg13g2_decap_8 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_4 FILLER_27_133 ();
 sg13g2_decap_4 FILLER_27_176 ();
 sg13g2_decap_8 FILLER_27_187 ();
 sg13g2_decap_8 FILLER_27_194 ();
 sg13g2_decap_4 FILLER_27_206 ();
 sg13g2_fill_1 FILLER_27_210 ();
 sg13g2_decap_4 FILLER_27_220 ();
 sg13g2_fill_1 FILLER_27_224 ();
 sg13g2_fill_1 FILLER_27_246 ();
 sg13g2_decap_8 FILLER_27_262 ();
 sg13g2_decap_8 FILLER_27_269 ();
 sg13g2_decap_8 FILLER_27_276 ();
 sg13g2_decap_8 FILLER_27_283 ();
 sg13g2_decap_8 FILLER_27_290 ();
 sg13g2_decap_8 FILLER_27_297 ();
 sg13g2_decap_8 FILLER_27_304 ();
 sg13g2_decap_8 FILLER_27_311 ();
 sg13g2_decap_4 FILLER_27_318 ();
 sg13g2_fill_1 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_332 ();
 sg13g2_decap_8 FILLER_27_339 ();
 sg13g2_decap_8 FILLER_27_346 ();
 sg13g2_decap_8 FILLER_27_353 ();
 sg13g2_decap_8 FILLER_27_360 ();
 sg13g2_decap_8 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_374 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_fill_2 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_128 ();
 sg13g2_decap_4 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_137 ();
 sg13g2_decap_4 FILLER_28_163 ();
 sg13g2_fill_2 FILLER_28_167 ();
 sg13g2_fill_2 FILLER_28_190 ();
 sg13g2_fill_1 FILLER_28_192 ();
 sg13g2_fill_2 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_240 ();
 sg13g2_decap_8 FILLER_28_247 ();
 sg13g2_decap_8 FILLER_28_263 ();
 sg13g2_decap_8 FILLER_28_270 ();
 sg13g2_decap_8 FILLER_28_277 ();
 sg13g2_decap_8 FILLER_28_284 ();
 sg13g2_decap_8 FILLER_28_291 ();
 sg13g2_fill_2 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_310 ();
 sg13g2_decap_4 FILLER_28_316 ();
 sg13g2_fill_2 FILLER_28_320 ();
 sg13g2_decap_4 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_351 ();
 sg13g2_fill_2 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_370 ();
 sg13g2_decap_4 FILLER_28_377 ();
 sg13g2_fill_2 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_4 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_fill_1 FILLER_29_166 ();
 sg13g2_decap_8 FILLER_29_170 ();
 sg13g2_decap_8 FILLER_29_188 ();
 sg13g2_decap_8 FILLER_29_209 ();
 sg13g2_decap_4 FILLER_29_216 ();
 sg13g2_fill_1 FILLER_29_220 ();
 sg13g2_fill_2 FILLER_29_226 ();
 sg13g2_decap_8 FILLER_29_236 ();
 sg13g2_decap_8 FILLER_29_268 ();
 sg13g2_decap_8 FILLER_29_275 ();
 sg13g2_fill_1 FILLER_29_306 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_29_326 ();
 sg13g2_decap_4 FILLER_29_353 ();
 sg13g2_decap_8 FILLER_29_374 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_119 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_fill_1 FILLER_30_198 ();
 sg13g2_decap_4 FILLER_30_219 ();
 sg13g2_fill_1 FILLER_30_263 ();
 sg13g2_decap_4 FILLER_30_282 ();
 sg13g2_fill_1 FILLER_30_286 ();
 sg13g2_fill_1 FILLER_30_300 ();
 sg13g2_fill_1 FILLER_30_310 ();
 sg13g2_fill_2 FILLER_30_321 ();
 sg13g2_fill_2 FILLER_30_338 ();
 sg13g2_decap_8 FILLER_30_344 ();
 sg13g2_fill_2 FILLER_30_351 ();
 sg13g2_decap_8 FILLER_30_368 ();
 sg13g2_fill_2 FILLER_30_384 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_4 FILLER_31_119 ();
 sg13g2_fill_1 FILLER_31_164 ();
 sg13g2_decap_4 FILLER_31_170 ();
 sg13g2_decap_4 FILLER_31_188 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_decap_4 FILLER_31_217 ();
 sg13g2_fill_2 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_240 ();
 sg13g2_fill_2 FILLER_31_246 ();
 sg13g2_fill_1 FILLER_31_248 ();
 sg13g2_fill_2 FILLER_31_264 ();
 sg13g2_decap_8 FILLER_31_275 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_fill_1 FILLER_31_290 ();
 sg13g2_decap_8 FILLER_31_296 ();
 sg13g2_decap_8 FILLER_31_303 ();
 sg13g2_fill_2 FILLER_31_310 ();
 sg13g2_fill_1 FILLER_31_312 ();
 sg13g2_fill_2 FILLER_31_317 ();
 sg13g2_fill_1 FILLER_31_319 ();
 sg13g2_fill_2 FILLER_31_329 ();
 sg13g2_fill_1 FILLER_31_331 ();
 sg13g2_decap_8 FILLER_31_342 ();
 sg13g2_fill_1 FILLER_31_354 ();
 sg13g2_decap_4 FILLER_31_363 ();
 sg13g2_fill_1 FILLER_31_367 ();
 sg13g2_decap_8 FILLER_31_373 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_fill_2 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_166 ();
 sg13g2_fill_2 FILLER_32_192 ();
 sg13g2_fill_2 FILLER_32_223 ();
 sg13g2_decap_8 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_decap_4 FILLER_32_280 ();
 sg13g2_fill_2 FILLER_32_284 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_fill_2 FILLER_32_311 ();
 sg13g2_fill_2 FILLER_32_331 ();
 sg13g2_fill_2 FILLER_32_337 ();
 sg13g2_fill_2 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_346 ();
 sg13g2_fill_2 FILLER_32_362 ();
 sg13g2_fill_1 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_383 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_4 FILLER_33_105 ();
 sg13g2_decap_4 FILLER_33_169 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_2 FILLER_33_180 ();
 sg13g2_decap_4 FILLER_33_199 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_fill_2 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_238 ();
 sg13g2_decap_4 FILLER_33_253 ();
 sg13g2_fill_1 FILLER_33_257 ();
 sg13g2_decap_8 FILLER_33_263 ();
 sg13g2_fill_2 FILLER_33_270 ();
 sg13g2_fill_1 FILLER_33_272 ();
 sg13g2_fill_1 FILLER_33_278 ();
 sg13g2_fill_1 FILLER_33_308 ();
 sg13g2_fill_1 FILLER_33_319 ();
 sg13g2_fill_2 FILLER_33_326 ();
 sg13g2_fill_1 FILLER_33_328 ();
 sg13g2_decap_4 FILLER_33_334 ();
 sg13g2_fill_2 FILLER_33_338 ();
 sg13g2_fill_2 FILLER_33_345 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_decap_4 FILLER_33_356 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_decap_4 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_4 FILLER_34_119 ();
 sg13g2_fill_1 FILLER_34_123 ();
 sg13g2_fill_1 FILLER_34_132 ();
 sg13g2_decap_4 FILLER_34_168 ();
 sg13g2_decap_4 FILLER_34_217 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_decap_8 FILLER_34_228 ();
 sg13g2_fill_2 FILLER_34_235 ();
 sg13g2_fill_1 FILLER_34_237 ();
 sg13g2_decap_4 FILLER_34_248 ();
 sg13g2_decap_8 FILLER_34_272 ();
 sg13g2_fill_2 FILLER_34_279 ();
 sg13g2_fill_1 FILLER_34_281 ();
 sg13g2_fill_2 FILLER_34_302 ();
 sg13g2_fill_1 FILLER_34_304 ();
 sg13g2_fill_2 FILLER_34_308 ();
 sg13g2_fill_1 FILLER_34_349 ();
 sg13g2_fill_2 FILLER_34_355 ();
 sg13g2_fill_2 FILLER_34_367 ();
 sg13g2_fill_2 FILLER_34_378 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_fill_2 FILLER_34_390 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_120 ();
 sg13g2_fill_1 FILLER_35_122 ();
 sg13g2_fill_2 FILLER_35_130 ();
 sg13g2_fill_2 FILLER_35_149 ();
 sg13g2_decap_4 FILLER_35_161 ();
 sg13g2_fill_1 FILLER_35_165 ();
 sg13g2_fill_2 FILLER_35_169 ();
 sg13g2_fill_1 FILLER_35_171 ();
 sg13g2_decap_4 FILLER_35_190 ();
 sg13g2_decap_4 FILLER_35_233 ();
 sg13g2_decap_4 FILLER_35_248 ();
 sg13g2_decap_8 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_270 ();
 sg13g2_decap_8 FILLER_35_304 ();
 sg13g2_fill_2 FILLER_35_311 ();
 sg13g2_decap_8 FILLER_35_333 ();
 sg13g2_fill_1 FILLER_35_340 ();
 sg13g2_decap_8 FILLER_35_355 ();
 sg13g2_decap_8 FILLER_35_372 ();
 sg13g2_fill_2 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_395 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_4 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_4 FILLER_36_161 ();
 sg13g2_fill_2 FILLER_36_165 ();
 sg13g2_fill_2 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_174 ();
 sg13g2_decap_8 FILLER_36_205 ();
 sg13g2_decap_8 FILLER_36_212 ();
 sg13g2_decap_4 FILLER_36_255 ();
 sg13g2_fill_2 FILLER_36_262 ();
 sg13g2_fill_1 FILLER_36_264 ();
 sg13g2_decap_4 FILLER_36_268 ();
 sg13g2_fill_2 FILLER_36_272 ();
 sg13g2_decap_4 FILLER_36_284 ();
 sg13g2_decap_4 FILLER_36_293 ();
 sg13g2_fill_2 FILLER_36_297 ();
 sg13g2_fill_2 FILLER_36_310 ();
 sg13g2_fill_2 FILLER_36_317 ();
 sg13g2_fill_2 FILLER_36_329 ();
 sg13g2_fill_1 FILLER_36_331 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_fill_2 FILLER_36_380 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_decap_4 FILLER_36_393 ();
 sg13g2_fill_1 FILLER_36_397 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_fill_1 FILLER_37_175 ();
 sg13g2_decap_4 FILLER_37_181 ();
 sg13g2_fill_2 FILLER_37_185 ();
 sg13g2_decap_8 FILLER_37_214 ();
 sg13g2_fill_1 FILLER_37_221 ();
 sg13g2_decap_4 FILLER_37_233 ();
 sg13g2_fill_1 FILLER_37_237 ();
 sg13g2_fill_2 FILLER_37_278 ();
 sg13g2_fill_1 FILLER_37_280 ();
 sg13g2_decap_4 FILLER_37_332 ();
 sg13g2_fill_1 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_352 ();
 sg13g2_fill_2 FILLER_37_372 ();
 sg13g2_fill_1 FILLER_37_374 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_4 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_211 ();
 sg13g2_decap_8 FILLER_38_235 ();
 sg13g2_decap_8 FILLER_38_242 ();
 sg13g2_decap_4 FILLER_38_249 ();
 sg13g2_fill_1 FILLER_38_253 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_4 FILLER_38_266 ();
 sg13g2_fill_2 FILLER_38_270 ();
 sg13g2_fill_1 FILLER_38_286 ();
 sg13g2_fill_2 FILLER_38_312 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_decap_8 FILLER_38_353 ();
 sg13g2_decap_8 FILLER_38_360 ();
 sg13g2_decap_8 FILLER_38_367 ();
 sg13g2_fill_2 FILLER_38_374 ();
 sg13g2_decap_8 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 assign uio_oe[0] = net80;
 assign uio_oe[1] = net81;
 assign uio_oe[2] = net82;
 assign uio_oe[3] = net83;
 assign uio_oe[4] = net84;
 assign uio_oe[5] = net85;
 assign uio_oe[6] = net86;
 assign uio_oe[7] = net87;
 assign uio_out[0] = net88;
 assign uio_out[1] = net89;
 assign uio_out[2] = net90;
 assign uio_out[3] = net91;
 assign uio_out[4] = net92;
 assign uio_out[5] = net93;
 assign uio_out[6] = net94;
 assign uio_out[7] = net95;
endmodule

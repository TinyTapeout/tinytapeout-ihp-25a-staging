module tt_um_jmack2201 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire clknet_0_clk;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire \wrapper.h_count[0] ;
 wire \wrapper.h_count[1] ;
 wire \wrapper.h_count[2] ;
 wire \wrapper.h_count[3] ;
 wire \wrapper.h_count[4] ;
 wire \wrapper.h_count[5] ;
 wire \wrapper.h_count[6] ;
 wire \wrapper.h_count[7] ;
 wire \wrapper.h_count[8] ;
 wire \wrapper.h_count[9] ;
 wire \wrapper.hsync ;
 wire \wrapper.pixel.background_state[0] ;
 wire \wrapper.pixel.background_state[1] ;
 wire \wrapper.pixel.background_state[2] ;
 wire \wrapper.pixel.background_state[3] ;
 wire \wrapper.pixel.lfsr_reg[0] ;
 wire \wrapper.pixel.lfsr_reg[10] ;
 wire \wrapper.pixel.lfsr_reg[11] ;
 wire \wrapper.pixel.lfsr_reg[12] ;
 wire \wrapper.pixel.lfsr_reg[13] ;
 wire \wrapper.pixel.lfsr_reg[14] ;
 wire \wrapper.pixel.lfsr_reg[15] ;
 wire \wrapper.pixel.lfsr_reg[1] ;
 wire \wrapper.pixel.lfsr_reg[2] ;
 wire \wrapper.pixel.lfsr_reg[3] ;
 wire \wrapper.pixel.lfsr_reg[4] ;
 wire \wrapper.pixel.lfsr_reg[5] ;
 wire \wrapper.pixel.lfsr_reg[6] ;
 wire \wrapper.pixel.lfsr_reg[7] ;
 wire \wrapper.pixel.lfsr_reg[8] ;
 wire \wrapper.pixel.lfsr_reg[9] ;
 wire \wrapper.pixel.looping_background_count[0] ;
 wire \wrapper.pixel.looping_background_count[1] ;
 wire \wrapper.pixel.looping_background_count[2] ;
 wire \wrapper.pixel.looping_background_count[3] ;
 wire \wrapper.pixel.moving_counter[0] ;
 wire \wrapper.pixel.moving_counter[1] ;
 wire \wrapper.pixel.moving_counter[2] ;
 wire \wrapper.pixel.moving_counter[3] ;
 wire \wrapper.pixel.moving_counter[4] ;
 wire \wrapper.pixel.moving_counter[5] ;
 wire \wrapper.pixel.moving_counter[6] ;
 wire \wrapper.pixel.moving_counter[7] ;
 wire \wrapper.pixel.prev_y[0] ;
 wire \wrapper.pixel.prev_y[1] ;
 wire \wrapper.pixel.prev_y[2] ;
 wire \wrapper.pixel.prev_y[3] ;
 wire \wrapper.pixel.prev_y[4] ;
 wire \wrapper.pixel.prev_y[5] ;
 wire \wrapper.pixel.prev_y[6] ;
 wire \wrapper.pixel.prev_y[7] ;
 wire \wrapper.pixel.prev_y[8] ;
 wire \wrapper.pixel.prev_y[9] ;
 wire \wrapper.pixel.rom0.color_out[0] ;
 wire \wrapper.pixel.rom0.color_out[1] ;
 wire \wrapper.pixel.rom0.color_out[2] ;
 wire \wrapper.pixel.rom0.color_out[3] ;
 wire \wrapper.pixel.rom0.color_out[4] ;
 wire \wrapper.pixel.rom0.color_out[5] ;
 wire \wrapper.pixel.solid_color[0] ;
 wire \wrapper.pixel.solid_color[1] ;
 wire \wrapper.pixel.solid_color[2] ;
 wire \wrapper.pixel.solid_color[3] ;
 wire \wrapper.pixel.solid_color[4] ;
 wire \wrapper.pixel.solid_color[5] ;
 wire \wrapper.pixel.sprite_left[0] ;
 wire \wrapper.pixel.sprite_left[1] ;
 wire \wrapper.pixel.sprite_left[2] ;
 wire \wrapper.pixel.sprite_left[3] ;
 wire \wrapper.pixel.sprite_left[4] ;
 wire \wrapper.pixel.sprite_left[5] ;
 wire \wrapper.pixel.sprite_left[6] ;
 wire \wrapper.pixel.sprite_left[7] ;
 wire \wrapper.pixel.sprite_left[8] ;
 wire \wrapper.pixel.sprite_left[9] ;
 wire \wrapper.pixel.sprite_top[0] ;
 wire \wrapper.pixel.sprite_top[1] ;
 wire \wrapper.pixel.sprite_top[2] ;
 wire \wrapper.pixel.sprite_top[3] ;
 wire \wrapper.pixel.sprite_top[4] ;
 wire \wrapper.pixel.sprite_top[5] ;
 wire \wrapper.pixel.sprite_top[6] ;
 wire \wrapper.pixel.sprite_top[7] ;
 wire \wrapper.pixel.sprite_top[8] ;
 wire \wrapper.pixel.sprite_top[9] ;
 wire \wrapper.pixel.vpos[0] ;
 wire \wrapper.pixel.vpos[1] ;
 wire \wrapper.pixel.vpos[2] ;
 wire \wrapper.pixel.vpos[3] ;
 wire \wrapper.pixel.vpos[4] ;
 wire \wrapper.pixel.vpos[5] ;
 wire \wrapper.pixel.vpos[6] ;
 wire \wrapper.pixel.vpos[7] ;
 wire \wrapper.pixel.vpos[8] ;
 wire \wrapper.pixel.vpos[9] ;
 wire \wrapper.pixel.vsync ;
 wire \wrapper.pixel.x_mov ;
 wire \wrapper.pixel.y_mov ;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;

 sg13g2_inv_1 _1533_ (.Y(_0601_),
    .A(net219));
 sg13g2_inv_1 _1534_ (.Y(_0602_),
    .A(net218));
 sg13g2_inv_2 _1535_ (.Y(_0603_),
    .A(\wrapper.pixel.vpos[7] ));
 sg13g2_inv_4 _1536_ (.A(net541),
    .Y(_0604_));
 sg13g2_inv_2 _1537_ (.Y(_0605_),
    .A(net544));
 sg13g2_inv_1 _1538_ (.Y(_0606_),
    .A(net551));
 sg13g2_inv_2 _1539_ (.Y(_0607_),
    .A(net552));
 sg13g2_inv_2 _1540_ (.Y(_0608_),
    .A(net557));
 sg13g2_inv_1 _1541_ (.Y(_0609_),
    .A(\wrapper.pixel.sprite_top[7] ));
 sg13g2_inv_1 _1542_ (.Y(_0610_),
    .A(\wrapper.pixel.sprite_top[4] ));
 sg13g2_inv_1 _1543_ (.Y(_0611_),
    .A(net191));
 sg13g2_inv_1 _1544_ (.Y(_0612_),
    .A(\wrapper.pixel.sprite_top[1] ));
 sg13g2_inv_1 _1545_ (.Y(_0613_),
    .A(\wrapper.pixel.sprite_top[0] ));
 sg13g2_inv_1 _1546_ (.Y(_0614_),
    .A(\wrapper.pixel.sprite_left[7] ));
 sg13g2_inv_1 _1547_ (.Y(_0615_),
    .A(\wrapper.pixel.sprite_left[5] ));
 sg13g2_inv_1 _1548_ (.Y(_0616_),
    .A(\wrapper.pixel.sprite_left[4] ));
 sg13g2_inv_1 _1549_ (.Y(_0617_),
    .A(net215));
 sg13g2_inv_1 _1550_ (.Y(_0618_),
    .A(\wrapper.pixel.sprite_left[0] ));
 sg13g2_inv_1 _1551_ (.Y(_0619_),
    .A(net169));
 sg13g2_inv_1 _1552_ (.Y(_0620_),
    .A(net168));
 sg13g2_inv_1 _1553_ (.Y(_0621_),
    .A(net161));
 sg13g2_inv_1 _1554_ (.Y(_0622_),
    .A(net181));
 sg13g2_inv_1 _1555_ (.Y(_0623_),
    .A(net162));
 sg13g2_inv_1 _1556_ (.Y(_0624_),
    .A(net183));
 sg13g2_inv_1 _1557_ (.Y(_0625_),
    .A(\wrapper.pixel.background_state[0] ));
 sg13g2_inv_1 _1558_ (.Y(_0626_),
    .A(net156));
 sg13g2_inv_1 _1559_ (.Y(_0627_),
    .A(net177));
 sg13g2_inv_2 _1560_ (.Y(_0628_),
    .A(net579));
 sg13g2_inv_1 _1561_ (.Y(_0629_),
    .A(\wrapper.h_count[4] ));
 sg13g2_inv_1 _1562_ (.Y(_0630_),
    .A(\wrapper.pixel.prev_y[1] ));
 sg13g2_inv_1 _1563_ (.Y(_0631_),
    .A(net147));
 sg13g2_inv_1 _1564_ (.Y(_0632_),
    .A(\wrapper.pixel.prev_y[6] ));
 sg13g2_inv_1 _1565_ (.Y(_0633_),
    .A(_0007_));
 sg13g2_inv_1 _1566_ (.Y(_0634_),
    .A(\wrapper.pixel.moving_counter[4] ));
 sg13g2_inv_1 _1567_ (.Y(_0635_),
    .A(\wrapper.pixel.moving_counter[6] ));
 sg13g2_inv_1 _1568_ (.Y(_0636_),
    .A(_0019_));
 sg13g2_inv_1 _1569_ (.Y(_0637_),
    .A(_0020_));
 sg13g2_inv_1 _1570_ (.Y(_0638_),
    .A(\wrapper.pixel.rom0.color_out[1] ));
 sg13g2_nor2b_1 _1571_ (.A(\wrapper.pixel.vpos[8] ),
    .B_N(\wrapper.pixel.sprite_top[8] ),
    .Y(_0639_));
 sg13g2_xnor2_1 _1572_ (.Y(_0640_),
    .A(\wrapper.pixel.vpos[8] ),
    .B(\wrapper.pixel.sprite_top[8] ));
 sg13g2_nand2b_1 _1573_ (.Y(_0641_),
    .B(\wrapper.pixel.sprite_top[6] ),
    .A_N(net540));
 sg13g2_nand2b_1 _1574_ (.Y(_0642_),
    .B(net540),
    .A_N(\wrapper.pixel.sprite_top[6] ));
 sg13g2_inv_1 _1575_ (.Y(_0643_),
    .A(_0642_));
 sg13g2_nand2_1 _1576_ (.Y(_0644_),
    .A(_0641_),
    .B(_0642_));
 sg13g2_nand2_1 _1577_ (.Y(_0645_),
    .A(_0604_),
    .B(\wrapper.pixel.sprite_top[5] ));
 sg13g2_nor2_1 _1578_ (.A(_0604_),
    .B(\wrapper.pixel.sprite_top[5] ),
    .Y(_0646_));
 sg13g2_nor2b_1 _1579_ (.A(\wrapper.pixel.sprite_top[4] ),
    .B_N(net543),
    .Y(_0647_));
 sg13g2_nand2b_1 _1580_ (.Y(_0648_),
    .B(net544),
    .A_N(\wrapper.pixel.sprite_top[3] ));
 sg13g2_nor2b_1 _1581_ (.A(\wrapper.pixel.sprite_top[2] ),
    .B_N(net546),
    .Y(_0649_));
 sg13g2_xnor2_1 _1582_ (.Y(_0650_),
    .A(net546),
    .B(\wrapper.pixel.sprite_top[2] ));
 sg13g2_nand2_1 _1583_ (.Y(_0651_),
    .A(net548),
    .B(_0612_));
 sg13g2_xor2_1 _1584_ (.B(\wrapper.pixel.sprite_top[1] ),
    .A(net548),
    .X(_0652_));
 sg13g2_nor2_2 _1585_ (.A(net550),
    .B(_0613_),
    .Y(_0653_));
 sg13g2_o21ai_1 _1586_ (.B1(_0651_),
    .Y(_0654_),
    .A1(_0652_),
    .A2(_0653_));
 sg13g2_a21oi_2 _1587_ (.B1(_0649_),
    .Y(_0655_),
    .A2(_0654_),
    .A1(_0650_));
 sg13g2_xor2_1 _1588_ (.B(\wrapper.pixel.sprite_top[3] ),
    .A(net544),
    .X(_0656_));
 sg13g2_o21ai_1 _1589_ (.B1(_0648_),
    .Y(_0657_),
    .A1(_0655_),
    .A2(_0656_));
 sg13g2_xnor2_1 _1590_ (.Y(_0658_),
    .A(net543),
    .B(\wrapper.pixel.sprite_top[4] ));
 sg13g2_a21o_1 _1591_ (.A2(_0658_),
    .A1(_0657_),
    .B1(_0647_),
    .X(_0659_));
 sg13g2_a21o_1 _1592_ (.A2(_0659_),
    .A1(_0645_),
    .B1(_0646_),
    .X(_0660_));
 sg13g2_a221oi_1 _1593_ (.B2(_0660_),
    .C1(_0643_),
    .B1(_0641_),
    .A1(\wrapper.pixel.vpos[7] ),
    .Y(_0661_),
    .A2(_0609_));
 sg13g2_a21oi_1 _1594_ (.A1(_0603_),
    .A2(\wrapper.pixel.sprite_top[7] ),
    .Y(_0662_),
    .B1(_0661_));
 sg13g2_xnor2_1 _1595_ (.Y(_0663_),
    .A(_0640_),
    .B(_0662_));
 sg13g2_nand2b_1 _1596_ (.Y(_0664_),
    .B(\wrapper.pixel.sprite_left[8] ),
    .A_N(\wrapper.h_count[8] ));
 sg13g2_xnor2_1 _1597_ (.Y(_0665_),
    .A(\wrapper.pixel.sprite_left[8] ),
    .B(\wrapper.h_count[8] ));
 sg13g2_nor2_1 _1598_ (.A(_0614_),
    .B(net562),
    .Y(_0666_));
 sg13g2_nand2b_1 _1599_ (.Y(_0667_),
    .B(net563),
    .A_N(\wrapper.pixel.sprite_left[6] ));
 sg13g2_inv_1 _1600_ (.Y(_0668_),
    .A(_0667_));
 sg13g2_nand2b_1 _1601_ (.Y(_0669_),
    .B(\wrapper.pixel.sprite_left[6] ),
    .A_N(net563));
 sg13g2_nand2_1 _1602_ (.Y(_0670_),
    .A(_0667_),
    .B(_0669_));
 sg13g2_nor2_1 _1603_ (.A(_0615_),
    .B(net564),
    .Y(_0671_));
 sg13g2_nand2_1 _1604_ (.Y(_0672_),
    .A(_0615_),
    .B(net564));
 sg13g2_nor2_1 _1605_ (.A(\wrapper.pixel.sprite_left[4] ),
    .B(_0629_),
    .Y(_0673_));
 sg13g2_nand2b_1 _1606_ (.Y(_0674_),
    .B(\wrapper.h_count[3] ),
    .A_N(\wrapper.pixel.sprite_left[3] ));
 sg13g2_xor2_1 _1607_ (.B(\wrapper.h_count[3] ),
    .A(\wrapper.pixel.sprite_left[3] ),
    .X(_0675_));
 sg13g2_nor2b_1 _1608_ (.A(\wrapper.pixel.sprite_left[2] ),
    .B_N(net565),
    .Y(_0676_));
 sg13g2_nand2b_1 _1609_ (.Y(_0677_),
    .B(\wrapper.h_count[1] ),
    .A_N(\wrapper.pixel.sprite_left[1] ));
 sg13g2_xor2_1 _1610_ (.B(\wrapper.h_count[1] ),
    .A(\wrapper.pixel.sprite_left[1] ),
    .X(_0678_));
 sg13g2_nor2b_2 _1611_ (.A(net566),
    .B_N(\wrapper.pixel.sprite_left[0] ),
    .Y(_0679_));
 sg13g2_o21ai_1 _1612_ (.B1(_0677_),
    .Y(_0680_),
    .A1(_0678_),
    .A2(_0679_));
 sg13g2_xnor2_1 _1613_ (.Y(_0681_),
    .A(\wrapper.pixel.sprite_left[2] ),
    .B(net565));
 sg13g2_a21oi_2 _1614_ (.B1(_0676_),
    .Y(_0682_),
    .A2(_0681_),
    .A1(_0680_));
 sg13g2_o21ai_1 _1615_ (.B1(_0674_),
    .Y(_0683_),
    .A1(_0675_),
    .A2(_0682_));
 sg13g2_xnor2_1 _1616_ (.Y(_0684_),
    .A(\wrapper.pixel.sprite_left[4] ),
    .B(\wrapper.h_count[4] ));
 sg13g2_a21oi_2 _1617_ (.B1(_0673_),
    .Y(_0685_),
    .A2(_0684_),
    .A1(_0683_));
 sg13g2_o21ai_1 _1618_ (.B1(_0672_),
    .Y(_0686_),
    .A1(_0671_),
    .A2(_0685_));
 sg13g2_a221oi_1 _1619_ (.B2(_0686_),
    .C1(_0668_),
    .B1(_0669_),
    .A1(_0614_),
    .Y(_0687_),
    .A2(net561));
 sg13g2_or3_1 _1620_ (.A(_0665_),
    .B(_0666_),
    .C(_0687_),
    .X(_0688_));
 sg13g2_xnor2_1 _1621_ (.Y(_0689_),
    .A(_0670_),
    .B(_0686_));
 sg13g2_xnor2_1 _1622_ (.Y(_0690_),
    .A(_0644_),
    .B(_0660_));
 sg13g2_xor2_1 _1623_ (.B(\wrapper.pixel.sprite_top[9] ),
    .A(\wrapper.pixel.vpos[9] ),
    .X(_0691_));
 sg13g2_xnor2_1 _1624_ (.Y(_0692_),
    .A(_0639_),
    .B(_0691_));
 sg13g2_xnor2_1 _1625_ (.Y(_0693_),
    .A(\wrapper.pixel.sprite_left[9] ),
    .B(\wrapper.h_count[9] ));
 sg13g2_xnor2_1 _1626_ (.Y(_0694_),
    .A(_0664_),
    .B(_0693_));
 sg13g2_xnor2_1 _1627_ (.Y(_0695_),
    .A(\wrapper.pixel.vpos[7] ),
    .B(\wrapper.pixel.sprite_top[7] ));
 sg13g2_xnor2_1 _1628_ (.Y(_0696_),
    .A(_0641_),
    .B(_0695_));
 sg13g2_xnor2_1 _1629_ (.Y(_0697_),
    .A(\wrapper.pixel.sprite_left[7] ),
    .B(net561));
 sg13g2_xnor2_1 _1630_ (.Y(_0698_),
    .A(_0669_),
    .B(_0697_));
 sg13g2_nand4_1 _1631_ (.B(_0694_),
    .C(_0696_),
    .A(_0692_),
    .Y(_0699_),
    .D(_0698_));
 sg13g2_nor3_1 _1632_ (.A(_0689_),
    .B(_0690_),
    .C(_0699_),
    .Y(_0700_));
 sg13g2_o21ai_1 _1633_ (.B1(_0665_),
    .Y(_0701_),
    .A1(_0666_),
    .A2(_0687_));
 sg13g2_and4_2 _1634_ (.A(_0663_),
    .B(_0688_),
    .C(_0700_),
    .D(_0701_),
    .X(_0702_));
 sg13g2_inv_1 _1635_ (.Y(_0703_),
    .A(_0702_));
 sg13g2_nor2_2 _1636_ (.A(net560),
    .B(\wrapper.pixel.background_state[0] ),
    .Y(_0704_));
 sg13g2_nor2_2 _1637_ (.A(\wrapper.pixel.background_state[3] ),
    .B(\wrapper.pixel.background_state[2] ),
    .Y(_0705_));
 sg13g2_and2_2 _1638_ (.A(_0704_),
    .B(_0705_),
    .X(_0706_));
 sg13g2_nand2_2 _1639_ (.Y(_0707_),
    .A(_0704_),
    .B(_0705_));
 sg13g2_nand2_1 _1640_ (.Y(_0708_),
    .A(_0620_),
    .B(_0706_));
 sg13g2_nand2_2 _1641_ (.Y(_0709_),
    .A(net560),
    .B(\wrapper.pixel.background_state[0] ));
 sg13g2_nand2_2 _1642_ (.Y(_0710_),
    .A(net558),
    .B(net559));
 sg13g2_nor2_2 _1643_ (.A(_0709_),
    .B(_0710_),
    .Y(_0711_));
 sg13g2_nor2b_1 _1644_ (.A(\wrapper.pixel.background_state[0] ),
    .B_N(net560),
    .Y(_0712_));
 sg13g2_nand2b_1 _1645_ (.Y(_0713_),
    .B(net560),
    .A_N(\wrapper.pixel.background_state[0] ));
 sg13g2_nor2_2 _1646_ (.A(_0710_),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_nor2_1 _1647_ (.A(net560),
    .B(_0625_),
    .Y(_0715_));
 sg13g2_nand2b_2 _1648_ (.Y(_0716_),
    .B(\wrapper.pixel.background_state[0] ),
    .A_N(net560));
 sg13g2_nor2b_1 _1649_ (.A(net559),
    .B_N(net558),
    .Y(_0717_));
 sg13g2_nand2b_1 _1650_ (.Y(_0718_),
    .B(net558),
    .A_N(net559));
 sg13g2_nor2b_2 _1651_ (.A(net558),
    .B_N(net559),
    .Y(_0719_));
 sg13g2_nand3b_1 _1652_ (.B(net559),
    .C(net560),
    .Y(_0720_),
    .A_N(net558));
 sg13g2_a22oi_1 _1653_ (.Y(_0721_),
    .B1(_0718_),
    .B2(_0720_),
    .A2(_0716_),
    .A1(_0713_));
 sg13g2_nor2_1 _1654_ (.A(\wrapper.pixel.moving_counter[0] ),
    .B(\wrapper.pixel.moving_counter[1] ),
    .Y(_0722_));
 sg13g2_nor3_1 _1655_ (.A(\wrapper.pixel.moving_counter[2] ),
    .B(\wrapper.pixel.moving_counter[0] ),
    .C(\wrapper.pixel.moving_counter[1] ),
    .Y(_0723_));
 sg13g2_nor2b_1 _1656_ (.A(\wrapper.pixel.moving_counter[3] ),
    .B_N(_0723_),
    .Y(_0724_));
 sg13g2_nand2_1 _1657_ (.Y(_0725_),
    .A(_0634_),
    .B(_0724_));
 sg13g2_xnor2_1 _1658_ (.Y(_0726_),
    .A(\wrapper.pixel.moving_counter[4] ),
    .B(_0724_));
 sg13g2_nand2_1 _1659_ (.Y(_0727_),
    .A(_0009_),
    .B(net525));
 sg13g2_o21ai_1 _1660_ (.B1(_0727_),
    .Y(_0728_),
    .A1(net524),
    .A2(_0726_));
 sg13g2_and2_1 _1661_ (.A(\wrapper.pixel.vpos[4] ),
    .B(_0728_),
    .X(_0729_));
 sg13g2_xnor2_1 _1662_ (.Y(_0730_),
    .A(net543),
    .B(_0728_));
 sg13g2_xnor2_1 _1663_ (.Y(_0731_),
    .A(\wrapper.pixel.moving_counter[3] ),
    .B(_0723_));
 sg13g2_nand2_1 _1664_ (.Y(_0732_),
    .A(_0010_),
    .B(net524));
 sg13g2_o21ai_1 _1665_ (.B1(_0732_),
    .Y(_0733_),
    .A1(net524),
    .A2(_0731_));
 sg13g2_nor2_1 _1666_ (.A(net545),
    .B(_0733_),
    .Y(_0734_));
 sg13g2_xnor2_1 _1667_ (.Y(_0735_),
    .A(\wrapper.pixel.moving_counter[2] ),
    .B(_0722_));
 sg13g2_nand2_1 _1668_ (.Y(_0736_),
    .A(_0011_),
    .B(net524));
 sg13g2_o21ai_1 _1669_ (.B1(_0736_),
    .Y(_0737_),
    .A1(net524),
    .A2(_0735_));
 sg13g2_and2_1 _1670_ (.A(net547),
    .B(_0737_),
    .X(_0738_));
 sg13g2_nand2_1 _1671_ (.Y(_0739_),
    .A(\wrapper.pixel.moving_counter[0] ),
    .B(\wrapper.pixel.moving_counter[1] ));
 sg13g2_nand2b_1 _1672_ (.Y(_0740_),
    .B(_0739_),
    .A_N(_0722_));
 sg13g2_mux2_1 _1673_ (.A0(_0740_),
    .A1(_0012_),
    .S(net524),
    .X(_0741_));
 sg13g2_nand2_1 _1674_ (.Y(_0742_),
    .A(net549),
    .B(_0741_));
 sg13g2_nor2b_1 _1675_ (.A(net551),
    .B_N(\wrapper.pixel.moving_counter[0] ),
    .Y(_0743_));
 sg13g2_xnor2_1 _1676_ (.Y(_0744_),
    .A(net549),
    .B(_0741_));
 sg13g2_o21ai_1 _1677_ (.B1(_0742_),
    .Y(_0745_),
    .A1(_0743_),
    .A2(_0744_));
 sg13g2_xor2_1 _1678_ (.B(_0737_),
    .A(net547),
    .X(_0746_));
 sg13g2_a21oi_1 _1679_ (.A1(_0745_),
    .A2(_0746_),
    .Y(_0747_),
    .B1(_0738_));
 sg13g2_a221oi_1 _1680_ (.B2(_0746_),
    .C1(_0738_),
    .B1(_0745_),
    .A1(net545),
    .Y(_0748_),
    .A2(_0733_));
 sg13g2_nor3_2 _1681_ (.A(_0730_),
    .B(_0734_),
    .C(_0748_),
    .Y(_0749_));
 sg13g2_o21ai_1 _1682_ (.B1(_0730_),
    .Y(_0750_),
    .A1(_0734_),
    .A2(_0748_));
 sg13g2_nand2b_1 _1683_ (.Y(_0751_),
    .B(_0750_),
    .A_N(_0749_));
 sg13g2_a22oi_1 _1684_ (.Y(_0752_),
    .B1(_0719_),
    .B2(_0704_),
    .A2(_0717_),
    .A1(_0625_));
 sg13g2_nor2_1 _1685_ (.A(_0010_),
    .B(net522),
    .Y(_0753_));
 sg13g2_a21oi_2 _1686_ (.B1(_0753_),
    .Y(_0754_),
    .A2(net522),
    .A1(_0731_));
 sg13g2_nor2_1 _1687_ (.A(\wrapper.h_count[3] ),
    .B(_0754_),
    .Y(_0755_));
 sg13g2_nor2_1 _1688_ (.A(_0011_),
    .B(net522),
    .Y(_0756_));
 sg13g2_a21oi_1 _1689_ (.A1(_0735_),
    .A2(net522),
    .Y(_0757_),
    .B1(_0756_));
 sg13g2_and2_1 _1690_ (.A(\wrapper.h_count[2] ),
    .B(_0757_),
    .X(_0758_));
 sg13g2_mux2_1 _1691_ (.A0(_0012_),
    .A1(_0740_),
    .S(net522),
    .X(_0759_));
 sg13g2_nand2_1 _1692_ (.Y(_0760_),
    .A(\wrapper.h_count[1] ),
    .B(_0759_));
 sg13g2_nor2b_1 _1693_ (.A(\wrapper.h_count[0] ),
    .B_N(\wrapper.pixel.moving_counter[0] ),
    .Y(_0761_));
 sg13g2_xnor2_1 _1694_ (.Y(_0762_),
    .A(\wrapper.h_count[1] ),
    .B(_0759_));
 sg13g2_o21ai_1 _1695_ (.B1(_0760_),
    .Y(_0763_),
    .A1(_0761_),
    .A2(_0762_));
 sg13g2_xor2_1 _1696_ (.B(_0757_),
    .A(net565),
    .X(_0764_));
 sg13g2_a21oi_1 _1697_ (.A1(_0763_),
    .A2(_0764_),
    .Y(_0765_),
    .B1(_0758_));
 sg13g2_a221oi_1 _1698_ (.B2(_0764_),
    .C1(_0758_),
    .B1(_0763_),
    .A1(\wrapper.h_count[3] ),
    .Y(_0766_),
    .A2(_0754_));
 sg13g2_nor2_1 _1699_ (.A(_0009_),
    .B(net522),
    .Y(_0767_));
 sg13g2_a21oi_1 _1700_ (.A1(_0726_),
    .A2(net523),
    .Y(_0768_),
    .B1(_0767_));
 sg13g2_xor2_1 _1701_ (.B(_0768_),
    .A(_0008_),
    .X(_0769_));
 sg13g2_nor3_2 _1702_ (.A(_0755_),
    .B(_0766_),
    .C(_0769_),
    .Y(_0770_));
 sg13g2_o21ai_1 _1703_ (.B1(_0769_),
    .Y(_0771_),
    .A1(_0755_),
    .A2(_0766_));
 sg13g2_nand2b_1 _1704_ (.Y(_0772_),
    .B(_0771_),
    .A_N(_0770_));
 sg13g2_nand3b_1 _1705_ (.B(_0751_),
    .C(_0772_),
    .Y(_0773_),
    .A_N(net543));
 sg13g2_a21oi_1 _1706_ (.A1(_0714_),
    .A2(_0773_),
    .Y(_0774_),
    .B1(_0711_));
 sg13g2_or2_1 _1707_ (.X(_0775_),
    .B(_0772_),
    .A(_0751_));
 sg13g2_nand3_1 _1708_ (.B(_0751_),
    .C(_0772_),
    .A(_0714_),
    .Y(_0776_));
 sg13g2_nand3_1 _1709_ (.B(_0775_),
    .C(_0776_),
    .A(net543),
    .Y(_0777_));
 sg13g2_o21ai_1 _1710_ (.B1(_0777_),
    .Y(_0778_),
    .A1(net543),
    .A2(_0775_));
 sg13g2_xnor2_1 _1711_ (.Y(_0779_),
    .A(_0763_),
    .B(_0764_));
 sg13g2_nand2_1 _1712_ (.Y(_0780_),
    .A(_0709_),
    .B(_0718_));
 sg13g2_o21ai_1 _1713_ (.B1(_0780_),
    .Y(_0781_),
    .A1(_0709_),
    .A2(_0719_));
 sg13g2_nor3_1 _1714_ (.A(net558),
    .B(net559),
    .C(_0709_),
    .Y(_0782_));
 sg13g2_a21o_1 _1715_ (.A2(_0719_),
    .A1(_0704_),
    .B1(_0782_),
    .X(_0783_));
 sg13g2_o21ai_1 _1716_ (.B1(_0719_),
    .Y(_0784_),
    .A1(_0712_),
    .A2(_0715_));
 sg13g2_nor2b_1 _1717_ (.A(_0783_),
    .B_N(_0784_),
    .Y(_0785_));
 sg13g2_nor3_2 _1718_ (.A(net558),
    .B(net559),
    .C(_0716_),
    .Y(_0786_));
 sg13g2_nand2_2 _1719_ (.Y(_0787_),
    .A(_0705_),
    .B(_0712_));
 sg13g2_inv_1 _1720_ (.Y(_0788_),
    .A(_0787_));
 sg13g2_o21ai_1 _1721_ (.B1(_0707_),
    .Y(_0789_),
    .A1(_0013_),
    .A2(_0785_));
 sg13g2_a221oi_1 _1722_ (.B2(\wrapper.h_count[1] ),
    .C1(_0789_),
    .B1(_0788_),
    .A1(net549),
    .Y(_0790_),
    .A2(_0786_));
 sg13g2_o21ai_1 _1723_ (.B1(_0790_),
    .Y(_0791_),
    .A1(_0779_),
    .A2(_0781_));
 sg13g2_inv_1 _1724_ (.Y(_0792_),
    .A(_0791_));
 sg13g2_nor3_1 _1725_ (.A(net560),
    .B(\wrapper.pixel.background_state[0] ),
    .C(_0710_),
    .Y(_0793_));
 sg13g2_nand3_1 _1726_ (.B(net559),
    .C(_0704_),
    .A(net558),
    .Y(_0794_));
 sg13g2_xor2_1 _1727_ (.B(\wrapper.h_count[4] ),
    .A(net543),
    .X(_0795_));
 sg13g2_xnor2_1 _1728_ (.Y(_0796_),
    .A(\wrapper.pixel.lfsr_reg[14] ),
    .B(_0795_));
 sg13g2_nor2_2 _1729_ (.A(_0709_),
    .B(_0718_),
    .Y(_0797_));
 sg13g2_nor2_2 _1730_ (.A(_0710_),
    .B(_0716_),
    .Y(_0798_));
 sg13g2_a22oi_1 _1731_ (.Y(_0799_),
    .B1(_0798_),
    .B2(_0795_),
    .A2(_0797_),
    .A1(\wrapper.pixel.lfsr_reg[14] ));
 sg13g2_o21ai_1 _1732_ (.B1(_0799_),
    .Y(_0800_),
    .A1(_0794_),
    .A2(_0796_));
 sg13g2_nor2_1 _1733_ (.A(_0791_),
    .B(_0800_),
    .Y(_0801_));
 sg13g2_o21ai_1 _1734_ (.B1(_0801_),
    .Y(_0802_),
    .A1(_0774_),
    .A2(_0778_));
 sg13g2_a21oi_1 _1735_ (.A1(_0708_),
    .A2(_0802_),
    .Y(_0803_),
    .B1(_0702_));
 sg13g2_nor2_1 _1736_ (.A(_0603_),
    .B(_0604_),
    .Y(_0804_));
 sg13g2_nand3_1 _1737_ (.B(net540),
    .C(_0804_),
    .A(\wrapper.pixel.vpos[8] ),
    .Y(_0805_));
 sg13g2_o21ai_1 _1738_ (.B1(_0633_),
    .Y(_0806_),
    .A1(net561),
    .A2(\wrapper.h_count[8] ));
 sg13g2_nand3_1 _1739_ (.B(_0805_),
    .C(_0806_),
    .A(_0601_),
    .Y(_0807_));
 sg13g2_nor2_1 _1740_ (.A(\wrapper.pixel.rom0.color_out[4] ),
    .B(_0703_),
    .Y(_0808_));
 sg13g2_nor3_2 _1741_ (.A(_0803_),
    .B(_0807_),
    .C(_0808_),
    .Y(uo_out[4]));
 sg13g2_and2_1 _1742_ (.A(\wrapper.h_count[4] ),
    .B(_0768_),
    .X(_0809_));
 sg13g2_nor2_1 _1743_ (.A(_0015_),
    .B(net523),
    .Y(_0810_));
 sg13g2_xor2_1 _1744_ (.B(_0725_),
    .A(\wrapper.pixel.moving_counter[5] ),
    .X(_0811_));
 sg13g2_a21oi_1 _1745_ (.A1(net522),
    .A2(_0811_),
    .Y(_0812_),
    .B1(_0810_));
 sg13g2_xnor2_1 _1746_ (.Y(_0813_),
    .A(_0014_),
    .B(_0812_));
 sg13g2_o21ai_1 _1747_ (.B1(_0813_),
    .Y(_0814_),
    .A1(_0770_),
    .A2(_0809_));
 sg13g2_or3_1 _1748_ (.A(_0770_),
    .B(_0809_),
    .C(_0813_),
    .X(_0815_));
 sg13g2_and2_1 _1749_ (.A(_0814_),
    .B(_0815_),
    .X(_0816_));
 sg13g2_nor2_1 _1750_ (.A(_0729_),
    .B(_0749_),
    .Y(_0817_));
 sg13g2_nand2_1 _1751_ (.Y(_0818_),
    .A(_0015_),
    .B(net525));
 sg13g2_o21ai_1 _1752_ (.B1(_0818_),
    .Y(_0819_),
    .A1(net525),
    .A2(_0811_));
 sg13g2_nand2_1 _1753_ (.Y(_0820_),
    .A(\wrapper.pixel.vpos[5] ),
    .B(_0819_));
 sg13g2_xnor2_1 _1754_ (.Y(_0821_),
    .A(net541),
    .B(_0819_));
 sg13g2_inv_1 _1755_ (.Y(_0822_),
    .A(_0821_));
 sg13g2_o21ai_1 _1756_ (.B1(_0822_),
    .Y(_0823_),
    .A1(_0729_),
    .A2(_0749_));
 sg13g2_xnor2_1 _1757_ (.Y(_0824_),
    .A(_0817_),
    .B(_0822_));
 sg13g2_nand2_1 _1758_ (.Y(_0825_),
    .A(_0816_),
    .B(_0824_));
 sg13g2_xor2_1 _1759_ (.B(_0824_),
    .A(_0816_),
    .X(_0826_));
 sg13g2_xnor2_1 _1760_ (.Y(_0827_),
    .A(_0604_),
    .B(_0826_));
 sg13g2_xnor2_1 _1761_ (.Y(_0828_),
    .A(_0604_),
    .B(_0825_));
 sg13g2_nand2_1 _1762_ (.Y(_0829_),
    .A(_0781_),
    .B(_0784_));
 sg13g2_xor2_1 _1763_ (.B(\wrapper.h_count[5] ),
    .A(net541),
    .X(_0830_));
 sg13g2_xor2_1 _1764_ (.B(_0830_),
    .A(\wrapper.pixel.lfsr_reg[15] ),
    .X(_0831_));
 sg13g2_nand2b_1 _1765_ (.Y(_0832_),
    .B(_0786_),
    .A_N(_0014_));
 sg13g2_nand2_1 _1766_ (.Y(_0833_),
    .A(_0783_),
    .B(_0816_));
 sg13g2_a221oi_1 _1767_ (.B2(_0830_),
    .C1(_0706_),
    .B1(_0798_),
    .A1(\wrapper.pixel.lfsr_reg[15] ),
    .Y(_0834_),
    .A2(_0797_));
 sg13g2_o21ai_1 _1768_ (.B1(_0832_),
    .Y(_0835_),
    .A1(_0016_),
    .A2(_0787_));
 sg13g2_a221oi_1 _1769_ (.B2(_0793_),
    .C1(_0835_),
    .B1(_0831_),
    .A1(_0824_),
    .Y(_0836_),
    .A2(_0829_));
 sg13g2_nand3_1 _1770_ (.B(_0834_),
    .C(_0836_),
    .A(_0833_),
    .Y(_0837_));
 sg13g2_a221oi_1 _1771_ (.B2(_0711_),
    .C1(_0837_),
    .B1(_0828_),
    .A1(_0714_),
    .Y(_0838_),
    .A2(_0827_));
 sg13g2_a21oi_1 _1772_ (.A1(_0619_),
    .A2(_0706_),
    .Y(_0839_),
    .B1(_0702_));
 sg13g2_nand2b_1 _1773_ (.Y(_0840_),
    .B(_0839_),
    .A_N(_0838_));
 sg13g2_nand2_1 _1774_ (.Y(_0841_),
    .A(\wrapper.pixel.rom0.color_out[5] ),
    .B(_0702_));
 sg13g2_a21oi_2 _1775_ (.B1(_0807_),
    .Y(uo_out[0]),
    .A2(_0841_),
    .A1(_0840_));
 sg13g2_xnor2_1 _1776_ (.Y(_0842_),
    .A(_0745_),
    .B(_0746_));
 sg13g2_nand3b_1 _1777_ (.B(_0779_),
    .C(_0842_),
    .Y(_0843_),
    .A_N(net547));
 sg13g2_a21oi_1 _1778_ (.A1(_0714_),
    .A2(_0843_),
    .Y(_0844_),
    .B1(_0711_));
 sg13g2_nor3_1 _1779_ (.A(net547),
    .B(_0779_),
    .C(_0842_),
    .Y(_0845_));
 sg13g2_nand3_1 _1780_ (.B(_0779_),
    .C(_0842_),
    .A(_0714_),
    .Y(_0846_));
 sg13g2_o21ai_1 _1781_ (.B1(net547),
    .Y(_0847_),
    .A1(_0779_),
    .A2(_0842_));
 sg13g2_nor2b_1 _1782_ (.A(_0847_),
    .B_N(_0846_),
    .Y(_0848_));
 sg13g2_nor3_2 _1783_ (.A(_0844_),
    .B(_0845_),
    .C(_0848_),
    .Y(_0849_));
 sg13g2_xor2_1 _1784_ (.B(net565),
    .A(net547),
    .X(_0850_));
 sg13g2_xnor2_1 _1785_ (.Y(_0851_),
    .A(\wrapper.pixel.lfsr_reg[12] ),
    .B(_0850_));
 sg13g2_a22oi_1 _1786_ (.Y(_0852_),
    .B1(_0798_),
    .B2(_0850_),
    .A2(_0797_),
    .A1(\wrapper.pixel.lfsr_reg[12] ));
 sg13g2_o21ai_1 _1787_ (.B1(_0852_),
    .Y(_0853_),
    .A1(_0794_),
    .A2(_0851_));
 sg13g2_nor2_1 _1788_ (.A(_0849_),
    .B(_0853_),
    .Y(_0854_));
 sg13g2_a22oi_1 _1789_ (.Y(_0855_),
    .B1(_0792_),
    .B2(_0854_),
    .A2(_0706_),
    .A1(_0622_));
 sg13g2_nand2_1 _1790_ (.Y(_0856_),
    .A(_0703_),
    .B(_0855_));
 sg13g2_nand2_1 _1791_ (.Y(_0857_),
    .A(\wrapper.pixel.rom0.color_out[2] ),
    .B(_0702_));
 sg13g2_a21oi_2 _1792_ (.B1(_0807_),
    .Y(uo_out[5]),
    .A2(_0857_),
    .A1(_0856_));
 sg13g2_nand2_1 _1793_ (.Y(_0858_),
    .A(_0621_),
    .B(_0706_));
 sg13g2_nor3_1 _1794_ (.A(\wrapper.pixel.moving_counter[5] ),
    .B(\wrapper.pixel.moving_counter[6] ),
    .C(_0725_),
    .Y(_0859_));
 sg13g2_o21ai_1 _1795_ (.B1(\wrapper.pixel.moving_counter[6] ),
    .Y(_0860_),
    .A1(\wrapper.pixel.moving_counter[5] ),
    .A2(_0725_));
 sg13g2_nor2b_1 _1796_ (.A(_0859_),
    .B_N(_0860_),
    .Y(_0861_));
 sg13g2_nand2_1 _1797_ (.Y(_0862_),
    .A(_0017_),
    .B(net525));
 sg13g2_o21ai_1 _1798_ (.B1(_0862_),
    .Y(_0863_),
    .A1(net525),
    .A2(_0861_));
 sg13g2_nand2_1 _1799_ (.Y(_0864_),
    .A(\wrapper.pixel.vpos[6] ),
    .B(_0863_));
 sg13g2_xnor2_1 _1800_ (.Y(_0865_),
    .A(\wrapper.pixel.vpos[6] ),
    .B(_0863_));
 sg13g2_a21o_1 _1801_ (.A2(_0823_),
    .A1(_0820_),
    .B1(_0865_),
    .X(_0866_));
 sg13g2_nand3_1 _1802_ (.B(_0823_),
    .C(_0865_),
    .A(_0820_),
    .Y(_0867_));
 sg13g2_nand3_1 _1803_ (.B(_0866_),
    .C(_0867_),
    .A(_0829_),
    .Y(_0868_));
 sg13g2_xnor2_1 _1804_ (.Y(_0869_),
    .A(net545),
    .B(_0733_));
 sg13g2_xnor2_1 _1805_ (.Y(_0870_),
    .A(_0747_),
    .B(_0869_));
 sg13g2_xnor2_1 _1806_ (.Y(_0871_),
    .A(\wrapper.h_count[3] ),
    .B(_0754_));
 sg13g2_xnor2_1 _1807_ (.Y(_0872_),
    .A(_0765_),
    .B(_0871_));
 sg13g2_nor2_1 _1808_ (.A(_0870_),
    .B(_0872_),
    .Y(_0873_));
 sg13g2_xnor2_1 _1809_ (.Y(_0874_),
    .A(net545),
    .B(_0873_));
 sg13g2_xor2_1 _1810_ (.B(_0872_),
    .A(_0870_),
    .X(_0875_));
 sg13g2_xnor2_1 _1811_ (.Y(_0876_),
    .A(_0605_),
    .B(_0875_));
 sg13g2_xnor2_1 _1812_ (.Y(_0877_),
    .A(net544),
    .B(\wrapper.h_count[3] ));
 sg13g2_xor2_1 _1813_ (.B(_0877_),
    .A(\wrapper.pixel.lfsr_reg[13] ),
    .X(_0878_));
 sg13g2_nor3_1 _1814_ (.A(_0710_),
    .B(_0716_),
    .C(_0877_),
    .Y(_0879_));
 sg13g2_o21ai_1 _1815_ (.B1(_0707_),
    .Y(_0880_),
    .A1(_0018_),
    .A2(_0787_));
 sg13g2_nor2_1 _1816_ (.A(_0879_),
    .B(_0880_),
    .Y(_0881_));
 sg13g2_o21ai_1 _1817_ (.B1(_0881_),
    .Y(_0882_),
    .A1(_0794_),
    .A2(_0878_));
 sg13g2_a221oi_1 _1818_ (.B2(\wrapper.pixel.lfsr_reg[13] ),
    .C1(_0882_),
    .B1(_0797_),
    .A1(_0636_),
    .Y(_0883_),
    .A2(_0786_));
 sg13g2_a22oi_1 _1819_ (.Y(_0884_),
    .B1(_0876_),
    .B2(_0714_),
    .A2(_0874_),
    .A1(_0711_));
 sg13g2_nand2_1 _1820_ (.Y(_0885_),
    .A(net564),
    .B(_0812_));
 sg13g2_nor2_1 _1821_ (.A(_0017_),
    .B(net523),
    .Y(_0886_));
 sg13g2_a21oi_2 _1822_ (.B1(_0886_),
    .Y(_0887_),
    .A2(_0861_),
    .A1(net522));
 sg13g2_nand2_1 _1823_ (.Y(_0888_),
    .A(\wrapper.h_count[6] ),
    .B(_0887_));
 sg13g2_xnor2_1 _1824_ (.Y(_0889_),
    .A(net563),
    .B(_0887_));
 sg13g2_nand3_1 _1825_ (.B(_0885_),
    .C(_0889_),
    .A(_0814_),
    .Y(_0890_));
 sg13g2_a21o_1 _1826_ (.A2(_0885_),
    .A1(_0814_),
    .B1(_0889_),
    .X(_0891_));
 sg13g2_nand3_1 _1827_ (.B(_0890_),
    .C(_0891_),
    .A(_0783_),
    .Y(_0892_));
 sg13g2_nand4_1 _1828_ (.B(_0883_),
    .C(_0884_),
    .A(_0868_),
    .Y(_0893_),
    .D(_0892_));
 sg13g2_a21oi_1 _1829_ (.A1(_0858_),
    .A2(_0893_),
    .Y(_0894_),
    .B1(_0702_));
 sg13g2_nor2_1 _1830_ (.A(\wrapper.pixel.rom0.color_out[3] ),
    .B(_0703_),
    .Y(_0895_));
 sg13g2_nor3_2 _1831_ (.A(_0807_),
    .B(_0894_),
    .C(_0895_),
    .Y(uo_out[1]));
 sg13g2_nand2_1 _1832_ (.Y(_0896_),
    .A(_0606_),
    .B(\wrapper.h_count[0] ));
 sg13g2_xor2_1 _1833_ (.B(net566),
    .A(net550),
    .X(_0897_));
 sg13g2_xnor2_1 _1834_ (.Y(_0898_),
    .A(\wrapper.pixel.lfsr_reg[10] ),
    .B(_0897_));
 sg13g2_o21ai_1 _1835_ (.B1(_0711_),
    .Y(_0899_),
    .A1(_0606_),
    .A2(net566));
 sg13g2_a21oi_2 _1836_ (.B1(_0899_),
    .Y(_0900_),
    .A2(_0896_),
    .A1(\wrapper.pixel.moving_counter[0] ));
 sg13g2_a221oi_1 _1837_ (.B2(_0637_),
    .C1(_0900_),
    .B1(_0797_),
    .A1(net566),
    .Y(_0901_),
    .A2(_0714_));
 sg13g2_o21ai_1 _1838_ (.B1(_0901_),
    .Y(_0902_),
    .A1(_0794_),
    .A2(_0898_));
 sg13g2_a21oi_1 _1839_ (.A1(_0798_),
    .A2(_0897_),
    .Y(_0903_),
    .B1(_0902_));
 sg13g2_a22oi_1 _1840_ (.Y(_0904_),
    .B1(_0792_),
    .B2(_0903_),
    .A2(_0706_),
    .A1(_0624_));
 sg13g2_mux2_1 _1841_ (.A0(_0904_),
    .A1(\wrapper.pixel.rom0.color_out[0] ),
    .S(_0702_),
    .X(_0905_));
 sg13g2_nor2b_2 _1842_ (.A(_0807_),
    .B_N(_0905_),
    .Y(uo_out[6]));
 sg13g2_nand2_1 _1843_ (.Y(_0906_),
    .A(_0864_),
    .B(_0866_));
 sg13g2_xnor2_1 _1844_ (.Y(_0907_),
    .A(\wrapper.pixel.moving_counter[7] ),
    .B(_0859_));
 sg13g2_nand2_1 _1845_ (.Y(_0908_),
    .A(_0021_),
    .B(net524));
 sg13g2_o21ai_1 _1846_ (.B1(_0908_),
    .Y(_0909_),
    .A1(net524),
    .A2(_0907_));
 sg13g2_xnor2_1 _1847_ (.Y(_0910_),
    .A(\wrapper.pixel.vpos[7] ),
    .B(_0909_));
 sg13g2_xnor2_1 _1848_ (.Y(_0911_),
    .A(_0906_),
    .B(_0910_));
 sg13g2_nand2_1 _1849_ (.Y(_0912_),
    .A(_0888_),
    .B(_0891_));
 sg13g2_nor2_1 _1850_ (.A(_0021_),
    .B(net523),
    .Y(_0913_));
 sg13g2_a21oi_1 _1851_ (.A1(net523),
    .A2(_0907_),
    .Y(_0914_),
    .B1(_0913_));
 sg13g2_xnor2_1 _1852_ (.Y(_0915_),
    .A(net562),
    .B(_0914_));
 sg13g2_xnor2_1 _1853_ (.Y(_0916_),
    .A(_0912_),
    .B(_0915_));
 sg13g2_xor2_1 _1854_ (.B(_0744_),
    .A(_0743_),
    .X(_0917_));
 sg13g2_xor2_1 _1855_ (.B(_0762_),
    .A(_0761_),
    .X(_0918_));
 sg13g2_nand2_1 _1856_ (.Y(_0919_),
    .A(_0917_),
    .B(_0918_));
 sg13g2_xnor2_1 _1857_ (.Y(_0920_),
    .A(_0917_),
    .B(_0918_));
 sg13g2_xnor2_1 _1858_ (.Y(_0921_),
    .A(net549),
    .B(_0920_));
 sg13g2_xor2_1 _1859_ (.B(\wrapper.h_count[1] ),
    .A(net549),
    .X(_0922_));
 sg13g2_xor2_1 _1860_ (.B(_0922_),
    .A(\wrapper.pixel.lfsr_reg[11] ),
    .X(_0923_));
 sg13g2_a21oi_1 _1861_ (.A1(_0798_),
    .A2(_0922_),
    .Y(_0924_),
    .B1(_0706_));
 sg13g2_a22oi_1 _1862_ (.Y(_0925_),
    .B1(_0797_),
    .B2(\wrapper.pixel.lfsr_reg[11] ),
    .A2(_0786_),
    .A1(net562));
 sg13g2_o21ai_1 _1863_ (.B1(_0925_),
    .Y(_0926_),
    .A1(_0022_),
    .A2(_0787_));
 sg13g2_a21oi_1 _1864_ (.A1(_0793_),
    .A2(_0923_),
    .Y(_0927_),
    .B1(_0926_));
 sg13g2_xor2_1 _1865_ (.B(_0919_),
    .A(net549),
    .X(_0928_));
 sg13g2_a22oi_1 _1866_ (.Y(_0929_),
    .B1(_0928_),
    .B2(_0711_),
    .A2(_0921_),
    .A1(_0714_));
 sg13g2_nand3_1 _1867_ (.B(_0927_),
    .C(_0929_),
    .A(_0924_),
    .Y(_0930_));
 sg13g2_a221oi_1 _1868_ (.B2(_0783_),
    .C1(_0930_),
    .B1(_0916_),
    .A1(_0829_),
    .Y(_0931_),
    .A2(_0911_));
 sg13g2_nor2_1 _1869_ (.A(\wrapper.pixel.solid_color[1] ),
    .B(_0707_),
    .Y(_0932_));
 sg13g2_o21ai_1 _1870_ (.B1(_0703_),
    .Y(_0933_),
    .A1(_0931_),
    .A2(_0932_));
 sg13g2_a21oi_1 _1871_ (.A1(_0638_),
    .A2(_0702_),
    .Y(_0934_),
    .B1(_0807_));
 sg13g2_and2_2 _1872_ (.A(_0933_),
    .B(_0934_),
    .X(uo_out[2]));
 sg13g2_xnor2_1 _1873_ (.Y(_0935_),
    .A(_0657_),
    .B(_0658_));
 sg13g2_inv_2 _1874_ (.Y(_0936_),
    .A(net458));
 sg13g2_xor2_1 _1875_ (.B(_0684_),
    .A(_0683_),
    .X(_0937_));
 sg13g2_xnor2_1 _1876_ (.Y(_0938_),
    .A(_0683_),
    .B(_0684_));
 sg13g2_xor2_1 _1877_ (.B(_0682_),
    .A(_0675_),
    .X(_0939_));
 sg13g2_xnor2_1 _1878_ (.Y(_0940_),
    .A(_0675_),
    .B(_0682_));
 sg13g2_nor2_2 _1879_ (.A(net476),
    .B(net501),
    .Y(_0941_));
 sg13g2_nand2_1 _1880_ (.Y(_0942_),
    .A(net469),
    .B(net495));
 sg13g2_nor2b_1 _1881_ (.A(_0671_),
    .B_N(_0672_),
    .Y(_0943_));
 sg13g2_xnor2_1 _1882_ (.Y(_0944_),
    .A(_0685_),
    .B(_0943_));
 sg13g2_xor2_1 _1883_ (.B(_0943_),
    .A(_0685_),
    .X(_0945_));
 sg13g2_xor2_1 _1884_ (.B(_0679_),
    .A(_0678_),
    .X(_0946_));
 sg13g2_xnor2_1 _1885_ (.Y(_0947_),
    .A(_0678_),
    .B(_0679_));
 sg13g2_xnor2_1 _1886_ (.Y(_0948_),
    .A(\wrapper.pixel.sprite_left[0] ),
    .B(net566));
 sg13g2_xor2_1 _1887_ (.B(net566),
    .A(\wrapper.pixel.sprite_left[0] ),
    .X(_0949_));
 sg13g2_xor2_1 _1888_ (.B(_0681_),
    .A(_0680_),
    .X(_0950_));
 sg13g2_xnor2_1 _1889_ (.Y(_0951_),
    .A(_0680_),
    .B(_0681_));
 sg13g2_nand2_2 _1890_ (.Y(_0952_),
    .A(net538),
    .B(net519));
 sg13g2_nor2_2 _1891_ (.A(_0946_),
    .B(_0948_),
    .Y(_0953_));
 sg13g2_nand2_2 _1892_ (.Y(_0954_),
    .A(_0947_),
    .B(net538));
 sg13g2_nor2_1 _1893_ (.A(net517),
    .B(_0954_),
    .Y(_0955_));
 sg13g2_nand2_2 _1894_ (.Y(_0956_),
    .A(_0950_),
    .B(_0953_));
 sg13g2_nand2_2 _1895_ (.Y(_0957_),
    .A(net469),
    .B(_0956_));
 sg13g2_nand3_1 _1896_ (.B(net446),
    .C(_0957_),
    .A(_0942_),
    .Y(_0958_));
 sg13g2_and2_2 _1897_ (.A(_0678_),
    .B(_0948_),
    .X(_0959_));
 sg13g2_nand2_2 _1898_ (.Y(_0960_),
    .A(_0678_),
    .B(_0948_));
 sg13g2_nor2_2 _1899_ (.A(net494),
    .B(net516),
    .Y(_0961_));
 sg13g2_nand2_2 _1900_ (.Y(_0962_),
    .A(net502),
    .B(net520));
 sg13g2_nor2_1 _1901_ (.A(net518),
    .B(_0960_),
    .Y(_0963_));
 sg13g2_nand2_2 _1902_ (.Y(_0964_),
    .A(net519),
    .B(_0959_));
 sg13g2_nand2_1 _1903_ (.Y(_0965_),
    .A(net505),
    .B(_0963_));
 sg13g2_a21oi_1 _1904_ (.A1(net479),
    .A2(_0965_),
    .Y(_0966_),
    .B1(_0958_));
 sg13g2_nor2_2 _1905_ (.A(net538),
    .B(net519),
    .Y(_0967_));
 sg13g2_nor2_2 _1906_ (.A(_0678_),
    .B(_0949_),
    .Y(_0968_));
 sg13g2_nand2b_2 _1907_ (.Y(_0969_),
    .B(_0948_),
    .A_N(_0678_));
 sg13g2_nor2_2 _1908_ (.A(_0950_),
    .B(_0969_),
    .Y(_0970_));
 sg13g2_nand2_1 _1909_ (.Y(_0971_),
    .A(net518),
    .B(_0968_));
 sg13g2_nor2_2 _1910_ (.A(net503),
    .B(net520),
    .Y(_0972_));
 sg13g2_nand2_2 _1911_ (.Y(_0973_),
    .A(net495),
    .B(net516));
 sg13g2_nor2_2 _1912_ (.A(net503),
    .B(net491),
    .Y(_0974_));
 sg13g2_nand2_2 _1913_ (.Y(_0975_),
    .A(net498),
    .B(_0970_));
 sg13g2_nor2_2 _1914_ (.A(net474),
    .B(net450),
    .Y(_0976_));
 sg13g2_xnor2_1 _1915_ (.Y(_0977_),
    .A(net550),
    .B(\wrapper.pixel.sprite_top[0] ));
 sg13g2_xor2_1 _1916_ (.B(\wrapper.pixel.sprite_top[0] ),
    .A(net550),
    .X(_0978_));
 sg13g2_xor2_1 _1917_ (.B(_0653_),
    .A(_0652_),
    .X(_0979_));
 sg13g2_xnor2_1 _1918_ (.Y(_0980_),
    .A(_0652_),
    .B(_0653_));
 sg13g2_nor2_2 _1919_ (.A(_0652_),
    .B(net527),
    .Y(_0981_));
 sg13g2_nand2_2 _1920_ (.Y(_0982_),
    .A(net532),
    .B(net508));
 sg13g2_nor2_1 _1921_ (.A(net484),
    .B(net450),
    .Y(_0983_));
 sg13g2_a221oi_1 _1922_ (.B2(_0959_),
    .C1(_0982_),
    .B1(net443),
    .A1(_0974_),
    .Y(_0984_),
    .A2(_0976_));
 sg13g2_nand2b_1 _1923_ (.Y(_0985_),
    .B(_0984_),
    .A_N(_0966_));
 sg13g2_nor2_2 _1924_ (.A(_0946_),
    .B(net520),
    .Y(_0986_));
 sg13g2_nand2_2 _1925_ (.Y(_0987_),
    .A(_0947_),
    .B(net516));
 sg13g2_nand2_2 _1926_ (.Y(_0988_),
    .A(net518),
    .B(_0953_));
 sg13g2_nand2_1 _1927_ (.Y(_0989_),
    .A(_0953_),
    .B(_0972_));
 sg13g2_a21oi_2 _1928_ (.B1(net470),
    .Y(_0990_),
    .A2(_0972_),
    .A1(_0953_));
 sg13g2_nor2_1 _1929_ (.A(net529),
    .B(net511),
    .Y(_0991_));
 sg13g2_nand2_2 _1930_ (.Y(_0992_),
    .A(_0652_),
    .B(net532));
 sg13g2_nor2_1 _1931_ (.A(net501),
    .B(net490),
    .Y(_0993_));
 sg13g2_nand2_2 _1932_ (.Y(_0994_),
    .A(net494),
    .B(_0986_));
 sg13g2_nor2_2 _1933_ (.A(net471),
    .B(_0993_),
    .Y(_0995_));
 sg13g2_nor2_2 _1934_ (.A(net445),
    .B(_0995_),
    .Y(_0996_));
 sg13g2_nand2_2 _1935_ (.Y(_0997_),
    .A(net495),
    .B(net490));
 sg13g2_nand3_1 _1936_ (.B(_0964_),
    .C(net490),
    .A(net494),
    .Y(_0998_));
 sg13g2_nor2_1 _1937_ (.A(_0947_),
    .B(_0948_),
    .Y(_0999_));
 sg13g2_nand2_2 _1938_ (.Y(_1000_),
    .A(_0946_),
    .B(net538));
 sg13g2_nor2_2 _1939_ (.A(net516),
    .B(_1000_),
    .Y(_1001_));
 sg13g2_nand2_2 _1940_ (.Y(_1002_),
    .A(net519),
    .B(net506));
 sg13g2_nand2_1 _1941_ (.Y(_1003_),
    .A(net501),
    .B(_1002_));
 sg13g2_nand3_1 _1942_ (.B(_0998_),
    .C(_1003_),
    .A(_0996_),
    .Y(_1004_));
 sg13g2_o21ai_1 _1943_ (.B1(_1004_),
    .Y(_1005_),
    .A1(_0958_),
    .A2(_0990_));
 sg13g2_xor2_1 _1944_ (.B(_0656_),
    .A(_0655_),
    .X(_1006_));
 sg13g2_xnor2_1 _1945_ (.Y(_1007_),
    .A(_0655_),
    .B(_0656_));
 sg13g2_xor2_1 _1946_ (.B(_0654_),
    .A(_0650_),
    .X(_1008_));
 sg13g2_xnor2_1 _1947_ (.Y(_1009_),
    .A(_0650_),
    .B(_0654_));
 sg13g2_nor2_2 _1948_ (.A(_1007_),
    .B(_1009_),
    .Y(_1010_));
 sg13g2_nand2_1 _1949_ (.Y(_1011_),
    .A(_1006_),
    .B(net488));
 sg13g2_o21ai_1 _1950_ (.B1(_1010_),
    .Y(_1012_),
    .A1(net521),
    .A2(_1005_));
 sg13g2_nor2_1 _1951_ (.A(net536),
    .B(net510),
    .Y(_1013_));
 sg13g2_nand2_1 _1952_ (.Y(_1014_),
    .A(net527),
    .B(net512));
 sg13g2_nand2_1 _1953_ (.Y(_1015_),
    .A(net498),
    .B(net491));
 sg13g2_nand3_1 _1954_ (.B(_0964_),
    .C(net492),
    .A(net499),
    .Y(_1016_));
 sg13g2_nand2_2 _1955_ (.Y(_1017_),
    .A(net503),
    .B(net491));
 sg13g2_nand3_1 _1956_ (.B(_1016_),
    .C(_1017_),
    .A(net443),
    .Y(_1018_));
 sg13g2_nor2_2 _1957_ (.A(net533),
    .B(net513),
    .Y(_1019_));
 sg13g2_nor2_2 _1958_ (.A(net503),
    .B(net518),
    .Y(_1020_));
 sg13g2_nand2_1 _1959_ (.Y(_1021_),
    .A(net493),
    .B(net519));
 sg13g2_o21ai_1 _1960_ (.B1(net453),
    .Y(_1022_),
    .A1(_0942_),
    .A2(_0964_));
 sg13g2_nand3_1 _1961_ (.B(net516),
    .C(net506),
    .A(net493),
    .Y(_1023_));
 sg13g2_nor2_1 _1962_ (.A(net469),
    .B(_1023_),
    .Y(_1024_));
 sg13g2_nor2_2 _1963_ (.A(net499),
    .B(net520),
    .Y(_1025_));
 sg13g2_nand2_2 _1964_ (.Y(_1026_),
    .A(net505),
    .B(net517));
 sg13g2_nand3_1 _1965_ (.B(net507),
    .C(_1025_),
    .A(net480),
    .Y(_1027_));
 sg13g2_nand2_1 _1966_ (.Y(_1028_),
    .A(net446),
    .B(_1027_));
 sg13g2_o21ai_1 _1967_ (.B1(_1028_),
    .Y(_1029_),
    .A1(_1022_),
    .A2(_1024_));
 sg13g2_a221oi_1 _1968_ (.B2(_1029_),
    .C1(_1012_),
    .B1(_1019_),
    .A1(net486),
    .Y(_1030_),
    .A2(_1018_));
 sg13g2_nand2_1 _1969_ (.Y(_1031_),
    .A(_0949_),
    .B(_0961_));
 sg13g2_a21oi_1 _1970_ (.A1(net469),
    .A2(_1031_),
    .Y(_1032_),
    .B1(_0990_));
 sg13g2_nor2b_1 _1971_ (.A(_1032_),
    .B_N(_0966_),
    .Y(_1033_));
 sg13g2_a21o_1 _1972_ (.A2(_1032_),
    .A1(net453),
    .B1(_0982_),
    .X(_1034_));
 sg13g2_nand2_2 _1973_ (.Y(_1035_),
    .A(net497),
    .B(_0967_));
 sg13g2_a21oi_1 _1974_ (.A1(net479),
    .A2(net468),
    .Y(_1036_),
    .B1(net446));
 sg13g2_o21ai_1 _1975_ (.B1(net469),
    .Y(_1037_),
    .A1(net502),
    .A2(_0960_));
 sg13g2_nor2_1 _1976_ (.A(net473),
    .B(net454),
    .Y(_1038_));
 sg13g2_nand2_2 _1977_ (.Y(_1039_),
    .A(net484),
    .B(net450));
 sg13g2_nor2_2 _1978_ (.A(net518),
    .B(_0968_),
    .Y(_1040_));
 sg13g2_nand2_2 _1979_ (.Y(_1041_),
    .A(net520),
    .B(_0969_));
 sg13g2_nor2_2 _1980_ (.A(_0997_),
    .B(_1040_),
    .Y(_1042_));
 sg13g2_a221oi_1 _1981_ (.B2(_1042_),
    .C1(_1014_),
    .B1(net440),
    .A1(_1036_),
    .Y(_1043_),
    .A2(_1037_));
 sg13g2_nor2_2 _1982_ (.A(net495),
    .B(_0988_),
    .Y(_1044_));
 sg13g2_nor2_1 _1983_ (.A(net470),
    .B(_1044_),
    .Y(_1045_));
 sg13g2_a21oi_1 _1984_ (.A1(net507),
    .A2(_1025_),
    .Y(_1046_),
    .B1(net480));
 sg13g2_o21ai_1 _1985_ (.B1(net446),
    .Y(_1047_),
    .A1(_1045_),
    .A2(_1046_));
 sg13g2_a21oi_1 _1986_ (.A1(_1022_),
    .A2(_1047_),
    .Y(_1048_),
    .B1(net521));
 sg13g2_nor2_2 _1987_ (.A(_1007_),
    .B(net488),
    .Y(_1049_));
 sg13g2_nand2_2 _1988_ (.Y(_1050_),
    .A(_1006_),
    .B(_1009_));
 sg13g2_o21ai_1 _1989_ (.B1(net504),
    .Y(_1051_),
    .A1(net517),
    .A2(_0969_));
 sg13g2_nand2_1 _1990_ (.Y(_1052_),
    .A(net497),
    .B(_0956_));
 sg13g2_o21ai_1 _1991_ (.B1(_1051_),
    .Y(_1053_),
    .A1(_0955_),
    .A2(_1015_));
 sg13g2_a21oi_1 _1992_ (.A1(net470),
    .A2(_1053_),
    .Y(_1054_),
    .B1(_0990_));
 sg13g2_nor2_2 _1993_ (.A(net453),
    .B(_0962_),
    .Y(_1055_));
 sg13g2_nand2_1 _1994_ (.Y(_1056_),
    .A(_0968_),
    .B(_1055_));
 sg13g2_o21ai_1 _1995_ (.B1(_1019_),
    .Y(_1057_),
    .A1(_1054_),
    .A2(_1056_));
 sg13g2_a21oi_1 _1996_ (.A1(net452),
    .A2(_1054_),
    .Y(_1058_),
    .B1(_1057_));
 sg13g2_nor4_1 _1997_ (.A(_1043_),
    .B(_1048_),
    .C(_1050_),
    .D(_1058_),
    .Y(_1059_));
 sg13g2_o21ai_1 _1998_ (.B1(_1059_),
    .Y(_1060_),
    .A1(_1033_),
    .A2(_1034_));
 sg13g2_nor2_2 _1999_ (.A(_0947_),
    .B(net516),
    .Y(_1061_));
 sg13g2_nand2_2 _2000_ (.Y(_1062_),
    .A(_0946_),
    .B(net519));
 sg13g2_nor2_1 _2001_ (.A(_0986_),
    .B(_1061_),
    .Y(_1063_));
 sg13g2_nor2_2 _2002_ (.A(net520),
    .B(_0960_),
    .Y(_1064_));
 sg13g2_nand2_2 _2003_ (.Y(_1065_),
    .A(net517),
    .B(_0959_));
 sg13g2_nand2_2 _2004_ (.Y(_1066_),
    .A(net500),
    .B(_1065_));
 sg13g2_a221oi_1 _2005_ (.B2(net502),
    .C1(net532),
    .B1(_1065_),
    .A1(net479),
    .Y(_1067_),
    .A2(net468));
 sg13g2_o21ai_1 _2006_ (.B1(_1067_),
    .Y(_1068_),
    .A1(_0948_),
    .A2(_1063_));
 sg13g2_nor2_1 _2007_ (.A(net502),
    .B(_1065_),
    .Y(_1069_));
 sg13g2_nand2b_2 _2008_ (.Y(_1070_),
    .B(net479),
    .A_N(_1069_));
 sg13g2_nor2_2 _2009_ (.A(net493),
    .B(_0953_),
    .Y(_1071_));
 sg13g2_nor2_1 _2010_ (.A(net526),
    .B(_1071_),
    .Y(_1072_));
 sg13g2_nor2_1 _2011_ (.A(net517),
    .B(net506),
    .Y(_1073_));
 sg13g2_nor2_2 _2012_ (.A(net520),
    .B(_0968_),
    .Y(_1074_));
 sg13g2_nor2_2 _2013_ (.A(_0970_),
    .B(_1001_),
    .Y(_1075_));
 sg13g2_nand2_1 _2014_ (.Y(_1076_),
    .A(net502),
    .B(_0988_));
 sg13g2_nand4_1 _2015_ (.B(_1070_),
    .C(_1075_),
    .A(net532),
    .Y(_1077_),
    .D(_1076_));
 sg13g2_nand2_1 _2016_ (.Y(_1078_),
    .A(_1068_),
    .B(_1077_));
 sg13g2_o21ai_1 _2017_ (.B1(net469),
    .Y(_1079_),
    .A1(_0997_),
    .A2(_1061_));
 sg13g2_nor2_1 _2018_ (.A(_0982_),
    .B(_0990_),
    .Y(_1080_));
 sg13g2_nand4_1 _2019_ (.B(net490),
    .C(_1019_),
    .A(net495),
    .Y(_1081_),
    .D(_1070_));
 sg13g2_nand2_1 _2020_ (.Y(_1082_),
    .A(net488),
    .B(_1081_));
 sg13g2_a221oi_1 _2021_ (.B2(_1080_),
    .C1(_1082_),
    .B1(_1079_),
    .A1(net513),
    .Y(_1083_),
    .A2(_1078_));
 sg13g2_nand2_1 _2022_ (.Y(_1084_),
    .A(net495),
    .B(_1001_));
 sg13g2_nand2_2 _2023_ (.Y(_1085_),
    .A(_0969_),
    .B(_1000_));
 sg13g2_nor2_1 _2024_ (.A(_0968_),
    .B(net507),
    .Y(_1086_));
 sg13g2_nor2_2 _2025_ (.A(net517),
    .B(_1085_),
    .Y(_1087_));
 sg13g2_a21oi_2 _2026_ (.B1(net478),
    .Y(_1088_),
    .A2(_1087_),
    .A1(net500));
 sg13g2_a21oi_1 _2027_ (.A1(_1084_),
    .A2(_1088_),
    .Y(_1089_),
    .B1(net521));
 sg13g2_nand2_2 _2028_ (.Y(_1090_),
    .A(net517),
    .B(_1085_));
 sg13g2_nor2_2 _2029_ (.A(net475),
    .B(_0972_),
    .Y(_1091_));
 sg13g2_nand2_1 _2030_ (.Y(_1092_),
    .A(net495),
    .B(_1061_));
 sg13g2_o21ai_1 _2031_ (.B1(net479),
    .Y(_1093_),
    .A1(_0948_),
    .A2(_0973_));
 sg13g2_a221oi_1 _2032_ (.B2(net469),
    .C1(net512),
    .B1(_1092_),
    .A1(net532),
    .Y(_1094_),
    .A2(_1090_));
 sg13g2_nand2_2 _2033_ (.Y(_1095_),
    .A(net516),
    .B(_1000_));
 sg13g2_nor2_1 _2034_ (.A(net519),
    .B(net506),
    .Y(_1096_));
 sg13g2_nor2_2 _2035_ (.A(net504),
    .B(_1096_),
    .Y(_1097_));
 sg13g2_nand3_1 _2036_ (.B(net486),
    .C(_1097_),
    .A(_0952_),
    .Y(_1098_));
 sg13g2_o21ai_1 _2037_ (.B1(_1009_),
    .Y(_1099_),
    .A1(net480),
    .A2(_1098_));
 sg13g2_a221oi_1 _2038_ (.B2(_1094_),
    .C1(_1099_),
    .B1(_1093_),
    .A1(_1070_),
    .Y(_1100_),
    .A2(_1089_));
 sg13g2_nor4_1 _2039_ (.A(net446),
    .B(_1006_),
    .C(_1083_),
    .D(_1100_),
    .Y(_1101_));
 sg13g2_a21oi_1 _2040_ (.A1(_0985_),
    .A2(_1030_),
    .Y(_1102_),
    .B1(_1101_));
 sg13g2_a21oi_1 _2041_ (.A1(_1060_),
    .A2(_1102_),
    .Y(_1103_),
    .B1(net457));
 sg13g2_xnor2_1 _2042_ (.Y(_1104_),
    .A(net541),
    .B(\wrapper.pixel.sprite_top[5] ));
 sg13g2_xnor2_1 _2043_ (.Y(_1105_),
    .A(_0659_),
    .B(_1104_));
 sg13g2_xor2_1 _2044_ (.B(_1104_),
    .A(_0659_),
    .X(_1106_));
 sg13g2_nand4_1 _2045_ (.B(_1006_),
    .C(net487),
    .A(net443),
    .Y(_1107_),
    .D(_1044_));
 sg13g2_a21o_1 _2046_ (.A2(_1107_),
    .A1(_1011_),
    .B1(_0936_),
    .X(_1108_));
 sg13g2_nand2_1 _2047_ (.Y(_1109_),
    .A(net503),
    .B(_1064_));
 sg13g2_nor2_1 _2048_ (.A(net509),
    .B(_1109_),
    .Y(_1110_));
 sg13g2_a21oi_1 _2049_ (.A1(net442),
    .A2(_1110_),
    .Y(_1111_),
    .B1(_1009_));
 sg13g2_o21ai_1 _2050_ (.B1(_1105_),
    .Y(_1112_),
    .A1(_1108_),
    .A2(_1111_));
 sg13g2_nand2_2 _2051_ (.Y(_1113_),
    .A(_0941_),
    .B(net455));
 sg13g2_o21ai_1 _2052_ (.B1(net536),
    .Y(_1114_),
    .A1(net491),
    .A2(_1113_));
 sg13g2_nor2_2 _2053_ (.A(_0947_),
    .B(net519),
    .Y(_1115_));
 sg13g2_nand2b_2 _2054_ (.Y(_1116_),
    .B(net500),
    .A_N(_1115_));
 sg13g2_nor3_2 _2055_ (.A(net493),
    .B(_0953_),
    .C(_1115_),
    .Y(_1117_));
 sg13g2_a21oi_2 _2056_ (.B1(_1117_),
    .Y(_1118_),
    .A2(_0964_),
    .A1(net494));
 sg13g2_a21oi_1 _2057_ (.A1(net441),
    .A2(_1118_),
    .Y(_1119_),
    .B1(_1114_));
 sg13g2_a21o_1 _2058_ (.A2(net490),
    .A1(_0954_),
    .B1(_1113_),
    .X(_1120_));
 sg13g2_o21ai_1 _2059_ (.B1(net441),
    .Y(_1121_),
    .A1(_0974_),
    .A2(_1044_));
 sg13g2_nand3_1 _2060_ (.B(_1120_),
    .C(_1121_),
    .A(net529),
    .Y(_1122_));
 sg13g2_nor2_1 _2061_ (.A(net509),
    .B(_1119_),
    .Y(_1123_));
 sg13g2_nor2_2 _2062_ (.A(net501),
    .B(_1001_),
    .Y(_1124_));
 sg13g2_nand2_2 _2063_ (.Y(_1125_),
    .A(net494),
    .B(_1002_));
 sg13g2_a221oi_1 _2064_ (.B2(net492),
    .C1(net533),
    .B1(_1124_),
    .A1(net500),
    .Y(_1126_),
    .A2(_1065_));
 sg13g2_a21oi_1 _2065_ (.A1(_0965_),
    .A2(_0994_),
    .Y(_1127_),
    .B1(net526));
 sg13g2_o21ai_1 _2066_ (.B1(net443),
    .Y(_1128_),
    .A1(_1126_),
    .A2(_1127_));
 sg13g2_o21ai_1 _2067_ (.B1(_1023_),
    .Y(_1129_),
    .A1(_1026_),
    .A2(_1085_));
 sg13g2_a22oi_1 _2068_ (.Y(_1130_),
    .B1(_1129_),
    .B2(net530),
    .A2(_1072_),
    .A1(_1016_));
 sg13g2_o21ai_1 _2069_ (.B1(_1128_),
    .Y(_1131_),
    .A1(_1039_),
    .A2(_1130_));
 sg13g2_nor2_2 _2070_ (.A(_1006_),
    .B(net488),
    .Y(_1132_));
 sg13g2_nand2_2 _2071_ (.Y(_1133_),
    .A(_1007_),
    .B(_1009_));
 sg13g2_a221oi_1 _2072_ (.B2(net509),
    .C1(_1133_),
    .B1(_1131_),
    .A1(_1122_),
    .Y(_1134_),
    .A2(_1123_));
 sg13g2_nand2_2 _2073_ (.Y(_1135_),
    .A(_1007_),
    .B(net488));
 sg13g2_nor2_2 _2074_ (.A(net497),
    .B(_0967_),
    .Y(_1136_));
 sg13g2_nand2_2 _2075_ (.Y(_1137_),
    .A(net503),
    .B(_1095_));
 sg13g2_nand2_2 _2076_ (.Y(_1138_),
    .A(_0973_),
    .B(_1137_));
 sg13g2_nor2_2 _2077_ (.A(net476),
    .B(net531),
    .Y(_1139_));
 sg13g2_nand3_1 _2078_ (.B(_1069_),
    .C(_1139_),
    .A(net452),
    .Y(_1140_));
 sg13g2_nand2_2 _2079_ (.Y(_1141_),
    .A(_0998_),
    .B(_1035_));
 sg13g2_nand3_1 _2080_ (.B(_0988_),
    .C(_1002_),
    .A(net500),
    .Y(_1142_));
 sg13g2_nand3_1 _2081_ (.B(net526),
    .C(_1090_),
    .A(net493),
    .Y(_1143_));
 sg13g2_nand2_1 _2082_ (.Y(_1144_),
    .A(net531),
    .B(_1141_));
 sg13g2_nand4_1 _2083_ (.B(_1142_),
    .C(_1143_),
    .A(net440),
    .Y(_1145_),
    .D(_1144_));
 sg13g2_a22oi_1 _2084_ (.Y(_1146_),
    .B1(_1140_),
    .B2(_1145_),
    .A2(_1138_),
    .A1(net513));
 sg13g2_nand3_1 _2085_ (.B(_0968_),
    .C(_1091_),
    .A(_0962_),
    .Y(_1147_));
 sg13g2_o21ai_1 _2086_ (.B1(_0988_),
    .Y(_1148_),
    .A1(net538),
    .A2(net518));
 sg13g2_a21oi_1 _2087_ (.A1(net480),
    .A2(_1148_),
    .Y(_1149_),
    .B1(_0982_));
 sg13g2_o21ai_1 _2088_ (.B1(net470),
    .Y(_1150_),
    .A1(net538),
    .A2(_0962_));
 sg13g2_nand2b_1 _2089_ (.Y(_1151_),
    .B(_1150_),
    .A_N(_1045_));
 sg13g2_a221oi_1 _2090_ (.B2(net489),
    .C1(_1149_),
    .B1(_1151_),
    .A1(net486),
    .Y(_1152_),
    .A2(_1147_));
 sg13g2_o21ai_1 _2091_ (.B1(net457),
    .Y(_1153_),
    .A1(_1050_),
    .A2(_1152_));
 sg13g2_nor2_1 _2092_ (.A(net476),
    .B(net526),
    .Y(_1154_));
 sg13g2_nand2_2 _2093_ (.Y(_1155_),
    .A(net471),
    .B(net533));
 sg13g2_nor3_2 _2094_ (.A(net511),
    .B(net506),
    .C(_1115_),
    .Y(_1156_));
 sg13g2_nor2_1 _2095_ (.A(_1155_),
    .B(_1156_),
    .Y(_1157_));
 sg13g2_nor2_1 _2096_ (.A(net504),
    .B(_1064_),
    .Y(_1158_));
 sg13g2_a221oi_1 _2097_ (.B2(net502),
    .C1(_1009_),
    .B1(_1157_),
    .A1(net479),
    .Y(_1159_),
    .A2(_1069_));
 sg13g2_nand3_1 _2098_ (.B(net538),
    .C(_1062_),
    .A(net479),
    .Y(_1160_));
 sg13g2_a21oi_1 _2099_ (.A1(net469),
    .A2(_1061_),
    .Y(_1161_),
    .B1(net532));
 sg13g2_a221oi_1 _2100_ (.B2(_1161_),
    .C1(net495),
    .B1(_1160_),
    .A1(_0956_),
    .Y(_1162_),
    .A2(net488));
 sg13g2_o21ai_1 _2101_ (.B1(net446),
    .Y(_1163_),
    .A1(net513),
    .A2(_1162_));
 sg13g2_o21ai_1 _2102_ (.B1(_1006_),
    .Y(_1164_),
    .A1(_1159_),
    .A2(_1163_));
 sg13g2_o21ai_1 _2103_ (.B1(_1164_),
    .Y(_1165_),
    .A1(_1135_),
    .A2(_1146_));
 sg13g2_nor3_1 _2104_ (.A(_1134_),
    .B(_1153_),
    .C(_1165_),
    .Y(_1166_));
 sg13g2_nor2_1 _2105_ (.A(net458),
    .B(_1133_),
    .Y(_1167_));
 sg13g2_nor2_2 _2106_ (.A(net498),
    .B(net491),
    .Y(_1168_));
 sg13g2_nand2_2 _2107_ (.Y(_1169_),
    .A(net503),
    .B(_0970_));
 sg13g2_nand3_1 _2108_ (.B(_0963_),
    .C(_1019_),
    .A(net496),
    .Y(_1170_));
 sg13g2_o21ai_1 _2109_ (.B1(_1170_),
    .Y(_1171_),
    .A1(net521),
    .A2(_1084_));
 sg13g2_a21oi_1 _2110_ (.A1(_0981_),
    .A2(_1168_),
    .Y(_1172_),
    .B1(_1171_));
 sg13g2_nor4_1 _2111_ (.A(net457),
    .B(_1039_),
    .C(_1133_),
    .D(_1172_),
    .Y(_1173_));
 sg13g2_or3_1 _2112_ (.A(_1105_),
    .B(_1166_),
    .C(_1173_),
    .X(_1174_));
 sg13g2_o21ai_1 _2113_ (.B1(_1174_),
    .Y(_0000_),
    .A1(_1103_),
    .A2(_1112_));
 sg13g2_o21ai_1 _2114_ (.B1(_0954_),
    .Y(_1175_),
    .A1(_0949_),
    .A2(net510));
 sg13g2_nand3_1 _2115_ (.B(_1025_),
    .C(_1175_),
    .A(net442),
    .Y(_1176_));
 sg13g2_a21o_1 _2116_ (.A2(net489),
    .A1(_0946_),
    .B1(_1176_),
    .X(_1177_));
 sg13g2_o21ai_1 _2117_ (.B1(net458),
    .Y(_1178_),
    .A1(net444),
    .A2(_1177_));
 sg13g2_and2_1 _2118_ (.A(_1105_),
    .B(_1178_),
    .X(_1179_));
 sg13g2_a21oi_1 _2119_ (.A1(_0954_),
    .A2(_1158_),
    .Y(_1180_),
    .B1(_1168_));
 sg13g2_nor3_1 _2120_ (.A(net482),
    .B(net449),
    .C(_1180_),
    .Y(_1181_));
 sg13g2_nand2b_1 _2121_ (.Y(_1182_),
    .B(net442),
    .A_N(_1180_));
 sg13g2_nor2_2 _2122_ (.A(net494),
    .B(_1062_),
    .Y(_1183_));
 sg13g2_nand2_2 _2123_ (.Y(_1184_),
    .A(net501),
    .B(_1061_));
 sg13g2_nand2_1 _2124_ (.Y(_1185_),
    .A(_1095_),
    .B(_1124_));
 sg13g2_nand2_1 _2125_ (.Y(_1186_),
    .A(_1184_),
    .B(_1185_));
 sg13g2_nor2_2 _2126_ (.A(net493),
    .B(_1041_),
    .Y(_1187_));
 sg13g2_nor2_1 _2127_ (.A(net478),
    .B(_0961_),
    .Y(_1188_));
 sg13g2_nor2_2 _2128_ (.A(net481),
    .B(_1187_),
    .Y(_1189_));
 sg13g2_or2_1 _2129_ (.X(_1190_),
    .B(_1188_),
    .A(net452));
 sg13g2_nor2_1 _2130_ (.A(net454),
    .B(_1189_),
    .Y(_1191_));
 sg13g2_or2_1 _2131_ (.X(_1192_),
    .B(_1189_),
    .A(net454));
 sg13g2_a21oi_1 _2132_ (.A1(net498),
    .A2(_1041_),
    .Y(_1193_),
    .B1(net473));
 sg13g2_nand2b_1 _2133_ (.Y(_1194_),
    .B(net454),
    .A_N(_1193_));
 sg13g2_a221oi_1 _2134_ (.B2(_1194_),
    .C1(net534),
    .B1(_1192_),
    .A1(net440),
    .Y(_1195_),
    .A2(_1186_));
 sg13g2_a221oi_1 _2135_ (.B2(net447),
    .C1(net529),
    .B1(_1189_),
    .A1(net440),
    .Y(_1196_),
    .A2(_1183_));
 sg13g2_a21oi_2 _2136_ (.B1(net478),
    .Y(_1197_),
    .A2(_1142_),
    .A1(_1052_));
 sg13g2_nand2_1 _2137_ (.Y(_1198_),
    .A(net498),
    .B(_1074_));
 sg13g2_a22oi_1 _2138_ (.Y(_1199_),
    .B1(_1198_),
    .B2(_0976_),
    .A2(_1197_),
    .A1(net455));
 sg13g2_a221oi_1 _2139_ (.B2(_1199_),
    .C1(net514),
    .B1(_1196_),
    .A1(_1182_),
    .Y(_1200_),
    .A2(_1195_));
 sg13g2_nor2_2 _2140_ (.A(net482),
    .B(_1183_),
    .Y(_1201_));
 sg13g2_nand2_1 _2141_ (.Y(_1202_),
    .A(net473),
    .B(_1184_));
 sg13g2_a21oi_1 _2142_ (.A1(_0954_),
    .A2(net490),
    .Y(_1203_),
    .B1(_1074_));
 sg13g2_nand2_2 _2143_ (.Y(_1204_),
    .A(net493),
    .B(_0988_));
 sg13g2_o21ai_1 _2144_ (.B1(net483),
    .Y(_1205_),
    .A1(_1064_),
    .A2(_1204_));
 sg13g2_nor2_1 _2145_ (.A(_1203_),
    .B(_1205_),
    .Y(_1206_));
 sg13g2_nand2_2 _2146_ (.Y(_1207_),
    .A(net448),
    .B(_1201_));
 sg13g2_a22oi_1 _2147_ (.Y(_1208_),
    .B1(_1206_),
    .B2(net447),
    .A2(_1125_),
    .A1(_0976_));
 sg13g2_nand3_1 _2148_ (.B(_1207_),
    .C(_1208_),
    .A(_1182_),
    .Y(_1209_));
 sg13g2_nand2_1 _2149_ (.Y(_1210_),
    .A(net487),
    .B(_1209_));
 sg13g2_nor2_2 _2150_ (.A(net455),
    .B(_1201_),
    .Y(_1211_));
 sg13g2_nand2_2 _2151_ (.Y(_1212_),
    .A(net449),
    .B(_1202_));
 sg13g2_nor2_2 _2152_ (.A(net505),
    .B(_1061_),
    .Y(_1213_));
 sg13g2_nand2_2 _2153_ (.Y(_1214_),
    .A(net494),
    .B(_1062_));
 sg13g2_a21oi_1 _2154_ (.A1(net482),
    .A2(_1214_),
    .Y(_1215_),
    .B1(net447));
 sg13g2_a221oi_1 _2155_ (.B2(_0976_),
    .C1(_1181_),
    .B1(_1214_),
    .A1(net448),
    .Y(_1216_),
    .A2(_1201_));
 sg13g2_a22oi_1 _2156_ (.Y(_1217_),
    .B1(_1136_),
    .B2(_0946_),
    .A2(_1075_),
    .A1(net497));
 sg13g2_o21ai_1 _2157_ (.B1(_1216_),
    .Y(_1218_),
    .A1(_1039_),
    .A2(_1217_));
 sg13g2_a21oi_1 _2158_ (.A1(net489),
    .A2(_1218_),
    .Y(_1219_),
    .B1(_1200_));
 sg13g2_a21oi_1 _2159_ (.A1(_1210_),
    .A2(_1219_),
    .Y(_1220_),
    .B1(net444));
 sg13g2_and3_2 _2160_ (.X(_1221_),
    .A(net476),
    .B(_0994_),
    .C(net468));
 sg13g2_nand3_1 _2161_ (.B(_0994_),
    .C(net468),
    .A(net476),
    .Y(_1222_));
 sg13g2_nand3_1 _2162_ (.B(_1184_),
    .C(_1214_),
    .A(_0988_),
    .Y(_1223_));
 sg13g2_a21oi_1 _2163_ (.A1(_1222_),
    .A2(_1223_),
    .Y(_1224_),
    .B1(_1000_));
 sg13g2_nand2_1 _2164_ (.Y(_1225_),
    .A(net448),
    .B(net535));
 sg13g2_nor2_2 _2165_ (.A(net445),
    .B(_1221_),
    .Y(_1226_));
 sg13g2_a221oi_1 _2166_ (.B2(_1223_),
    .C1(net526),
    .B1(_1226_),
    .A1(_1055_),
    .Y(_1227_),
    .A2(_1224_));
 sg13g2_a221oi_1 _2167_ (.B2(_1071_),
    .C1(net445),
    .B1(_1062_),
    .A1(_0995_),
    .Y(_1228_),
    .A2(net468));
 sg13g2_a221oi_1 _2168_ (.B2(_1021_),
    .C1(net531),
    .B1(_1228_),
    .A1(net440),
    .Y(_1229_),
    .A2(_1187_));
 sg13g2_o21ai_1 _2169_ (.B1(net508),
    .Y(_1230_),
    .A1(_1227_),
    .A2(_1229_));
 sg13g2_nor2_1 _2170_ (.A(net446),
    .B(_1091_),
    .Y(_1231_));
 sg13g2_nand2_1 _2171_ (.Y(_1232_),
    .A(net452),
    .B(_1093_));
 sg13g2_o21ai_1 _2172_ (.B1(_1232_),
    .Y(_1233_),
    .A1(_1042_),
    .A2(_1190_));
 sg13g2_nand3_1 _2173_ (.B(_0975_),
    .C(_1197_),
    .A(net453),
    .Y(_1234_));
 sg13g2_a21oi_1 _2174_ (.A1(_1233_),
    .A2(_1234_),
    .Y(_1235_),
    .B1(_1014_));
 sg13g2_nand2_1 _2175_ (.Y(_1236_),
    .A(_0954_),
    .B(_1020_));
 sg13g2_and2_1 _2176_ (.A(_1023_),
    .B(_1236_),
    .X(_1237_));
 sg13g2_a21oi_1 _2177_ (.A1(_0964_),
    .A2(_1071_),
    .Y(_1238_),
    .B1(_1221_));
 sg13g2_a21oi_1 _2178_ (.A1(_1237_),
    .A2(_1238_),
    .Y(_1239_),
    .B1(net445));
 sg13g2_nor3_2 _2179_ (.A(net472),
    .B(net497),
    .C(_0986_),
    .Y(_1240_));
 sg13g2_nor2_2 _2180_ (.A(net456),
    .B(_1240_),
    .Y(_1241_));
 sg13g2_o21ai_1 _2181_ (.B1(_1056_),
    .Y(_1242_),
    .A1(_1239_),
    .A2(_1241_));
 sg13g2_o21ai_1 _2182_ (.B1(_1230_),
    .Y(_1243_),
    .A1(net521),
    .A2(_1242_));
 sg13g2_o21ai_1 _2183_ (.B1(_1049_),
    .Y(_1244_),
    .A1(_1235_),
    .A2(_1243_));
 sg13g2_nor3_1 _2184_ (.A(net476),
    .B(net526),
    .C(_1214_),
    .Y(_1245_));
 sg13g2_a21oi_1 _2185_ (.A1(_0941_),
    .A2(_1041_),
    .Y(_1246_),
    .B1(_1245_));
 sg13g2_a21oi_1 _2186_ (.A1(_1226_),
    .A2(_1246_),
    .Y(_1247_),
    .B1(net508));
 sg13g2_nor2_1 _2187_ (.A(net488),
    .B(_1247_),
    .Y(_1248_));
 sg13g2_a21oi_1 _2188_ (.A1(_1125_),
    .A2(_1184_),
    .Y(_1249_),
    .B1(net476));
 sg13g2_o21ai_1 _2189_ (.B1(net531),
    .Y(_1250_),
    .A1(_0961_),
    .A2(_1124_));
 sg13g2_nand2_1 _2190_ (.Y(_1251_),
    .A(net452),
    .B(_1250_));
 sg13g2_nor2_1 _2191_ (.A(_1249_),
    .B(_1251_),
    .Y(_1252_));
 sg13g2_a21oi_1 _2192_ (.A1(_1070_),
    .A2(_1252_),
    .Y(_1253_),
    .B1(net512));
 sg13g2_nor2b_1 _2193_ (.A(_1253_),
    .B_N(_1248_),
    .Y(_1254_));
 sg13g2_nor3_1 _2194_ (.A(net471),
    .B(net531),
    .C(_0993_),
    .Y(_1255_));
 sg13g2_nor3_1 _2195_ (.A(net445),
    .B(_1221_),
    .C(_1255_),
    .Y(_1256_));
 sg13g2_nor2_1 _2196_ (.A(net497),
    .B(_1074_),
    .Y(_1257_));
 sg13g2_or2_2 _2197_ (.X(_1258_),
    .B(_1074_),
    .A(_1051_));
 sg13g2_nand2_1 _2198_ (.Y(_1259_),
    .A(_0994_),
    .B(_1258_));
 sg13g2_nor2_1 _2199_ (.A(_1155_),
    .B(_1258_),
    .Y(_1260_));
 sg13g2_nor2_1 _2200_ (.A(net504),
    .B(_1073_),
    .Y(_1261_));
 sg13g2_or2_1 _2201_ (.X(_1262_),
    .B(_1073_),
    .A(net504));
 sg13g2_o21ai_1 _2202_ (.B1(net493),
    .Y(_1263_),
    .A1(_0986_),
    .A2(_1001_));
 sg13g2_nand2b_1 _2203_ (.Y(_1264_),
    .B(_1263_),
    .A_N(_1117_));
 sg13g2_a221oi_1 _2204_ (.B2(_1139_),
    .C1(net512),
    .B1(_1264_),
    .A1(_1154_),
    .Y(_1265_),
    .A2(_1259_));
 sg13g2_nand3_1 _2205_ (.B(_0956_),
    .C(_1065_),
    .A(net500),
    .Y(_1266_));
 sg13g2_nand2_1 _2206_ (.Y(_1267_),
    .A(_1263_),
    .B(_1266_));
 sg13g2_a22oi_1 _2207_ (.Y(_1268_),
    .B1(net492),
    .B2(_1213_),
    .A2(_0961_),
    .A1(net538));
 sg13g2_a221oi_1 _2208_ (.B2(_1139_),
    .C1(net508),
    .B1(_1268_),
    .A1(_1154_),
    .Y(_1269_),
    .A2(_1267_));
 sg13g2_a22oi_1 _2209_ (.Y(_1270_),
    .B1(_1269_),
    .B2(_0996_),
    .A2(_1265_),
    .A1(_1256_));
 sg13g2_o21ai_1 _2210_ (.B1(_1007_),
    .Y(_1271_),
    .A1(_1009_),
    .A2(_1270_));
 sg13g2_o21ai_1 _2211_ (.B1(_1244_),
    .Y(_1272_),
    .A1(_1254_),
    .A2(_1271_));
 sg13g2_o21ai_1 _2212_ (.B1(_0936_),
    .Y(_1273_),
    .A1(_1220_),
    .A2(_1272_));
 sg13g2_o21ai_1 _2213_ (.B1(net509),
    .Y(_1274_),
    .A1(_0969_),
    .A2(net536));
 sg13g2_o21ai_1 _2214_ (.B1(_1274_),
    .Y(_1275_),
    .A1(_0960_),
    .A2(net529));
 sg13g2_nand4_1 _2215_ (.B(net441),
    .C(_1132_),
    .A(_1020_),
    .Y(_1276_),
    .D(_1275_));
 sg13g2_a21oi_2 _2216_ (.B1(_1105_),
    .Y(_1277_),
    .A2(_1276_),
    .A1(_0936_));
 sg13g2_nand2_1 _2217_ (.Y(_1278_),
    .A(_0960_),
    .B(_1020_));
 sg13g2_a221oi_1 _2218_ (.B2(_0947_),
    .C1(_1212_),
    .B1(_1025_),
    .A1(_0960_),
    .Y(_1279_),
    .A2(_1020_));
 sg13g2_o21ai_1 _2219_ (.B1(net515),
    .Y(_1280_),
    .A1(net536),
    .A2(_1279_));
 sg13g2_a21oi_1 _2220_ (.A1(_1138_),
    .A2(_1211_),
    .Y(_1281_),
    .B1(_1114_));
 sg13g2_a21oi_1 _2221_ (.A1(_0972_),
    .A2(net442),
    .Y(_1282_),
    .B1(_1211_));
 sg13g2_a21oi_1 _2222_ (.A1(_1015_),
    .A2(_1266_),
    .Y(_1283_),
    .B1(_1039_));
 sg13g2_nor3_1 _2223_ (.A(_0982_),
    .B(_1282_),
    .C(_1283_),
    .Y(_1284_));
 sg13g2_o21ai_1 _2224_ (.B1(_1212_),
    .Y(_1285_),
    .A1(_0987_),
    .A2(_1113_));
 sg13g2_nor2_1 _2225_ (.A(_0959_),
    .B(_1026_),
    .Y(_1286_));
 sg13g2_o21ai_1 _2226_ (.B1(net450),
    .Y(_1287_),
    .A1(_1097_),
    .A2(_1286_));
 sg13g2_nand3_1 _2227_ (.B(_1285_),
    .C(_1287_),
    .A(_1019_),
    .Y(_1288_));
 sg13g2_nor2b_1 _2228_ (.A(_1284_),
    .B_N(_1288_),
    .Y(_1289_));
 sg13g2_o21ai_1 _2229_ (.B1(_1289_),
    .Y(_1290_),
    .A1(_1280_),
    .A2(_1281_));
 sg13g2_nand2b_1 _2230_ (.Y(_1291_),
    .B(_1290_),
    .A_N(_1135_));
 sg13g2_a21oi_2 _2231_ (.B1(net482),
    .Y(_1292_),
    .A2(net490),
    .A1(net504));
 sg13g2_nor3_1 _2232_ (.A(net537),
    .B(_1240_),
    .C(_1292_),
    .Y(_1293_));
 sg13g2_nor2_1 _2233_ (.A(net474),
    .B(_1137_),
    .Y(_1294_));
 sg13g2_nand2_2 _2234_ (.Y(_1295_),
    .A(net474),
    .B(_1137_));
 sg13g2_nor2_1 _2235_ (.A(net529),
    .B(_1294_),
    .Y(_1296_));
 sg13g2_a21oi_1 _2236_ (.A1(_1295_),
    .A2(_1296_),
    .Y(_1297_),
    .B1(_1293_));
 sg13g2_o21ai_1 _2237_ (.B1(net510),
    .Y(_1298_),
    .A1(net456),
    .A2(_1297_));
 sg13g2_nor3_1 _2238_ (.A(net537),
    .B(_1097_),
    .C(_1168_),
    .Y(_1299_));
 sg13g2_or2_1 _2239_ (.X(_1300_),
    .B(_1044_),
    .A(net484));
 sg13g2_nand3b_1 _2240_ (.B(_1300_),
    .C(_1241_),
    .Y(_1301_),
    .A_N(_1299_));
 sg13g2_a21oi_1 _2241_ (.A1(net514),
    .A2(_1301_),
    .Y(_1302_),
    .B1(net444));
 sg13g2_o21ai_1 _2242_ (.B1(_1266_),
    .Y(_1303_),
    .A1(net501),
    .A2(_0963_));
 sg13g2_inv_1 _2243_ (.Y(_1304_),
    .A(_1303_));
 sg13g2_nand3_1 _2244_ (.B(net492),
    .C(_1041_),
    .A(_0941_),
    .Y(_1305_));
 sg13g2_a22oi_1 _2245_ (.Y(_1306_),
    .B1(_1305_),
    .B2(net452),
    .A2(_1303_),
    .A1(net478));
 sg13g2_o21ai_1 _2246_ (.B1(net513),
    .Y(_1307_),
    .A1(net531),
    .A2(_1306_));
 sg13g2_nor2_2 _2247_ (.A(net500),
    .B(_1087_),
    .Y(_1308_));
 sg13g2_o21ai_1 _2248_ (.B1(net497),
    .Y(_1309_),
    .A1(net517),
    .A2(_1085_));
 sg13g2_a21o_1 _2249_ (.A2(_1309_),
    .A1(_1066_),
    .B1(net472),
    .X(_1310_));
 sg13g2_a22oi_1 _2250_ (.Y(_1311_),
    .B1(_1310_),
    .B2(net449),
    .A2(net491),
    .A1(_0941_));
 sg13g2_a21o_1 _2251_ (.A2(_1311_),
    .A1(net535),
    .B1(_1307_),
    .X(_1312_));
 sg13g2_nand2_1 _2252_ (.Y(_1313_),
    .A(_1066_),
    .B(_1262_));
 sg13g2_nand3_1 _2253_ (.B(net447),
    .C(_1313_),
    .A(net482),
    .Y(_1314_));
 sg13g2_nand2_1 _2254_ (.Y(_1315_),
    .A(_1085_),
    .B(_1213_));
 sg13g2_a21oi_1 _2255_ (.A1(_1292_),
    .A2(_1315_),
    .Y(_1316_),
    .B1(net448));
 sg13g2_nor2_1 _2256_ (.A(net534),
    .B(_1316_),
    .Y(_1317_));
 sg13g2_nand2_1 _2257_ (.Y(_1318_),
    .A(_1201_),
    .B(_1315_));
 sg13g2_nand2_1 _2258_ (.Y(_1319_),
    .A(net468),
    .B(_1263_));
 sg13g2_nand3_1 _2259_ (.B(_1066_),
    .C(_1263_),
    .A(_1035_),
    .Y(_1320_));
 sg13g2_nand3_1 _2260_ (.B(net447),
    .C(_1320_),
    .A(net482),
    .Y(_1321_));
 sg13g2_a21oi_1 _2261_ (.A1(net454),
    .A2(_1318_),
    .Y(_1322_),
    .B1(net529));
 sg13g2_a22oi_1 _2262_ (.Y(_1323_),
    .B1(_1321_),
    .B2(_1322_),
    .A2(_1317_),
    .A1(_1314_));
 sg13g2_o21ai_1 _2263_ (.B1(_1312_),
    .Y(_1324_),
    .A1(net514),
    .A2(_1323_));
 sg13g2_nand3_1 _2264_ (.B(_1207_),
    .C(_1324_),
    .A(_1132_),
    .Y(_1325_));
 sg13g2_nor2_1 _2265_ (.A(net455),
    .B(_1088_),
    .Y(_1326_));
 sg13g2_nor2_1 _2266_ (.A(_1051_),
    .B(_1115_),
    .Y(_1327_));
 sg13g2_o21ai_1 _2267_ (.B1(net481),
    .Y(_1328_),
    .A1(_1261_),
    .A2(_1327_));
 sg13g2_a21oi_1 _2268_ (.A1(_1326_),
    .A2(_1328_),
    .Y(_1329_),
    .B1(net528));
 sg13g2_o21ai_1 _2269_ (.B1(net481),
    .Y(_1330_),
    .A1(_1257_),
    .A2(_1319_));
 sg13g2_o21ai_1 _2270_ (.B1(net472),
    .Y(_1331_),
    .A1(_0962_),
    .A2(net506));
 sg13g2_and3_1 _2271_ (.X(_1332_),
    .A(net447),
    .B(net514),
    .C(_1331_));
 sg13g2_a21oi_1 _2272_ (.A1(_1330_),
    .A2(_1332_),
    .Y(_1333_),
    .B1(_0991_));
 sg13g2_a21oi_1 _2273_ (.A1(_1116_),
    .A2(net467),
    .Y(_1334_),
    .B1(net471));
 sg13g2_a221oi_1 _2274_ (.B2(_1309_),
    .C1(net472),
    .B1(_1116_),
    .A1(_0961_),
    .Y(_1335_),
    .A2(_0968_));
 sg13g2_nor2b_1 _2275_ (.A(_1335_),
    .B_N(_1019_),
    .Y(_1336_));
 sg13g2_o21ai_1 _2276_ (.B1(_1023_),
    .Y(_1337_),
    .A1(_0959_),
    .A2(_1021_));
 sg13g2_o21ai_1 _2277_ (.B1(net533),
    .Y(_1338_),
    .A1(net496),
    .A2(_1063_));
 sg13g2_o21ai_1 _2278_ (.B1(_1155_),
    .Y(_1339_),
    .A1(_1337_),
    .A2(_1338_));
 sg13g2_nor3_1 _2279_ (.A(net454),
    .B(net515),
    .C(_1189_),
    .Y(_1340_));
 sg13g2_a22oi_1 _2280_ (.Y(_1341_),
    .B1(_1339_),
    .B2(_1340_),
    .A2(_1336_),
    .A1(_1326_));
 sg13g2_o21ai_1 _2281_ (.B1(_1341_),
    .Y(_1342_),
    .A1(_1329_),
    .A2(_1333_));
 sg13g2_a221oi_1 _2282_ (.B2(_1049_),
    .C1(_0936_),
    .B1(_1342_),
    .A1(_1298_),
    .Y(_1343_),
    .A2(_1302_));
 sg13g2_nand3_1 _2283_ (.B(_1325_),
    .C(_1343_),
    .A(_1291_),
    .Y(_1344_));
 sg13g2_a22oi_1 _2284_ (.Y(_0001_),
    .B1(_1277_),
    .B2(_1344_),
    .A2(_1273_),
    .A1(_1179_));
 sg13g2_o21ai_1 _2285_ (.B1(_1207_),
    .Y(_1345_),
    .A1(_1044_),
    .A2(_1314_));
 sg13g2_a22oi_1 _2286_ (.Y(_1346_),
    .B1(_1295_),
    .B2(net528),
    .A2(_1097_),
    .A1(_1041_));
 sg13g2_nor2_1 _2287_ (.A(net448),
    .B(_1346_),
    .Y(_1347_));
 sg13g2_o21ai_1 _2288_ (.B1(_1225_),
    .Y(_1348_),
    .A1(_1345_),
    .A2(_1347_));
 sg13g2_or2_1 _2289_ (.X(_1349_),
    .B(_1348_),
    .A(net514));
 sg13g2_nor2_1 _2290_ (.A(_0953_),
    .B(_1066_),
    .Y(_1350_));
 sg13g2_nand2_2 _2291_ (.Y(_1351_),
    .A(_1065_),
    .B(_1071_));
 sg13g2_nand2_1 _2292_ (.Y(_1352_),
    .A(net467),
    .B(_1351_));
 sg13g2_a22oi_1 _2293_ (.Y(_1353_),
    .B1(_1352_),
    .B2(net441),
    .A2(_1212_),
    .A1(_1113_));
 sg13g2_a21oi_1 _2294_ (.A1(_1016_),
    .A2(_1351_),
    .Y(_1354_),
    .B1(_1039_));
 sg13g2_a21oi_1 _2295_ (.A1(net442),
    .A2(_1213_),
    .Y(_1355_),
    .B1(_1211_));
 sg13g2_o21ai_1 _2296_ (.B1(net487),
    .Y(_1356_),
    .A1(_1354_),
    .A2(_1355_));
 sg13g2_a21oi_2 _2297_ (.B1(net481),
    .Y(_1357_),
    .A2(net506),
    .A1(_0961_));
 sg13g2_nand2_1 _2298_ (.Y(_1358_),
    .A(_1207_),
    .B(_1321_));
 sg13g2_inv_1 _2299_ (.Y(_1359_),
    .A(_1358_));
 sg13g2_o21ai_1 _2300_ (.B1(_1359_),
    .Y(_0121_),
    .A1(net448),
    .A2(_1357_));
 sg13g2_o21ai_1 _2301_ (.B1(_1356_),
    .Y(_0122_),
    .A1(_0992_),
    .A2(_1353_));
 sg13g2_a21oi_1 _2302_ (.A1(_0981_),
    .A2(_0121_),
    .Y(_0123_),
    .B1(_0122_));
 sg13g2_a21oi_1 _2303_ (.A1(_1349_),
    .A2(_0123_),
    .Y(_0124_),
    .B1(_1133_));
 sg13g2_a21o_1 _2304_ (.A2(_1262_),
    .A1(_1258_),
    .B1(net473),
    .X(_0125_));
 sg13g2_nand3_1 _2305_ (.B(_1331_),
    .C(_0125_),
    .A(net447),
    .Y(_0126_));
 sg13g2_a21oi_1 _2306_ (.A1(net534),
    .A2(_0126_),
    .Y(_0127_),
    .B1(_1333_));
 sg13g2_nand3_1 _2307_ (.B(_1184_),
    .C(net467),
    .A(net491),
    .Y(_0128_));
 sg13g2_nand2_1 _2308_ (.Y(_0129_),
    .A(net482),
    .B(_0128_));
 sg13g2_a21oi_1 _2309_ (.A1(_1191_),
    .A2(_0129_),
    .Y(_0130_),
    .B1(net534));
 sg13g2_nor2_1 _2310_ (.A(net497),
    .B(_1075_),
    .Y(_0131_));
 sg13g2_o21ai_1 _2311_ (.B1(net481),
    .Y(_0132_),
    .A1(_1337_),
    .A2(_0131_));
 sg13g2_a21oi_1 _2312_ (.A1(_1340_),
    .A2(_0132_),
    .Y(_0133_),
    .B1(_1019_));
 sg13g2_nor2_1 _2313_ (.A(_0130_),
    .B(_0133_),
    .Y(_0134_));
 sg13g2_nor2_1 _2314_ (.A(_0127_),
    .B(_0134_),
    .Y(_0135_));
 sg13g2_nand3_1 _2315_ (.B(_0997_),
    .C(_1169_),
    .A(net529),
    .Y(_0136_));
 sg13g2_nand2_1 _2316_ (.Y(_0137_),
    .A(_1241_),
    .B(_0136_));
 sg13g2_nand3b_1 _2317_ (.B(_1090_),
    .C(net504),
    .Y(_0138_),
    .A_N(_1073_));
 sg13g2_a21oi_1 _2318_ (.A1(net475),
    .A2(_0138_),
    .Y(_0139_),
    .B1(_0137_));
 sg13g2_o21ai_1 _2319_ (.B1(_1298_),
    .Y(_0140_),
    .A1(net510),
    .A2(_0139_));
 sg13g2_a22oi_1 _2320_ (.Y(_0141_),
    .B1(_0140_),
    .B2(_1010_),
    .A2(_0135_),
    .A1(_1049_));
 sg13g2_nor2_1 _2321_ (.A(net498),
    .B(_1090_),
    .Y(_0142_));
 sg13g2_a21oi_2 _2322_ (.B1(_0142_),
    .Y(_0143_),
    .A2(_0961_),
    .A1(_0948_));
 sg13g2_a21oi_1 _2323_ (.A1(_0998_),
    .A2(_0143_),
    .Y(_0144_),
    .B1(_1039_));
 sg13g2_nand3_1 _2324_ (.B(_1211_),
    .C(_1278_),
    .A(_1169_),
    .Y(_0145_));
 sg13g2_or2_1 _2325_ (.X(_0146_),
    .B(_1136_),
    .A(_0972_));
 sg13g2_a221oi_1 _2326_ (.B2(_0146_),
    .C1(_0992_),
    .B1(_1211_),
    .A1(_0974_),
    .Y(_0147_),
    .A2(net442));
 sg13g2_o21ai_1 _2327_ (.B1(net451),
    .Y(_0148_),
    .A1(_1097_),
    .A2(_0142_));
 sg13g2_a21o_1 _2328_ (.A2(_0148_),
    .A1(_1285_),
    .B1(net536),
    .X(_0149_));
 sg13g2_o21ai_1 _2329_ (.B1(net536),
    .Y(_0150_),
    .A1(_1282_),
    .A2(_0144_));
 sg13g2_nand2_1 _2330_ (.Y(_0151_),
    .A(_0149_),
    .B(_0150_));
 sg13g2_a221oi_1 _2331_ (.B2(net510),
    .C1(_0147_),
    .B1(_0151_),
    .A1(net486),
    .Y(_0152_),
    .A2(_0145_));
 sg13g2_o21ai_1 _2332_ (.B1(_0141_),
    .Y(_0153_),
    .A1(_1135_),
    .A2(_0152_));
 sg13g2_o21ai_1 _2333_ (.B1(net457),
    .Y(_0154_),
    .A1(_0124_),
    .A2(_0153_));
 sg13g2_nand3_1 _2334_ (.B(_1017_),
    .C(_1085_),
    .A(net442),
    .Y(_0155_));
 sg13g2_nand2_1 _2335_ (.Y(_0156_),
    .A(_0954_),
    .B(_0972_));
 sg13g2_nand4_1 _2336_ (.B(_0988_),
    .C(_1062_),
    .A(net502),
    .Y(_0157_),
    .D(_1065_));
 sg13g2_o21ai_1 _2337_ (.B1(_0157_),
    .Y(_0158_),
    .A1(_0959_),
    .A2(_1052_));
 sg13g2_a22oi_1 _2338_ (.Y(_0159_),
    .B1(_0158_),
    .B2(net442),
    .A2(_0156_),
    .A1(_0976_));
 sg13g2_a221oi_1 _2339_ (.B2(_1196_),
    .C1(net514),
    .B1(_0159_),
    .A1(_1195_),
    .Y(_0160_),
    .A2(_0155_));
 sg13g2_nor2_2 _2340_ (.A(_1096_),
    .B(net467),
    .Y(_0161_));
 sg13g2_o21ai_1 _2341_ (.B1(net473),
    .Y(_0162_),
    .A1(_1168_),
    .A2(_0161_));
 sg13g2_or2_1 _2342_ (.X(_0163_),
    .B(_0162_),
    .A(net447));
 sg13g2_nand3_1 _2343_ (.B(_1208_),
    .C(_0163_),
    .A(_1207_),
    .Y(_0164_));
 sg13g2_a22oi_1 _2344_ (.Y(_0165_),
    .B1(_1136_),
    .B2(_0946_),
    .A2(_1124_),
    .A1(net490));
 sg13g2_o21ai_1 _2345_ (.B1(_1191_),
    .Y(_0166_),
    .A1(net472),
    .A2(_0165_));
 sg13g2_a21oi_1 _2346_ (.A1(_1215_),
    .A2(_0162_),
    .Y(_0167_),
    .B1(net521));
 sg13g2_a221oi_1 _2347_ (.B2(_0167_),
    .C1(_0160_),
    .B1(_0166_),
    .A1(net487),
    .Y(_0168_),
    .A2(_0164_));
 sg13g2_a221oi_1 _2348_ (.B2(_1236_),
    .C1(net531),
    .B1(_1228_),
    .A1(net440),
    .Y(_0169_),
    .A2(_1187_));
 sg13g2_o21ai_1 _2349_ (.B1(net508),
    .Y(_0170_),
    .A1(_1227_),
    .A2(_0169_));
 sg13g2_nor2_1 _2350_ (.A(_1040_),
    .B(_1137_),
    .Y(_0171_));
 sg13g2_or3_1 _2351_ (.A(net453),
    .B(_1240_),
    .C(_0171_),
    .X(_0172_));
 sg13g2_a221oi_1 _2352_ (.B2(_1308_),
    .C1(_1221_),
    .B1(_1095_),
    .A1(_0964_),
    .Y(_0173_),
    .A2(_1071_));
 sg13g2_o21ai_1 _2353_ (.B1(_0172_),
    .Y(_0174_),
    .A1(net445),
    .A2(_0173_));
 sg13g2_a21oi_1 _2354_ (.A1(_1142_),
    .A2(net467),
    .Y(_0175_),
    .B1(net477));
 sg13g2_nand2_1 _2355_ (.Y(_0176_),
    .A(net468),
    .B(_0175_));
 sg13g2_o21ai_1 _2356_ (.B1(net486),
    .Y(_0177_),
    .A1(net452),
    .A2(_1188_));
 sg13g2_a21oi_1 _2357_ (.A1(_1231_),
    .A2(_0176_),
    .Y(_0178_),
    .B1(_0177_));
 sg13g2_a21oi_1 _2358_ (.A1(net489),
    .A2(_0174_),
    .Y(_0179_),
    .B1(_0178_));
 sg13g2_a21oi_1 _2359_ (.A1(_0170_),
    .A2(_0179_),
    .Y(_0180_),
    .B1(_1050_));
 sg13g2_o21ai_1 _2360_ (.B1(net479),
    .Y(_0181_),
    .A1(_0947_),
    .A2(_0973_));
 sg13g2_o21ai_1 _2361_ (.B1(net471),
    .Y(_0182_),
    .A1(_1183_),
    .A2(_1213_));
 sg13g2_nand2_1 _2362_ (.Y(_0183_),
    .A(_0181_),
    .B(_0182_));
 sg13g2_o21ai_1 _2363_ (.B1(net508),
    .Y(_0184_),
    .A1(_1251_),
    .A2(_0183_));
 sg13g2_a221oi_1 _2364_ (.B2(_1139_),
    .C1(_1260_),
    .B1(_1117_),
    .A1(_0941_),
    .Y(_0185_),
    .A2(_0986_));
 sg13g2_or2_1 _2365_ (.X(_0186_),
    .B(_0185_),
    .A(net512));
 sg13g2_nand2_1 _2366_ (.Y(_0187_),
    .A(_1263_),
    .B(_1351_));
 sg13g2_nor2_1 _2367_ (.A(net477),
    .B(net521),
    .Y(_0188_));
 sg13g2_o21ai_1 _2368_ (.B1(_1000_),
    .Y(_0189_),
    .A1(_0955_),
    .A2(_1116_));
 sg13g2_a21oi_1 _2369_ (.A1(net501),
    .A2(_1001_),
    .Y(_0190_),
    .B1(_1014_));
 sg13g2_nand2_1 _2370_ (.Y(_0191_),
    .A(net488),
    .B(_1226_));
 sg13g2_a221oi_1 _2371_ (.B2(_0190_),
    .C1(_0191_),
    .B1(_0189_),
    .A1(_0187_),
    .Y(_0192_),
    .A2(_0188_));
 sg13g2_a221oi_1 _2372_ (.B2(_0192_),
    .C1(_1006_),
    .B1(_0186_),
    .A1(_1248_),
    .Y(_0193_),
    .A2(_0184_));
 sg13g2_nor3_2 _2373_ (.A(net457),
    .B(_0180_),
    .C(_0193_),
    .Y(_0194_));
 sg13g2_o21ai_1 _2374_ (.B1(_0194_),
    .Y(_0195_),
    .A1(net444),
    .A2(_0168_));
 sg13g2_o21ai_1 _2375_ (.B1(_0195_),
    .Y(_0196_),
    .A1(_1108_),
    .A2(_1177_));
 sg13g2_a22oi_1 _2376_ (.Y(_0002_),
    .B1(_0196_),
    .B2(_1105_),
    .A2(_0154_),
    .A1(_1277_));
 sg13g2_a21oi_1 _2377_ (.A1(net516),
    .A2(_1071_),
    .Y(_0197_),
    .B1(net445));
 sg13g2_nand2b_1 _2378_ (.Y(_0198_),
    .B(_0990_),
    .A_N(_1069_));
 sg13g2_nand2_1 _2379_ (.Y(_0199_),
    .A(_1237_),
    .B(_0198_));
 sg13g2_a21oi_1 _2380_ (.A1(_1031_),
    .A2(_1040_),
    .Y(_0200_),
    .B1(_0990_));
 sg13g2_a21o_1 _2381_ (.A2(_1213_),
    .A1(net492),
    .B1(_1190_),
    .X(_0201_));
 sg13g2_nand3_1 _2382_ (.B(_1076_),
    .C(net467),
    .A(net443),
    .Y(_0202_));
 sg13g2_nand3_1 _2383_ (.B(_0201_),
    .C(_0202_),
    .A(net486),
    .Y(_0203_));
 sg13g2_nand3_1 _2384_ (.B(_0957_),
    .C(_1136_),
    .A(net446),
    .Y(_0204_));
 sg13g2_a22oi_1 _2385_ (.Y(_0205_),
    .B1(_1308_),
    .B2(net492),
    .A2(_1071_),
    .A1(_0964_));
 sg13g2_or2_1 _2386_ (.X(_0206_),
    .B(_0205_),
    .A(net477));
 sg13g2_a21oi_1 _2387_ (.A1(_1036_),
    .A2(_0206_),
    .Y(_0207_),
    .B1(net521));
 sg13g2_a22oi_1 _2388_ (.Y(_0208_),
    .B1(_0197_),
    .B2(_0200_),
    .A2(_1183_),
    .A1(net440));
 sg13g2_nand2_1 _2389_ (.Y(_0209_),
    .A(net532),
    .B(_0208_));
 sg13g2_mux2_1 _2390_ (.A0(_0197_),
    .A1(_1055_),
    .S(_0199_),
    .X(_0210_));
 sg13g2_o21ai_1 _2391_ (.B1(_0209_),
    .Y(_0211_),
    .A1(net532),
    .A2(_0210_));
 sg13g2_a22oi_1 _2392_ (.Y(_0212_),
    .B1(_0211_),
    .B2(net508),
    .A2(_0207_),
    .A1(_0204_));
 sg13g2_a21oi_1 _2393_ (.A1(_0203_),
    .A2(_0212_),
    .Y(_0213_),
    .B1(_1050_));
 sg13g2_o21ai_1 _2394_ (.B1(_1190_),
    .Y(_0214_),
    .A1(_1232_),
    .A2(_0175_));
 sg13g2_nand3_1 _2395_ (.B(net440),
    .C(net467),
    .A(_1003_),
    .Y(_0215_));
 sg13g2_nand3_1 _2396_ (.B(_0214_),
    .C(_0215_),
    .A(_0981_),
    .Y(_0216_));
 sg13g2_nand2b_1 _2397_ (.Y(_0217_),
    .B(_1136_),
    .A_N(_1087_));
 sg13g2_nand2_1 _2398_ (.Y(_0218_),
    .A(_0952_),
    .B(_0969_));
 sg13g2_xnor2_1 _2399_ (.Y(_0219_),
    .A(_0217_),
    .B(_0218_));
 sg13g2_nor2_1 _2400_ (.A(net528),
    .B(_1189_),
    .Y(_0220_));
 sg13g2_o21ai_1 _2401_ (.B1(_0220_),
    .Y(_0221_),
    .A1(net472),
    .A2(_0219_));
 sg13g2_nor2_1 _2402_ (.A(net534),
    .B(_1201_),
    .Y(_0222_));
 sg13g2_a21oi_1 _2403_ (.A1(_1205_),
    .A2(_0222_),
    .Y(_0223_),
    .B1(net454));
 sg13g2_o21ai_1 _2404_ (.B1(net535),
    .Y(_0224_),
    .A1(_1168_),
    .A2(_1193_));
 sg13g2_o21ai_1 _2405_ (.B1(_0224_),
    .Y(_0225_),
    .A1(_0957_),
    .A2(_0998_));
 sg13g2_nand3_1 _2406_ (.B(net528),
    .C(_1214_),
    .A(_0976_),
    .Y(_0226_));
 sg13g2_a221oi_1 _2407_ (.B2(net454),
    .C1(net509),
    .B1(_0225_),
    .A1(_0221_),
    .Y(_0227_),
    .A2(_0223_));
 sg13g2_o21ai_1 _2408_ (.B1(_0941_),
    .Y(_0228_),
    .A1(net506),
    .A2(_1115_));
 sg13g2_o21ai_1 _2409_ (.B1(_0228_),
    .Y(_0229_),
    .A1(net481),
    .A2(_0969_));
 sg13g2_o21ai_1 _2410_ (.B1(net482),
    .Y(_0230_),
    .A1(_1124_),
    .A2(_1183_));
 sg13g2_o21ai_1 _2411_ (.B1(_1191_),
    .Y(_0231_),
    .A1(_0986_),
    .A2(_0230_));
 sg13g2_o21ai_1 _2412_ (.B1(_0231_),
    .Y(_0232_),
    .A1(_1194_),
    .A2(_0229_));
 sg13g2_a221oi_1 _2413_ (.B2(_1019_),
    .C1(net444),
    .B1(_0232_),
    .A1(_0226_),
    .Y(_0233_),
    .A2(_0227_));
 sg13g2_nor3_1 _2414_ (.A(net477),
    .B(_0961_),
    .C(_1124_),
    .Y(_0234_));
 sg13g2_nor3_1 _2415_ (.A(net527),
    .B(_1024_),
    .C(_0234_),
    .Y(_0235_));
 sg13g2_nand2_2 _2416_ (.Y(_0236_),
    .A(net500),
    .B(_0952_));
 sg13g2_nand3_1 _2417_ (.B(_1092_),
    .C(_0236_),
    .A(net471),
    .Y(_0237_));
 sg13g2_a21oi_1 _2418_ (.A1(_0198_),
    .A2(_0237_),
    .Y(_0238_),
    .B1(net531));
 sg13g2_nor3_1 _2419_ (.A(net445),
    .B(_0235_),
    .C(_0238_),
    .Y(_0239_));
 sg13g2_o21ai_1 _2420_ (.B1(_1248_),
    .Y(_0240_),
    .A1(net513),
    .A2(_0239_));
 sg13g2_o21ai_1 _2421_ (.B1(net471),
    .Y(_0241_),
    .A1(_1141_),
    .A2(_1350_));
 sg13g2_nand2_1 _2422_ (.Y(_0242_),
    .A(_1204_),
    .B(_1266_));
 sg13g2_a21oi_1 _2423_ (.A1(_1139_),
    .A2(_0242_),
    .Y(_0243_),
    .B1(_1255_));
 sg13g2_a21oi_1 _2424_ (.A1(_0241_),
    .A2(_0243_),
    .Y(_0244_),
    .B1(net508));
 sg13g2_o21ai_1 _2425_ (.B1(net471),
    .Y(_0245_),
    .A1(_1257_),
    .A2(_1308_));
 sg13g2_nor2_1 _2426_ (.A(net526),
    .B(_0995_),
    .Y(_0246_));
 sg13g2_a21oi_2 _2427_ (.B1(net484),
    .Y(_0247_),
    .A2(_1086_),
    .A1(_1025_));
 sg13g2_nand2_1 _2428_ (.Y(_0248_),
    .A(_1092_),
    .B(_0247_));
 sg13g2_a221oi_1 _2429_ (.B2(net526),
    .C1(net512),
    .B1(_0248_),
    .A1(_0245_),
    .Y(_0249_),
    .A2(_0246_));
 sg13g2_nor3_1 _2430_ (.A(_0191_),
    .B(_0244_),
    .C(_0249_),
    .Y(_0250_));
 sg13g2_nor2_1 _2431_ (.A(_1006_),
    .B(_0250_),
    .Y(_0251_));
 sg13g2_a221oi_1 _2432_ (.B2(_0251_),
    .C1(net457),
    .B1(_0240_),
    .A1(_0216_),
    .Y(_0252_),
    .A2(_0233_));
 sg13g2_nor2b_2 _2433_ (.A(_0213_),
    .B_N(_0252_),
    .Y(_0253_));
 sg13g2_nand2b_1 _2434_ (.Y(_0254_),
    .B(_0982_),
    .A_N(_1176_));
 sg13g2_o21ai_1 _2435_ (.B1(_1105_),
    .Y(_0255_),
    .A1(_1108_),
    .A2(_0254_));
 sg13g2_o21ai_1 _2436_ (.B1(_1155_),
    .Y(_0256_),
    .A1(_1042_),
    .A2(_1295_));
 sg13g2_nand3_1 _2437_ (.B(_0952_),
    .C(_0988_),
    .A(net496),
    .Y(_0257_));
 sg13g2_a21o_1 _2438_ (.A2(_0257_),
    .A1(_1031_),
    .B1(net527),
    .X(_0258_));
 sg13g2_nand3_1 _2439_ (.B(_0256_),
    .C(_0258_),
    .A(net452),
    .Y(_0259_));
 sg13g2_a21oi_1 _2440_ (.A1(_1090_),
    .A2(_1261_),
    .Y(_0260_),
    .B1(net528));
 sg13g2_a21oi_1 _2441_ (.A1(_1351_),
    .A2(_0260_),
    .Y(_0261_),
    .B1(net472));
 sg13g2_nand4_1 _2442_ (.B(_1035_),
    .C(_1263_),
    .A(net528),
    .Y(_0262_),
    .D(_1266_));
 sg13g2_a221oi_1 _2443_ (.B2(_0262_),
    .C1(net515),
    .B1(_0261_),
    .A1(_1212_),
    .Y(_0263_),
    .A2(_0259_));
 sg13g2_o21ai_1 _2444_ (.B1(net467),
    .Y(_0264_),
    .A1(_0955_),
    .A2(_1116_));
 sg13g2_nand2_1 _2445_ (.Y(_0265_),
    .A(net478),
    .B(_0264_));
 sg13g2_nor3_1 _2446_ (.A(net481),
    .B(_0967_),
    .C(_1125_),
    .Y(_0266_));
 sg13g2_o21ai_1 _2447_ (.B1(_0265_),
    .Y(_0267_),
    .A1(net449),
    .A2(_0266_));
 sg13g2_a221oi_1 _2448_ (.B2(net535),
    .C1(_1307_),
    .B1(_0267_),
    .A1(net449),
    .Y(_0268_),
    .A2(_1357_));
 sg13g2_o21ai_1 _2449_ (.B1(_1007_),
    .Y(_0269_),
    .A1(_0263_),
    .A2(_0268_));
 sg13g2_o21ai_1 _2450_ (.B1(net481),
    .Y(_0270_),
    .A1(_1141_),
    .A2(_1327_));
 sg13g2_nor2_1 _2451_ (.A(net535),
    .B(_1189_),
    .Y(_0271_));
 sg13g2_a22oi_1 _2452_ (.Y(_0272_),
    .B1(_0270_),
    .B2(_0271_),
    .A2(_1339_),
    .A1(_1202_));
 sg13g2_nand3_1 _2453_ (.B(_1026_),
    .C(_1185_),
    .A(net483),
    .Y(_0273_));
 sg13g2_nand2_1 _2454_ (.Y(_0274_),
    .A(_1331_),
    .B(_0273_));
 sg13g2_o21ai_1 _2455_ (.B1(net489),
    .Y(_0275_),
    .A1(_1188_),
    .A2(_1334_));
 sg13g2_nand2_1 _2456_ (.Y(_0276_),
    .A(_1049_),
    .B(_0275_));
 sg13g2_a221oi_1 _2457_ (.B2(net487),
    .C1(_0276_),
    .B1(_0274_),
    .A1(net509),
    .Y(_0277_),
    .A2(_0272_));
 sg13g2_a22oi_1 _2458_ (.Y(_0278_),
    .B1(_1137_),
    .B2(_0975_),
    .A2(_1075_),
    .A1(net474));
 sg13g2_o21ai_1 _2459_ (.B1(net536),
    .Y(_0279_),
    .A1(_0974_),
    .A2(_1295_));
 sg13g2_nor2_1 _2460_ (.A(_0278_),
    .B(_0279_),
    .Y(_0280_));
 sg13g2_a21oi_1 _2461_ (.A1(_1109_),
    .A2(_1293_),
    .Y(_0281_),
    .B1(_0280_));
 sg13g2_a22oi_1 _2462_ (.Y(_0282_),
    .B1(_1017_),
    .B2(_0975_),
    .A2(net507),
    .A1(net474));
 sg13g2_a21oi_1 _2463_ (.A1(_1015_),
    .A2(_1169_),
    .Y(_0283_),
    .B1(net484));
 sg13g2_nor3_1 _2464_ (.A(_1299_),
    .B(_0282_),
    .C(_0283_),
    .Y(_0284_));
 sg13g2_o21ai_1 _2465_ (.B1(_1008_),
    .Y(_0285_),
    .A1(net509),
    .A2(_0284_));
 sg13g2_a21oi_1 _2466_ (.A1(net509),
    .A2(_0281_),
    .Y(_0286_),
    .B1(_0285_));
 sg13g2_o21ai_1 _2467_ (.B1(net450),
    .Y(_0287_),
    .A1(_0277_),
    .A2(_0286_));
 sg13g2_and3_1 _2468_ (.X(_0288_),
    .A(_1135_),
    .B(_0269_),
    .C(_0287_));
 sg13g2_and3_1 _2469_ (.X(_0289_),
    .A(net450),
    .B(_1026_),
    .C(_1278_));
 sg13g2_o21ai_1 _2470_ (.B1(_1207_),
    .Y(_0290_),
    .A1(_1114_),
    .A2(_0289_));
 sg13g2_nor2_1 _2471_ (.A(_1095_),
    .B(_1113_),
    .Y(_0291_));
 sg13g2_o21ai_1 _2472_ (.B1(_1021_),
    .Y(_0292_),
    .A1(_0959_),
    .A2(_0236_));
 sg13g2_nor3_1 _2473_ (.A(net535),
    .B(_1212_),
    .C(_0292_),
    .Y(_0293_));
 sg13g2_a21oi_1 _2474_ (.A1(_1016_),
    .A2(_1266_),
    .Y(_0294_),
    .B1(net472));
 sg13g2_nor4_1 _2475_ (.A(net455),
    .B(net528),
    .C(_1357_),
    .D(_0294_),
    .Y(_0295_));
 sg13g2_nor4_1 _2476_ (.A(net515),
    .B(_0291_),
    .C(_0293_),
    .D(_0295_),
    .Y(_0296_));
 sg13g2_o21ai_1 _2477_ (.B1(_1091_),
    .Y(_0297_),
    .A1(_1001_),
    .A2(_1017_));
 sg13g2_nand2_1 _2478_ (.Y(_0298_),
    .A(net450),
    .B(_0297_));
 sg13g2_a221oi_1 _2479_ (.B2(net486),
    .C1(_0296_),
    .B1(_0298_),
    .A1(net515),
    .Y(_0299_),
    .A2(_0290_));
 sg13g2_o21ai_1 _2480_ (.B1(net458),
    .Y(_0300_),
    .A1(_1135_),
    .A2(_0299_));
 sg13g2_nand3_1 _2481_ (.B(_0946_),
    .C(net489),
    .A(net498),
    .Y(_0301_));
 sg13g2_a22oi_1 _2482_ (.Y(_0302_),
    .B1(_1274_),
    .B2(_0301_),
    .A2(net491),
    .A1(net503));
 sg13g2_nand4_1 _2483_ (.B(_1091_),
    .C(_1167_),
    .A(net450),
    .Y(_0303_),
    .D(_0302_));
 sg13g2_and2_1 _2484_ (.A(_1106_),
    .B(_0303_),
    .X(_0304_));
 sg13g2_o21ai_1 _2485_ (.B1(_0304_),
    .Y(_0305_),
    .A1(_0288_),
    .A2(_0300_));
 sg13g2_o21ai_1 _2486_ (.B1(_0305_),
    .Y(_0003_),
    .A1(_0253_),
    .A2(_0255_));
 sg13g2_a21oi_1 _2487_ (.A1(_0997_),
    .A2(_0143_),
    .Y(_0306_),
    .B1(_1039_));
 sg13g2_o21ai_1 _2488_ (.B1(net536),
    .Y(_0307_),
    .A1(_1282_),
    .A2(_0306_));
 sg13g2_nand3_1 _2489_ (.B(_0149_),
    .C(_0307_),
    .A(net510),
    .Y(_0308_));
 sg13g2_a21oi_1 _2490_ (.A1(_1280_),
    .A2(_0308_),
    .Y(_0309_),
    .B1(_0147_));
 sg13g2_nor2_1 _2491_ (.A(_1135_),
    .B(_0309_),
    .Y(_0310_));
 sg13g2_nor3_1 _2492_ (.A(net534),
    .B(_1316_),
    .C(_1345_),
    .Y(_0311_));
 sg13g2_a21oi_1 _2493_ (.A1(_1041_),
    .A2(_1097_),
    .Y(_0312_),
    .B1(_1202_));
 sg13g2_o21ai_1 _2494_ (.B1(net534),
    .Y(_0313_),
    .A1(net448),
    .A2(_0312_));
 sg13g2_o21ai_1 _2495_ (.B1(net510),
    .Y(_0314_),
    .A1(_1358_),
    .A2(_0313_));
 sg13g2_nor2_1 _2496_ (.A(_0311_),
    .B(_0314_),
    .Y(_0315_));
 sg13g2_o21ai_1 _2497_ (.B1(_1086_),
    .Y(_0316_),
    .A1(_1020_),
    .A2(_1025_));
 sg13g2_a22oi_1 _2498_ (.Y(_0317_),
    .B1(_0316_),
    .B2(net441),
    .A2(_1212_),
    .A1(_1113_));
 sg13g2_o21ai_1 _2499_ (.B1(_1356_),
    .Y(_0318_),
    .A1(_0992_),
    .A2(_0317_));
 sg13g2_o21ai_1 _2500_ (.B1(_1132_),
    .Y(_0319_),
    .A1(_0315_),
    .A2(_0318_));
 sg13g2_o21ai_1 _2501_ (.B1(net514),
    .Y(_0320_),
    .A1(_0137_),
    .A2(_0247_));
 sg13g2_a21o_1 _2502_ (.A2(_0320_),
    .A1(_1298_),
    .B1(net444),
    .X(_0321_));
 sg13g2_a21oi_1 _2503_ (.A1(_1326_),
    .A2(_0125_),
    .Y(_0322_),
    .B1(net528));
 sg13g2_a21oi_1 _2504_ (.A1(_1326_),
    .A2(_0129_),
    .Y(_0323_),
    .B1(net534));
 sg13g2_nor2_1 _2505_ (.A(_0133_),
    .B(_0323_),
    .Y(_0324_));
 sg13g2_nor2_1 _2506_ (.A(_1050_),
    .B(_0324_),
    .Y(_0325_));
 sg13g2_o21ai_1 _2507_ (.B1(_0325_),
    .Y(_0326_),
    .A1(_1333_),
    .A2(_0322_));
 sg13g2_nand3_1 _2508_ (.B(_0321_),
    .C(_0326_),
    .A(_0319_),
    .Y(_0327_));
 sg13g2_o21ai_1 _2509_ (.B1(net457),
    .Y(_0328_),
    .A1(_0310_),
    .A2(_0327_));
 sg13g2_nand3_1 _2510_ (.B(_0956_),
    .C(_1158_),
    .A(net474),
    .Y(_0329_));
 sg13g2_o21ai_1 _2511_ (.B1(_0329_),
    .Y(_0330_),
    .A1(net483),
    .A2(_0157_));
 sg13g2_o21ai_1 _2512_ (.B1(net455),
    .Y(_0331_),
    .A1(_1091_),
    .A2(_0330_));
 sg13g2_a221oi_1 _2513_ (.B2(_0331_),
    .C1(net514),
    .B1(_1196_),
    .A1(_1182_),
    .Y(_0332_),
    .A2(_1195_));
 sg13g2_nor3_1 _2514_ (.A(net473),
    .B(net455),
    .C(_0165_),
    .Y(_0333_));
 sg13g2_nand2b_1 _2515_ (.Y(_0334_),
    .B(_1216_),
    .A_N(_0333_));
 sg13g2_a21oi_1 _2516_ (.A1(_0991_),
    .A2(_0334_),
    .Y(_0335_),
    .B1(_0332_));
 sg13g2_a21oi_1 _2517_ (.A1(_1210_),
    .A2(_0335_),
    .Y(_0336_),
    .B1(net444));
 sg13g2_a21oi_1 _2518_ (.A1(_1252_),
    .A2(_0181_),
    .Y(_0337_),
    .B1(net512));
 sg13g2_o21ai_1 _2519_ (.B1(_1132_),
    .Y(_0338_),
    .A1(_1247_),
    .A2(_0337_));
 sg13g2_nor2b_1 _2520_ (.A(_1118_),
    .B_N(_1139_),
    .Y(_0339_));
 sg13g2_nor3_1 _2521_ (.A(_1245_),
    .B(_1260_),
    .C(_0339_),
    .Y(_0340_));
 sg13g2_a21oi_1 _2522_ (.A1(_1256_),
    .A2(_0340_),
    .Y(_0341_),
    .B1(net512));
 sg13g2_nand3b_1 _2523_ (.B(_0236_),
    .C(_1226_),
    .Y(_0342_),
    .A_N(_0161_));
 sg13g2_o21ai_1 _2524_ (.B1(_0996_),
    .Y(_0343_),
    .A1(net476),
    .A2(_1304_));
 sg13g2_a221oi_1 _2525_ (.B2(net489),
    .C1(_0341_),
    .B1(_0343_),
    .A1(net486),
    .Y(_0344_),
    .A2(_0342_));
 sg13g2_o21ai_1 _2526_ (.B1(_0338_),
    .Y(_0345_),
    .A1(_1135_),
    .A2(_0344_));
 sg13g2_nand2b_1 _2527_ (.Y(_0346_),
    .B(_0172_),
    .A_N(_1239_));
 sg13g2_nand2_1 _2528_ (.Y(_0347_),
    .A(net468),
    .B(_1197_));
 sg13g2_a21oi_1 _2529_ (.A1(_1231_),
    .A2(_0347_),
    .Y(_0348_),
    .B1(_0177_));
 sg13g2_a21oi_1 _2530_ (.A1(net489),
    .A2(_0346_),
    .Y(_0349_),
    .B1(_0348_));
 sg13g2_a21oi_2 _2531_ (.B1(_1050_),
    .Y(_0350_),
    .A2(_0349_),
    .A1(_1230_));
 sg13g2_nor3_1 _2532_ (.A(_0336_),
    .B(_0345_),
    .C(_0350_),
    .Y(_0351_));
 sg13g2_nand2b_1 _2533_ (.Y(_0352_),
    .B(_0936_),
    .A_N(_0351_));
 sg13g2_a22oi_1 _2534_ (.Y(_0004_),
    .B1(_0352_),
    .B2(_1179_),
    .A2(_0328_),
    .A1(_1277_));
 sg13g2_and2_1 _2535_ (.A(net566),
    .B(\wrapper.h_count[1] ),
    .X(_0353_));
 sg13g2_nand3_1 _2536_ (.B(net565),
    .C(_0353_),
    .A(\wrapper.h_count[3] ),
    .Y(_0354_));
 sg13g2_inv_1 _2537_ (.Y(_0355_),
    .A(_0354_));
 sg13g2_nor4_1 _2538_ (.A(net564),
    .B(_0629_),
    .C(net561),
    .D(net563),
    .Y(_0356_));
 sg13g2_nand4_1 _2539_ (.B(\wrapper.h_count[9] ),
    .C(_0355_),
    .A(\wrapper.h_count[8] ),
    .Y(_0357_),
    .D(_0356_));
 sg13g2_and2_1 _2540_ (.A(net577),
    .B(_0357_),
    .X(_0358_));
 sg13g2_nand2_2 _2541_ (.Y(_0359_),
    .A(net579),
    .B(_0357_));
 sg13g2_and2_1 _2542_ (.A(net123),
    .B(net466),
    .X(_0028_));
 sg13g2_nor2_1 _2543_ (.A(net566),
    .B(net221),
    .Y(_0360_));
 sg13g2_nor3_1 _2544_ (.A(_0628_),
    .B(_0353_),
    .C(net222),
    .Y(_0029_));
 sg13g2_o21ai_1 _2545_ (.B1(net577),
    .Y(_0361_),
    .A1(net565),
    .A2(_0353_));
 sg13g2_a21oi_1 _2546_ (.A1(net565),
    .A2(_0353_),
    .Y(_0030_),
    .B1(_0361_));
 sg13g2_a21oi_1 _2547_ (.A1(net565),
    .A2(_0353_),
    .Y(_0362_),
    .B1(net205));
 sg13g2_nor3_1 _2548_ (.A(net571),
    .B(_0355_),
    .C(net206),
    .Y(_0031_));
 sg13g2_xnor2_1 _2549_ (.Y(_0363_),
    .A(_0629_),
    .B(_0354_));
 sg13g2_nor2_1 _2550_ (.A(_0359_),
    .B(_0363_),
    .Y(_0032_));
 sg13g2_nor2_1 _2551_ (.A(net179),
    .B(_0354_),
    .Y(_0364_));
 sg13g2_xnor2_1 _2552_ (.Y(_0365_),
    .A(net564),
    .B(_0364_));
 sg13g2_nor2_1 _2553_ (.A(_0359_),
    .B(net180),
    .Y(_0033_));
 sg13g2_nand2_1 _2554_ (.Y(_0366_),
    .A(net564),
    .B(\wrapper.h_count[4] ));
 sg13g2_nor2_1 _2555_ (.A(_0354_),
    .B(_0366_),
    .Y(_0367_));
 sg13g2_o21ai_1 _2556_ (.B1(net466),
    .Y(_0368_),
    .A1(net563),
    .A2(_0367_));
 sg13g2_a21oi_1 _2557_ (.A1(net563),
    .A2(_0367_),
    .Y(_0034_),
    .B1(_0368_));
 sg13g2_nor3_1 _2558_ (.A(net195),
    .B(_0354_),
    .C(_0366_),
    .Y(_0369_));
 sg13g2_o21ai_1 _2559_ (.B1(_0358_),
    .Y(_0370_),
    .A1(net561),
    .A2(_0369_));
 sg13g2_a21oi_1 _2560_ (.A1(net561),
    .A2(_0369_),
    .Y(_0035_),
    .B1(_0370_));
 sg13g2_nand4_1 _2561_ (.B(\wrapper.h_count[4] ),
    .C(net561),
    .A(net564),
    .Y(_0371_),
    .D(net563));
 sg13g2_nor2_1 _2562_ (.A(_0354_),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_nor2_1 _2563_ (.A(net208),
    .B(_0372_),
    .Y(_0373_));
 sg13g2_and2_1 _2564_ (.A(net208),
    .B(_0372_),
    .X(_0374_));
 sg13g2_nor3_1 _2565_ (.A(_0359_),
    .B(_0373_),
    .C(_0374_),
    .Y(_0036_));
 sg13g2_o21ai_1 _2566_ (.B1(_0358_),
    .Y(_0375_),
    .A1(net190),
    .A2(_0374_));
 sg13g2_a21oi_1 _2567_ (.A1(net190),
    .A2(_0374_),
    .Y(_0037_),
    .B1(_0375_));
 sg13g2_xor2_1 _2568_ (.B(\wrapper.pixel.prev_y[9] ),
    .A(\wrapper.pixel.vpos[9] ),
    .X(_0376_));
 sg13g2_nand2b_1 _2569_ (.Y(_0377_),
    .B(\wrapper.pixel.prev_y[6] ),
    .A_N(net540));
 sg13g2_nor2_1 _2570_ (.A(net548),
    .B(_0630_),
    .Y(_0378_));
 sg13g2_nand2b_1 _2571_ (.Y(_0379_),
    .B(net551),
    .A_N(\wrapper.pixel.prev_y[0] ));
 sg13g2_nand2b_1 _2572_ (.Y(_0380_),
    .B(net544),
    .A_N(\wrapper.pixel.prev_y[3] ));
 sg13g2_o21ai_1 _2573_ (.B1(_0377_),
    .Y(_0381_),
    .A1(_0602_),
    .A2(\wrapper.pixel.prev_y[8] ));
 sg13g2_xor2_1 _2574_ (.B(\wrapper.pixel.prev_y[7] ),
    .A(\wrapper.pixel.vpos[7] ),
    .X(_0382_));
 sg13g2_xor2_1 _2575_ (.B(\wrapper.pixel.prev_y[2] ),
    .A(net546),
    .X(_0383_));
 sg13g2_nor4_1 _2576_ (.A(_0378_),
    .B(_0381_),
    .C(_0382_),
    .D(_0383_),
    .Y(_0384_));
 sg13g2_xor2_1 _2577_ (.B(\wrapper.pixel.prev_y[4] ),
    .A(net542),
    .X(_0385_));
 sg13g2_a22oi_1 _2578_ (.Y(_0386_),
    .B1(_0632_),
    .B2(net540),
    .A2(\wrapper.pixel.prev_y[0] ),
    .A1(_0606_));
 sg13g2_o21ai_1 _2579_ (.B1(_0386_),
    .Y(_0387_),
    .A1(_0604_),
    .A2(\wrapper.pixel.prev_y[5] ));
 sg13g2_a22oi_1 _2580_ (.Y(_0388_),
    .B1(\wrapper.pixel.prev_y[5] ),
    .B2(_0604_),
    .A2(_0630_),
    .A1(net548));
 sg13g2_a22oi_1 _2581_ (.Y(_0389_),
    .B1(\wrapper.pixel.prev_y[8] ),
    .B2(_0602_),
    .A2(\wrapper.pixel.prev_y[3] ),
    .A1(_0605_));
 sg13g2_nand4_1 _2582_ (.B(_0380_),
    .C(_0388_),
    .A(_0379_),
    .Y(_0390_),
    .D(_0389_));
 sg13g2_nor4_1 _2583_ (.A(_0376_),
    .B(_0385_),
    .C(_0387_),
    .D(_0390_),
    .Y(_0391_));
 sg13g2_nor4_1 _2584_ (.A(\wrapper.pixel.vpos[7] ),
    .B(net540),
    .C(net541),
    .D(net542),
    .Y(_0392_));
 sg13g2_nor2_1 _2585_ (.A(net548),
    .B(net551),
    .Y(_0393_));
 sg13g2_nor4_1 _2586_ (.A(\wrapper.pixel.vpos[9] ),
    .B(\wrapper.pixel.vpos[8] ),
    .C(net544),
    .D(net546),
    .Y(_0394_));
 sg13g2_nand3_1 _2587_ (.B(_0393_),
    .C(_0394_),
    .A(_0392_),
    .Y(_0395_));
 sg13g2_a21o_1 _2588_ (.A2(_0391_),
    .A1(_0384_),
    .B1(_0395_),
    .X(_0396_));
 sg13g2_nor4_1 _2589_ (.A(\wrapper.pixel.sprite_top[9] ),
    .B(\wrapper.pixel.sprite_top[6] ),
    .C(\wrapper.pixel.sprite_top[5] ),
    .D(_0613_),
    .Y(_0397_));
 sg13g2_nor2_1 _2590_ (.A(net553),
    .B(\wrapper.pixel.sprite_top[8] ),
    .Y(_0398_));
 sg13g2_or2_1 _2591_ (.X(_0399_),
    .B(\wrapper.pixel.sprite_top[2] ),
    .A(\wrapper.pixel.sprite_top[3] ));
 sg13g2_nor3_1 _2592_ (.A(\wrapper.pixel.sprite_top[7] ),
    .B(\wrapper.pixel.sprite_top[1] ),
    .C(_0399_),
    .Y(_0400_));
 sg13g2_nand3_1 _2593_ (.B(_0398_),
    .C(_0400_),
    .A(_0610_),
    .Y(_0401_));
 sg13g2_nand3_1 _2594_ (.B(\wrapper.pixel.sprite_top[2] ),
    .C(\wrapper.pixel.sprite_top[1] ),
    .A(\wrapper.pixel.sprite_top[3] ),
    .Y(_0402_));
 sg13g2_nand4_1 _2595_ (.B(\wrapper.pixel.sprite_top[8] ),
    .C(\wrapper.pixel.sprite_top[7] ),
    .A(net554),
    .Y(_0403_),
    .D(\wrapper.pixel.sprite_top[4] ));
 sg13g2_o21ai_1 _2596_ (.B1(_0401_),
    .Y(_0404_),
    .A1(_0402_),
    .A2(_0403_));
 sg13g2_nand3b_1 _2597_ (.B(_0397_),
    .C(_0404_),
    .Y(_0405_),
    .A_N(net461));
 sg13g2_inv_2 _2598_ (.Y(_0406_),
    .A(_0405_));
 sg13g2_or3_1 _2599_ (.A(\wrapper.pixel.sprite_left[8] ),
    .B(\wrapper.pixel.sprite_left[7] ),
    .C(\wrapper.pixel.sprite_left[6] ),
    .X(_0407_));
 sg13g2_or2_1 _2600_ (.X(_0408_),
    .B(\wrapper.pixel.sprite_left[2] ),
    .A(\wrapper.pixel.sprite_left[3] ));
 sg13g2_nor3_1 _2601_ (.A(\wrapper.pixel.sprite_left[5] ),
    .B(\wrapper.pixel.sprite_left[4] ),
    .C(\wrapper.pixel.sprite_left[1] ),
    .Y(_0409_));
 sg13g2_nor3_1 _2602_ (.A(net557),
    .B(\wrapper.pixel.sprite_left[9] ),
    .C(_0408_),
    .Y(_0410_));
 sg13g2_nand4_1 _2603_ (.B(\wrapper.pixel.sprite_left[5] ),
    .C(\wrapper.pixel.sprite_left[3] ),
    .A(\wrapper.pixel.sprite_left[9] ),
    .Y(_0411_),
    .D(\wrapper.pixel.sprite_left[1] ));
 sg13g2_nor3_1 _2604_ (.A(_0608_),
    .B(_0616_),
    .C(_0411_),
    .Y(_0412_));
 sg13g2_a22oi_1 _2605_ (.Y(_0413_),
    .B1(_0412_),
    .B2(\wrapper.pixel.sprite_left[2] ),
    .A2(_0410_),
    .A1(_0409_));
 sg13g2_nor4_2 _2606_ (.A(_0618_),
    .B(net464),
    .C(_0407_),
    .Y(_0414_),
    .D(_0413_));
 sg13g2_nor2_2 _2607_ (.A(_0406_),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_o21ai_1 _2608_ (.B1(net583),
    .Y(_0416_),
    .A1(net134),
    .A2(_0415_));
 sg13g2_a21oi_1 _2609_ (.A1(_0627_),
    .A2(_0415_),
    .Y(_0038_),
    .B1(_0416_));
 sg13g2_nor2_1 _2610_ (.A(_0627_),
    .B(_0415_),
    .Y(_0417_));
 sg13g2_o21ai_1 _2611_ (.B1(net583),
    .Y(_0418_),
    .A1(net189),
    .A2(_0417_));
 sg13g2_nand2_1 _2612_ (.Y(_0419_),
    .A(net189),
    .B(_0417_));
 sg13g2_nor2b_1 _2613_ (.A(_0418_),
    .B_N(_0419_),
    .Y(_0039_));
 sg13g2_nand2b_1 _2614_ (.Y(_0420_),
    .B(_0419_),
    .A_N(net186));
 sg13g2_nand3_1 _2615_ (.B(net189),
    .C(_0417_),
    .A(net186),
    .Y(_0421_));
 sg13g2_and3_1 _2616_ (.X(_0040_),
    .A(net582),
    .B(_0420_),
    .C(_0421_));
 sg13g2_o21ai_1 _2617_ (.B1(net582),
    .Y(_0422_),
    .A1(_0626_),
    .A2(_0421_));
 sg13g2_a21oi_1 _2618_ (.A1(_0626_),
    .A2(_0421_),
    .Y(_0041_),
    .B1(_0422_));
 sg13g2_xor2_1 _2619_ (.B(net184),
    .A(net175),
    .X(_0423_));
 sg13g2_xor2_1 _2620_ (.B(net163),
    .A(\wrapper.pixel.lfsr_reg[15] ),
    .X(_0424_));
 sg13g2_a21oi_1 _2621_ (.A1(_0423_),
    .A2(_0424_),
    .Y(_0425_),
    .B1(net571));
 sg13g2_o21ai_1 _2622_ (.B1(_0425_),
    .Y(_0042_),
    .A1(_0423_),
    .A2(_0424_));
 sg13g2_and2_1 _2623_ (.A(net582),
    .B(net126),
    .X(_0043_));
 sg13g2_and2_1 _2624_ (.A(net583),
    .B(net131),
    .X(_0044_));
 sg13g2_and2_1 _2625_ (.A(net583),
    .B(net129),
    .X(_0045_));
 sg13g2_and2_1 _2626_ (.A(net583),
    .B(net124),
    .X(_0046_));
 sg13g2_and2_1 _2627_ (.A(net580),
    .B(net125),
    .X(_0047_));
 sg13g2_and2_1 _2628_ (.A(net580),
    .B(net132),
    .X(_0048_));
 sg13g2_and2_1 _2629_ (.A(net580),
    .B(net130),
    .X(_0049_));
 sg13g2_and2_1 _2630_ (.A(net580),
    .B(net133),
    .X(_0050_));
 sg13g2_and2_1 _2631_ (.A(net580),
    .B(net128),
    .X(_0051_));
 sg13g2_and2_1 _2632_ (.A(net580),
    .B(net127),
    .X(_0052_));
 sg13g2_and2_1 _2633_ (.A(net581),
    .B(net140),
    .X(_0053_));
 sg13g2_and2_1 _2634_ (.A(net581),
    .B(net149),
    .X(_0054_));
 sg13g2_and2_1 _2635_ (.A(net581),
    .B(net163),
    .X(_0055_));
 sg13g2_and2_1 _2636_ (.A(net584),
    .B(net175),
    .X(_0056_));
 sg13g2_and2_1 _2637_ (.A(net582),
    .B(net160),
    .X(_0057_));
 sg13g2_o21ai_1 _2638_ (.B1(net582),
    .Y(_0426_),
    .A1(\wrapper.pixel.background_state[0] ),
    .A2(net572));
 sg13g2_nor2b_1 _2639_ (.A(net573),
    .B_N(net1),
    .Y(_0427_));
 sg13g2_a21oi_1 _2640_ (.A1(net177),
    .A2(net7),
    .Y(_0428_),
    .B1(_0427_));
 sg13g2_a21oi_1 _2641_ (.A1(net572),
    .A2(_0428_),
    .Y(_0058_),
    .B1(_0426_));
 sg13g2_o21ai_1 _2642_ (.B1(net582),
    .Y(_0429_),
    .A1(net173),
    .A2(net572));
 sg13g2_nor2b_1 _2643_ (.A(net573),
    .B_N(net2),
    .Y(_0430_));
 sg13g2_a21oi_1 _2644_ (.A1(\wrapper.pixel.looping_background_count[1] ),
    .A2(net573),
    .Y(_0431_),
    .B1(_0430_));
 sg13g2_a21oi_1 _2645_ (.A1(net572),
    .A2(_0431_),
    .Y(_0059_),
    .B1(_0429_));
 sg13g2_o21ai_1 _2646_ (.B1(net582),
    .Y(_0432_),
    .A1(\wrapper.pixel.background_state[2] ),
    .A2(net572));
 sg13g2_nor2b_1 _2647_ (.A(net573),
    .B_N(net3),
    .Y(_0433_));
 sg13g2_a21oi_1 _2648_ (.A1(net186),
    .A2(net573),
    .Y(_0434_),
    .B1(_0433_));
 sg13g2_a21oi_1 _2649_ (.A1(net572),
    .A2(_0434_),
    .Y(_0060_),
    .B1(_0432_));
 sg13g2_o21ai_1 _2650_ (.B1(net582),
    .Y(_0435_),
    .A1(net182),
    .A2(net572));
 sg13g2_nor2b_1 _2651_ (.A(net573),
    .B_N(net4),
    .Y(_0436_));
 sg13g2_a21oi_1 _2652_ (.A1(net156),
    .A2(net573),
    .Y(_0437_),
    .B1(_0436_));
 sg13g2_a21oi_1 _2653_ (.A1(net572),
    .A2(_0437_),
    .Y(_0061_),
    .B1(_0435_));
 sg13g2_nor2_1 _2654_ (.A(net573),
    .B(net8),
    .Y(_0438_));
 sg13g2_a21oi_1 _2655_ (.A1(net1),
    .A2(net568),
    .Y(_0439_),
    .B1(net571));
 sg13g2_o21ai_1 _2656_ (.B1(_0439_),
    .Y(_0062_),
    .A1(_0624_),
    .A2(net568));
 sg13g2_a21oi_1 _2657_ (.A1(net2),
    .A2(net568),
    .Y(_0440_),
    .B1(net571));
 sg13g2_o21ai_1 _2658_ (.B1(_0440_),
    .Y(_0063_),
    .A1(_0623_),
    .A2(net567));
 sg13g2_a21oi_1 _2659_ (.A1(net3),
    .A2(net567),
    .Y(_0441_),
    .B1(net570));
 sg13g2_o21ai_1 _2660_ (.B1(_0441_),
    .Y(_0064_),
    .A1(_0622_),
    .A2(net568));
 sg13g2_a21oi_1 _2661_ (.A1(net4),
    .A2(net567),
    .Y(_0442_),
    .B1(net570));
 sg13g2_o21ai_1 _2662_ (.B1(_0442_),
    .Y(_0065_),
    .A1(_0621_),
    .A2(net567));
 sg13g2_a21oi_1 _2663_ (.A1(net5),
    .A2(net567),
    .Y(_0443_),
    .B1(net570));
 sg13g2_o21ai_1 _2664_ (.B1(_0443_),
    .Y(_0066_),
    .A1(_0620_),
    .A2(net567));
 sg13g2_a21oi_1 _2665_ (.A1(net6),
    .A2(net567),
    .Y(_0444_),
    .B1(net570));
 sg13g2_o21ai_1 _2666_ (.B1(_0444_),
    .Y(_0067_),
    .A1(_0619_),
    .A2(net567));
 sg13g2_o21ai_1 _2667_ (.B1(net579),
    .Y(_0445_),
    .A1(net164),
    .A2(net464));
 sg13g2_a21oi_1 _2668_ (.A1(_0618_),
    .A2(net464),
    .Y(_0068_),
    .B1(_0445_));
 sg13g2_xor2_1 _2669_ (.B(\wrapper.pixel.sprite_left[1] ),
    .A(net557),
    .X(_0446_));
 sg13g2_xnor2_1 _2670_ (.Y(_0447_),
    .A(net164),
    .B(_0446_));
 sg13g2_a21oi_1 _2671_ (.A1(net172),
    .A2(net465),
    .Y(_0448_),
    .B1(net571));
 sg13g2_o21ai_1 _2672_ (.B1(_0448_),
    .Y(_0069_),
    .A1(net465),
    .A2(_0447_));
 sg13g2_xor2_1 _2673_ (.B(\wrapper.pixel.sprite_left[2] ),
    .A(net555),
    .X(_0449_));
 sg13g2_a21o_1 _2674_ (.A2(\wrapper.pixel.sprite_left[1] ),
    .A1(_0608_),
    .B1(\wrapper.pixel.sprite_left[0] ),
    .X(_0450_));
 sg13g2_o21ai_1 _2675_ (.B1(_0450_),
    .Y(_0451_),
    .A1(_0608_),
    .A2(\wrapper.pixel.sprite_left[1] ));
 sg13g2_nor2_1 _2676_ (.A(_0449_),
    .B(_0451_),
    .Y(_0452_));
 sg13g2_xor2_1 _2677_ (.B(_0451_),
    .A(_0449_),
    .X(_0453_));
 sg13g2_o21ai_1 _2678_ (.B1(net579),
    .Y(_0454_),
    .A1(net462),
    .A2(_0453_));
 sg13g2_a21oi_1 _2679_ (.A1(_0617_),
    .A2(net462),
    .Y(_0070_),
    .B1(_0454_));
 sg13g2_nand2b_1 _2680_ (.Y(_0455_),
    .B(net555),
    .A_N(\wrapper.pixel.sprite_left[3] ));
 sg13g2_xor2_1 _2681_ (.B(\wrapper.pixel.sprite_left[3] ),
    .A(net555),
    .X(_0456_));
 sg13g2_a21oi_1 _2682_ (.A1(_0608_),
    .A2(\wrapper.pixel.sprite_left[2] ),
    .Y(_0457_),
    .B1(_0452_));
 sg13g2_xnor2_1 _2683_ (.Y(_0458_),
    .A(_0456_),
    .B(_0457_));
 sg13g2_a21oi_1 _2684_ (.A1(net223),
    .A2(net462),
    .Y(_0459_),
    .B1(net570));
 sg13g2_o21ai_1 _2685_ (.B1(_0459_),
    .Y(_0071_),
    .A1(net462),
    .A2(_0458_));
 sg13g2_xor2_1 _2686_ (.B(\wrapper.pixel.sprite_left[4] ),
    .A(net555),
    .X(_0460_));
 sg13g2_a22oi_1 _2687_ (.Y(_0461_),
    .B1(_0452_),
    .B2(_0455_),
    .A2(_0408_),
    .A1(_0608_));
 sg13g2_or2_1 _2688_ (.X(_0462_),
    .B(_0461_),
    .A(_0460_));
 sg13g2_a21oi_1 _2689_ (.A1(_0460_),
    .A2(_0461_),
    .Y(_0463_),
    .B1(net462));
 sg13g2_a22oi_1 _2690_ (.Y(_0464_),
    .B1(_0462_),
    .B2(_0463_),
    .A2(net462),
    .A1(net220));
 sg13g2_nand2_1 _2691_ (.Y(_0072_),
    .A(net584),
    .B(_0464_));
 sg13g2_a21oi_1 _2692_ (.A1(net200),
    .A2(net462),
    .Y(_0465_),
    .B1(net570));
 sg13g2_xor2_1 _2693_ (.B(\wrapper.pixel.sprite_left[5] ),
    .A(net556),
    .X(_0466_));
 sg13g2_o21ai_1 _2694_ (.B1(_0462_),
    .Y(_0467_),
    .A1(net556),
    .A2(_0616_));
 sg13g2_xor2_1 _2695_ (.B(_0467_),
    .A(_0466_),
    .X(_0468_));
 sg13g2_o21ai_1 _2696_ (.B1(_0465_),
    .Y(_0073_),
    .A1(net462),
    .A2(_0468_));
 sg13g2_nand2_1 _2697_ (.Y(_0469_),
    .A(_0608_),
    .B(\wrapper.pixel.sprite_left[6] ));
 sg13g2_xor2_1 _2698_ (.B(\wrapper.pixel.sprite_left[6] ),
    .A(net555),
    .X(_0470_));
 sg13g2_nor2_1 _2699_ (.A(_0462_),
    .B(_0466_),
    .Y(_0471_));
 sg13g2_a21oi_1 _2700_ (.A1(_0615_),
    .A2(_0616_),
    .Y(_0472_),
    .B1(net557));
 sg13g2_nor2_1 _2701_ (.A(_0471_),
    .B(_0472_),
    .Y(_0473_));
 sg13g2_nand2_1 _2702_ (.Y(_0474_),
    .A(net207),
    .B(net463));
 sg13g2_a21oi_1 _2703_ (.A1(_0470_),
    .A2(_0473_),
    .Y(_0475_),
    .B1(net463));
 sg13g2_o21ai_1 _2704_ (.B1(_0475_),
    .Y(_0476_),
    .A1(_0470_),
    .A2(_0473_));
 sg13g2_nand3_1 _2705_ (.B(_0474_),
    .C(_0476_),
    .A(net579),
    .Y(_0074_));
 sg13g2_a21oi_1 _2706_ (.A1(net201),
    .A2(net463),
    .Y(_0477_),
    .B1(net570));
 sg13g2_xor2_1 _2707_ (.B(\wrapper.pixel.sprite_left[7] ),
    .A(net555),
    .X(_0478_));
 sg13g2_o21ai_1 _2708_ (.B1(_0469_),
    .Y(_0479_),
    .A1(_0470_),
    .A2(_0473_));
 sg13g2_xor2_1 _2709_ (.B(_0479_),
    .A(_0478_),
    .X(_0480_));
 sg13g2_o21ai_1 _2710_ (.B1(_0477_),
    .Y(_0075_),
    .A1(net463),
    .A2(_0480_));
 sg13g2_nor4_1 _2711_ (.A(_0462_),
    .B(_0466_),
    .C(_0470_),
    .D(_0478_),
    .Y(_0481_));
 sg13g2_o21ai_1 _2712_ (.B1(_0469_),
    .Y(_0482_),
    .A1(net557),
    .A2(_0614_));
 sg13g2_nor3_2 _2713_ (.A(_0472_),
    .B(_0481_),
    .C(_0482_),
    .Y(_0483_));
 sg13g2_xnor2_1 _2714_ (.Y(_0484_),
    .A(net555),
    .B(\wrapper.pixel.sprite_left[8] ));
 sg13g2_xnor2_1 _2715_ (.Y(_0485_),
    .A(_0483_),
    .B(_0484_));
 sg13g2_nand2b_1 _2716_ (.Y(_0486_),
    .B(net463),
    .A_N(net226));
 sg13g2_o21ai_1 _2717_ (.B1(_0486_),
    .Y(_0487_),
    .A1(net463),
    .A2(_0485_));
 sg13g2_nor2_1 _2718_ (.A(net570),
    .B(_0487_),
    .Y(_0076_));
 sg13g2_a21oi_1 _2719_ (.A1(net556),
    .A2(\wrapper.pixel.sprite_left[8] ),
    .Y(_0488_),
    .B1(_0483_));
 sg13g2_o21ai_1 _2720_ (.B1(_0483_),
    .Y(_0489_),
    .A1(net556),
    .A2(\wrapper.pixel.sprite_left[8] ));
 sg13g2_inv_1 _2721_ (.Y(_0490_),
    .A(_0489_));
 sg13g2_nor3_1 _2722_ (.A(net463),
    .B(_0488_),
    .C(_0490_),
    .Y(_0491_));
 sg13g2_o21ai_1 _2723_ (.B1(net579),
    .Y(_0492_),
    .A1(net188),
    .A2(_0491_));
 sg13g2_a21oi_1 _2724_ (.A1(net188),
    .A2(_0491_),
    .Y(_0077_),
    .B1(_0492_));
 sg13g2_o21ai_1 _2725_ (.B1(net576),
    .Y(_0493_),
    .A1(net166),
    .A2(net461));
 sg13g2_a21oi_1 _2726_ (.A1(_0613_),
    .A2(net461),
    .Y(_0078_),
    .B1(_0493_));
 sg13g2_xor2_1 _2727_ (.B(\wrapper.pixel.sprite_top[1] ),
    .A(net554),
    .X(_0494_));
 sg13g2_xnor2_1 _2728_ (.Y(_0495_),
    .A(net166),
    .B(_0494_));
 sg13g2_a21oi_1 _2729_ (.A1(net176),
    .A2(net461),
    .Y(_0496_),
    .B1(net569));
 sg13g2_o21ai_1 _2730_ (.B1(_0496_),
    .Y(_0079_),
    .A1(net461),
    .A2(_0495_));
 sg13g2_xor2_1 _2731_ (.B(\wrapper.pixel.sprite_top[2] ),
    .A(net552),
    .X(_0497_));
 sg13g2_o21ai_1 _2732_ (.B1(_0613_),
    .Y(_0498_),
    .A1(net554),
    .A2(_0612_));
 sg13g2_o21ai_1 _2733_ (.B1(_0498_),
    .Y(_0499_),
    .A1(_0607_),
    .A2(\wrapper.pixel.sprite_top[1] ));
 sg13g2_nor2_1 _2734_ (.A(_0497_),
    .B(_0499_),
    .Y(_0500_));
 sg13g2_xor2_1 _2735_ (.B(_0499_),
    .A(_0497_),
    .X(_0501_));
 sg13g2_o21ai_1 _2736_ (.B1(net576),
    .Y(_0502_),
    .A1(net459),
    .A2(_0501_));
 sg13g2_a21oi_1 _2737_ (.A1(_0611_),
    .A2(net459),
    .Y(_0080_),
    .B1(_0502_));
 sg13g2_nand2b_1 _2738_ (.Y(_0503_),
    .B(net552),
    .A_N(\wrapper.pixel.sprite_top[3] ));
 sg13g2_xor2_1 _2739_ (.B(\wrapper.pixel.sprite_top[3] ),
    .A(net552),
    .X(_0504_));
 sg13g2_a21oi_1 _2740_ (.A1(_0607_),
    .A2(\wrapper.pixel.sprite_top[2] ),
    .Y(_0505_),
    .B1(_0500_));
 sg13g2_xnor2_1 _2741_ (.Y(_0506_),
    .A(_0504_),
    .B(_0505_));
 sg13g2_a21oi_1 _2742_ (.A1(net210),
    .A2(net459),
    .Y(_0507_),
    .B1(net569));
 sg13g2_o21ai_1 _2743_ (.B1(_0507_),
    .Y(_0081_),
    .A1(net459),
    .A2(_0506_));
 sg13g2_xnor2_1 _2744_ (.Y(_0508_),
    .A(net552),
    .B(\wrapper.pixel.sprite_top[4] ));
 sg13g2_inv_1 _2745_ (.Y(_0509_),
    .A(_0508_));
 sg13g2_a22oi_1 _2746_ (.Y(_0510_),
    .B1(_0500_),
    .B2(_0503_),
    .A2(_0399_),
    .A1(_0607_));
 sg13g2_nand2b_1 _2747_ (.Y(_0511_),
    .B(_0508_),
    .A_N(_0510_));
 sg13g2_a21oi_1 _2748_ (.A1(_0509_),
    .A2(_0510_),
    .Y(_0512_),
    .B1(net459));
 sg13g2_a22oi_1 _2749_ (.Y(_0513_),
    .B1(_0511_),
    .B2(_0512_),
    .A2(net459),
    .A1(net217));
 sg13g2_nand2_1 _2750_ (.Y(_0082_),
    .A(net576),
    .B(_0513_));
 sg13g2_a21oi_1 _2751_ (.A1(net224),
    .A2(net459),
    .Y(_0514_),
    .B1(net569));
 sg13g2_xor2_1 _2752_ (.B(\wrapper.pixel.sprite_top[5] ),
    .A(net552),
    .X(_0515_));
 sg13g2_o21ai_1 _2753_ (.B1(_0511_),
    .Y(_0516_),
    .A1(net552),
    .A2(_0610_));
 sg13g2_xor2_1 _2754_ (.B(_0516_),
    .A(_0515_),
    .X(_0517_));
 sg13g2_o21ai_1 _2755_ (.B1(_0514_),
    .Y(_0083_),
    .A1(net459),
    .A2(_0517_));
 sg13g2_nand2_1 _2756_ (.Y(_0518_),
    .A(_0607_),
    .B(\wrapper.pixel.sprite_top[6] ));
 sg13g2_xor2_1 _2757_ (.B(\wrapper.pixel.sprite_top[6] ),
    .A(net553),
    .X(_0519_));
 sg13g2_or2_1 _2758_ (.X(_0520_),
    .B(_0515_),
    .A(_0511_));
 sg13g2_o21ai_1 _2759_ (.B1(_0607_),
    .Y(_0521_),
    .A1(\wrapper.pixel.sprite_top[5] ),
    .A2(\wrapper.pixel.sprite_top[4] ));
 sg13g2_and2_1 _2760_ (.A(_0520_),
    .B(_0521_),
    .X(_0522_));
 sg13g2_nand2_1 _2761_ (.Y(_0523_),
    .A(net212),
    .B(net460));
 sg13g2_a21oi_1 _2762_ (.A1(_0519_),
    .A2(_0522_),
    .Y(_0524_),
    .B1(net460));
 sg13g2_o21ai_1 _2763_ (.B1(_0524_),
    .Y(_0525_),
    .A1(_0519_),
    .A2(_0522_));
 sg13g2_nand3_1 _2764_ (.B(_0523_),
    .C(_0525_),
    .A(net576),
    .Y(_0084_));
 sg13g2_a21oi_1 _2765_ (.A1(net216),
    .A2(net460),
    .Y(_0526_),
    .B1(net569));
 sg13g2_xor2_1 _2766_ (.B(\wrapper.pixel.sprite_top[7] ),
    .A(net553),
    .X(_0527_));
 sg13g2_o21ai_1 _2767_ (.B1(_0518_),
    .Y(_0528_),
    .A1(_0519_),
    .A2(_0522_));
 sg13g2_xor2_1 _2768_ (.B(_0528_),
    .A(_0527_),
    .X(_0529_));
 sg13g2_o21ai_1 _2769_ (.B1(_0526_),
    .Y(_0085_),
    .A1(net460),
    .A2(_0529_));
 sg13g2_nor3_1 _2770_ (.A(_0519_),
    .B(_0520_),
    .C(_0527_),
    .Y(_0530_));
 sg13g2_o21ai_1 _2771_ (.B1(_0607_),
    .Y(_0531_),
    .A1(\wrapper.pixel.sprite_top[7] ),
    .A2(\wrapper.pixel.sprite_top[6] ));
 sg13g2_nand2_1 _2772_ (.Y(_0532_),
    .A(_0521_),
    .B(_0531_));
 sg13g2_nor2_1 _2773_ (.A(_0530_),
    .B(_0532_),
    .Y(_0533_));
 sg13g2_xnor2_1 _2774_ (.Y(_0534_),
    .A(net553),
    .B(\wrapper.pixel.sprite_top[8] ));
 sg13g2_xnor2_1 _2775_ (.Y(_0535_),
    .A(_0533_),
    .B(_0534_));
 sg13g2_nand2b_1 _2776_ (.Y(_0536_),
    .B(net460),
    .A_N(net225));
 sg13g2_o21ai_1 _2777_ (.B1(_0536_),
    .Y(_0537_),
    .A1(net460),
    .A2(_0535_));
 sg13g2_nor2_1 _2778_ (.A(net569),
    .B(_0537_),
    .Y(_0086_));
 sg13g2_nor3_1 _2779_ (.A(_0398_),
    .B(_0530_),
    .C(_0532_),
    .Y(_0538_));
 sg13g2_a21oi_1 _2780_ (.A1(net552),
    .A2(\wrapper.pixel.sprite_top[8] ),
    .Y(_0539_),
    .B1(_0533_));
 sg13g2_nor3_1 _2781_ (.A(net460),
    .B(_0538_),
    .C(_0539_),
    .Y(_0540_));
 sg13g2_o21ai_1 _2782_ (.B1(net576),
    .Y(_0541_),
    .A1(net155),
    .A2(_0540_));
 sg13g2_a21oi_1 _2783_ (.A1(net155),
    .A2(_0540_),
    .Y(_0087_),
    .B1(_0541_));
 sg13g2_nand2b_1 _2784_ (.Y(_0542_),
    .B(net555),
    .A_N(_0414_));
 sg13g2_nand3_1 _2785_ (.B(net146),
    .C(_0414_),
    .A(_0608_),
    .Y(_0543_));
 sg13g2_nand3_1 _2786_ (.B(_0542_),
    .C(_0543_),
    .A(net579),
    .Y(_0088_));
 sg13g2_a21oi_1 _2787_ (.A1(_0607_),
    .A2(net136),
    .Y(_0544_),
    .B1(_0405_));
 sg13g2_o21ai_1 _2788_ (.B1(net576),
    .Y(_0545_),
    .A1(net554),
    .A2(_0406_));
 sg13g2_nor2_1 _2789_ (.A(_0544_),
    .B(_0545_),
    .Y(_0089_));
 sg13g2_and2_1 _2790_ (.A(net585),
    .B(_0023_),
    .X(_0090_));
 sg13g2_nor2_1 _2791_ (.A(net569),
    .B(_0740_),
    .Y(_0091_));
 sg13g2_xor2_1 _2792_ (.B(_0739_),
    .A(\wrapper.pixel.moving_counter[2] ),
    .X(_0546_));
 sg13g2_nor2_1 _2793_ (.A(net569),
    .B(_0546_),
    .Y(_0092_));
 sg13g2_nor2_1 _2794_ (.A(_0011_),
    .B(_0739_),
    .Y(_0547_));
 sg13g2_o21ai_1 _2795_ (.B1(net578),
    .Y(_0548_),
    .A1(\wrapper.pixel.moving_counter[3] ),
    .A2(_0547_));
 sg13g2_a21oi_1 _2796_ (.A1(\wrapper.pixel.moving_counter[3] ),
    .A2(_0547_),
    .Y(_0093_),
    .B1(_0548_));
 sg13g2_nand4_1 _2797_ (.B(\wrapper.pixel.moving_counter[2] ),
    .C(\wrapper.pixel.moving_counter[0] ),
    .A(\wrapper.pixel.moving_counter[3] ),
    .Y(_0549_),
    .D(\wrapper.pixel.moving_counter[1] ));
 sg13g2_inv_1 _2798_ (.Y(_0550_),
    .A(_0549_));
 sg13g2_o21ai_1 _2799_ (.B1(net578),
    .Y(_0551_),
    .A1(_0634_),
    .A2(_0549_));
 sg13g2_a21oi_1 _2800_ (.A1(_0634_),
    .A2(_0549_),
    .Y(_0094_),
    .B1(_0551_));
 sg13g2_nor2_1 _2801_ (.A(_0009_),
    .B(_0549_),
    .Y(_0552_));
 sg13g2_o21ai_1 _2802_ (.B1(net578),
    .Y(_0553_),
    .A1(\wrapper.pixel.moving_counter[5] ),
    .A2(_0552_));
 sg13g2_a21oi_1 _2803_ (.A1(\wrapper.pixel.moving_counter[5] ),
    .A2(_0552_),
    .Y(_0095_),
    .B1(_0553_));
 sg13g2_nand3_1 _2804_ (.B(\wrapper.pixel.moving_counter[5] ),
    .C(_0550_),
    .A(\wrapper.pixel.moving_counter[4] ),
    .Y(_0554_));
 sg13g2_o21ai_1 _2805_ (.B1(net580),
    .Y(_0555_),
    .A1(_0635_),
    .A2(_0554_));
 sg13g2_a21oi_1 _2806_ (.A1(_0635_),
    .A2(_0554_),
    .Y(_0096_),
    .B1(_0555_));
 sg13g2_nor2_1 _2807_ (.A(_0017_),
    .B(_0554_),
    .Y(_0556_));
 sg13g2_o21ai_1 _2808_ (.B1(net580),
    .Y(_0557_),
    .A1(\wrapper.pixel.moving_counter[7] ),
    .A2(_0556_));
 sg13g2_a21oi_1 _2809_ (.A1(\wrapper.pixel.moving_counter[7] ),
    .A2(_0556_),
    .Y(_0097_),
    .B1(_0557_));
 sg13g2_nor4_1 _2810_ (.A(net457),
    .B(_0982_),
    .C(_0989_),
    .D(net444),
    .Y(_0558_));
 sg13g2_nand3_1 _2811_ (.B(_1105_),
    .C(_0558_),
    .A(_0976_),
    .Y(_0098_));
 sg13g2_mux2_1 _2812_ (.A0(net158),
    .A1(net551),
    .S(net578),
    .X(_0099_));
 sg13g2_mux2_1 _2813_ (.A0(net145),
    .A1(net548),
    .S(net578),
    .X(_0100_));
 sg13g2_nand2_1 _2814_ (.Y(_0559_),
    .A(net546),
    .B(net578));
 sg13g2_o21ai_1 _2815_ (.B1(_0559_),
    .Y(_0101_),
    .A1(net578),
    .A2(_0631_));
 sg13g2_nor2_1 _2816_ (.A(net575),
    .B(net151),
    .Y(_0560_));
 sg13g2_a21oi_1 _2817_ (.A1(_0605_),
    .A2(net575),
    .Y(_0102_),
    .B1(_0560_));
 sg13g2_mux2_1 _2818_ (.A0(net154),
    .A1(net542),
    .S(net574),
    .X(_0103_));
 sg13g2_mux2_1 _2819_ (.A0(net170),
    .A1(net541),
    .S(net575),
    .X(_0104_));
 sg13g2_mux2_1 _2820_ (.A0(net150),
    .A1(net540),
    .S(net578),
    .X(_0105_));
 sg13g2_nor2_1 _2821_ (.A(net575),
    .B(net153),
    .Y(_0561_));
 sg13g2_a21oi_1 _2822_ (.A1(_0603_),
    .A2(net574),
    .Y(_0106_),
    .B1(_0561_));
 sg13g2_nor2_1 _2823_ (.A(net574),
    .B(net143),
    .Y(_0562_));
 sg13g2_a21oi_1 _2824_ (.A1(_0602_),
    .A2(net574),
    .Y(_0107_),
    .B1(_0562_));
 sg13g2_nor2_1 _2825_ (.A(net574),
    .B(net141),
    .Y(_0563_));
 sg13g2_a21oi_1 _2826_ (.A1(_0601_),
    .A2(net574),
    .Y(_0108_),
    .B1(_0563_));
 sg13g2_nand4_1 _2827_ (.B(net546),
    .C(_0392_),
    .A(\wrapper.pixel.vpos[9] ),
    .Y(_0564_),
    .D(_0393_));
 sg13g2_nor3_1 _2828_ (.A(\wrapper.pixel.vpos[8] ),
    .B(_0605_),
    .C(_0564_),
    .Y(_0565_));
 sg13g2_nor3_2 _2829_ (.A(net569),
    .B(_0357_),
    .C(_0565_),
    .Y(_0566_));
 sg13g2_nor2_1 _2830_ (.A(net550),
    .B(_0566_),
    .Y(_0567_));
 sg13g2_a21oi_1 _2831_ (.A1(net550),
    .A2(_0359_),
    .Y(_0109_),
    .B1(_0567_));
 sg13g2_a21oi_1 _2832_ (.A1(net550),
    .A2(_0359_),
    .Y(_0568_),
    .B1(net138));
 sg13g2_nand2_1 _2833_ (.Y(_0569_),
    .A(net549),
    .B(net550));
 sg13g2_o21ai_1 _2834_ (.B1(net577),
    .Y(_0570_),
    .A1(_0357_),
    .A2(_0569_));
 sg13g2_nor2_1 _2835_ (.A(net139),
    .B(_0570_),
    .Y(_0110_));
 sg13g2_xor2_1 _2836_ (.B(_0569_),
    .A(net202),
    .X(_0571_));
 sg13g2_a22oi_1 _2837_ (.Y(_0572_),
    .B1(_0566_),
    .B2(_0571_),
    .A2(net466),
    .A1(net547));
 sg13g2_inv_1 _2838_ (.Y(_0111_),
    .A(net203));
 sg13g2_nand3_1 _2839_ (.B(net548),
    .C(net551),
    .A(net546),
    .Y(_0573_));
 sg13g2_nor2_1 _2840_ (.A(_0605_),
    .B(_0573_),
    .Y(_0574_));
 sg13g2_xnor2_1 _2841_ (.Y(_0575_),
    .A(net544),
    .B(_0573_));
 sg13g2_a22oi_1 _2842_ (.Y(_0576_),
    .B1(_0566_),
    .B2(_0575_),
    .A2(net466),
    .A1(net544));
 sg13g2_inv_1 _2843_ (.Y(_0112_),
    .A(_0576_));
 sg13g2_nor2b_1 _2844_ (.A(_0357_),
    .B_N(_0574_),
    .Y(_0577_));
 sg13g2_and2_2 _2845_ (.A(net542),
    .B(_0574_),
    .X(_0578_));
 sg13g2_o21ai_1 _2846_ (.B1(net574),
    .Y(_0579_),
    .A1(net542),
    .A2(_0577_));
 sg13g2_a21oi_1 _2847_ (.A1(net542),
    .A2(_0577_),
    .Y(_0113_),
    .B1(_0579_));
 sg13g2_xnor2_1 _2848_ (.Y(_0580_),
    .A(net198),
    .B(_0578_));
 sg13g2_a22oi_1 _2849_ (.Y(_0581_),
    .B1(_0566_),
    .B2(_0580_),
    .A2(net466),
    .A1(net541));
 sg13g2_inv_1 _2850_ (.Y(_0114_),
    .A(net199));
 sg13g2_nand2_1 _2851_ (.Y(_0582_),
    .A(net541),
    .B(_0578_));
 sg13g2_or2_1 _2852_ (.X(_0583_),
    .B(_0582_),
    .A(_0018_));
 sg13g2_nand2_1 _2853_ (.Y(_0584_),
    .A(_0566_),
    .B(_0583_));
 sg13g2_a21oi_1 _2854_ (.A1(_0018_),
    .A2(_0582_),
    .Y(_0585_),
    .B1(_0584_));
 sg13g2_a21o_1 _2855_ (.A2(net466),
    .A1(net196),
    .B1(_0585_),
    .X(_0115_));
 sg13g2_xor2_1 _2856_ (.B(_0583_),
    .A(net192),
    .X(_0586_));
 sg13g2_a22oi_1 _2857_ (.Y(_0587_),
    .B1(_0566_),
    .B2(net193),
    .A2(net466),
    .A1(\wrapper.pixel.vpos[7] ));
 sg13g2_inv_1 _2858_ (.Y(_0116_),
    .A(net194));
 sg13g2_nand4_1 _2859_ (.B(net542),
    .C(_0804_),
    .A(net540),
    .Y(_0588_),
    .D(_0577_));
 sg13g2_nand2b_1 _2860_ (.Y(_0589_),
    .B(_0578_),
    .A_N(_0805_));
 sg13g2_o21ai_1 _2861_ (.B1(net574),
    .Y(_0590_),
    .A1(_0357_),
    .A2(_0589_));
 sg13g2_a21oi_1 _2862_ (.A1(_0602_),
    .A2(_0588_),
    .Y(_0117_),
    .B1(_0590_));
 sg13g2_a21oi_1 _2863_ (.A1(_0566_),
    .A2(_0589_),
    .Y(_0591_),
    .B1(net466));
 sg13g2_nor2_1 _2864_ (.A(net219),
    .B(_0805_),
    .Y(_0592_));
 sg13g2_nand3_1 _2865_ (.B(_0578_),
    .C(_0592_),
    .A(_0566_),
    .Y(_0593_));
 sg13g2_o21ai_1 _2866_ (.B1(_0593_),
    .Y(_0118_),
    .A1(_0601_),
    .A2(_0591_));
 sg13g2_nor3_1 _2867_ (.A(net542),
    .B(_0605_),
    .C(net546),
    .Y(_0594_));
 sg13g2_nand3_1 _2868_ (.B(_0592_),
    .C(_0594_),
    .A(net548),
    .Y(_0595_));
 sg13g2_nand2_1 _2869_ (.Y(_0119_),
    .A(net577),
    .B(_0595_));
 sg13g2_nor3_1 _2870_ (.A(net564),
    .B(\wrapper.h_count[4] ),
    .C(net563),
    .Y(_0596_));
 sg13g2_nor2b_1 _2871_ (.A(_0596_),
    .B_N(\wrapper.h_count[9] ),
    .Y(_0597_));
 sg13g2_a22oi_1 _2872_ (.Y(_0598_),
    .B1(_0597_),
    .B2(net561),
    .A2(\wrapper.h_count[9] ),
    .A1(\wrapper.h_count[8] ));
 sg13g2_nor2b_1 _2873_ (.A(\wrapper.h_count[8] ),
    .B_N(\wrapper.h_count[9] ),
    .Y(_0599_));
 sg13g2_a21oi_1 _2874_ (.A1(_0371_),
    .A2(_0599_),
    .Y(_0600_),
    .B1(net204));
 sg13g2_o21ai_1 _2875_ (.B1(net579),
    .Y(_0120_),
    .A1(_0598_),
    .A2(_0600_));
 sg13g2_dfrbp_1 _2876_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net35),
    .D(_0028_),
    .Q_N(_0027_),
    .Q(\wrapper.h_count[0] ));
 sg13g2_dfrbp_1 _2877_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net76),
    .D(_0029_),
    .Q_N(_1430_),
    .Q(\wrapper.h_count[1] ));
 sg13g2_dfrbp_1 _2878_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net75),
    .D(_0030_),
    .Q_N(_1429_),
    .Q(\wrapper.h_count[2] ));
 sg13g2_dfrbp_1 _2879_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net74),
    .D(_0031_),
    .Q_N(_1428_),
    .Q(\wrapper.h_count[3] ));
 sg13g2_dfrbp_1 _2880_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net73),
    .D(_0032_),
    .Q_N(_0008_),
    .Q(\wrapper.h_count[4] ));
 sg13g2_dfrbp_1 _2881_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net72),
    .D(_0033_),
    .Q_N(_0014_),
    .Q(\wrapper.h_count[5] ));
 sg13g2_dfrbp_1 _2882_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net71),
    .D(_0034_),
    .Q_N(_0019_),
    .Q(\wrapper.h_count[6] ));
 sg13g2_dfrbp_1 _2883_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net70),
    .D(_0035_),
    .Q_N(_1427_),
    .Q(\wrapper.h_count[7] ));
 sg13g2_dfrbp_1 _2884_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net69),
    .D(_0036_),
    .Q_N(_1426_),
    .Q(\wrapper.h_count[8] ));
 sg13g2_dfrbp_1 _2885_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net36),
    .D(_0037_),
    .Q_N(_0007_),
    .Q(\wrapper.h_count[9] ));
 sg13g2_dfrbp_1 _2886_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net37),
    .D(_0000_),
    .Q_N(_1431_),
    .Q(\wrapper.pixel.rom0.color_out[0] ));
 sg13g2_dfrbp_1 _2887_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net38),
    .D(_0001_),
    .Q_N(_1432_),
    .Q(\wrapper.pixel.rom0.color_out[1] ));
 sg13g2_dfrbp_1 _2888_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net39),
    .D(_0002_),
    .Q_N(_1433_),
    .Q(\wrapper.pixel.rom0.color_out[2] ));
 sg13g2_dfrbp_1 _2889_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net95),
    .D(_0003_),
    .Q_N(_1434_),
    .Q(\wrapper.pixel.rom0.color_out[4] ));
 sg13g2_dfrbp_1 _2890_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net68),
    .D(_0004_),
    .Q_N(_1425_),
    .Q(\wrapper.pixel.rom0.color_out[5] ));
 sg13g2_dfrbp_1 _2891_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net67),
    .D(net135),
    .Q_N(_0026_),
    .Q(\wrapper.pixel.looping_background_count[0] ));
 sg13g2_dfrbp_1 _2892_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net65),
    .D(_0039_),
    .Q_N(_1424_),
    .Q(\wrapper.pixel.looping_background_count[1] ));
 sg13g2_dfrbp_1 _2893_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net63),
    .D(_0040_),
    .Q_N(_1423_),
    .Q(\wrapper.pixel.looping_background_count[2] ));
 sg13g2_dfrbp_1 _2894_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net61),
    .D(net157),
    .Q_N(_1422_),
    .Q(\wrapper.pixel.looping_background_count[3] ));
 sg13g2_dfrbp_1 _2895_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net59),
    .D(net185),
    .Q_N(_1421_),
    .Q(\wrapper.pixel.lfsr_reg[0] ));
 sg13g2_dfrbp_1 _2896_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net58),
    .D(_0043_),
    .Q_N(_1420_),
    .Q(\wrapper.pixel.lfsr_reg[1] ));
 sg13g2_dfrbp_1 _2897_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net57),
    .D(_0044_),
    .Q_N(_1419_),
    .Q(\wrapper.pixel.lfsr_reg[2] ));
 sg13g2_dfrbp_1 _2898_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net56),
    .D(_0045_),
    .Q_N(_1418_),
    .Q(\wrapper.pixel.lfsr_reg[3] ));
 sg13g2_dfrbp_1 _2899_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net55),
    .D(_0046_),
    .Q_N(_1417_),
    .Q(\wrapper.pixel.lfsr_reg[4] ));
 sg13g2_dfrbp_1 _2900_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net54),
    .D(_0047_),
    .Q_N(_1416_),
    .Q(\wrapper.pixel.lfsr_reg[5] ));
 sg13g2_dfrbp_1 _2901_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net53),
    .D(_0048_),
    .Q_N(_1415_),
    .Q(\wrapper.pixel.lfsr_reg[6] ));
 sg13g2_dfrbp_1 _2902_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net52),
    .D(_0049_),
    .Q_N(_1414_),
    .Q(\wrapper.pixel.lfsr_reg[7] ));
 sg13g2_dfrbp_1 _2903_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net51),
    .D(_0050_),
    .Q_N(_1413_),
    .Q(\wrapper.pixel.lfsr_reg[8] ));
 sg13g2_dfrbp_1 _2904_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net50),
    .D(_0051_),
    .Q_N(_1412_),
    .Q(\wrapper.pixel.lfsr_reg[9] ));
 sg13g2_dfrbp_1 _2905_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net49),
    .D(_0052_),
    .Q_N(_0020_),
    .Q(\wrapper.pixel.lfsr_reg[10] ));
 sg13g2_dfrbp_1 _2906_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net48),
    .D(_0053_),
    .Q_N(_1411_),
    .Q(\wrapper.pixel.lfsr_reg[11] ));
 sg13g2_dfrbp_1 _2907_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net47),
    .D(_0054_),
    .Q_N(_1410_),
    .Q(\wrapper.pixel.lfsr_reg[12] ));
 sg13g2_dfrbp_1 _2908_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net46),
    .D(_0055_),
    .Q_N(_1409_),
    .Q(\wrapper.pixel.lfsr_reg[13] ));
 sg13g2_dfrbp_1 _2909_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net45),
    .D(_0056_),
    .Q_N(_1408_),
    .Q(\wrapper.pixel.lfsr_reg[14] ));
 sg13g2_dfrbp_1 _2910_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net44),
    .D(_0057_),
    .Q_N(_1407_),
    .Q(\wrapper.pixel.lfsr_reg[15] ));
 sg13g2_dfrbp_1 _2911_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net43),
    .D(net178),
    .Q_N(_1406_),
    .Q(\wrapper.pixel.background_state[0] ));
 sg13g2_dfrbp_1 _2912_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net41),
    .D(net174),
    .Q_N(_1405_),
    .Q(\wrapper.pixel.background_state[1] ));
 sg13g2_dfrbp_1 _2913_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net34),
    .D(net187),
    .Q_N(_1404_),
    .Q(\wrapper.pixel.background_state[2] ));
 sg13g2_dfrbp_1 _2914_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net32),
    .D(_0061_),
    .Q_N(_1403_),
    .Q(\wrapper.pixel.background_state[3] ));
 sg13g2_dfrbp_1 _2915_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net30),
    .D(_0062_),
    .Q_N(_1402_),
    .Q(\wrapper.pixel.solid_color[0] ));
 sg13g2_dfrbp_1 _2916_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net28),
    .D(_0063_),
    .Q_N(_1401_),
    .Q(\wrapper.pixel.solid_color[1] ));
 sg13g2_dfrbp_1 _2917_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net26),
    .D(_0064_),
    .Q_N(_1400_),
    .Q(\wrapper.pixel.solid_color[2] ));
 sg13g2_dfrbp_1 _2918_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net122),
    .D(_0065_),
    .Q_N(_1399_),
    .Q(\wrapper.pixel.solid_color[3] ));
 sg13g2_dfrbp_1 _2919_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net120),
    .D(_0066_),
    .Q_N(_1398_),
    .Q(\wrapper.pixel.solid_color[4] ));
 sg13g2_dfrbp_1 _2920_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net118),
    .D(_0067_),
    .Q_N(_1397_),
    .Q(\wrapper.pixel.solid_color[5] ));
 sg13g2_dfrbp_1 _2921_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net116),
    .D(net165),
    .Q_N(_0025_),
    .Q(\wrapper.pixel.sprite_left[0] ));
 sg13g2_dfrbp_1 _2922_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net114),
    .D(_0069_),
    .Q_N(_1396_),
    .Q(\wrapper.pixel.sprite_left[1] ));
 sg13g2_dfrbp_1 _2923_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net112),
    .D(_0070_),
    .Q_N(_1395_),
    .Q(\wrapper.pixel.sprite_left[2] ));
 sg13g2_dfrbp_1 _2924_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net110),
    .D(_0071_),
    .Q_N(_1394_),
    .Q(\wrapper.pixel.sprite_left[3] ));
 sg13g2_dfrbp_1 _2925_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net108),
    .D(_0072_),
    .Q_N(_1393_),
    .Q(\wrapper.pixel.sprite_left[4] ));
 sg13g2_dfrbp_1 _2926_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net106),
    .D(_0073_),
    .Q_N(_1392_),
    .Q(\wrapper.pixel.sprite_left[5] ));
 sg13g2_dfrbp_1 _2927_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net104),
    .D(_0074_),
    .Q_N(_1391_),
    .Q(\wrapper.pixel.sprite_left[6] ));
 sg13g2_dfrbp_1 _2928_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net102),
    .D(_0075_),
    .Q_N(_1390_),
    .Q(\wrapper.pixel.sprite_left[7] ));
 sg13g2_dfrbp_1 _2929_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net100),
    .D(_0076_),
    .Q_N(_1389_),
    .Q(\wrapper.pixel.sprite_left[8] ));
 sg13g2_dfrbp_1 _2930_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net98),
    .D(_0077_),
    .Q_N(_1388_),
    .Q(\wrapper.pixel.sprite_left[9] ));
 sg13g2_dfrbp_1 _2931_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net96),
    .D(net167),
    .Q_N(_0024_),
    .Q(\wrapper.pixel.sprite_top[0] ));
 sg13g2_dfrbp_1 _2932_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net94),
    .D(_0079_),
    .Q_N(_1387_),
    .Q(\wrapper.pixel.sprite_top[1] ));
 sg13g2_dfrbp_1 _2933_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net92),
    .D(_0080_),
    .Q_N(_1386_),
    .Q(\wrapper.pixel.sprite_top[2] ));
 sg13g2_dfrbp_1 _2934_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net90),
    .D(_0081_),
    .Q_N(_1385_),
    .Q(\wrapper.pixel.sprite_top[3] ));
 sg13g2_dfrbp_1 _2935_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net88),
    .D(_0082_),
    .Q_N(_1384_),
    .Q(\wrapper.pixel.sprite_top[4] ));
 sg13g2_dfrbp_1 _2936_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net86),
    .D(_0083_),
    .Q_N(_1383_),
    .Q(\wrapper.pixel.sprite_top[5] ));
 sg13g2_dfrbp_1 _2937_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net84),
    .D(_0084_),
    .Q_N(_1382_),
    .Q(\wrapper.pixel.sprite_top[6] ));
 sg13g2_dfrbp_1 _2938_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net82),
    .D(_0085_),
    .Q_N(_1381_),
    .Q(\wrapper.pixel.sprite_top[7] ));
 sg13g2_dfrbp_1 _2939_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net80),
    .D(_0086_),
    .Q_N(_1380_),
    .Q(\wrapper.pixel.sprite_top[8] ));
 sg13g2_dfrbp_1 _2940_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net78),
    .D(_0087_),
    .Q_N(_1379_),
    .Q(\wrapper.pixel.sprite_top[9] ));
 sg13g2_dfrbp_1 _2941_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net66),
    .D(_0088_),
    .Q_N(_0006_),
    .Q(\wrapper.pixel.x_mov ));
 sg13g2_dfrbp_1 _2942_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net62),
    .D(net137),
    .Q_N(_0005_),
    .Q(\wrapper.pixel.y_mov ));
 sg13g2_dfrbp_1 _2943_ (.CLK(net539),
    .RESET_B(net42),
    .D(_0090_),
    .Q_N(_0023_),
    .Q(\wrapper.pixel.moving_counter[0] ));
 sg13g2_dfrbp_1 _2944_ (.CLK(net539),
    .RESET_B(net40),
    .D(_0091_),
    .Q_N(_0012_),
    .Q(\wrapper.pixel.moving_counter[1] ));
 sg13g2_dfrbp_1 _2945_ (.CLK(net539),
    .RESET_B(net33),
    .D(_0092_),
    .Q_N(_0011_),
    .Q(\wrapper.pixel.moving_counter[2] ));
 sg13g2_dfrbp_1 _2946_ (.CLK(net539),
    .RESET_B(net31),
    .D(_0093_),
    .Q_N(_0010_),
    .Q(\wrapper.pixel.moving_counter[3] ));
 sg13g2_dfrbp_1 _2947_ (.CLK(net539),
    .RESET_B(net29),
    .D(_0094_),
    .Q_N(_0009_),
    .Q(\wrapper.pixel.moving_counter[4] ));
 sg13g2_dfrbp_1 _2948_ (.CLK(\wrapper.pixel.vsync ),
    .RESET_B(net27),
    .D(_0095_),
    .Q_N(_0015_),
    .Q(\wrapper.pixel.moving_counter[5] ));
 sg13g2_dfrbp_1 _2949_ (.CLK(net539),
    .RESET_B(net25),
    .D(_0096_),
    .Q_N(_0017_),
    .Q(\wrapper.pixel.moving_counter[6] ));
 sg13g2_dfrbp_1 _2950_ (.CLK(net539),
    .RESET_B(net121),
    .D(_0097_),
    .Q_N(_0021_),
    .Q(\wrapper.pixel.moving_counter[7] ));
 sg13g2_dfrbp_1 _2951_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net119),
    .D(_0098_),
    .Q_N(_1378_),
    .Q(\wrapper.pixel.rom0.color_out[3] ));
 sg13g2_dfrbp_1 _2952_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net117),
    .D(net159),
    .Q_N(_1377_),
    .Q(\wrapper.pixel.prev_y[0] ));
 sg13g2_dfrbp_1 _2953_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net115),
    .D(_0100_),
    .Q_N(_1376_),
    .Q(\wrapper.pixel.prev_y[1] ));
 sg13g2_dfrbp_1 _2954_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net113),
    .D(net148),
    .Q_N(_1375_),
    .Q(\wrapper.pixel.prev_y[2] ));
 sg13g2_dfrbp_1 _2955_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net111),
    .D(net152),
    .Q_N(_1374_),
    .Q(\wrapper.pixel.prev_y[3] ));
 sg13g2_dfrbp_1 _2956_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net109),
    .D(_0103_),
    .Q_N(_1373_),
    .Q(\wrapper.pixel.prev_y[4] ));
 sg13g2_dfrbp_1 _2957_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net107),
    .D(net171),
    .Q_N(_1372_),
    .Q(\wrapper.pixel.prev_y[5] ));
 sg13g2_dfrbp_1 _2958_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net105),
    .D(_0105_),
    .Q_N(_1371_),
    .Q(\wrapper.pixel.prev_y[6] ));
 sg13g2_dfrbp_1 _2959_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net103),
    .D(_0106_),
    .Q_N(_1370_),
    .Q(\wrapper.pixel.prev_y[7] ));
 sg13g2_dfrbp_1 _2960_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net101),
    .D(net144),
    .Q_N(_1369_),
    .Q(\wrapper.pixel.prev_y[8] ));
 sg13g2_dfrbp_1 _2961_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net99),
    .D(net142),
    .Q_N(_1368_),
    .Q(\wrapper.pixel.prev_y[9] ));
 sg13g2_dfrbp_1 _2962_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net97),
    .D(_0109_),
    .Q_N(_1367_),
    .Q(\wrapper.pixel.vpos[0] ));
 sg13g2_dfrbp_1 _2963_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net93),
    .D(_0110_),
    .Q_N(_1366_),
    .Q(\wrapper.pixel.vpos[1] ));
 sg13g2_dfrbp_1 _2964_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net89),
    .D(_0111_),
    .Q_N(_0013_),
    .Q(\wrapper.pixel.vpos[2] ));
 sg13g2_dfrbp_1 _2965_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net85),
    .D(_0112_),
    .Q_N(_1365_),
    .Q(\wrapper.pixel.vpos[3] ));
 sg13g2_dfrbp_1 _2966_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net81),
    .D(_0113_),
    .Q_N(_1364_),
    .Q(\wrapper.pixel.vpos[4] ));
 sg13g2_dfrbp_1 _2967_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net77),
    .D(_0114_),
    .Q_N(_0016_),
    .Q(\wrapper.pixel.vpos[5] ));
 sg13g2_dfrbp_1 _2968_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net60),
    .D(net197),
    .Q_N(_0018_),
    .Q(\wrapper.pixel.vpos[6] ));
 sg13g2_dfrbp_1 _2969_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net91),
    .D(_0116_),
    .Q_N(_0022_),
    .Q(\wrapper.pixel.vpos[7] ));
 sg13g2_dfrbp_1 _2970_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net83),
    .D(_0117_),
    .Q_N(_1363_),
    .Q(\wrapper.pixel.vpos[8] ));
 sg13g2_dfrbp_1 _2971_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net64),
    .D(_0118_),
    .Q_N(_1362_),
    .Q(\wrapper.pixel.vpos[9] ));
 sg13g2_dfrbp_1 _2972_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net87),
    .D(_0119_),
    .Q_N(_1361_),
    .Q(\wrapper.pixel.vsync ));
 sg13g2_dfrbp_1 _2973_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net79),
    .D(_0120_),
    .Q_N(_1360_),
    .Q(\wrapper.hsync ));
 sg13g2_tiehi _2917__26 (.L_HI(net26));
 sg13g2_tiehi _2948__27 (.L_HI(net27));
 sg13g2_tiehi _2916__28 (.L_HI(net28));
 sg13g2_tiehi _2947__29 (.L_HI(net29));
 sg13g2_tiehi _2915__30 (.L_HI(net30));
 sg13g2_tiehi _2946__31 (.L_HI(net31));
 sg13g2_tiehi _2914__32 (.L_HI(net32));
 sg13g2_tiehi _2945__33 (.L_HI(net33));
 sg13g2_tiehi _2913__34 (.L_HI(net34));
 sg13g2_tiehi _2876__35 (.L_HI(net35));
 sg13g2_tiehi _2885__36 (.L_HI(net36));
 sg13g2_tiehi _2886__37 (.L_HI(net37));
 sg13g2_tiehi _2887__38 (.L_HI(net38));
 sg13g2_tiehi _2888__39 (.L_HI(net39));
 sg13g2_tiehi _2944__40 (.L_HI(net40));
 sg13g2_tiehi _2912__41 (.L_HI(net41));
 sg13g2_tiehi _2943__42 (.L_HI(net42));
 sg13g2_tiehi _2911__43 (.L_HI(net43));
 sg13g2_tiehi _2910__44 (.L_HI(net44));
 sg13g2_tiehi _2909__45 (.L_HI(net45));
 sg13g2_tiehi _2908__46 (.L_HI(net46));
 sg13g2_tiehi _2907__47 (.L_HI(net47));
 sg13g2_tiehi _2906__48 (.L_HI(net48));
 sg13g2_tiehi _2905__49 (.L_HI(net49));
 sg13g2_tiehi _2904__50 (.L_HI(net50));
 sg13g2_tiehi _2903__51 (.L_HI(net51));
 sg13g2_tiehi _2902__52 (.L_HI(net52));
 sg13g2_tiehi _2901__53 (.L_HI(net53));
 sg13g2_tiehi _2900__54 (.L_HI(net54));
 sg13g2_tiehi _2899__55 (.L_HI(net55));
 sg13g2_tiehi _2898__56 (.L_HI(net56));
 sg13g2_tiehi _2897__57 (.L_HI(net57));
 sg13g2_tiehi _2896__58 (.L_HI(net58));
 sg13g2_tiehi _2895__59 (.L_HI(net59));
 sg13g2_tiehi _2968__60 (.L_HI(net60));
 sg13g2_tiehi _2894__61 (.L_HI(net61));
 sg13g2_tiehi _2942__62 (.L_HI(net62));
 sg13g2_tiehi _2893__63 (.L_HI(net63));
 sg13g2_tiehi _2971__64 (.L_HI(net64));
 sg13g2_tiehi _2892__65 (.L_HI(net65));
 sg13g2_tiehi _2941__66 (.L_HI(net66));
 sg13g2_tiehi _2891__67 (.L_HI(net67));
 sg13g2_tiehi _2890__68 (.L_HI(net68));
 sg13g2_tiehi _2884__69 (.L_HI(net69));
 sg13g2_tiehi _2883__70 (.L_HI(net70));
 sg13g2_tiehi _2882__71 (.L_HI(net71));
 sg13g2_tiehi _2881__72 (.L_HI(net72));
 sg13g2_tiehi _2880__73 (.L_HI(net73));
 sg13g2_tiehi _2879__74 (.L_HI(net74));
 sg13g2_tiehi _2878__75 (.L_HI(net75));
 sg13g2_tiehi _2877__76 (.L_HI(net76));
 sg13g2_tiehi _2967__77 (.L_HI(net77));
 sg13g2_tiehi _2940__78 (.L_HI(net78));
 sg13g2_tiehi _2973__79 (.L_HI(net79));
 sg13g2_tiehi _2939__80 (.L_HI(net80));
 sg13g2_tiehi _2966__81 (.L_HI(net81));
 sg13g2_tiehi _2938__82 (.L_HI(net82));
 sg13g2_tiehi _2970__83 (.L_HI(net83));
 sg13g2_tiehi _2937__84 (.L_HI(net84));
 sg13g2_tiehi _2965__85 (.L_HI(net85));
 sg13g2_tiehi _2936__86 (.L_HI(net86));
 sg13g2_tiehi _2972__87 (.L_HI(net87));
 sg13g2_tiehi _2935__88 (.L_HI(net88));
 sg13g2_tiehi _2964__89 (.L_HI(net89));
 sg13g2_tiehi _2934__90 (.L_HI(net90));
 sg13g2_tiehi _2969__91 (.L_HI(net91));
 sg13g2_tiehi _2933__92 (.L_HI(net92));
 sg13g2_tiehi _2963__93 (.L_HI(net93));
 sg13g2_tiehi _2932__94 (.L_HI(net94));
 sg13g2_tiehi _2889__95 (.L_HI(net95));
 sg13g2_tiehi _2931__96 (.L_HI(net96));
 sg13g2_tiehi _2962__97 (.L_HI(net97));
 sg13g2_tiehi _2930__98 (.L_HI(net98));
 sg13g2_tiehi _2961__99 (.L_HI(net99));
 sg13g2_tiehi _2929__100 (.L_HI(net100));
 sg13g2_tiehi _2960__101 (.L_HI(net101));
 sg13g2_tiehi _2928__102 (.L_HI(net102));
 sg13g2_tiehi _2959__103 (.L_HI(net103));
 sg13g2_tiehi _2927__104 (.L_HI(net104));
 sg13g2_tiehi _2958__105 (.L_HI(net105));
 sg13g2_tiehi _2926__106 (.L_HI(net106));
 sg13g2_tiehi _2957__107 (.L_HI(net107));
 sg13g2_tiehi _2925__108 (.L_HI(net108));
 sg13g2_tiehi _2956__109 (.L_HI(net109));
 sg13g2_tiehi _2924__110 (.L_HI(net110));
 sg13g2_tiehi _2955__111 (.L_HI(net111));
 sg13g2_tiehi _2923__112 (.L_HI(net112));
 sg13g2_tiehi _2954__113 (.L_HI(net113));
 sg13g2_tiehi _2922__114 (.L_HI(net114));
 sg13g2_tiehi _2953__115 (.L_HI(net115));
 sg13g2_tiehi _2921__116 (.L_HI(net116));
 sg13g2_tiehi _2952__117 (.L_HI(net117));
 sg13g2_tiehi _2920__118 (.L_HI(net118));
 sg13g2_tiehi _2951__119 (.L_HI(net119));
 sg13g2_tiehi _2919__120 (.L_HI(net120));
 sg13g2_tiehi _2950__121 (.L_HI(net121));
 sg13g2_tiehi _2918__122 (.L_HI(net122));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_jmack2201_10 (.L_LO(net10));
 sg13g2_tielo tt_um_jmack2201_11 (.L_LO(net11));
 sg13g2_tielo tt_um_jmack2201_12 (.L_LO(net12));
 sg13g2_tielo tt_um_jmack2201_13 (.L_LO(net13));
 sg13g2_tielo tt_um_jmack2201_14 (.L_LO(net14));
 sg13g2_tielo tt_um_jmack2201_15 (.L_LO(net15));
 sg13g2_tielo tt_um_jmack2201_16 (.L_LO(net16));
 sg13g2_tielo tt_um_jmack2201_17 (.L_LO(net17));
 sg13g2_tielo tt_um_jmack2201_18 (.L_LO(net18));
 sg13g2_tielo tt_um_jmack2201_19 (.L_LO(net19));
 sg13g2_tielo tt_um_jmack2201_20 (.L_LO(net20));
 sg13g2_tielo tt_um_jmack2201_21 (.L_LO(net21));
 sg13g2_tielo tt_um_jmack2201_22 (.L_LO(net22));
 sg13g2_tielo tt_um_jmack2201_23 (.L_LO(net23));
 sg13g2_tielo tt_um_jmack2201_24 (.L_LO(net24));
 sg13g2_tiehi _2949__25 (.L_HI(net25));
 sg13g2_buf_4 _3088_ (.X(uo_out[3]),
    .A(net539));
 sg13g2_buf_1 _3089_ (.A(\wrapper.hsync ),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout440 (.X(net440),
    .A(_1038_));
 sg13g2_buf_2 fanout441 (.A(_1038_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(net443),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_0983_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_1011_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(net451),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(net451),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(net449),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(net451),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(net451),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_0945_),
    .X(net451));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(net456));
 sg13g2_buf_2 fanout453 (.A(net456),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(net455),
    .X(net454));
 sg13g2_buf_4 fanout455 (.X(net455),
    .A(net456));
 sg13g2_buf_2 fanout456 (.A(_0944_),
    .X(net456));
 sg13g2_buf_4 fanout457 (.X(net457),
    .A(_0935_));
 sg13g2_buf_2 fanout458 (.A(_0935_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(net461),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(net461),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(net465),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(net464),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(net464),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(net465),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_0396_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_0358_),
    .X(net466));
 sg13g2_buf_4 fanout467 (.X(net467),
    .A(_1309_));
 sg13g2_buf_4 fanout468 (.X(net468),
    .A(_1035_));
 sg13g2_buf_2 fanout469 (.A(net475),
    .X(net469));
 sg13g2_buf_1 fanout470 (.A(net475),
    .X(net470));
 sg13g2_buf_4 fanout471 (.X(net471),
    .A(net475));
 sg13g2_buf_2 fanout472 (.A(net474),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(net474),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net475),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_0938_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(net478),
    .X(net476));
 sg13g2_buf_1 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_4 fanout478 (.X(net478),
    .A(net485));
 sg13g2_buf_2 fanout479 (.A(net485),
    .X(net479));
 sg13g2_buf_1 fanout480 (.A(net485),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(net483),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(net483),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(net484),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(net485),
    .X(net484));
 sg13g2_buf_1 fanout485 (.A(_0937_),
    .X(net485));
 sg13g2_buf_4 fanout486 (.X(net486),
    .A(_1013_));
 sg13g2_buf_2 fanout487 (.A(_1013_),
    .X(net487));
 sg13g2_buf_4 fanout488 (.X(net488),
    .A(_1008_));
 sg13g2_buf_4 fanout489 (.X(net489),
    .A(_0991_));
 sg13g2_buf_4 fanout490 (.X(net490),
    .A(_0987_));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(net492));
 sg13g2_buf_2 fanout492 (.A(_0971_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(net494),
    .X(net493));
 sg13g2_buf_4 fanout494 (.X(net494),
    .A(net496));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(net496));
 sg13g2_buf_2 fanout496 (.A(net499),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(net498),
    .X(net497));
 sg13g2_buf_4 fanout498 (.X(net498),
    .A(net499));
 sg13g2_buf_2 fanout499 (.A(_0940_),
    .X(net499));
 sg13g2_buf_4 fanout500 (.X(net500),
    .A(net501));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(net502));
 sg13g2_buf_2 fanout502 (.A(net505),
    .X(net502));
 sg13g2_buf_4 fanout503 (.X(net503),
    .A(net504));
 sg13g2_buf_4 fanout504 (.X(net504),
    .A(net505));
 sg13g2_buf_2 fanout505 (.A(_0939_),
    .X(net505));
 sg13g2_buf_4 fanout506 (.X(net506),
    .A(_0999_));
 sg13g2_buf_1 fanout507 (.A(_0999_),
    .X(net507));
 sg13g2_buf_4 fanout508 (.X(net508),
    .A(net511));
 sg13g2_buf_2 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(net511),
    .X(net510));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(_0980_));
 sg13g2_buf_2 fanout512 (.A(net513),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_0979_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(net515),
    .X(net514));
 sg13g2_buf_4 fanout515 (.X(net515),
    .A(_0979_));
 sg13g2_buf_4 fanout516 (.X(net516),
    .A(net518));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(net518));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(_0951_));
 sg13g2_buf_4 fanout519 (.X(net519),
    .A(net520));
 sg13g2_buf_4 fanout520 (.X(net520),
    .A(_0950_));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(_0992_));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(_0752_));
 sg13g2_buf_1 fanout523 (.A(_0752_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_0721_),
    .X(net524));
 sg13g2_buf_1 fanout525 (.A(_0721_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(net530),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(net530),
    .X(net527));
 sg13g2_buf_4 fanout528 (.X(net528),
    .A(net529));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(net530));
 sg13g2_buf_2 fanout530 (.A(_0978_),
    .X(net530));
 sg13g2_buf_4 fanout531 (.X(net531),
    .A(net533));
 sg13g2_buf_2 fanout532 (.A(net533),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_0977_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net535),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(net537),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(net537),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_0977_),
    .X(net537));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(_0949_));
 sg13g2_buf_2 fanout539 (.A(\wrapper.pixel.vsync ),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(\wrapper.pixel.vpos[6] ),
    .X(net540));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(\wrapper.pixel.vpos[5] ));
 sg13g2_buf_2 fanout542 (.A(net543),
    .X(net542));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(\wrapper.pixel.vpos[4] ));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(net213));
 sg13g2_buf_2 fanout545 (.A(\wrapper.pixel.vpos[3] ),
    .X(net545));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(net227));
 sg13g2_buf_2 fanout547 (.A(\wrapper.pixel.vpos[2] ),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net549),
    .X(net548));
 sg13g2_buf_4 fanout549 (.X(net549),
    .A(\wrapper.pixel.vpos[1] ));
 sg13g2_buf_4 fanout550 (.X(net550),
    .A(net214));
 sg13g2_buf_2 fanout551 (.A(\wrapper.pixel.vpos[0] ),
    .X(net551));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(net554));
 sg13g2_buf_2 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(\wrapper.pixel.y_mov ),
    .X(net554));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(net557));
 sg13g2_buf_1 fanout556 (.A(net557),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(\wrapper.pixel.x_mov ),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(\wrapper.pixel.background_state[3] ),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(\wrapper.pixel.background_state[2] ),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(\wrapper.pixel.background_state[1] ),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net562),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(\wrapper.h_count[7] ),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(net211),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(\wrapper.h_count[5] ),
    .X(net564));
 sg13g2_buf_4 fanout565 (.X(net565),
    .A(net209));
 sg13g2_buf_4 fanout566 (.X(net566),
    .A(\wrapper.h_count[0] ));
 sg13g2_buf_2 fanout567 (.A(_0438_),
    .X(net567));
 sg13g2_buf_1 fanout568 (.A(_0438_),
    .X(net568));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(_0628_));
 sg13g2_buf_2 fanout570 (.A(net571),
    .X(net570));
 sg13g2_buf_4 fanout571 (.X(net571),
    .A(_0628_));
 sg13g2_buf_2 fanout572 (.A(net8),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(net7),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net576),
    .X(net574));
 sg13g2_buf_1 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_4 fanout576 (.X(net576),
    .A(net577));
 sg13g2_buf_2 fanout577 (.A(net585),
    .X(net577));
 sg13g2_buf_4 fanout578 (.X(net578),
    .A(net585));
 sg13g2_buf_4 fanout579 (.X(net579),
    .A(net584));
 sg13g2_buf_2 fanout580 (.A(net581),
    .X(net580));
 sg13g2_buf_1 fanout581 (.A(net584),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(net584),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(net584),
    .X(net583));
 sg13g2_buf_4 fanout584 (.X(net584),
    .A(net585));
 sg13g2_buf_1 fanout585 (.A(rst_n),
    .X(net585));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_jmack2201_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0027_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold2 (.A(\wrapper.pixel.lfsr_reg[3] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold3 (.A(\wrapper.pixel.lfsr_reg[4] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold4 (.A(\wrapper.pixel.lfsr_reg[0] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold5 (.A(\wrapper.pixel.lfsr_reg[9] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold6 (.A(\wrapper.pixel.lfsr_reg[8] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold7 (.A(\wrapper.pixel.lfsr_reg[2] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold8 (.A(\wrapper.pixel.lfsr_reg[6] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold9 (.A(\wrapper.pixel.lfsr_reg[1] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold10 (.A(\wrapper.pixel.lfsr_reg[5] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold11 (.A(\wrapper.pixel.lfsr_reg[7] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0026_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0038_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0005_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0089_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold16 (.A(\wrapper.pixel.vpos[1] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0568_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold18 (.A(\wrapper.pixel.lfsr_reg[10] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold19 (.A(\wrapper.pixel.prev_y[9] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0108_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold21 (.A(\wrapper.pixel.prev_y[8] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0107_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold23 (.A(\wrapper.pixel.prev_y[1] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0006_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold25 (.A(\wrapper.pixel.prev_y[2] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0101_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold27 (.A(\wrapper.pixel.lfsr_reg[11] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold28 (.A(\wrapper.pixel.prev_y[6] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold29 (.A(\wrapper.pixel.prev_y[3] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0102_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold31 (.A(\wrapper.pixel.prev_y[7] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold32 (.A(\wrapper.pixel.prev_y[4] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold33 (.A(\wrapper.pixel.sprite_top[9] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold34 (.A(\wrapper.pixel.looping_background_count[3] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0041_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold36 (.A(\wrapper.pixel.prev_y[0] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0099_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold38 (.A(\wrapper.pixel.lfsr_reg[14] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold39 (.A(\wrapper.pixel.solid_color[3] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold40 (.A(\wrapper.pixel.solid_color[1] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold41 (.A(\wrapper.pixel.lfsr_reg[12] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0025_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0068_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0024_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0078_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold46 (.A(\wrapper.pixel.solid_color[4] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold47 (.A(\wrapper.pixel.solid_color[5] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold48 (.A(\wrapper.pixel.prev_y[5] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0104_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold50 (.A(\wrapper.pixel.sprite_left[1] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold51 (.A(\wrapper.pixel.background_state[1] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0059_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold53 (.A(\wrapper.pixel.lfsr_reg[13] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold54 (.A(\wrapper.pixel.sprite_top[1] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold55 (.A(\wrapper.pixel.looping_background_count[0] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0058_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0008_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0365_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold59 (.A(\wrapper.pixel.solid_color[2] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold60 (.A(\wrapper.pixel.background_state[3] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold61 (.A(\wrapper.pixel.solid_color[0] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0020_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0042_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold64 (.A(\wrapper.pixel.looping_background_count[2] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0060_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold66 (.A(\wrapper.pixel.sprite_left[9] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold67 (.A(\wrapper.pixel.looping_background_count[1] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold68 (.A(\wrapper.h_count[9] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold69 (.A(\wrapper.pixel.sprite_top[2] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0022_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0586_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0587_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0019_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold74 (.A(\wrapper.pixel.vpos[6] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0115_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0016_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0581_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold78 (.A(\wrapper.pixel.sprite_left[5] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold79 (.A(\wrapper.pixel.sprite_left[7] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0013_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0572_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0007_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold83 (.A(\wrapper.h_count[3] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0362_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold85 (.A(\wrapper.pixel.sprite_left[6] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold86 (.A(\wrapper.h_count[8] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold87 (.A(\wrapper.h_count[2] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold88 (.A(\wrapper.pixel.sprite_top[3] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold89 (.A(\wrapper.h_count[6] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold90 (.A(\wrapper.pixel.sprite_top[6] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold91 (.A(\wrapper.pixel.vpos[3] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold92 (.A(\wrapper.pixel.vpos[0] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold93 (.A(\wrapper.pixel.sprite_left[2] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold94 (.A(\wrapper.pixel.sprite_top[7] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold95 (.A(\wrapper.pixel.sprite_top[4] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold96 (.A(\wrapper.pixel.vpos[8] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold97 (.A(\wrapper.pixel.vpos[9] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold98 (.A(\wrapper.pixel.sprite_left[4] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold99 (.A(\wrapper.h_count[1] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0360_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold101 (.A(\wrapper.pixel.sprite_left[3] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold102 (.A(\wrapper.pixel.sprite_top[5] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold103 (.A(\wrapper.pixel.sprite_top[8] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold104 (.A(\wrapper.pixel.sprite_left[8] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold105 (.A(\wrapper.pixel.vpos[2] ),
    .X(net227));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_fill_2 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_267 ();
 sg13g2_decap_8 FILLER_24_274 ();
 sg13g2_decap_8 FILLER_24_281 ();
 sg13g2_decap_8 FILLER_24_288 ();
 sg13g2_decap_8 FILLER_24_295 ();
 sg13g2_decap_8 FILLER_24_302 ();
 sg13g2_decap_8 FILLER_24_309 ();
 sg13g2_decap_8 FILLER_24_316 ();
 sg13g2_decap_8 FILLER_24_323 ();
 sg13g2_decap_8 FILLER_24_330 ();
 sg13g2_decap_8 FILLER_24_337 ();
 sg13g2_decap_8 FILLER_24_344 ();
 sg13g2_decap_8 FILLER_24_351 ();
 sg13g2_decap_8 FILLER_24_358 ();
 sg13g2_decap_8 FILLER_24_365 ();
 sg13g2_decap_8 FILLER_24_372 ();
 sg13g2_decap_8 FILLER_24_379 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_fill_2 FILLER_25_168 ();
 sg13g2_fill_1 FILLER_25_170 ();
 sg13g2_decap_8 FILLER_25_197 ();
 sg13g2_decap_8 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_211 ();
 sg13g2_decap_8 FILLER_25_218 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_232 ();
 sg13g2_fill_2 FILLER_25_259 ();
 sg13g2_fill_2 FILLER_25_265 ();
 sg13g2_decap_8 FILLER_25_293 ();
 sg13g2_decap_8 FILLER_25_300 ();
 sg13g2_decap_8 FILLER_25_307 ();
 sg13g2_decap_8 FILLER_25_314 ();
 sg13g2_decap_8 FILLER_25_321 ();
 sg13g2_decap_8 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_decap_8 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_349 ();
 sg13g2_decap_8 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_4 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_165 ();
 sg13g2_fill_1 FILLER_26_192 ();
 sg13g2_decap_8 FILLER_26_197 ();
 sg13g2_decap_4 FILLER_26_204 ();
 sg13g2_decap_8 FILLER_26_212 ();
 sg13g2_decap_8 FILLER_26_219 ();
 sg13g2_decap_4 FILLER_26_226 ();
 sg13g2_fill_2 FILLER_26_230 ();
 sg13g2_fill_1 FILLER_26_251 ();
 sg13g2_decap_8 FILLER_26_300 ();
 sg13g2_decap_8 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_314 ();
 sg13g2_decap_8 FILLER_26_321 ();
 sg13g2_decap_8 FILLER_26_328 ();
 sg13g2_decap_8 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_decap_8 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_4 FILLER_27_154 ();
 sg13g2_fill_2 FILLER_27_158 ();
 sg13g2_fill_1 FILLER_27_196 ();
 sg13g2_fill_1 FILLER_27_223 ();
 sg13g2_fill_1 FILLER_27_255 ();
 sg13g2_fill_1 FILLER_27_261 ();
 sg13g2_fill_1 FILLER_27_276 ();
 sg13g2_decap_8 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_decap_8 FILLER_27_309 ();
 sg13g2_decap_8 FILLER_27_316 ();
 sg13g2_decap_8 FILLER_27_323 ();
 sg13g2_decap_8 FILLER_27_330 ();
 sg13g2_decap_8 FILLER_27_337 ();
 sg13g2_decap_8 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_fill_2 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_fill_1 FILLER_28_186 ();
 sg13g2_fill_1 FILLER_28_204 ();
 sg13g2_fill_1 FILLER_28_235 ();
 sg13g2_decap_8 FILLER_28_307 ();
 sg13g2_decap_8 FILLER_28_314 ();
 sg13g2_decap_8 FILLER_28_321 ();
 sg13g2_decap_8 FILLER_28_328 ();
 sg13g2_decap_8 FILLER_28_335 ();
 sg13g2_decap_8 FILLER_28_342 ();
 sg13g2_decap_8 FILLER_28_349 ();
 sg13g2_decap_8 FILLER_28_356 ();
 sg13g2_decap_8 FILLER_28_363 ();
 sg13g2_decap_8 FILLER_28_370 ();
 sg13g2_decap_8 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_fill_2 FILLER_29_161 ();
 sg13g2_fill_2 FILLER_29_184 ();
 sg13g2_fill_1 FILLER_29_207 ();
 sg13g2_fill_2 FILLER_29_240 ();
 sg13g2_fill_1 FILLER_29_260 ();
 sg13g2_fill_1 FILLER_29_282 ();
 sg13g2_decap_8 FILLER_29_309 ();
 sg13g2_decap_8 FILLER_29_316 ();
 sg13g2_decap_8 FILLER_29_323 ();
 sg13g2_decap_8 FILLER_29_330 ();
 sg13g2_decap_8 FILLER_29_337 ();
 sg13g2_decap_8 FILLER_29_344 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_4 FILLER_30_168 ();
 sg13g2_fill_2 FILLER_30_209 ();
 sg13g2_fill_1 FILLER_30_211 ();
 sg13g2_fill_1 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_decap_8 FILLER_30_319 ();
 sg13g2_decap_8 FILLER_30_326 ();
 sg13g2_decap_8 FILLER_30_333 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_decap_8 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_354 ();
 sg13g2_decap_8 FILLER_30_361 ();
 sg13g2_decap_8 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_fill_2 FILLER_31_147 ();
 sg13g2_fill_1 FILLER_31_149 ();
 sg13g2_fill_1 FILLER_31_181 ();
 sg13g2_fill_1 FILLER_31_189 ();
 sg13g2_fill_1 FILLER_31_195 ();
 sg13g2_decap_8 FILLER_31_200 ();
 sg13g2_decap_8 FILLER_31_207 ();
 sg13g2_decap_4 FILLER_31_214 ();
 sg13g2_fill_2 FILLER_31_240 ();
 sg13g2_fill_1 FILLER_31_259 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_306 ();
 sg13g2_decap_8 FILLER_31_313 ();
 sg13g2_decap_8 FILLER_31_320 ();
 sg13g2_decap_8 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_334 ();
 sg13g2_decap_8 FILLER_31_341 ();
 sg13g2_decap_8 FILLER_31_348 ();
 sg13g2_decap_8 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_362 ();
 sg13g2_decap_8 FILLER_31_369 ();
 sg13g2_decap_8 FILLER_31_376 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_4 FILLER_32_147 ();
 sg13g2_fill_1 FILLER_32_151 ();
 sg13g2_decap_4 FILLER_32_186 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_fill_2 FILLER_32_213 ();
 sg13g2_fill_1 FILLER_32_215 ();
 sg13g2_fill_2 FILLER_32_266 ();
 sg13g2_fill_1 FILLER_32_289 ();
 sg13g2_decap_8 FILLER_32_316 ();
 sg13g2_decap_8 FILLER_32_323 ();
 sg13g2_decap_8 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_decap_8 FILLER_32_351 ();
 sg13g2_decap_8 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_4 FILLER_33_161 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_decap_4 FILLER_33_169 ();
 sg13g2_fill_1 FILLER_33_173 ();
 sg13g2_decap_8 FILLER_33_179 ();
 sg13g2_fill_1 FILLER_33_229 ();
 sg13g2_decap_8 FILLER_33_260 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_fill_2 FILLER_34_167 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_fill_1 FILLER_34_203 ();
 sg13g2_fill_2 FILLER_34_209 ();
 sg13g2_fill_2 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_231 ();
 sg13g2_fill_1 FILLER_34_240 ();
 sg13g2_decap_8 FILLER_34_256 ();
 sg13g2_decap_8 FILLER_34_263 ();
 sg13g2_decap_4 FILLER_34_270 ();
 sg13g2_fill_2 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_282 ();
 sg13g2_decap_8 FILLER_34_307 ();
 sg13g2_decap_8 FILLER_34_314 ();
 sg13g2_decap_8 FILLER_34_321 ();
 sg13g2_decap_8 FILLER_34_328 ();
 sg13g2_decap_8 FILLER_34_335 ();
 sg13g2_decap_8 FILLER_34_342 ();
 sg13g2_decap_8 FILLER_34_349 ();
 sg13g2_decap_8 FILLER_34_356 ();
 sg13g2_decap_8 FILLER_34_363 ();
 sg13g2_decap_8 FILLER_34_370 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_189 ();
 sg13g2_fill_1 FILLER_35_208 ();
 sg13g2_decap_8 FILLER_35_213 ();
 sg13g2_decap_4 FILLER_35_220 ();
 sg13g2_fill_1 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_270 ();
 sg13g2_fill_2 FILLER_35_277 ();
 sg13g2_fill_1 FILLER_35_286 ();
 sg13g2_fill_2 FILLER_35_291 ();
 sg13g2_decap_4 FILLER_35_306 ();
 sg13g2_fill_2 FILLER_35_310 ();
 sg13g2_decap_8 FILLER_35_316 ();
 sg13g2_decap_8 FILLER_35_323 ();
 sg13g2_decap_8 FILLER_35_330 ();
 sg13g2_decap_8 FILLER_35_337 ();
 sg13g2_decap_8 FILLER_35_344 ();
 sg13g2_decap_8 FILLER_35_351 ();
 sg13g2_decap_8 FILLER_35_358 ();
 sg13g2_decap_8 FILLER_35_365 ();
 sg13g2_decap_8 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_4 FILLER_36_154 ();
 sg13g2_fill_2 FILLER_36_158 ();
 sg13g2_fill_1 FILLER_36_170 ();
 sg13g2_decap_8 FILLER_36_201 ();
 sg13g2_decap_4 FILLER_36_208 ();
 sg13g2_fill_2 FILLER_36_237 ();
 sg13g2_fill_1 FILLER_36_239 ();
 sg13g2_fill_2 FILLER_36_275 ();
 sg13g2_fill_1 FILLER_36_290 ();
 sg13g2_decap_8 FILLER_36_325 ();
 sg13g2_decap_8 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_339 ();
 sg13g2_decap_8 FILLER_36_346 ();
 sg13g2_decap_8 FILLER_36_353 ();
 sg13g2_decap_8 FILLER_36_360 ();
 sg13g2_decap_8 FILLER_36_367 ();
 sg13g2_decap_8 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_fill_2 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_93 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_fill_2 FILLER_37_154 ();
 sg13g2_fill_1 FILLER_37_156 ();
 sg13g2_decap_4 FILLER_37_165 ();
 sg13g2_decap_4 FILLER_37_174 ();
 sg13g2_decap_4 FILLER_37_183 ();
 sg13g2_fill_1 FILLER_37_187 ();
 sg13g2_decap_8 FILLER_37_193 ();
 sg13g2_fill_1 FILLER_37_200 ();
 sg13g2_fill_2 FILLER_37_211 ();
 sg13g2_fill_1 FILLER_37_247 ();
 sg13g2_fill_2 FILLER_37_259 ();
 sg13g2_fill_1 FILLER_37_271 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_56 ();
 sg13g2_fill_1 FILLER_38_58 ();
 sg13g2_decap_4 FILLER_38_69 ();
 sg13g2_fill_2 FILLER_38_73 ();
 sg13g2_fill_2 FILLER_38_83 ();
 sg13g2_fill_1 FILLER_38_85 ();
 sg13g2_fill_2 FILLER_38_101 ();
 sg13g2_fill_2 FILLER_38_117 ();
 sg13g2_fill_1 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_fill_2 FILLER_38_161 ();
 sg13g2_fill_1 FILLER_38_163 ();
 sg13g2_fill_2 FILLER_38_197 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_fill_1 FILLER_38_291 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_352 ();
 sg13g2_decap_8 FILLER_38_359 ();
 sg13g2_decap_8 FILLER_38_366 ();
 sg13g2_decap_8 FILLER_38_373 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_fill_1 FILLER_39_49 ();
 sg13g2_fill_2 FILLER_39_73 ();
 sg13g2_fill_2 FILLER_39_122 ();
 sg13g2_fill_2 FILLER_39_146 ();
 sg13g2_fill_1 FILLER_39_148 ();
 sg13g2_fill_1 FILLER_39_165 ();
 sg13g2_fill_2 FILLER_39_174 ();
 sg13g2_fill_1 FILLER_39_186 ();
 sg13g2_fill_2 FILLER_39_213 ();
 sg13g2_decap_4 FILLER_39_233 ();
 sg13g2_fill_1 FILLER_39_237 ();
 sg13g2_fill_1 FILLER_39_309 ();
 sg13g2_fill_1 FILLER_39_318 ();
 sg13g2_fill_2 FILLER_39_324 ();
 sg13g2_fill_1 FILLER_39_326 ();
 sg13g2_decap_8 FILLER_39_344 ();
 sg13g2_decap_8 FILLER_39_351 ();
 sg13g2_decap_8 FILLER_39_358 ();
 sg13g2_decap_8 FILLER_39_365 ();
 sg13g2_decap_8 FILLER_39_372 ();
 sg13g2_decap_8 FILLER_39_379 ();
 sg13g2_decap_8 FILLER_39_386 ();
 sg13g2_decap_8 FILLER_39_393 ();
 sg13g2_decap_8 FILLER_39_400 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_fill_2 FILLER_40_49 ();
 sg13g2_fill_1 FILLER_40_51 ();
 sg13g2_fill_1 FILLER_40_58 ();
 sg13g2_fill_1 FILLER_40_69 ();
 sg13g2_fill_1 FILLER_40_88 ();
 sg13g2_fill_1 FILLER_40_104 ();
 sg13g2_fill_1 FILLER_40_118 ();
 sg13g2_fill_2 FILLER_40_131 ();
 sg13g2_fill_1 FILLER_40_133 ();
 sg13g2_fill_2 FILLER_40_164 ();
 sg13g2_fill_1 FILLER_40_166 ();
 sg13g2_fill_2 FILLER_40_178 ();
 sg13g2_fill_1 FILLER_40_180 ();
 sg13g2_fill_2 FILLER_40_200 ();
 sg13g2_fill_1 FILLER_40_202 ();
 sg13g2_decap_8 FILLER_40_218 ();
 sg13g2_decap_4 FILLER_40_225 ();
 sg13g2_fill_2 FILLER_40_229 ();
 sg13g2_decap_4 FILLER_40_235 ();
 sg13g2_fill_1 FILLER_40_248 ();
 sg13g2_fill_2 FILLER_40_270 ();
 sg13g2_fill_1 FILLER_40_272 ();
 sg13g2_decap_4 FILLER_40_286 ();
 sg13g2_decap_8 FILLER_40_295 ();
 sg13g2_fill_2 FILLER_40_302 ();
 sg13g2_fill_1 FILLER_40_312 ();
 sg13g2_decap_8 FILLER_40_317 ();
 sg13g2_decap_4 FILLER_40_324 ();
 sg13g2_decap_8 FILLER_40_332 ();
 sg13g2_decap_8 FILLER_40_339 ();
 sg13g2_decap_8 FILLER_40_346 ();
 sg13g2_decap_8 FILLER_40_353 ();
 sg13g2_decap_8 FILLER_40_360 ();
 sg13g2_decap_8 FILLER_40_367 ();
 sg13g2_decap_8 FILLER_40_374 ();
 sg13g2_decap_8 FILLER_40_381 ();
 sg13g2_decap_8 FILLER_40_388 ();
 sg13g2_decap_8 FILLER_40_395 ();
 sg13g2_decap_8 FILLER_40_402 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_4 FILLER_41_42 ();
 sg13g2_fill_2 FILLER_41_46 ();
 sg13g2_fill_1 FILLER_41_62 ();
 sg13g2_decap_4 FILLER_41_69 ();
 sg13g2_fill_2 FILLER_41_78 ();
 sg13g2_fill_1 FILLER_41_80 ();
 sg13g2_fill_2 FILLER_41_127 ();
 sg13g2_fill_1 FILLER_41_129 ();
 sg13g2_fill_2 FILLER_41_160 ();
 sg13g2_fill_1 FILLER_41_162 ();
 sg13g2_fill_1 FILLER_41_171 ();
 sg13g2_fill_2 FILLER_41_189 ();
 sg13g2_fill_1 FILLER_41_191 ();
 sg13g2_decap_8 FILLER_41_209 ();
 sg13g2_decap_4 FILLER_41_216 ();
 sg13g2_fill_1 FILLER_41_220 ();
 sg13g2_fill_1 FILLER_41_271 ();
 sg13g2_fill_2 FILLER_41_310 ();
 sg13g2_fill_1 FILLER_41_312 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_fill_2 FILLER_42_35 ();
 sg13g2_fill_2 FILLER_42_66 ();
 sg13g2_fill_2 FILLER_42_74 ();
 sg13g2_fill_1 FILLER_42_76 ();
 sg13g2_fill_1 FILLER_42_93 ();
 sg13g2_decap_4 FILLER_42_98 ();
 sg13g2_fill_2 FILLER_42_102 ();
 sg13g2_fill_1 FILLER_42_118 ();
 sg13g2_decap_4 FILLER_42_199 ();
 sg13g2_fill_2 FILLER_42_203 ();
 sg13g2_fill_2 FILLER_42_254 ();
 sg13g2_fill_1 FILLER_42_290 ();
 sg13g2_fill_1 FILLER_42_325 ();
 sg13g2_decap_8 FILLER_42_352 ();
 sg13g2_decap_8 FILLER_42_359 ();
 sg13g2_decap_8 FILLER_42_366 ();
 sg13g2_decap_8 FILLER_42_373 ();
 sg13g2_decap_8 FILLER_42_380 ();
 sg13g2_decap_8 FILLER_42_387 ();
 sg13g2_decap_8 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_fill_1 FILLER_43_88 ();
 sg13g2_fill_1 FILLER_43_104 ();
 sg13g2_fill_2 FILLER_43_119 ();
 sg13g2_fill_1 FILLER_43_121 ();
 sg13g2_fill_2 FILLER_43_126 ();
 sg13g2_fill_1 FILLER_43_128 ();
 sg13g2_decap_4 FILLER_43_137 ();
 sg13g2_fill_2 FILLER_43_141 ();
 sg13g2_decap_8 FILLER_43_151 ();
 sg13g2_fill_1 FILLER_43_193 ();
 sg13g2_fill_2 FILLER_43_202 ();
 sg13g2_fill_2 FILLER_43_240 ();
 sg13g2_fill_2 FILLER_43_269 ();
 sg13g2_fill_1 FILLER_43_271 ();
 sg13g2_fill_2 FILLER_43_286 ();
 sg13g2_fill_1 FILLER_43_296 ();
 sg13g2_fill_1 FILLER_43_321 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_4 FILLER_44_69 ();
 sg13g2_fill_1 FILLER_44_89 ();
 sg13g2_fill_2 FILLER_44_100 ();
 sg13g2_fill_1 FILLER_44_115 ();
 sg13g2_decap_4 FILLER_44_122 ();
 sg13g2_fill_1 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_132 ();
 sg13g2_decap_4 FILLER_44_139 ();
 sg13g2_decap_8 FILLER_44_155 ();
 sg13g2_decap_8 FILLER_44_162 ();
 sg13g2_fill_2 FILLER_44_173 ();
 sg13g2_fill_2 FILLER_44_178 ();
 sg13g2_decap_8 FILLER_44_194 ();
 sg13g2_decap_4 FILLER_44_201 ();
 sg13g2_decap_4 FILLER_44_208 ();
 sg13g2_decap_8 FILLER_44_225 ();
 sg13g2_fill_2 FILLER_44_257 ();
 sg13g2_fill_2 FILLER_44_296 ();
 sg13g2_fill_1 FILLER_44_298 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_decap_4 FILLER_44_315 ();
 sg13g2_fill_1 FILLER_44_319 ();
 sg13g2_decap_4 FILLER_44_324 ();
 sg13g2_fill_2 FILLER_44_337 ();
 sg13g2_decap_8 FILLER_44_354 ();
 sg13g2_decap_8 FILLER_44_361 ();
 sg13g2_decap_8 FILLER_44_368 ();
 sg13g2_decap_8 FILLER_44_375 ();
 sg13g2_decap_8 FILLER_44_382 ();
 sg13g2_decap_8 FILLER_44_389 ();
 sg13g2_decap_8 FILLER_44_396 ();
 sg13g2_decap_4 FILLER_44_403 ();
 sg13g2_fill_2 FILLER_44_407 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_fill_2 FILLER_45_56 ();
 sg13g2_fill_2 FILLER_45_71 ();
 sg13g2_fill_1 FILLER_45_73 ();
 sg13g2_fill_1 FILLER_45_81 ();
 sg13g2_fill_2 FILLER_45_114 ();
 sg13g2_fill_1 FILLER_45_127 ();
 sg13g2_decap_8 FILLER_45_137 ();
 sg13g2_fill_1 FILLER_45_144 ();
 sg13g2_decap_4 FILLER_45_156 ();
 sg13g2_fill_1 FILLER_45_160 ();
 sg13g2_fill_2 FILLER_45_169 ();
 sg13g2_fill_1 FILLER_45_171 ();
 sg13g2_fill_1 FILLER_45_192 ();
 sg13g2_decap_8 FILLER_45_219 ();
 sg13g2_decap_4 FILLER_45_226 ();
 sg13g2_fill_1 FILLER_45_230 ();
 sg13g2_fill_1 FILLER_45_307 ();
 sg13g2_fill_2 FILLER_45_316 ();
 sg13g2_fill_1 FILLER_45_332 ();
 sg13g2_decap_8 FILLER_45_351 ();
 sg13g2_decap_8 FILLER_45_358 ();
 sg13g2_decap_8 FILLER_45_365 ();
 sg13g2_decap_8 FILLER_45_372 ();
 sg13g2_decap_8 FILLER_45_379 ();
 sg13g2_decap_8 FILLER_45_386 ();
 sg13g2_decap_8 FILLER_45_393 ();
 sg13g2_decap_8 FILLER_45_400 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_fill_2 FILLER_46_42 ();
 sg13g2_fill_2 FILLER_46_52 ();
 sg13g2_fill_1 FILLER_46_54 ();
 sg13g2_fill_1 FILLER_46_73 ();
 sg13g2_decap_8 FILLER_46_78 ();
 sg13g2_decap_8 FILLER_46_85 ();
 sg13g2_decap_4 FILLER_46_92 ();
 sg13g2_fill_1 FILLER_46_96 ();
 sg13g2_fill_1 FILLER_46_106 ();
 sg13g2_fill_2 FILLER_46_119 ();
 sg13g2_fill_1 FILLER_46_121 ();
 sg13g2_fill_1 FILLER_46_130 ();
 sg13g2_fill_2 FILLER_46_150 ();
 sg13g2_fill_1 FILLER_46_157 ();
 sg13g2_decap_4 FILLER_46_171 ();
 sg13g2_fill_2 FILLER_46_183 ();
 sg13g2_fill_1 FILLER_46_205 ();
 sg13g2_decap_4 FILLER_46_219 ();
 sg13g2_fill_1 FILLER_46_223 ();
 sg13g2_decap_8 FILLER_46_229 ();
 sg13g2_fill_1 FILLER_46_236 ();
 sg13g2_fill_2 FILLER_46_331 ();
 sg13g2_decap_8 FILLER_46_359 ();
 sg13g2_decap_8 FILLER_46_366 ();
 sg13g2_decap_8 FILLER_46_373 ();
 sg13g2_decap_8 FILLER_46_380 ();
 sg13g2_decap_8 FILLER_46_387 ();
 sg13g2_decap_8 FILLER_46_394 ();
 sg13g2_decap_8 FILLER_46_401 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_fill_2 FILLER_47_49 ();
 sg13g2_fill_2 FILLER_47_63 ();
 sg13g2_fill_2 FILLER_47_70 ();
 sg13g2_fill_2 FILLER_47_80 ();
 sg13g2_decap_4 FILLER_47_91 ();
 sg13g2_fill_2 FILLER_47_95 ();
 sg13g2_fill_2 FILLER_47_101 ();
 sg13g2_fill_1 FILLER_47_103 ();
 sg13g2_fill_2 FILLER_47_109 ();
 sg13g2_fill_1 FILLER_47_111 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_162 ();
 sg13g2_fill_2 FILLER_47_177 ();
 sg13g2_fill_1 FILLER_47_179 ();
 sg13g2_fill_2 FILLER_47_188 ();
 sg13g2_fill_1 FILLER_47_201 ();
 sg13g2_fill_1 FILLER_47_304 ();
 sg13g2_fill_1 FILLER_47_338 ();
 sg13g2_decap_8 FILLER_47_348 ();
 sg13g2_decap_8 FILLER_47_355 ();
 sg13g2_decap_8 FILLER_47_362 ();
 sg13g2_decap_8 FILLER_47_369 ();
 sg13g2_decap_8 FILLER_47_376 ();
 sg13g2_decap_8 FILLER_47_383 ();
 sg13g2_decap_8 FILLER_47_390 ();
 sg13g2_decap_8 FILLER_47_397 ();
 sg13g2_decap_4 FILLER_47_404 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_fill_2 FILLER_48_42 ();
 sg13g2_fill_1 FILLER_48_44 ();
 sg13g2_fill_1 FILLER_48_60 ();
 sg13g2_fill_2 FILLER_48_74 ();
 sg13g2_fill_1 FILLER_48_76 ();
 sg13g2_fill_1 FILLER_48_95 ();
 sg13g2_fill_2 FILLER_48_108 ();
 sg13g2_fill_2 FILLER_48_124 ();
 sg13g2_fill_1 FILLER_48_126 ();
 sg13g2_fill_2 FILLER_48_136 ();
 sg13g2_decap_4 FILLER_48_144 ();
 sg13g2_fill_2 FILLER_48_148 ();
 sg13g2_fill_2 FILLER_48_163 ();
 sg13g2_decap_8 FILLER_48_181 ();
 sg13g2_decap_8 FILLER_48_188 ();
 sg13g2_fill_1 FILLER_48_195 ();
 sg13g2_fill_2 FILLER_48_209 ();
 sg13g2_fill_1 FILLER_48_211 ();
 sg13g2_decap_4 FILLER_48_257 ();
 sg13g2_fill_1 FILLER_48_261 ();
 sg13g2_fill_1 FILLER_48_311 ();
 sg13g2_decap_8 FILLER_48_316 ();
 sg13g2_decap_8 FILLER_48_327 ();
 sg13g2_decap_4 FILLER_48_334 ();
 sg13g2_fill_1 FILLER_48_338 ();
 sg13g2_decap_8 FILLER_48_344 ();
 sg13g2_decap_8 FILLER_48_351 ();
 sg13g2_decap_8 FILLER_48_358 ();
 sg13g2_decap_8 FILLER_48_365 ();
 sg13g2_decap_8 FILLER_48_372 ();
 sg13g2_decap_8 FILLER_48_379 ();
 sg13g2_decap_8 FILLER_48_386 ();
 sg13g2_decap_8 FILLER_48_393 ();
 sg13g2_decap_8 FILLER_48_400 ();
 sg13g2_fill_2 FILLER_48_407 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_4 FILLER_49_35 ();
 sg13g2_fill_2 FILLER_49_67 ();
 sg13g2_fill_1 FILLER_49_98 ();
 sg13g2_fill_2 FILLER_49_106 ();
 sg13g2_fill_1 FILLER_49_108 ();
 sg13g2_fill_2 FILLER_49_117 ();
 sg13g2_fill_1 FILLER_49_119 ();
 sg13g2_fill_1 FILLER_49_125 ();
 sg13g2_decap_4 FILLER_49_146 ();
 sg13g2_decap_4 FILLER_49_156 ();
 sg13g2_fill_2 FILLER_49_160 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_200 ();
 sg13g2_decap_8 FILLER_49_207 ();
 sg13g2_fill_1 FILLER_49_233 ();
 sg13g2_fill_2 FILLER_49_246 ();
 sg13g2_fill_1 FILLER_49_248 ();
 sg13g2_decap_4 FILLER_49_257 ();
 sg13g2_fill_1 FILLER_49_261 ();
 sg13g2_decap_8 FILLER_49_307 ();
 sg13g2_decap_8 FILLER_49_314 ();
 sg13g2_fill_2 FILLER_49_321 ();
 sg13g2_fill_2 FILLER_49_327 ();
 sg13g2_decap_8 FILLER_49_359 ();
 sg13g2_decap_8 FILLER_49_366 ();
 sg13g2_decap_8 FILLER_49_373 ();
 sg13g2_decap_8 FILLER_49_380 ();
 sg13g2_decap_8 FILLER_49_387 ();
 sg13g2_decap_8 FILLER_49_394 ();
 sg13g2_decap_8 FILLER_49_401 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_fill_2 FILLER_50_42 ();
 sg13g2_fill_2 FILLER_50_59 ();
 sg13g2_fill_1 FILLER_50_61 ();
 sg13g2_decap_4 FILLER_50_73 ();
 sg13g2_fill_2 FILLER_50_113 ();
 sg13g2_fill_2 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_165 ();
 sg13g2_decap_8 FILLER_50_172 ();
 sg13g2_decap_4 FILLER_50_179 ();
 sg13g2_fill_2 FILLER_50_183 ();
 sg13g2_decap_8 FILLER_50_266 ();
 sg13g2_fill_2 FILLER_50_273 ();
 sg13g2_decap_8 FILLER_50_284 ();
 sg13g2_fill_1 FILLER_50_291 ();
 sg13g2_fill_2 FILLER_50_302 ();
 sg13g2_fill_1 FILLER_50_304 ();
 sg13g2_fill_1 FILLER_50_327 ();
 sg13g2_decap_8 FILLER_50_359 ();
 sg13g2_decap_8 FILLER_50_366 ();
 sg13g2_decap_8 FILLER_50_373 ();
 sg13g2_decap_8 FILLER_50_380 ();
 sg13g2_decap_8 FILLER_50_387 ();
 sg13g2_decap_8 FILLER_50_394 ();
 sg13g2_decap_8 FILLER_50_401 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_4 FILLER_51_42 ();
 sg13g2_fill_1 FILLER_51_46 ();
 sg13g2_fill_2 FILLER_51_53 ();
 sg13g2_fill_1 FILLER_51_55 ();
 sg13g2_fill_1 FILLER_51_75 ();
 sg13g2_decap_4 FILLER_51_82 ();
 sg13g2_fill_1 FILLER_51_86 ();
 sg13g2_decap_4 FILLER_51_119 ();
 sg13g2_fill_2 FILLER_51_123 ();
 sg13g2_fill_2 FILLER_51_144 ();
 sg13g2_fill_2 FILLER_51_151 ();
 sg13g2_decap_4 FILLER_51_167 ();
 sg13g2_fill_1 FILLER_51_184 ();
 sg13g2_fill_2 FILLER_51_190 ();
 sg13g2_fill_1 FILLER_51_224 ();
 sg13g2_fill_2 FILLER_51_255 ();
 sg13g2_fill_1 FILLER_51_275 ();
 sg13g2_decap_8 FILLER_51_290 ();
 sg13g2_fill_1 FILLER_51_297 ();
 sg13g2_fill_1 FILLER_51_316 ();
 sg13g2_decap_8 FILLER_51_361 ();
 sg13g2_decap_8 FILLER_51_368 ();
 sg13g2_decap_8 FILLER_51_375 ();
 sg13g2_decap_8 FILLER_51_382 ();
 sg13g2_decap_8 FILLER_51_389 ();
 sg13g2_decap_8 FILLER_51_396 ();
 sg13g2_decap_4 FILLER_51_403 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_4 FILLER_52_35 ();
 sg13g2_fill_2 FILLER_52_56 ();
 sg13g2_fill_1 FILLER_52_58 ();
 sg13g2_fill_1 FILLER_52_67 ();
 sg13g2_fill_1 FILLER_52_74 ();
 sg13g2_decap_8 FILLER_52_80 ();
 sg13g2_fill_2 FILLER_52_87 ();
 sg13g2_fill_1 FILLER_52_89 ();
 sg13g2_decap_8 FILLER_52_94 ();
 sg13g2_decap_4 FILLER_52_101 ();
 sg13g2_decap_8 FILLER_52_127 ();
 sg13g2_fill_1 FILLER_52_143 ();
 sg13g2_decap_4 FILLER_52_148 ();
 sg13g2_fill_2 FILLER_52_152 ();
 sg13g2_fill_2 FILLER_52_158 ();
 sg13g2_fill_1 FILLER_52_160 ();
 sg13g2_fill_2 FILLER_52_191 ();
 sg13g2_fill_1 FILLER_52_236 ();
 sg13g2_fill_2 FILLER_52_245 ();
 sg13g2_fill_1 FILLER_52_247 ();
 sg13g2_fill_2 FILLER_52_296 ();
 sg13g2_fill_1 FILLER_52_333 ();
 sg13g2_decap_8 FILLER_52_353 ();
 sg13g2_decap_8 FILLER_52_360 ();
 sg13g2_decap_8 FILLER_52_367 ();
 sg13g2_decap_8 FILLER_52_374 ();
 sg13g2_decap_8 FILLER_52_381 ();
 sg13g2_decap_8 FILLER_52_388 ();
 sg13g2_decap_8 FILLER_52_395 ();
 sg13g2_decap_8 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_fill_2 FILLER_53_35 ();
 sg13g2_fill_1 FILLER_53_37 ();
 sg13g2_decap_4 FILLER_53_95 ();
 sg13g2_fill_1 FILLER_53_99 ();
 sg13g2_fill_2 FILLER_53_111 ();
 sg13g2_fill_2 FILLER_53_137 ();
 sg13g2_fill_1 FILLER_53_139 ();
 sg13g2_fill_2 FILLER_53_145 ();
 sg13g2_fill_2 FILLER_53_152 ();
 sg13g2_fill_2 FILLER_53_185 ();
 sg13g2_fill_1 FILLER_53_187 ();
 sg13g2_fill_2 FILLER_53_206 ();
 sg13g2_fill_1 FILLER_53_208 ();
 sg13g2_fill_1 FILLER_53_220 ();
 sg13g2_fill_2 FILLER_53_255 ();
 sg13g2_fill_1 FILLER_53_257 ();
 sg13g2_fill_1 FILLER_53_278 ();
 sg13g2_decap_8 FILLER_53_289 ();
 sg13g2_decap_8 FILLER_53_296 ();
 sg13g2_fill_2 FILLER_53_303 ();
 sg13g2_fill_1 FILLER_53_305 ();
 sg13g2_decap_4 FILLER_53_318 ();
 sg13g2_fill_2 FILLER_53_322 ();
 sg13g2_decap_8 FILLER_53_332 ();
 sg13g2_decap_8 FILLER_53_339 ();
 sg13g2_decap_8 FILLER_53_346 ();
 sg13g2_decap_8 FILLER_53_353 ();
 sg13g2_decap_8 FILLER_53_360 ();
 sg13g2_decap_8 FILLER_53_367 ();
 sg13g2_decap_8 FILLER_53_374 ();
 sg13g2_decap_8 FILLER_53_381 ();
 sg13g2_decap_8 FILLER_53_388 ();
 sg13g2_decap_8 FILLER_53_395 ();
 sg13g2_decap_8 FILLER_53_402 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_4 FILLER_54_35 ();
 sg13g2_fill_1 FILLER_54_39 ();
 sg13g2_fill_2 FILLER_54_63 ();
 sg13g2_fill_1 FILLER_54_65 ();
 sg13g2_fill_2 FILLER_54_90 ();
 sg13g2_fill_1 FILLER_54_92 ();
 sg13g2_fill_1 FILLER_54_121 ();
 sg13g2_fill_2 FILLER_54_145 ();
 sg13g2_fill_2 FILLER_54_155 ();
 sg13g2_fill_2 FILLER_54_183 ();
 sg13g2_decap_8 FILLER_54_201 ();
 sg13g2_fill_1 FILLER_54_208 ();
 sg13g2_fill_2 FILLER_54_212 ();
 sg13g2_fill_1 FILLER_54_219 ();
 sg13g2_fill_2 FILLER_54_229 ();
 sg13g2_fill_1 FILLER_54_231 ();
 sg13g2_fill_2 FILLER_54_236 ();
 sg13g2_fill_2 FILLER_54_252 ();
 sg13g2_decap_8 FILLER_54_286 ();
 sg13g2_decap_8 FILLER_54_293 ();
 sg13g2_fill_1 FILLER_54_300 ();
 sg13g2_fill_2 FILLER_54_308 ();
 sg13g2_decap_8 FILLER_54_322 ();
 sg13g2_decap_8 FILLER_54_329 ();
 sg13g2_decap_4 FILLER_54_336 ();
 sg13g2_fill_2 FILLER_54_340 ();
 sg13g2_decap_8 FILLER_54_350 ();
 sg13g2_decap_8 FILLER_54_357 ();
 sg13g2_decap_8 FILLER_54_364 ();
 sg13g2_decap_8 FILLER_54_371 ();
 sg13g2_decap_8 FILLER_54_378 ();
 sg13g2_decap_8 FILLER_54_385 ();
 sg13g2_decap_8 FILLER_54_392 ();
 sg13g2_decap_8 FILLER_54_399 ();
 sg13g2_fill_2 FILLER_54_406 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_fill_2 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_60 ();
 sg13g2_decap_8 FILLER_55_67 ();
 sg13g2_decap_4 FILLER_55_74 ();
 sg13g2_fill_2 FILLER_55_78 ();
 sg13g2_fill_1 FILLER_55_90 ();
 sg13g2_fill_2 FILLER_55_104 ();
 sg13g2_decap_4 FILLER_55_121 ();
 sg13g2_fill_2 FILLER_55_135 ();
 sg13g2_fill_2 FILLER_55_142 ();
 sg13g2_fill_1 FILLER_55_144 ();
 sg13g2_fill_2 FILLER_55_150 ();
 sg13g2_fill_1 FILLER_55_152 ();
 sg13g2_decap_8 FILLER_55_165 ();
 sg13g2_decap_4 FILLER_55_172 ();
 sg13g2_decap_8 FILLER_55_181 ();
 sg13g2_fill_2 FILLER_55_188 ();
 sg13g2_fill_1 FILLER_55_190 ();
 sg13g2_decap_4 FILLER_55_211 ();
 sg13g2_decap_8 FILLER_55_231 ();
 sg13g2_fill_1 FILLER_55_250 ();
 sg13g2_decap_4 FILLER_55_294 ();
 sg13g2_decap_4 FILLER_55_303 ();
 sg13g2_fill_2 FILLER_55_307 ();
 sg13g2_decap_4 FILLER_55_313 ();
 sg13g2_fill_1 FILLER_55_317 ();
 sg13g2_fill_2 FILLER_55_327 ();
 sg13g2_decap_8 FILLER_55_356 ();
 sg13g2_decap_8 FILLER_55_363 ();
 sg13g2_decap_8 FILLER_55_370 ();
 sg13g2_decap_8 FILLER_55_377 ();
 sg13g2_decap_8 FILLER_55_384 ();
 sg13g2_decap_8 FILLER_55_391 ();
 sg13g2_decap_8 FILLER_55_398 ();
 sg13g2_decap_4 FILLER_55_405 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_4 FILLER_56_35 ();
 sg13g2_fill_2 FILLER_56_39 ();
 sg13g2_fill_2 FILLER_56_61 ();
 sg13g2_fill_2 FILLER_56_73 ();
 sg13g2_fill_1 FILLER_56_81 ();
 sg13g2_decap_8 FILLER_56_111 ();
 sg13g2_decap_4 FILLER_56_123 ();
 sg13g2_fill_2 FILLER_56_146 ();
 sg13g2_fill_1 FILLER_56_148 ();
 sg13g2_fill_2 FILLER_56_159 ();
 sg13g2_fill_1 FILLER_56_161 ();
 sg13g2_fill_1 FILLER_56_168 ();
 sg13g2_decap_8 FILLER_56_177 ();
 sg13g2_decap_4 FILLER_56_194 ();
 sg13g2_fill_1 FILLER_56_198 ();
 sg13g2_fill_1 FILLER_56_204 ();
 sg13g2_decap_4 FILLER_56_213 ();
 sg13g2_decap_8 FILLER_56_222 ();
 sg13g2_decap_4 FILLER_56_229 ();
 sg13g2_fill_2 FILLER_56_233 ();
 sg13g2_fill_2 FILLER_56_261 ();
 sg13g2_fill_2 FILLER_56_272 ();
 sg13g2_fill_1 FILLER_56_279 ();
 sg13g2_fill_2 FILLER_56_329 ();
 sg13g2_fill_1 FILLER_56_331 ();
 sg13g2_decap_8 FILLER_56_363 ();
 sg13g2_decap_8 FILLER_56_370 ();
 sg13g2_decap_8 FILLER_56_377 ();
 sg13g2_decap_8 FILLER_56_384 ();
 sg13g2_decap_8 FILLER_56_391 ();
 sg13g2_decap_8 FILLER_56_398 ();
 sg13g2_decap_4 FILLER_56_405 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_4 FILLER_57_78 ();
 sg13g2_fill_2 FILLER_57_82 ();
 sg13g2_decap_4 FILLER_57_88 ();
 sg13g2_decap_8 FILLER_57_97 ();
 sg13g2_fill_1 FILLER_57_139 ();
 sg13g2_fill_2 FILLER_57_150 ();
 sg13g2_fill_1 FILLER_57_152 ();
 sg13g2_fill_1 FILLER_57_183 ();
 sg13g2_fill_2 FILLER_57_213 ();
 sg13g2_fill_1 FILLER_57_260 ();
 sg13g2_fill_1 FILLER_57_325 ();
 sg13g2_decap_8 FILLER_57_360 ();
 sg13g2_decap_8 FILLER_57_367 ();
 sg13g2_decap_8 FILLER_57_374 ();
 sg13g2_decap_8 FILLER_57_381 ();
 sg13g2_decap_8 FILLER_57_388 ();
 sg13g2_decap_8 FILLER_57_395 ();
 sg13g2_decap_8 FILLER_57_402 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_4 FILLER_58_35 ();
 sg13g2_fill_2 FILLER_58_39 ();
 sg13g2_fill_2 FILLER_58_61 ();
 sg13g2_fill_2 FILLER_58_73 ();
 sg13g2_fill_1 FILLER_58_75 ();
 sg13g2_fill_1 FILLER_58_84 ();
 sg13g2_fill_2 FILLER_58_109 ();
 sg13g2_fill_1 FILLER_58_125 ();
 sg13g2_fill_2 FILLER_58_137 ();
 sg13g2_decap_4 FILLER_58_156 ();
 sg13g2_fill_1 FILLER_58_160 ();
 sg13g2_decap_8 FILLER_58_173 ();
 sg13g2_decap_8 FILLER_58_190 ();
 sg13g2_fill_2 FILLER_58_197 ();
 sg13g2_fill_1 FILLER_58_214 ();
 sg13g2_fill_1 FILLER_58_220 ();
 sg13g2_decap_8 FILLER_58_250 ();
 sg13g2_fill_1 FILLER_58_257 ();
 sg13g2_fill_2 FILLER_58_336 ();
 sg13g2_decap_8 FILLER_58_348 ();
 sg13g2_decap_8 FILLER_58_355 ();
 sg13g2_decap_8 FILLER_58_362 ();
 sg13g2_decap_8 FILLER_58_369 ();
 sg13g2_decap_8 FILLER_58_376 ();
 sg13g2_decap_8 FILLER_58_383 ();
 sg13g2_decap_8 FILLER_58_390 ();
 sg13g2_decap_8 FILLER_58_397 ();
 sg13g2_decap_4 FILLER_58_404 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_fill_1 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_55 ();
 sg13g2_fill_2 FILLER_59_62 ();
 sg13g2_fill_1 FILLER_59_73 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_fill_2 FILLER_59_91 ();
 sg13g2_fill_1 FILLER_59_108 ();
 sg13g2_fill_2 FILLER_59_117 ();
 sg13g2_decap_4 FILLER_59_143 ();
 sg13g2_decap_8 FILLER_59_161 ();
 sg13g2_decap_4 FILLER_59_168 ();
 sg13g2_fill_2 FILLER_59_172 ();
 sg13g2_decap_8 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_196 ();
 sg13g2_decap_4 FILLER_59_203 ();
 sg13g2_fill_1 FILLER_59_207 ();
 sg13g2_decap_8 FILLER_59_242 ();
 sg13g2_decap_8 FILLER_59_249 ();
 sg13g2_decap_8 FILLER_59_256 ();
 sg13g2_decap_4 FILLER_59_263 ();
 sg13g2_fill_1 FILLER_59_267 ();
 sg13g2_decap_8 FILLER_59_289 ();
 sg13g2_decap_8 FILLER_59_310 ();
 sg13g2_decap_8 FILLER_59_329 ();
 sg13g2_decap_8 FILLER_59_336 ();
 sg13g2_decap_8 FILLER_59_343 ();
 sg13g2_decap_8 FILLER_59_350 ();
 sg13g2_decap_8 FILLER_59_357 ();
 sg13g2_decap_8 FILLER_59_364 ();
 sg13g2_decap_8 FILLER_59_371 ();
 sg13g2_decap_8 FILLER_59_378 ();
 sg13g2_decap_8 FILLER_59_385 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_decap_8 FILLER_59_399 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_4 FILLER_60_42 ();
 sg13g2_fill_1 FILLER_60_46 ();
 sg13g2_fill_2 FILLER_60_52 ();
 sg13g2_decap_8 FILLER_60_64 ();
 sg13g2_decap_4 FILLER_60_76 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_4 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_115 ();
 sg13g2_decap_8 FILLER_60_122 ();
 sg13g2_decap_8 FILLER_60_129 ();
 sg13g2_decap_4 FILLER_60_141 ();
 sg13g2_fill_1 FILLER_60_158 ();
 sg13g2_fill_2 FILLER_60_169 ();
 sg13g2_fill_2 FILLER_60_197 ();
 sg13g2_fill_1 FILLER_60_199 ();
 sg13g2_decap_8 FILLER_60_205 ();
 sg13g2_fill_1 FILLER_60_212 ();
 sg13g2_fill_1 FILLER_60_229 ();
 sg13g2_fill_2 FILLER_60_235 ();
 sg13g2_fill_1 FILLER_60_237 ();
 sg13g2_decap_8 FILLER_60_260 ();
 sg13g2_fill_1 FILLER_60_272 ();
 sg13g2_decap_8 FILLER_60_277 ();
 sg13g2_decap_8 FILLER_60_284 ();
 sg13g2_decap_8 FILLER_60_291 ();
 sg13g2_decap_8 FILLER_60_298 ();
 sg13g2_fill_2 FILLER_60_305 ();
 sg13g2_decap_8 FILLER_60_322 ();
 sg13g2_decap_8 FILLER_60_329 ();
 sg13g2_decap_8 FILLER_60_336 ();
 sg13g2_decap_8 FILLER_60_343 ();
 sg13g2_decap_8 FILLER_60_350 ();
 sg13g2_decap_8 FILLER_60_357 ();
 sg13g2_decap_8 FILLER_60_364 ();
 sg13g2_decap_8 FILLER_60_371 ();
 sg13g2_decap_8 FILLER_60_378 ();
 sg13g2_decap_8 FILLER_60_385 ();
 sg13g2_decap_8 FILLER_60_392 ();
 sg13g2_decap_8 FILLER_60_399 ();
 sg13g2_fill_2 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_4 FILLER_61_35 ();
 sg13g2_fill_2 FILLER_61_51 ();
 sg13g2_fill_1 FILLER_61_53 ();
 sg13g2_fill_1 FILLER_61_85 ();
 sg13g2_fill_2 FILLER_61_91 ();
 sg13g2_fill_1 FILLER_61_93 ();
 sg13g2_fill_1 FILLER_61_98 ();
 sg13g2_decap_4 FILLER_61_104 ();
 sg13g2_fill_1 FILLER_61_108 ();
 sg13g2_fill_2 FILLER_61_140 ();
 sg13g2_fill_1 FILLER_61_142 ();
 sg13g2_decap_4 FILLER_61_169 ();
 sg13g2_fill_2 FILLER_61_173 ();
 sg13g2_decap_8 FILLER_61_213 ();
 sg13g2_decap_8 FILLER_61_220 ();
 sg13g2_decap_8 FILLER_61_227 ();
 sg13g2_fill_2 FILLER_61_234 ();
 sg13g2_decap_4 FILLER_61_257 ();
 sg13g2_fill_2 FILLER_61_291 ();
 sg13g2_fill_1 FILLER_61_293 ();
 sg13g2_decap_8 FILLER_61_356 ();
 sg13g2_decap_8 FILLER_61_363 ();
 sg13g2_decap_8 FILLER_61_370 ();
 sg13g2_decap_8 FILLER_61_377 ();
 sg13g2_decap_8 FILLER_61_384 ();
 sg13g2_decap_8 FILLER_61_391 ();
 sg13g2_decap_8 FILLER_61_398 ();
 sg13g2_decap_4 FILLER_61_405 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_4 FILLER_62_28 ();
 sg13g2_fill_1 FILLER_62_32 ();
 sg13g2_fill_2 FILLER_62_62 ();
 sg13g2_fill_1 FILLER_62_64 ();
 sg13g2_fill_2 FILLER_62_87 ();
 sg13g2_decap_4 FILLER_62_109 ();
 sg13g2_fill_2 FILLER_62_124 ();
 sg13g2_fill_2 FILLER_62_146 ();
 sg13g2_fill_1 FILLER_62_148 ();
 sg13g2_decap_8 FILLER_62_155 ();
 sg13g2_decap_8 FILLER_62_162 ();
 sg13g2_decap_8 FILLER_62_169 ();
 sg13g2_decap_8 FILLER_62_176 ();
 sg13g2_fill_2 FILLER_62_183 ();
 sg13g2_fill_1 FILLER_62_185 ();
 sg13g2_decap_4 FILLER_62_209 ();
 sg13g2_fill_2 FILLER_62_213 ();
 sg13g2_decap_8 FILLER_62_223 ();
 sg13g2_decap_8 FILLER_62_230 ();
 sg13g2_decap_4 FILLER_62_237 ();
 sg13g2_fill_2 FILLER_62_262 ();
 sg13g2_fill_1 FILLER_62_264 ();
 sg13g2_fill_1 FILLER_62_294 ();
 sg13g2_decap_8 FILLER_62_352 ();
 sg13g2_decap_8 FILLER_62_359 ();
 sg13g2_decap_8 FILLER_62_366 ();
 sg13g2_decap_8 FILLER_62_373 ();
 sg13g2_decap_8 FILLER_62_380 ();
 sg13g2_decap_8 FILLER_62_387 ();
 sg13g2_decap_8 FILLER_62_394 ();
 sg13g2_decap_8 FILLER_62_401 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_fill_1 FILLER_63_57 ();
 sg13g2_fill_2 FILLER_63_133 ();
 sg13g2_fill_2 FILLER_63_143 ();
 sg13g2_fill_2 FILLER_63_157 ();
 sg13g2_decap_8 FILLER_63_203 ();
 sg13g2_decap_8 FILLER_63_210 ();
 sg13g2_decap_8 FILLER_63_217 ();
 sg13g2_fill_1 FILLER_63_231 ();
 sg13g2_fill_2 FILLER_63_262 ();
 sg13g2_fill_1 FILLER_63_316 ();
 sg13g2_fill_1 FILLER_63_328 ();
 sg13g2_decap_8 FILLER_63_356 ();
 sg13g2_decap_8 FILLER_63_363 ();
 sg13g2_decap_8 FILLER_63_370 ();
 sg13g2_decap_8 FILLER_63_377 ();
 sg13g2_decap_8 FILLER_63_384 ();
 sg13g2_decap_8 FILLER_63_391 ();
 sg13g2_decap_8 FILLER_63_398 ();
 sg13g2_decap_4 FILLER_63_405 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_4 FILLER_64_42 ();
 sg13g2_decap_4 FILLER_64_66 ();
 sg13g2_decap_4 FILLER_64_75 ();
 sg13g2_fill_1 FILLER_64_79 ();
 sg13g2_decap_4 FILLER_64_110 ();
 sg13g2_decap_4 FILLER_64_127 ();
 sg13g2_fill_1 FILLER_64_131 ();
 sg13g2_fill_1 FILLER_64_136 ();
 sg13g2_fill_2 FILLER_64_151 ();
 sg13g2_decap_8 FILLER_64_173 ();
 sg13g2_fill_1 FILLER_64_188 ();
 sg13g2_fill_2 FILLER_64_211 ();
 sg13g2_fill_1 FILLER_64_213 ();
 sg13g2_fill_2 FILLER_64_240 ();
 sg13g2_fill_2 FILLER_64_266 ();
 sg13g2_fill_1 FILLER_64_268 ();
 sg13g2_fill_1 FILLER_64_274 ();
 sg13g2_fill_1 FILLER_64_319 ();
 sg13g2_fill_1 FILLER_64_324 ();
 sg13g2_fill_2 FILLER_64_334 ();
 sg13g2_fill_1 FILLER_64_336 ();
 sg13g2_decap_8 FILLER_64_351 ();
 sg13g2_decap_8 FILLER_64_358 ();
 sg13g2_decap_8 FILLER_64_365 ();
 sg13g2_decap_8 FILLER_64_372 ();
 sg13g2_decap_8 FILLER_64_379 ();
 sg13g2_decap_8 FILLER_64_386 ();
 sg13g2_decap_8 FILLER_64_393 ();
 sg13g2_decap_8 FILLER_64_400 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_fill_2 FILLER_65_42 ();
 sg13g2_decap_4 FILLER_65_64 ();
 sg13g2_fill_1 FILLER_65_76 ();
 sg13g2_decap_8 FILLER_65_81 ();
 sg13g2_fill_1 FILLER_65_88 ();
 sg13g2_decap_4 FILLER_65_94 ();
 sg13g2_fill_2 FILLER_65_102 ();
 sg13g2_fill_1 FILLER_65_109 ();
 sg13g2_fill_2 FILLER_65_118 ();
 sg13g2_decap_4 FILLER_65_138 ();
 sg13g2_fill_2 FILLER_65_169 ();
 sg13g2_fill_2 FILLER_65_197 ();
 sg13g2_fill_2 FILLER_65_216 ();
 sg13g2_decap_4 FILLER_65_230 ();
 sg13g2_fill_2 FILLER_65_237 ();
 sg13g2_decap_8 FILLER_65_260 ();
 sg13g2_decap_4 FILLER_65_271 ();
 sg13g2_decap_8 FILLER_65_278 ();
 sg13g2_decap_8 FILLER_65_285 ();
 sg13g2_fill_1 FILLER_65_292 ();
 sg13g2_fill_2 FILLER_65_299 ();
 sg13g2_fill_1 FILLER_65_301 ();
 sg13g2_decap_4 FILLER_65_313 ();
 sg13g2_decap_8 FILLER_65_357 ();
 sg13g2_decap_8 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_371 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_decap_8 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_399 ();
 sg13g2_fill_2 FILLER_65_406 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_fill_1 FILLER_66_42 ();
 sg13g2_fill_1 FILLER_66_71 ();
 sg13g2_fill_2 FILLER_66_86 ();
 sg13g2_fill_1 FILLER_66_88 ();
 sg13g2_decap_4 FILLER_66_106 ();
 sg13g2_fill_1 FILLER_66_110 ();
 sg13g2_fill_2 FILLER_66_120 ();
 sg13g2_fill_2 FILLER_66_131 ();
 sg13g2_decap_4 FILLER_66_142 ();
 sg13g2_fill_1 FILLER_66_146 ();
 sg13g2_fill_2 FILLER_66_156 ();
 sg13g2_decap_8 FILLER_66_163 ();
 sg13g2_decap_8 FILLER_66_170 ();
 sg13g2_decap_8 FILLER_66_177 ();
 sg13g2_fill_2 FILLER_66_196 ();
 sg13g2_fill_2 FILLER_66_242 ();
 sg13g2_fill_1 FILLER_66_244 ();
 sg13g2_decap_8 FILLER_66_264 ();
 sg13g2_fill_1 FILLER_66_271 ();
 sg13g2_decap_8 FILLER_66_288 ();
 sg13g2_decap_8 FILLER_66_295 ();
 sg13g2_fill_2 FILLER_66_302 ();
 sg13g2_decap_8 FILLER_66_374 ();
 sg13g2_decap_8 FILLER_66_381 ();
 sg13g2_decap_8 FILLER_66_388 ();
 sg13g2_decap_8 FILLER_66_395 ();
 sg13g2_decap_8 FILLER_66_402 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_4 FILLER_67_42 ();
 sg13g2_fill_1 FILLER_67_56 ();
 sg13g2_fill_2 FILLER_67_62 ();
 sg13g2_fill_1 FILLER_67_64 ();
 sg13g2_fill_2 FILLER_67_81 ();
 sg13g2_fill_1 FILLER_67_83 ();
 sg13g2_fill_2 FILLER_67_103 ();
 sg13g2_fill_2 FILLER_67_114 ();
 sg13g2_fill_1 FILLER_67_116 ();
 sg13g2_fill_1 FILLER_67_134 ();
 sg13g2_fill_1 FILLER_67_143 ();
 sg13g2_fill_2 FILLER_67_157 ();
 sg13g2_fill_1 FILLER_67_159 ();
 sg13g2_fill_2 FILLER_67_171 ();
 sg13g2_fill_1 FILLER_67_173 ();
 sg13g2_fill_2 FILLER_67_232 ();
 sg13g2_fill_1 FILLER_67_296 ();
 sg13g2_decap_8 FILLER_67_311 ();
 sg13g2_decap_4 FILLER_67_318 ();
 sg13g2_fill_1 FILLER_67_322 ();
 sg13g2_decap_8 FILLER_67_361 ();
 sg13g2_decap_8 FILLER_67_368 ();
 sg13g2_decap_8 FILLER_67_375 ();
 sg13g2_decap_8 FILLER_67_382 ();
 sg13g2_decap_8 FILLER_67_389 ();
 sg13g2_decap_8 FILLER_67_396 ();
 sg13g2_decap_4 FILLER_67_403 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_4 FILLER_68_49 ();
 sg13g2_fill_1 FILLER_68_53 ();
 sg13g2_decap_4 FILLER_68_58 ();
 sg13g2_fill_1 FILLER_68_62 ();
 sg13g2_fill_2 FILLER_68_73 ();
 sg13g2_fill_1 FILLER_68_85 ();
 sg13g2_decap_4 FILLER_68_92 ();
 sg13g2_fill_2 FILLER_68_96 ();
 sg13g2_fill_2 FILLER_68_108 ();
 sg13g2_fill_2 FILLER_68_121 ();
 sg13g2_fill_2 FILLER_68_141 ();
 sg13g2_fill_1 FILLER_68_143 ();
 sg13g2_decap_4 FILLER_68_169 ();
 sg13g2_fill_1 FILLER_68_249 ();
 sg13g2_fill_1 FILLER_68_341 ();
 sg13g2_fill_2 FILLER_68_351 ();
 sg13g2_fill_1 FILLER_68_353 ();
 sg13g2_decap_8 FILLER_68_363 ();
 sg13g2_decap_8 FILLER_68_370 ();
 sg13g2_decap_8 FILLER_68_377 ();
 sg13g2_decap_8 FILLER_68_384 ();
 sg13g2_decap_8 FILLER_68_391 ();
 sg13g2_decap_8 FILLER_68_398 ();
 sg13g2_decap_4 FILLER_68_405 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_fill_2 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_64 ();
 sg13g2_fill_2 FILLER_69_71 ();
 sg13g2_decap_8 FILLER_69_78 ();
 sg13g2_decap_4 FILLER_69_85 ();
 sg13g2_fill_2 FILLER_69_89 ();
 sg13g2_fill_2 FILLER_69_145 ();
 sg13g2_fill_1 FILLER_69_147 ();
 sg13g2_fill_1 FILLER_69_153 ();
 sg13g2_fill_1 FILLER_69_165 ();
 sg13g2_fill_1 FILLER_69_200 ();
 sg13g2_fill_1 FILLER_69_211 ();
 sg13g2_fill_2 FILLER_69_225 ();
 sg13g2_fill_1 FILLER_69_227 ();
 sg13g2_fill_2 FILLER_69_237 ();
 sg13g2_fill_2 FILLER_69_269 ();
 sg13g2_fill_2 FILLER_69_276 ();
 sg13g2_fill_1 FILLER_69_278 ();
 sg13g2_fill_2 FILLER_69_301 ();
 sg13g2_fill_1 FILLER_69_334 ();
 sg13g2_decap_8 FILLER_69_361 ();
 sg13g2_decap_8 FILLER_69_368 ();
 sg13g2_decap_8 FILLER_69_375 ();
 sg13g2_decap_8 FILLER_69_382 ();
 sg13g2_decap_8 FILLER_69_389 ();
 sg13g2_decap_8 FILLER_69_396 ();
 sg13g2_decap_4 FILLER_69_403 ();
 sg13g2_fill_2 FILLER_69_407 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_fill_1 FILLER_70_42 ();
 sg13g2_fill_2 FILLER_70_67 ();
 sg13g2_fill_1 FILLER_70_89 ();
 sg13g2_decap_8 FILLER_70_94 ();
 sg13g2_fill_1 FILLER_70_101 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_fill_2 FILLER_70_140 ();
 sg13g2_fill_2 FILLER_70_153 ();
 sg13g2_decap_8 FILLER_70_170 ();
 sg13g2_fill_2 FILLER_70_181 ();
 sg13g2_fill_1 FILLER_70_183 ();
 sg13g2_fill_1 FILLER_70_188 ();
 sg13g2_decap_4 FILLER_70_194 ();
 sg13g2_fill_2 FILLER_70_198 ();
 sg13g2_decap_4 FILLER_70_209 ();
 sg13g2_decap_4 FILLER_70_221 ();
 sg13g2_decap_8 FILLER_70_239 ();
 sg13g2_fill_1 FILLER_70_246 ();
 sg13g2_fill_2 FILLER_70_273 ();
 sg13g2_fill_1 FILLER_70_275 ();
 sg13g2_decap_4 FILLER_70_280 ();
 sg13g2_fill_1 FILLER_70_284 ();
 sg13g2_fill_2 FILLER_70_353 ();
 sg13g2_decap_8 FILLER_70_368 ();
 sg13g2_decap_8 FILLER_70_375 ();
 sg13g2_decap_8 FILLER_70_382 ();
 sg13g2_decap_8 FILLER_70_389 ();
 sg13g2_decap_8 FILLER_70_396 ();
 sg13g2_decap_4 FILLER_70_403 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_fill_1 FILLER_71_49 ();
 sg13g2_fill_2 FILLER_71_60 ();
 sg13g2_fill_1 FILLER_71_62 ();
 sg13g2_fill_1 FILLER_71_97 ();
 sg13g2_decap_8 FILLER_71_103 ();
 sg13g2_decap_8 FILLER_71_110 ();
 sg13g2_decap_4 FILLER_71_117 ();
 sg13g2_fill_1 FILLER_71_121 ();
 sg13g2_decap_8 FILLER_71_137 ();
 sg13g2_decap_8 FILLER_71_144 ();
 sg13g2_fill_1 FILLER_71_151 ();
 sg13g2_decap_8 FILLER_71_162 ();
 sg13g2_decap_8 FILLER_71_169 ();
 sg13g2_decap_8 FILLER_71_176 ();
 sg13g2_decap_8 FILLER_71_183 ();
 sg13g2_decap_8 FILLER_71_190 ();
 sg13g2_decap_8 FILLER_71_197 ();
 sg13g2_decap_8 FILLER_71_216 ();
 sg13g2_decap_4 FILLER_71_223 ();
 sg13g2_fill_1 FILLER_71_227 ();
 sg13g2_decap_8 FILLER_71_240 ();
 sg13g2_decap_8 FILLER_71_247 ();
 sg13g2_decap_8 FILLER_71_262 ();
 sg13g2_fill_2 FILLER_71_269 ();
 sg13g2_fill_1 FILLER_71_271 ();
 sg13g2_fill_2 FILLER_71_322 ();
 sg13g2_fill_1 FILLER_71_324 ();
 sg13g2_decap_8 FILLER_71_373 ();
 sg13g2_decap_8 FILLER_71_380 ();
 sg13g2_decap_8 FILLER_71_387 ();
 sg13g2_decap_8 FILLER_71_394 ();
 sg13g2_decap_8 FILLER_71_401 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_fill_2 FILLER_72_49 ();
 sg13g2_fill_1 FILLER_72_51 ();
 sg13g2_fill_1 FILLER_72_70 ();
 sg13g2_decap_4 FILLER_72_109 ();
 sg13g2_fill_2 FILLER_72_113 ();
 sg13g2_decap_8 FILLER_72_120 ();
 sg13g2_fill_1 FILLER_72_127 ();
 sg13g2_decap_8 FILLER_72_138 ();
 sg13g2_decap_4 FILLER_72_145 ();
 sg13g2_fill_2 FILLER_72_149 ();
 sg13g2_fill_1 FILLER_72_163 ();
 sg13g2_fill_1 FILLER_72_205 ();
 sg13g2_fill_2 FILLER_72_219 ();
 sg13g2_decap_4 FILLER_72_244 ();
 sg13g2_decap_4 FILLER_72_265 ();
 sg13g2_fill_1 FILLER_72_278 ();
 sg13g2_fill_2 FILLER_72_288 ();
 sg13g2_fill_1 FILLER_72_290 ();
 sg13g2_decap_8 FILLER_72_366 ();
 sg13g2_decap_8 FILLER_72_373 ();
 sg13g2_decap_8 FILLER_72_380 ();
 sg13g2_decap_8 FILLER_72_387 ();
 sg13g2_decap_8 FILLER_72_394 ();
 sg13g2_decap_8 FILLER_72_401 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_fill_1 FILLER_73_56 ();
 sg13g2_fill_1 FILLER_73_61 ();
 sg13g2_fill_2 FILLER_73_67 ();
 sg13g2_decap_8 FILLER_73_111 ();
 sg13g2_fill_2 FILLER_73_118 ();
 sg13g2_fill_2 FILLER_73_141 ();
 sg13g2_fill_1 FILLER_73_143 ();
 sg13g2_fill_2 FILLER_73_149 ();
 sg13g2_fill_1 FILLER_73_151 ();
 sg13g2_fill_2 FILLER_73_170 ();
 sg13g2_fill_1 FILLER_73_172 ();
 sg13g2_fill_2 FILLER_73_197 ();
 sg13g2_fill_2 FILLER_73_205 ();
 sg13g2_fill_2 FILLER_73_324 ();
 sg13g2_decap_8 FILLER_73_370 ();
 sg13g2_decap_8 FILLER_73_377 ();
 sg13g2_decap_8 FILLER_73_384 ();
 sg13g2_decap_8 FILLER_73_391 ();
 sg13g2_decap_8 FILLER_73_398 ();
 sg13g2_decap_4 FILLER_73_405 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_fill_1 FILLER_74_60 ();
 sg13g2_fill_2 FILLER_74_77 ();
 sg13g2_fill_1 FILLER_74_98 ();
 sg13g2_fill_2 FILLER_74_109 ();
 sg13g2_fill_1 FILLER_74_111 ();
 sg13g2_fill_2 FILLER_74_117 ();
 sg13g2_fill_1 FILLER_74_119 ();
 sg13g2_fill_1 FILLER_74_186 ();
 sg13g2_fill_1 FILLER_74_221 ();
 sg13g2_fill_1 FILLER_74_237 ();
 sg13g2_fill_2 FILLER_74_247 ();
 sg13g2_fill_1 FILLER_74_249 ();
 sg13g2_fill_2 FILLER_74_276 ();
 sg13g2_fill_1 FILLER_74_283 ();
 sg13g2_decap_8 FILLER_74_362 ();
 sg13g2_decap_8 FILLER_74_369 ();
 sg13g2_decap_8 FILLER_74_376 ();
 sg13g2_decap_8 FILLER_74_383 ();
 sg13g2_decap_8 FILLER_74_390 ();
 sg13g2_decap_8 FILLER_74_397 ();
 sg13g2_decap_4 FILLER_74_404 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_fill_1 FILLER_75_49 ();
 sg13g2_decap_4 FILLER_75_78 ();
 sg13g2_fill_2 FILLER_75_82 ();
 sg13g2_fill_1 FILLER_75_93 ();
 sg13g2_fill_2 FILLER_75_99 ();
 sg13g2_fill_1 FILLER_75_101 ();
 sg13g2_decap_4 FILLER_75_165 ();
 sg13g2_fill_2 FILLER_75_169 ();
 sg13g2_fill_1 FILLER_75_216 ();
 sg13g2_decap_4 FILLER_75_252 ();
 sg13g2_fill_1 FILLER_75_268 ();
 sg13g2_fill_2 FILLER_75_297 ();
 sg13g2_fill_1 FILLER_75_299 ();
 sg13g2_fill_2 FILLER_75_327 ();
 sg13g2_fill_1 FILLER_75_329 ();
 sg13g2_decap_8 FILLER_75_343 ();
 sg13g2_decap_8 FILLER_75_350 ();
 sg13g2_decap_8 FILLER_75_357 ();
 sg13g2_decap_8 FILLER_75_364 ();
 sg13g2_decap_8 FILLER_75_371 ();
 sg13g2_decap_8 FILLER_75_378 ();
 sg13g2_decap_8 FILLER_75_385 ();
 sg13g2_decap_8 FILLER_75_392 ();
 sg13g2_decap_8 FILLER_75_399 ();
 sg13g2_fill_2 FILLER_75_406 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_fill_2 FILLER_76_42 ();
 sg13g2_fill_2 FILLER_76_88 ();
 sg13g2_fill_1 FILLER_76_90 ();
 sg13g2_decap_8 FILLER_76_100 ();
 sg13g2_fill_1 FILLER_76_107 ();
 sg13g2_fill_2 FILLER_76_128 ();
 sg13g2_fill_1 FILLER_76_130 ();
 sg13g2_decap_8 FILLER_76_145 ();
 sg13g2_decap_8 FILLER_76_152 ();
 sg13g2_fill_1 FILLER_76_159 ();
 sg13g2_fill_2 FILLER_76_207 ();
 sg13g2_fill_2 FILLER_76_231 ();
 sg13g2_decap_4 FILLER_76_247 ();
 sg13g2_fill_2 FILLER_76_251 ();
 sg13g2_fill_2 FILLER_76_256 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_392 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_fill_2 FILLER_76_406 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_4 FILLER_77_49 ();
 sg13g2_fill_2 FILLER_77_79 ();
 sg13g2_fill_1 FILLER_77_81 ();
 sg13g2_fill_2 FILLER_77_88 ();
 sg13g2_fill_1 FILLER_77_90 ();
 sg13g2_fill_2 FILLER_77_101 ();
 sg13g2_fill_1 FILLER_77_103 ();
 sg13g2_fill_1 FILLER_77_139 ();
 sg13g2_decap_8 FILLER_77_145 ();
 sg13g2_decap_8 FILLER_77_152 ();
 sg13g2_decap_8 FILLER_77_159 ();
 sg13g2_decap_4 FILLER_77_166 ();
 sg13g2_fill_1 FILLER_77_170 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_4 FILLER_77_182 ();
 sg13g2_fill_1 FILLER_77_186 ();
 sg13g2_fill_2 FILLER_77_229 ();
 sg13g2_fill_1 FILLER_77_231 ();
 sg13g2_decap_4 FILLER_77_236 ();
 sg13g2_fill_1 FILLER_77_240 ();
 sg13g2_fill_2 FILLER_77_254 ();
 sg13g2_fill_1 FILLER_77_266 ();
 sg13g2_fill_2 FILLER_77_271 ();
 sg13g2_fill_1 FILLER_77_309 ();
 sg13g2_decap_8 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_364 ();
 sg13g2_decap_8 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_fill_2 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_fill_2 FILLER_78_63 ();
 sg13g2_fill_1 FILLER_78_65 ();
 sg13g2_fill_1 FILLER_78_98 ();
 sg13g2_fill_2 FILLER_78_115 ();
 sg13g2_decap_8 FILLER_78_127 ();
 sg13g2_decap_8 FILLER_78_134 ();
 sg13g2_decap_8 FILLER_78_141 ();
 sg13g2_decap_8 FILLER_78_148 ();
 sg13g2_decap_8 FILLER_78_155 ();
 sg13g2_decap_8 FILLER_78_162 ();
 sg13g2_decap_8 FILLER_78_169 ();
 sg13g2_decap_8 FILLER_78_176 ();
 sg13g2_decap_4 FILLER_78_183 ();
 sg13g2_fill_2 FILLER_78_187 ();
 sg13g2_fill_2 FILLER_78_203 ();
 sg13g2_decap_4 FILLER_78_231 ();
 sg13g2_fill_2 FILLER_78_261 ();
 sg13g2_fill_1 FILLER_78_280 ();
 sg13g2_fill_2 FILLER_78_286 ();
 sg13g2_fill_1 FILLER_78_298 ();
 sg13g2_fill_2 FILLER_78_317 ();
 sg13g2_fill_1 FILLER_78_319 ();
 sg13g2_decap_8 FILLER_78_333 ();
 sg13g2_decap_8 FILLER_78_340 ();
 sg13g2_decap_8 FILLER_78_347 ();
 sg13g2_decap_8 FILLER_78_354 ();
 sg13g2_decap_8 FILLER_78_361 ();
 sg13g2_decap_8 FILLER_78_368 ();
 sg13g2_decap_8 FILLER_78_375 ();
 sg13g2_decap_8 FILLER_78_382 ();
 sg13g2_decap_8 FILLER_78_389 ();
 sg13g2_decap_8 FILLER_78_396 ();
 sg13g2_decap_4 FILLER_78_403 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_4 FILLER_79_75 ();
 sg13g2_fill_2 FILLER_79_79 ();
 sg13g2_fill_2 FILLER_79_90 ();
 sg13g2_fill_2 FILLER_79_96 ();
 sg13g2_decap_4 FILLER_79_107 ();
 sg13g2_fill_1 FILLER_79_111 ();
 sg13g2_decap_8 FILLER_79_117 ();
 sg13g2_decap_8 FILLER_79_124 ();
 sg13g2_decap_8 FILLER_79_131 ();
 sg13g2_decap_8 FILLER_79_138 ();
 sg13g2_decap_8 FILLER_79_145 ();
 sg13g2_decap_8 FILLER_79_152 ();
 sg13g2_decap_8 FILLER_79_159 ();
 sg13g2_decap_8 FILLER_79_166 ();
 sg13g2_decap_8 FILLER_79_173 ();
 sg13g2_decap_4 FILLER_79_180 ();
 sg13g2_fill_1 FILLER_79_184 ();
 sg13g2_fill_2 FILLER_79_211 ();
 sg13g2_fill_1 FILLER_79_213 ();
 sg13g2_fill_2 FILLER_79_218 ();
 sg13g2_fill_1 FILLER_79_220 ();
 sg13g2_decap_8 FILLER_79_329 ();
 sg13g2_decap_8 FILLER_79_336 ();
 sg13g2_decap_8 FILLER_79_343 ();
 sg13g2_decap_8 FILLER_79_350 ();
 sg13g2_decap_8 FILLER_79_357 ();
 sg13g2_decap_8 FILLER_79_364 ();
 sg13g2_decap_8 FILLER_79_371 ();
 sg13g2_decap_8 FILLER_79_378 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_fill_2 FILLER_79_406 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_fill_1 FILLER_80_84 ();
 sg13g2_fill_2 FILLER_80_93 ();
 sg13g2_fill_1 FILLER_80_103 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_fill_2 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_200 ();
 sg13g2_decap_8 FILLER_80_207 ();
 sg13g2_fill_2 FILLER_80_214 ();
 sg13g2_decap_8 FILLER_80_220 ();
 sg13g2_decap_4 FILLER_80_227 ();
 sg13g2_fill_1 FILLER_80_231 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_fill_1 FILLER_80_243 ();
 sg13g2_decap_4 FILLER_80_248 ();
 sg13g2_fill_1 FILLER_80_256 ();
 sg13g2_fill_1 FILLER_80_304 ();
 sg13g2_fill_1 FILLER_80_319 ();
 sg13g2_decap_4 FILLER_80_324 ();
 sg13g2_decap_4 FILLER_80_332 ();
 sg13g2_decap_4 FILLER_80_340 ();
 sg13g2_decap_4 FILLER_80_348 ();
 sg13g2_decap_4 FILLER_80_356 ();
 sg13g2_decap_4 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_372 ();
 sg13g2_decap_8 FILLER_80_379 ();
 sg13g2_decap_8 FILLER_80_386 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_8 FILLER_80_400 ();
 sg13g2_fill_2 FILLER_80_407 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule

module tt_um_DaDDS (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire net13;
 wire \top_level.adder.b[0] ;
 wire \top_level.adder.b[10] ;
 wire \top_level.adder.b[11] ;
 wire \top_level.adder.b[12] ;
 wire \top_level.adder.b[13] ;
 wire \top_level.adder.b[14] ;
 wire \top_level.adder.b[15] ;
 wire \top_level.adder.b[1] ;
 wire \top_level.adder.b[2] ;
 wire \top_level.adder.b[3] ;
 wire \top_level.adder.b[4] ;
 wire \top_level.adder.b[5] ;
 wire \top_level.adder.b[6] ;
 wire \top_level.adder.b[7] ;
 wire \top_level.adder.b[8] ;
 wire \top_level.adder.b[9] ;
 wire \top_level.adder.sum[0] ;
 wire \top_level.adder.sum[10] ;
 wire \top_level.adder.sum[11] ;
 wire \top_level.adder.sum[12] ;
 wire \top_level.adder.sum[13] ;
 wire \top_level.adder.sum[14] ;
 wire \top_level.adder.sum[15] ;
 wire \top_level.adder.sum[1] ;
 wire \top_level.adder.sum[2] ;
 wire \top_level.adder.sum[3] ;
 wire \top_level.adder.sum[4] ;
 wire \top_level.adder.sum[5] ;
 wire \top_level.adder.sum[6] ;
 wire \top_level.adder.sum[7] ;
 wire \top_level.adder.sum[8] ;
 wire \top_level.adder.sum[9] ;
 wire \top_level.freq0_reg_out[0] ;
 wire \top_level.freq0_reg_out[10] ;
 wire \top_level.freq0_reg_out[11] ;
 wire \top_level.freq0_reg_out[12] ;
 wire \top_level.freq0_reg_out[13] ;
 wire \top_level.freq0_reg_out[14] ;
 wire \top_level.freq0_reg_out[15] ;
 wire \top_level.freq0_reg_out[1] ;
 wire \top_level.freq0_reg_out[2] ;
 wire \top_level.freq0_reg_out[3] ;
 wire \top_level.freq0_reg_out[4] ;
 wire \top_level.freq0_reg_out[5] ;
 wire \top_level.freq0_reg_out[6] ;
 wire \top_level.freq0_reg_out[7] ;
 wire \top_level.freq0_reg_out[8] ;
 wire \top_level.freq0_reg_out[9] ;
 wire \top_level.freq1_reg_out[0] ;
 wire \top_level.freq1_reg_out[10] ;
 wire \top_level.freq1_reg_out[11] ;
 wire \top_level.freq1_reg_out[12] ;
 wire \top_level.freq1_reg_out[13] ;
 wire \top_level.freq1_reg_out[14] ;
 wire \top_level.freq1_reg_out[15] ;
 wire \top_level.freq1_reg_out[1] ;
 wire \top_level.freq1_reg_out[2] ;
 wire \top_level.freq1_reg_out[3] ;
 wire \top_level.freq1_reg_out[4] ;
 wire \top_level.freq1_reg_out[5] ;
 wire \top_level.freq1_reg_out[6] ;
 wire \top_level.freq1_reg_out[7] ;
 wire \top_level.freq1_reg_out[8] ;
 wire \top_level.freq1_reg_out[9] ;
 wire \top_level.uart.bit_index_reg[0] ;
 wire \top_level.uart.bit_index_reg[1] ;
 wire \top_level.uart.bit_index_reg[2] ;
 wire \top_level.uart.bit_index_reg[3] ;
 wire \top_level.uart.byte_number ;
 wire \top_level.uart.clk_count_reg[0] ;
 wire \top_level.uart.clk_count_reg[10] ;
 wire \top_level.uart.clk_count_reg[11] ;
 wire \top_level.uart.clk_count_reg[1] ;
 wire \top_level.uart.clk_count_reg[2] ;
 wire \top_level.uart.clk_count_reg[3] ;
 wire \top_level.uart.clk_count_reg[4] ;
 wire \top_level.uart.clk_count_reg[5] ;
 wire \top_level.uart.clk_count_reg[6] ;
 wire \top_level.uart.clk_count_reg[7] ;
 wire \top_level.uart.clk_count_reg[8] ;
 wire \top_level.uart.clk_count_reg[9] ;
 wire \top_level.uart.rx_data_reg ;
 wire \top_level.uart.state_reg[0] ;
 wire \top_level.uart.state_reg[1] ;
 wire \top_level.uart.state_reg[2] ;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;

 sg13g2_inv_1 _0569_ (.Y(_0065_),
    .A(\top_level.uart.clk_count_reg[9] ));
 sg13g2_inv_1 _0570_ (.Y(_0066_),
    .A(net74));
 sg13g2_inv_2 _0571_ (.Y(_0067_),
    .A(net156));
 sg13g2_inv_1 _0572_ (.Y(_0068_),
    .A(net105));
 sg13g2_inv_1 _0573_ (.Y(_0069_),
    .A(net160));
 sg13g2_nand2b_1 _0574_ (.Y(_0070_),
    .B(_0011_),
    .A_N(net161));
 sg13g2_nand2_1 _0575_ (.Y(_0071_),
    .A(net157),
    .B(_0011_));
 sg13g2_or2_1 _0576_ (.X(_0072_),
    .B(\top_level.adder.b[12] ),
    .A(net157));
 sg13g2_nand3_1 _0577_ (.B(_0071_),
    .C(_0072_),
    .A(net162),
    .Y(_0073_));
 sg13g2_nand2_2 _0578_ (.Y(_0074_),
    .A(_0070_),
    .B(_0073_));
 sg13g2_nand2b_2 _0579_ (.Y(_0075_),
    .B(_0012_),
    .A_N(net162));
 sg13g2_nand2_1 _0580_ (.Y(_0076_),
    .A(net157),
    .B(_0012_));
 sg13g2_or2_1 _0581_ (.X(_0077_),
    .B(\top_level.adder.b[13] ),
    .A(net157));
 sg13g2_nand3_1 _0582_ (.B(_0076_),
    .C(_0077_),
    .A(net162),
    .Y(_0078_));
 sg13g2_and2_1 _0583_ (.A(_0075_),
    .B(_0078_),
    .X(_0079_));
 sg13g2_nand2_2 _0584_ (.Y(_0080_),
    .A(_0075_),
    .B(_0078_));
 sg13g2_nor2_1 _0585_ (.A(_0074_),
    .B(_0080_),
    .Y(_0081_));
 sg13g2_nand4_1 _0586_ (.B(_0073_),
    .C(_0075_),
    .A(_0070_),
    .Y(_0082_),
    .D(_0078_));
 sg13g2_nor2b_1 _0587_ (.A(net161),
    .B_N(_0008_),
    .Y(_0083_));
 sg13g2_nand2_1 _0588_ (.Y(_0084_),
    .A(net159),
    .B(_0008_));
 sg13g2_or2_1 _0589_ (.X(_0085_),
    .B(\top_level.adder.b[9] ),
    .A(net159));
 sg13g2_nand3_1 _0590_ (.B(_0084_),
    .C(_0085_),
    .A(net161),
    .Y(_0086_));
 sg13g2_nor2b_1 _0591_ (.A(_0083_),
    .B_N(_0086_),
    .Y(_0087_));
 sg13g2_nand2b_1 _0592_ (.Y(_0088_),
    .B(_0086_),
    .A_N(_0083_));
 sg13g2_nand2b_1 _0593_ (.Y(_0089_),
    .B(_0010_),
    .A_N(net161));
 sg13g2_nand2_1 _0594_ (.Y(_0090_),
    .A(net157),
    .B(_0010_));
 sg13g2_or2_1 _0595_ (.X(_0091_),
    .B(\top_level.adder.b[11] ),
    .A(net158));
 sg13g2_nand3_1 _0596_ (.B(_0090_),
    .C(_0091_),
    .A(net162),
    .Y(_0092_));
 sg13g2_nand2b_1 _0597_ (.Y(_0093_),
    .B(\top_level.adder.b[10] ),
    .A_N(net161));
 sg13g2_nand2_1 _0598_ (.Y(_0094_),
    .A(net157),
    .B(\top_level.adder.b[10] ));
 sg13g2_or2_1 _0599_ (.X(_0095_),
    .B(_0009_),
    .A(net157));
 sg13g2_nand3_1 _0600_ (.B(_0094_),
    .C(_0095_),
    .A(net161),
    .Y(_0096_));
 sg13g2_a22oi_1 _0601_ (.Y(_0097_),
    .B1(_0093_),
    .B2(_0096_),
    .A2(_0092_),
    .A1(_0089_));
 sg13g2_inv_1 _0602_ (.Y(_0098_),
    .A(net143));
 sg13g2_nand2_2 _0603_ (.Y(_0099_),
    .A(net144),
    .B(net143));
 sg13g2_nand2b_1 _0604_ (.Y(_0100_),
    .B(_0009_),
    .A_N(net161));
 sg13g2_nand2_1 _0605_ (.Y(_0101_),
    .A(net157),
    .B(_0009_));
 sg13g2_or2_1 _0606_ (.X(_0102_),
    .B(\top_level.adder.b[10] ),
    .A(net158));
 sg13g2_nand3_1 _0607_ (.B(_0101_),
    .C(_0102_),
    .A(net161),
    .Y(_0103_));
 sg13g2_a22oi_1 _0608_ (.Y(_0104_),
    .B1(_0100_),
    .B2(_0103_),
    .A2(_0092_),
    .A1(_0089_));
 sg13g2_nor2b_1 _0609_ (.A(net162),
    .B_N(_0006_),
    .Y(_0105_));
 sg13g2_nand2_1 _0610_ (.Y(_0106_),
    .A(net158),
    .B(_0006_));
 sg13g2_or2_1 _0611_ (.X(_0107_),
    .B(\top_level.adder.b[8] ),
    .A(net158));
 sg13g2_nand3_1 _0612_ (.B(_0106_),
    .C(_0107_),
    .A(\top_level.adder.b[14] ),
    .Y(_0108_));
 sg13g2_nor2b_2 _0613_ (.A(_0105_),
    .B_N(_0108_),
    .Y(_0109_));
 sg13g2_nand2b_2 _0614_ (.Y(_0110_),
    .B(_0108_),
    .A_N(_0105_));
 sg13g2_nor2_1 _0615_ (.A(net145),
    .B(_0110_),
    .Y(_0111_));
 sg13g2_nand2_1 _0616_ (.Y(_0112_),
    .A(_0088_),
    .B(_0109_));
 sg13g2_a22oi_1 _0617_ (.Y(_0113_),
    .B1(_0104_),
    .B2(_0111_),
    .A2(net143),
    .A1(net144));
 sg13g2_nand4_1 _0618_ (.B(_0092_),
    .C(_0100_),
    .A(_0089_),
    .Y(_0114_),
    .D(_0103_));
 sg13g2_nand2_2 _0619_ (.Y(_0115_),
    .A(net144),
    .B(_0110_));
 sg13g2_nand4_1 _0620_ (.B(_0092_),
    .C(_0093_),
    .A(_0089_),
    .Y(_0116_),
    .D(_0096_));
 sg13g2_or2_1 _0621_ (.X(_0117_),
    .B(_0116_),
    .A(net144));
 sg13g2_o21ai_1 _0622_ (.B1(_0117_),
    .Y(_0118_),
    .A1(net142),
    .A2(_0115_));
 sg13g2_nand2b_1 _0623_ (.Y(_0119_),
    .B(_0080_),
    .A_N(_0074_));
 sg13g2_or2_1 _0624_ (.X(_0120_),
    .B(net141),
    .A(_0116_));
 sg13g2_or2_1 _0625_ (.X(_0121_),
    .B(net141),
    .A(_0117_));
 sg13g2_and2_2 _0626_ (.A(_0074_),
    .B(_0079_),
    .X(_0122_));
 sg13g2_nand2_2 _0627_ (.Y(_0123_),
    .A(_0074_),
    .B(_0079_));
 sg13g2_nand2b_1 _0628_ (.Y(_0124_),
    .B(_0122_),
    .A_N(_0099_));
 sg13g2_nand2_1 _0629_ (.Y(_0125_),
    .A(_0104_),
    .B(_0122_));
 sg13g2_nand2_1 _0630_ (.Y(_0126_),
    .A(net146),
    .B(_0104_));
 sg13g2_nand3_1 _0631_ (.B(_0104_),
    .C(_0110_),
    .A(net146),
    .Y(_0127_));
 sg13g2_inv_1 _0632_ (.Y(_0128_),
    .A(_0127_));
 sg13g2_nand2_1 _0633_ (.Y(_0129_),
    .A(net145),
    .B(net143));
 sg13g2_nand2_2 _0634_ (.Y(_0130_),
    .A(net145),
    .B(_0109_));
 sg13g2_nand3_1 _0635_ (.B(net143),
    .C(_0109_),
    .A(net145),
    .Y(_0131_));
 sg13g2_nand2_1 _0636_ (.Y(_0132_),
    .A(net145),
    .B(_0110_));
 sg13g2_nor2b_1 _0637_ (.A(_0082_),
    .B_N(_0104_),
    .Y(_0133_));
 sg13g2_a21oi_1 _0638_ (.A1(_0127_),
    .A2(_0131_),
    .Y(_0134_),
    .B1(_0082_));
 sg13g2_a22oi_1 _0639_ (.Y(_0135_),
    .B1(_0075_),
    .B2(_0078_),
    .A2(_0073_),
    .A1(_0070_));
 sg13g2_nand2_2 _0640_ (.Y(_0136_),
    .A(_0074_),
    .B(_0080_));
 sg13g2_or2_1 _0641_ (.X(_0137_),
    .B(_0130_),
    .A(net142));
 sg13g2_a21oi_1 _0642_ (.A1(_0098_),
    .A2(net142),
    .Y(_0138_),
    .B1(_0130_));
 sg13g2_a22oi_1 _0643_ (.Y(_0139_),
    .B1(_0135_),
    .B2(_0138_),
    .A2(_0128_),
    .A1(_0080_));
 sg13g2_nand2b_1 _0644_ (.Y(_0140_),
    .B(_0138_),
    .A_N(net141));
 sg13g2_nand2b_1 _0645_ (.Y(_0141_),
    .B(_0135_),
    .A_N(_0116_));
 sg13g2_o21ai_1 _0646_ (.B1(_0140_),
    .Y(_0142_),
    .A1(_0112_),
    .A2(_0141_));
 sg13g2_inv_1 _0647_ (.Y(_0143_),
    .A(_0142_));
 sg13g2_or2_1 _0648_ (.X(_0144_),
    .B(_0141_),
    .A(_0130_));
 sg13g2_nor3_1 _0649_ (.A(net142),
    .B(_0115_),
    .C(_0123_),
    .Y(_0145_));
 sg13g2_nor2_1 _0650_ (.A(_0123_),
    .B(_0129_),
    .Y(_0146_));
 sg13g2_or2_1 _0651_ (.X(_0147_),
    .B(_0114_),
    .A(_0112_));
 sg13g2_o21ai_1 _0652_ (.B1(_0137_),
    .Y(_0148_),
    .A1(_0115_),
    .A2(_0116_));
 sg13g2_nand3_1 _0653_ (.B(net144),
    .C(_0097_),
    .A(_0080_),
    .Y(_0149_));
 sg13g2_a21oi_1 _0654_ (.A1(_0099_),
    .A2(_0147_),
    .Y(_0150_),
    .B1(_0136_));
 sg13g2_nand2b_1 _0655_ (.Y(_0151_),
    .B(_0081_),
    .A_N(_0113_));
 sg13g2_o21ai_1 _0656_ (.B1(_0144_),
    .Y(_0152_),
    .A1(_0123_),
    .A2(_0129_));
 sg13g2_nor3_1 _0657_ (.A(_0099_),
    .B(_0109_),
    .C(net141),
    .Y(_0153_));
 sg13g2_nand4_1 _0658_ (.B(_0124_),
    .C(_0125_),
    .A(_0121_),
    .Y(_0154_),
    .D(_0151_));
 sg13g2_nor4_1 _0659_ (.A(_0134_),
    .B(_0145_),
    .C(_0150_),
    .D(_0152_),
    .Y(_0155_));
 sg13g2_nor2b_1 _0660_ (.A(_0154_),
    .B_N(_0155_),
    .Y(_0156_));
 sg13g2_a221oi_1 _0661_ (.B2(_0148_),
    .C1(_0153_),
    .B1(_0122_),
    .A1(_0081_),
    .Y(_0157_),
    .A2(_0118_));
 sg13g2_nand4_1 _0662_ (.B(_0143_),
    .C(_0156_),
    .A(_0139_),
    .Y(_0158_),
    .D(_0157_));
 sg13g2_or4_1 _0663_ (.A(\top_level.freq1_reg_out[2] ),
    .B(\top_level.freq1_reg_out[3] ),
    .C(\top_level.freq1_reg_out[4] ),
    .D(\top_level.freq1_reg_out[5] ),
    .X(_0159_));
 sg13g2_nor3_1 _0664_ (.A(\top_level.freq1_reg_out[0] ),
    .B(\top_level.freq1_reg_out[1] ),
    .C(_0159_),
    .Y(_0160_));
 sg13g2_nor3_1 _0665_ (.A(\top_level.freq1_reg_out[14] ),
    .B(\top_level.freq1_reg_out[15] ),
    .C(net163),
    .Y(_0161_));
 sg13g2_nor4_1 _0666_ (.A(\top_level.freq1_reg_out[10] ),
    .B(\top_level.freq1_reg_out[11] ),
    .C(\top_level.freq1_reg_out[12] ),
    .D(\top_level.freq1_reg_out[13] ),
    .Y(_0162_));
 sg13g2_nor4_1 _0667_ (.A(\top_level.freq1_reg_out[6] ),
    .B(\top_level.freq1_reg_out[7] ),
    .C(\top_level.freq1_reg_out[8] ),
    .D(\top_level.freq1_reg_out[9] ),
    .Y(_0163_));
 sg13g2_nand4_1 _0668_ (.B(_0161_),
    .C(_0162_),
    .A(_0160_),
    .Y(_0164_),
    .D(_0163_));
 sg13g2_nand3b_1 _0669_ (.B(net144),
    .C(_0104_),
    .Y(_0165_),
    .A_N(net141));
 sg13g2_nand2b_2 _0670_ (.Y(_0166_),
    .B(_0135_),
    .A_N(net142));
 sg13g2_nand3_1 _0671_ (.B(_0165_),
    .C(_0166_),
    .A(_0144_),
    .Y(_0167_));
 sg13g2_or2_1 _0672_ (.X(_0168_),
    .B(_0141_),
    .A(_0132_));
 sg13g2_nand3_1 _0673_ (.B(_0104_),
    .C(_0109_),
    .A(net146),
    .Y(_0169_));
 sg13g2_o21ai_1 _0674_ (.B1(_0168_),
    .Y(_0170_),
    .A1(_0136_),
    .A2(_0169_));
 sg13g2_nor2_1 _0675_ (.A(net146),
    .B(_0116_),
    .Y(_0171_));
 sg13g2_a21oi_1 _0676_ (.A1(net145),
    .A2(net143),
    .Y(_0172_),
    .B1(_0171_));
 sg13g2_nor2_1 _0677_ (.A(net141),
    .B(_0172_),
    .Y(_0173_));
 sg13g2_a21o_1 _0678_ (.A2(_0126_),
    .A1(_0099_),
    .B1(net141),
    .X(_0174_));
 sg13g2_o21ai_1 _0679_ (.B1(_0174_),
    .Y(_0175_),
    .A1(_0136_),
    .A2(_0172_));
 sg13g2_a21oi_1 _0680_ (.A1(_0113_),
    .A2(_0127_),
    .Y(_0176_),
    .B1(_0136_));
 sg13g2_nor2_1 _0681_ (.A(_0170_),
    .B(_0176_),
    .Y(_0177_));
 sg13g2_nor3_1 _0682_ (.A(_0167_),
    .B(_0173_),
    .C(_0175_),
    .Y(_0178_));
 sg13g2_and2_1 _0683_ (.A(_0118_),
    .B(_0122_),
    .X(_0179_));
 sg13g2_nor2_1 _0684_ (.A(_0123_),
    .B(_0172_),
    .Y(_0180_));
 sg13g2_a21oi_1 _0685_ (.A1(net142),
    .A2(_0116_),
    .Y(_0181_),
    .B1(_0082_));
 sg13g2_a21o_1 _0686_ (.A2(net143),
    .A1(_0081_),
    .B1(_0181_),
    .X(_0182_));
 sg13g2_a21o_1 _0687_ (.A2(_0110_),
    .A1(net144),
    .B1(net142),
    .X(_0183_));
 sg13g2_nor2_1 _0688_ (.A(_0123_),
    .B(_0183_),
    .Y(_0184_));
 sg13g2_or3_1 _0689_ (.A(_0133_),
    .B(_0182_),
    .C(_0184_),
    .X(_0185_));
 sg13g2_nor3_1 _0690_ (.A(_0179_),
    .B(_0180_),
    .C(_0185_),
    .Y(_0186_));
 sg13g2_or2_1 _0691_ (.X(_0187_),
    .B(_0119_),
    .A(_0114_));
 sg13g2_and4_1 _0692_ (.A(_0121_),
    .B(_0124_),
    .C(_0125_),
    .D(_0187_),
    .X(_0188_));
 sg13g2_nand4_1 _0693_ (.B(_0178_),
    .C(_0186_),
    .A(_0177_),
    .Y(_0189_),
    .D(_0188_));
 sg13g2_o21ai_1 _0694_ (.B1(_0164_),
    .Y(_0190_),
    .A1(_0069_),
    .A2(_0189_));
 sg13g2_and2_1 _0695_ (.A(_0069_),
    .B(_0189_),
    .X(_0191_));
 sg13g2_mux2_1 _0696_ (.A0(_0191_),
    .A1(net160),
    .S(_0158_),
    .X(_0192_));
 sg13g2_nor2_2 _0697_ (.A(_0190_),
    .B(_0192_),
    .Y(uo_out[0]));
 sg13g2_a21oi_1 _0698_ (.A1(_0113_),
    .A2(_0147_),
    .Y(_0193_),
    .B1(_0079_));
 sg13g2_o21ai_1 _0699_ (.B1(_0121_),
    .Y(_0194_),
    .A1(net144),
    .A2(_0166_));
 sg13g2_a21oi_1 _0700_ (.A1(_0120_),
    .A2(_0166_),
    .Y(_0195_),
    .B1(_0132_));
 sg13g2_o21ai_1 _0701_ (.B1(_0168_),
    .Y(_0196_),
    .A1(_0115_),
    .A2(_0120_));
 sg13g2_nor2_1 _0702_ (.A(_0082_),
    .B(_0183_),
    .Y(_0197_));
 sg13g2_nand2_1 _0703_ (.Y(_0198_),
    .A(net143),
    .B(net141));
 sg13g2_nor3_1 _0704_ (.A(_0122_),
    .B(_0132_),
    .C(_0198_),
    .Y(_0199_));
 sg13g2_nor3_1 _0705_ (.A(_0196_),
    .B(_0197_),
    .C(_0199_),
    .Y(_0200_));
 sg13g2_nor2b_1 _0706_ (.A(_0104_),
    .B_N(_0116_),
    .Y(_0201_));
 sg13g2_a21oi_1 _0707_ (.A1(_0098_),
    .A2(_0201_),
    .Y(_0202_),
    .B1(_0110_));
 sg13g2_nor2_1 _0708_ (.A(_0111_),
    .B(net142),
    .Y(_0203_));
 sg13g2_o21ai_1 _0709_ (.B1(_0122_),
    .Y(_0204_),
    .A1(_0202_),
    .A2(_0203_));
 sg13g2_nor4_1 _0710_ (.A(_0134_),
    .B(_0142_),
    .C(_0193_),
    .D(_0195_),
    .Y(_0205_));
 sg13g2_nand3_1 _0711_ (.B(_0204_),
    .C(_0205_),
    .A(_0200_),
    .Y(_0206_));
 sg13g2_mux2_1 _0712_ (.A0(_0191_),
    .A1(net159),
    .S(_0206_),
    .X(_0207_));
 sg13g2_nor2_2 _0713_ (.A(_0190_),
    .B(_0207_),
    .Y(uo_out[1]));
 sg13g2_nand2_1 _0714_ (.Y(_0208_),
    .A(_0125_),
    .B(_0187_));
 sg13g2_nand2_1 _0715_ (.Y(_0209_),
    .A(net145),
    .B(_0208_));
 sg13g2_nor2_1 _0716_ (.A(_0179_),
    .B(_0196_),
    .Y(_0210_));
 sg13g2_a21oi_1 _0717_ (.A1(_0121_),
    .A2(_0149_),
    .Y(_0211_),
    .B1(_0110_));
 sg13g2_nand2_1 _0718_ (.Y(_0212_),
    .A(_0130_),
    .B(_0133_));
 sg13g2_o21ai_1 _0719_ (.B1(_0212_),
    .Y(_0213_),
    .A1(net145),
    .A2(_0166_));
 sg13g2_nor4_1 _0720_ (.A(_0146_),
    .B(_0181_),
    .C(_0211_),
    .D(_0213_),
    .Y(_0214_));
 sg13g2_nand4_1 _0721_ (.B(_0209_),
    .C(_0210_),
    .A(_0139_),
    .Y(_0215_),
    .D(_0214_));
 sg13g2_mux2_1 _0722_ (.A0(_0191_),
    .A1(net159),
    .S(_0215_),
    .X(_0216_));
 sg13g2_nor2_1 _0723_ (.A(_0190_),
    .B(_0216_),
    .Y(uo_out[2]));
 sg13g2_or3_1 _0724_ (.A(_0179_),
    .B(_0182_),
    .C(_0194_),
    .X(_0217_));
 sg13g2_or2_1 _0725_ (.X(_0218_),
    .B(_0120_),
    .A(_0112_));
 sg13g2_nand2_1 _0726_ (.Y(_0219_),
    .A(_0074_),
    .B(_0171_));
 sg13g2_nand3_1 _0727_ (.B(_0218_),
    .C(_0219_),
    .A(_0125_),
    .Y(_0220_));
 sg13g2_o21ai_1 _0728_ (.B1(_0149_),
    .Y(_0221_),
    .A1(_0074_),
    .A2(_0169_));
 sg13g2_nor4_1 _0729_ (.A(_0170_),
    .B(_0217_),
    .C(_0220_),
    .D(_0221_),
    .Y(_0222_));
 sg13g2_mux2_1 _0730_ (.A0(net159),
    .A1(_0191_),
    .S(_0222_),
    .X(_0223_));
 sg13g2_nor2_2 _0731_ (.A(_0190_),
    .B(_0223_),
    .Y(uo_out[3]));
 sg13g2_nand2_1 _0732_ (.Y(_0224_),
    .A(_0165_),
    .B(_0168_));
 sg13g2_nor4_1 _0733_ (.A(_0175_),
    .B(_0185_),
    .C(_0208_),
    .D(_0224_),
    .Y(_0225_));
 sg13g2_mux2_1 _0734_ (.A0(net159),
    .A1(_0191_),
    .S(_0225_),
    .X(_0226_));
 sg13g2_nor2_1 _0735_ (.A(_0190_),
    .B(_0226_),
    .Y(uo_out[4]));
 sg13g2_nor2b_1 _0736_ (.A(_0167_),
    .B_N(_0124_),
    .Y(_0227_));
 sg13g2_and3_1 _0737_ (.X(_0228_),
    .A(_0174_),
    .B(_0186_),
    .C(_0227_));
 sg13g2_mux2_1 _0738_ (.A0(net159),
    .A1(_0191_),
    .S(_0228_),
    .X(_0229_));
 sg13g2_nor2_1 _0739_ (.A(_0190_),
    .B(_0229_),
    .Y(uo_out[5]));
 sg13g2_a21oi_1 _0740_ (.A1(_0177_),
    .A2(_0178_),
    .Y(_0230_),
    .B1(_0173_));
 sg13g2_xnor2_1 _0741_ (.Y(_0231_),
    .A(net159),
    .B(_0230_));
 sg13g2_and2_1 _0742_ (.A(_0164_),
    .B(_0231_),
    .X(uo_out[6]));
 sg13g2_or2_1 _0743_ (.X(uo_out[7]),
    .B(_0191_),
    .A(_0190_));
 sg13g2_mux2_1 _0744_ (.A0(net23),
    .A1(\top_level.freq1_reg_out[0] ),
    .S(net3),
    .X(_0232_));
 sg13g2_nand2_1 _0745_ (.Y(_0233_),
    .A(net34),
    .B(_0232_));
 sg13g2_mux2_1 _0746_ (.A0(\top_level.freq0_reg_out[1] ),
    .A1(\top_level.freq1_reg_out[1] ),
    .S(net165),
    .X(_0234_));
 sg13g2_nand2_1 _0747_ (.Y(_0235_),
    .A(net76),
    .B(_0234_));
 sg13g2_xnor2_1 _0748_ (.Y(_0236_),
    .A(net76),
    .B(_0234_));
 sg13g2_xor2_1 _0749_ (.B(_0236_),
    .A(_0233_),
    .X(\top_level.adder.sum[1] ));
 sg13g2_o21ai_1 _0750_ (.B1(_0235_),
    .Y(_0237_),
    .A1(_0233_),
    .A2(_0236_));
 sg13g2_mux2_1 _0751_ (.A0(\top_level.freq0_reg_out[2] ),
    .A1(\top_level.freq1_reg_out[2] ),
    .S(net165),
    .X(_0238_));
 sg13g2_and2_1 _0752_ (.A(net93),
    .B(_0238_),
    .X(_0239_));
 sg13g2_or2_1 _0753_ (.X(_0240_),
    .B(_0238_),
    .A(net93));
 sg13g2_nand2b_1 _0754_ (.Y(_0241_),
    .B(_0240_),
    .A_N(_0239_));
 sg13g2_xnor2_1 _0755_ (.Y(\top_level.adder.sum[2] ),
    .A(_0237_),
    .B(_0241_));
 sg13g2_mux2_1 _0756_ (.A0(\top_level.freq0_reg_out[3] ),
    .A1(\top_level.freq1_reg_out[3] ),
    .S(net165),
    .X(_0242_));
 sg13g2_nor2b_1 _0757_ (.A(net89),
    .B_N(_0242_),
    .Y(_0243_));
 sg13g2_xnor2_1 _0758_ (.Y(_0244_),
    .A(net89),
    .B(_0242_));
 sg13g2_a21o_1 _0759_ (.A2(_0240_),
    .A1(_0237_),
    .B1(_0239_),
    .X(_0245_));
 sg13g2_xor2_1 _0760_ (.B(_0245_),
    .A(_0244_),
    .X(\top_level.adder.sum[3] ));
 sg13g2_a21oi_2 _0761_ (.B1(_0243_),
    .Y(_0246_),
    .A2(_0245_),
    .A1(_0244_));
 sg13g2_mux2_1 _0762_ (.A0(\top_level.freq0_reg_out[4] ),
    .A1(\top_level.freq1_reg_out[4] ),
    .S(net165),
    .X(_0247_));
 sg13g2_and2_1 _0763_ (.A(\top_level.adder.b[4] ),
    .B(_0247_),
    .X(_0248_));
 sg13g2_xnor2_1 _0764_ (.Y(_0249_),
    .A(\top_level.adder.b[4] ),
    .B(_0247_));
 sg13g2_nor2_1 _0765_ (.A(_0246_),
    .B(_0249_),
    .Y(_0250_));
 sg13g2_xor2_1 _0766_ (.B(_0249_),
    .A(_0246_),
    .X(\top_level.adder.sum[4] ));
 sg13g2_nor2_1 _0767_ (.A(\top_level.freq0_reg_out[5] ),
    .B(net165),
    .Y(_0251_));
 sg13g2_nor2b_1 _0768_ (.A(\top_level.freq1_reg_out[5] ),
    .B_N(net165),
    .Y(_0252_));
 sg13g2_o21ai_1 _0769_ (.B1(net100),
    .Y(_0253_),
    .A1(_0251_),
    .A2(_0252_));
 sg13g2_inv_1 _0770_ (.Y(_0254_),
    .A(_0253_));
 sg13g2_nor3_1 _0771_ (.A(net100),
    .B(_0251_),
    .C(_0252_),
    .Y(_0255_));
 sg13g2_nor2_1 _0772_ (.A(_0254_),
    .B(_0255_),
    .Y(_0256_));
 sg13g2_nor2_1 _0773_ (.A(_0248_),
    .B(_0250_),
    .Y(_0257_));
 sg13g2_xnor2_1 _0774_ (.Y(\top_level.adder.sum[5] ),
    .A(_0256_),
    .B(_0257_));
 sg13g2_mux2_1 _0775_ (.A0(\top_level.freq0_reg_out[6] ),
    .A1(\top_level.freq1_reg_out[6] ),
    .S(net164),
    .X(_0258_));
 sg13g2_and2_1 _0776_ (.A(net115),
    .B(_0258_),
    .X(_0259_));
 sg13g2_or2_1 _0777_ (.X(_0260_),
    .B(_0258_),
    .A(net115));
 sg13g2_nand2b_1 _0778_ (.Y(_0261_),
    .B(_0260_),
    .A_N(_0259_));
 sg13g2_or4_2 _0779_ (.A(_0246_),
    .B(_0249_),
    .C(_0254_),
    .D(_0255_),
    .X(_0262_));
 sg13g2_a21oi_1 _0780_ (.A1(_0248_),
    .A2(_0253_),
    .Y(_0263_),
    .B1(_0255_));
 sg13g2_nand2_1 _0781_ (.Y(_0264_),
    .A(_0262_),
    .B(_0263_));
 sg13g2_xnor2_1 _0782_ (.Y(\top_level.adder.sum[6] ),
    .A(_0261_),
    .B(_0264_));
 sg13g2_nor2_1 _0783_ (.A(\top_level.freq0_reg_out[7] ),
    .B(net163),
    .Y(_0265_));
 sg13g2_nor2b_1 _0784_ (.A(\top_level.freq1_reg_out[7] ),
    .B_N(net164),
    .Y(_0266_));
 sg13g2_or3_1 _0785_ (.A(net95),
    .B(_0265_),
    .C(_0266_),
    .X(_0267_));
 sg13g2_inv_1 _0786_ (.Y(_0268_),
    .A(_0267_));
 sg13g2_o21ai_1 _0787_ (.B1(net95),
    .Y(_0269_),
    .A1(_0265_),
    .A2(_0266_));
 sg13g2_nand2_1 _0788_ (.Y(_0270_),
    .A(_0267_),
    .B(_0269_));
 sg13g2_a21oi_1 _0789_ (.A1(_0260_),
    .A2(_0264_),
    .Y(_0271_),
    .B1(_0259_));
 sg13g2_xor2_1 _0790_ (.B(_0271_),
    .A(_0270_),
    .X(\top_level.adder.sum[7] ));
 sg13g2_a21oi_1 _0791_ (.A1(_0259_),
    .A2(_0269_),
    .Y(_0272_),
    .B1(_0268_));
 sg13g2_and2_1 _0792_ (.A(_0263_),
    .B(_0272_),
    .X(_0273_));
 sg13g2_a21oi_1 _0793_ (.A1(_0260_),
    .A2(_0269_),
    .Y(_0274_),
    .B1(_0268_));
 sg13g2_a21oi_1 _0794_ (.A1(_0262_),
    .A2(_0273_),
    .Y(_0275_),
    .B1(_0274_));
 sg13g2_a21o_1 _0795_ (.A2(_0273_),
    .A1(_0262_),
    .B1(_0274_),
    .X(_0276_));
 sg13g2_mux2_1 _0796_ (.A0(\top_level.freq0_reg_out[8] ),
    .A1(\top_level.freq1_reg_out[8] ),
    .S(net164),
    .X(_0277_));
 sg13g2_xnor2_1 _0797_ (.Y(_0278_),
    .A(net94),
    .B(_0277_));
 sg13g2_inv_1 _0798_ (.Y(_0279_),
    .A(_0278_));
 sg13g2_xnor2_1 _0799_ (.Y(\top_level.adder.sum[8] ),
    .A(_0276_),
    .B(_0278_));
 sg13g2_mux2_1 _0800_ (.A0(\top_level.freq0_reg_out[9] ),
    .A1(\top_level.freq1_reg_out[9] ),
    .S(net164),
    .X(_0280_));
 sg13g2_nor2b_1 _0801_ (.A(_0280_),
    .B_N(_0008_),
    .Y(_0281_));
 sg13g2_nand2b_1 _0802_ (.Y(_0282_),
    .B(_0280_),
    .A_N(_0008_));
 sg13g2_nor2b_1 _0803_ (.A(_0281_),
    .B_N(_0282_),
    .Y(_0283_));
 sg13g2_nand2_1 _0804_ (.Y(_0284_),
    .A(net109),
    .B(_0277_));
 sg13g2_o21ai_1 _0805_ (.B1(_0284_),
    .Y(_0285_),
    .A1(_0276_),
    .A2(_0279_));
 sg13g2_xor2_1 _0806_ (.B(_0285_),
    .A(_0283_),
    .X(\top_level.adder.sum[9] ));
 sg13g2_o21ai_1 _0807_ (.B1(_0282_),
    .Y(_0286_),
    .A1(_0281_),
    .A2(_0284_));
 sg13g2_inv_1 _0808_ (.Y(_0287_),
    .A(_0286_));
 sg13g2_nand2_1 _0809_ (.Y(_0288_),
    .A(_0278_),
    .B(_0283_));
 sg13g2_o21ai_1 _0810_ (.B1(_0287_),
    .Y(_0289_),
    .A1(_0276_),
    .A2(_0288_));
 sg13g2_mux2_1 _0811_ (.A0(\top_level.freq0_reg_out[10] ),
    .A1(\top_level.freq1_reg_out[10] ),
    .S(net163),
    .X(_0290_));
 sg13g2_xnor2_1 _0812_ (.Y(_0291_),
    .A(net116),
    .B(_0290_));
 sg13g2_inv_1 _0813_ (.Y(_0292_),
    .A(_0291_));
 sg13g2_xnor2_1 _0814_ (.Y(\top_level.adder.sum[10] ),
    .A(_0289_),
    .B(_0292_));
 sg13g2_a22oi_1 _0815_ (.Y(_0293_),
    .B1(_0291_),
    .B2(_0289_),
    .A2(_0290_),
    .A1(net97));
 sg13g2_mux2_1 _0816_ (.A0(\top_level.freq0_reg_out[11] ),
    .A1(\top_level.freq1_reg_out[11] ),
    .S(net163),
    .X(_0294_));
 sg13g2_xor2_1 _0817_ (.B(_0294_),
    .A(_0010_),
    .X(_0295_));
 sg13g2_xor2_1 _0818_ (.B(_0295_),
    .A(net98),
    .X(\top_level.adder.sum[11] ));
 sg13g2_nor3_1 _0819_ (.A(_0288_),
    .B(_0292_),
    .C(_0295_),
    .Y(_0296_));
 sg13g2_a22oi_1 _0820_ (.Y(_0297_),
    .B1(_0291_),
    .B2(_0286_),
    .A2(_0290_),
    .A1(\top_level.adder.b[10] ));
 sg13g2_nor2_1 _0821_ (.A(_0295_),
    .B(_0297_),
    .Y(_0298_));
 sg13g2_a221oi_1 _0822_ (.B2(_0275_),
    .C1(_0298_),
    .B1(_0296_),
    .A1(\top_level.adder.b[11] ),
    .Y(_0299_),
    .A2(_0294_));
 sg13g2_inv_1 _0823_ (.Y(_0300_),
    .A(_0299_));
 sg13g2_mux2_1 _0824_ (.A0(\top_level.freq0_reg_out[12] ),
    .A1(\top_level.freq1_reg_out[12] ),
    .S(net163),
    .X(_0301_));
 sg13g2_xnor2_1 _0825_ (.Y(_0302_),
    .A(net107),
    .B(_0301_));
 sg13g2_xnor2_1 _0826_ (.Y(\top_level.adder.sum[12] ),
    .A(_0299_),
    .B(_0302_));
 sg13g2_mux2_1 _0827_ (.A0(\top_level.freq0_reg_out[13] ),
    .A1(\top_level.freq1_reg_out[13] ),
    .S(net163),
    .X(_0303_));
 sg13g2_xnor2_1 _0828_ (.Y(_0304_),
    .A(_0012_),
    .B(_0303_));
 sg13g2_and2_1 _0829_ (.A(net103),
    .B(_0301_),
    .X(_0305_));
 sg13g2_a21oi_1 _0830_ (.A1(_0300_),
    .A2(_0302_),
    .Y(_0306_),
    .B1(_0305_));
 sg13g2_nand2_1 _0831_ (.Y(_0307_),
    .A(_0302_),
    .B(_0304_));
 sg13g2_xnor2_1 _0832_ (.Y(\top_level.adder.sum[13] ),
    .A(_0304_),
    .B(_0306_));
 sg13g2_mux2_1 _0833_ (.A0(\top_level.freq0_reg_out[14] ),
    .A1(\top_level.freq1_reg_out[14] ),
    .S(net163),
    .X(_0308_));
 sg13g2_and2_1 _0834_ (.A(net162),
    .B(_0308_),
    .X(_0309_));
 sg13g2_xnor2_1 _0835_ (.Y(_0310_),
    .A(net162),
    .B(_0308_));
 sg13g2_inv_1 _0836_ (.Y(_0311_),
    .A(_0310_));
 sg13g2_a22oi_1 _0837_ (.Y(_0312_),
    .B1(_0304_),
    .B2(_0305_),
    .A2(_0303_),
    .A1(net113));
 sg13g2_o21ai_1 _0838_ (.B1(_0312_),
    .Y(_0313_),
    .A1(_0299_),
    .A2(_0307_));
 sg13g2_xnor2_1 _0839_ (.Y(\top_level.adder.sum[14] ),
    .A(_0310_),
    .B(_0313_));
 sg13g2_a21oi_1 _0840_ (.A1(_0311_),
    .A2(_0313_),
    .Y(_0314_),
    .B1(_0309_));
 sg13g2_mux2_1 _0841_ (.A0(net28),
    .A1(net49),
    .S(net163),
    .X(_0315_));
 sg13g2_xnor2_1 _0842_ (.Y(_0316_),
    .A(net68),
    .B(_0315_));
 sg13g2_xnor2_1 _0843_ (.Y(\top_level.adder.sum[15] ),
    .A(_0314_),
    .B(_0316_));
 sg13g2_xor2_1 _0844_ (.B(_0232_),
    .A(net34),
    .X(\top_level.adder.sum[0] ));
 sg13g2_nor4_2 _0845_ (.A(\top_level.uart.clk_count_reg[5] ),
    .B(\top_level.uart.clk_count_reg[4] ),
    .C(\top_level.uart.clk_count_reg[7] ),
    .Y(_0317_),
    .D(net50));
 sg13g2_nor2_1 _0846_ (.A(\top_level.uart.clk_count_reg[3] ),
    .B(\top_level.uart.clk_count_reg[8] ),
    .Y(_0318_));
 sg13g2_a21oi_1 _0847_ (.A1(_0317_),
    .A2(_0318_),
    .Y(_0319_),
    .B1(_0065_));
 sg13g2_nor3_2 _0848_ (.A(net74),
    .B(\top_level.uart.clk_count_reg[10] ),
    .C(_0319_),
    .Y(_0320_));
 sg13g2_or3_1 _0849_ (.A(\top_level.uart.clk_count_reg[11] ),
    .B(\top_level.uart.clk_count_reg[10] ),
    .C(_0319_),
    .X(_0321_));
 sg13g2_nand2_1 _0850_ (.Y(_0322_),
    .A(\top_level.uart.state_reg[0] ),
    .B(_0003_));
 sg13g2_nand2_1 _0851_ (.Y(_0323_),
    .A(\top_level.uart.state_reg[0] ),
    .B(\top_level.uart.state_reg[1] ));
 sg13g2_nand3_1 _0852_ (.B(\top_level.uart.state_reg[1] ),
    .C(net119),
    .A(\top_level.uart.state_reg[0] ),
    .Y(_0324_));
 sg13g2_nor2_2 _0853_ (.A(_0320_),
    .B(_0324_),
    .Y(_0325_));
 sg13g2_and2_1 _0854_ (.A(net2),
    .B(_0325_),
    .X(_0326_));
 sg13g2_nand2_1 _0855_ (.Y(_0327_),
    .A(net2),
    .B(_0325_));
 sg13g2_nor2_1 _0856_ (.A(net155),
    .B(net137),
    .Y(_0328_));
 sg13g2_nand2b_2 _0857_ (.Y(_0329_),
    .B(_0326_),
    .A_N(net154));
 sg13g2_nor2b_2 _0858_ (.A(\top_level.uart.bit_index_reg[1] ),
    .B_N(\top_level.uart.bit_index_reg[0] ),
    .Y(_0330_));
 sg13g2_nor2b_1 _0859_ (.A(net151),
    .B_N(_0330_),
    .Y(_0331_));
 sg13g2_nand2b_1 _0860_ (.Y(_0332_),
    .B(_0330_),
    .A_N(net150));
 sg13g2_nand2b_1 _0861_ (.Y(_0333_),
    .B(_0331_),
    .A_N(net148));
 sg13g2_o21ai_1 _0862_ (.B1(net62),
    .Y(_0334_),
    .A1(_0329_),
    .A2(_0333_));
 sg13g2_nor2_1 _0863_ (.A(\top_level.uart.bit_index_reg[1] ),
    .B(net152),
    .Y(_0335_));
 sg13g2_nor3_2 _0864_ (.A(\top_level.uart.bit_index_reg[1] ),
    .B(net152),
    .C(net151),
    .Y(_0336_));
 sg13g2_nand2_1 _0865_ (.Y(_0337_),
    .A(net148),
    .B(_0336_));
 sg13g2_nand2b_1 _0866_ (.Y(_0338_),
    .B(_0336_),
    .A_N(net149));
 sg13g2_nand2b_1 _0867_ (.Y(_0339_),
    .B(net149),
    .A_N(_0336_));
 sg13g2_nand3b_1 _0868_ (.B(_0338_),
    .C(_0339_),
    .Y(_0340_),
    .A_N(net155));
 sg13g2_nor2_2 _0869_ (.A(_0067_),
    .B(_0340_),
    .Y(_0341_));
 sg13g2_nand2_1 _0870_ (.Y(_0342_),
    .A(_0331_),
    .B(_0341_));
 sg13g2_o21ai_1 _0871_ (.B1(_0334_),
    .Y(_0013_),
    .A1(net137),
    .A2(_0342_));
 sg13g2_nor3_2 _0872_ (.A(_0068_),
    .B(net152),
    .C(net151),
    .Y(_0343_));
 sg13g2_nand2b_1 _0873_ (.Y(_0344_),
    .B(_0343_),
    .A_N(\top_level.uart.bit_index_reg[3] ));
 sg13g2_o21ai_1 _0874_ (.B1(net56),
    .Y(_0345_),
    .A1(_0329_),
    .A2(_0344_));
 sg13g2_nand2_1 _0875_ (.Y(_0346_),
    .A(_0341_),
    .B(_0343_));
 sg13g2_o21ai_1 _0876_ (.B1(net57),
    .Y(_0014_),
    .A1(net137),
    .A2(_0346_));
 sg13g2_and2_1 _0877_ (.A(\top_level.uart.bit_index_reg[1] ),
    .B(net152),
    .X(_0347_));
 sg13g2_nand2_1 _0878_ (.Y(_0348_),
    .A(\top_level.uart.bit_index_reg[1] ),
    .B(net152));
 sg13g2_nor2_2 _0879_ (.A(net150),
    .B(_0348_),
    .Y(_0349_));
 sg13g2_nand2b_1 _0880_ (.Y(_0350_),
    .B(_0349_),
    .A_N(net148));
 sg13g2_o21ai_1 _0881_ (.B1(net67),
    .Y(_0351_),
    .A1(_0329_),
    .A2(_0350_));
 sg13g2_nand2_1 _0882_ (.Y(_0352_),
    .A(_0341_),
    .B(_0349_));
 sg13g2_o21ai_1 _0883_ (.B1(_0351_),
    .Y(_0015_),
    .A1(net137),
    .A2(_0352_));
 sg13g2_nand2_2 _0884_ (.Y(_0353_),
    .A(net151),
    .B(_0335_));
 sg13g2_or2_1 _0885_ (.X(_0354_),
    .B(_0353_),
    .A(net148));
 sg13g2_o21ai_1 _0886_ (.B1(net54),
    .Y(_0355_),
    .A1(_0329_),
    .A2(_0354_));
 sg13g2_nand3_1 _0887_ (.B(_0335_),
    .C(_0341_),
    .A(net151),
    .Y(_0356_));
 sg13g2_o21ai_1 _0888_ (.B1(_0355_),
    .Y(_0016_),
    .A1(net137),
    .A2(_0356_));
 sg13g2_and2_1 _0889_ (.A(net150),
    .B(_0330_),
    .X(_0357_));
 sg13g2_nand2_1 _0890_ (.Y(_0358_),
    .A(net150),
    .B(_0330_));
 sg13g2_nand2b_1 _0891_ (.Y(_0359_),
    .B(_0357_),
    .A_N(net148));
 sg13g2_o21ai_1 _0892_ (.B1(net53),
    .Y(_0360_),
    .A1(_0329_),
    .A2(_0359_));
 sg13g2_nand2_1 _0893_ (.Y(_0361_),
    .A(_0341_),
    .B(_0357_));
 sg13g2_o21ai_1 _0894_ (.B1(_0360_),
    .Y(_0017_),
    .A1(net137),
    .A2(_0361_));
 sg13g2_nand3b_1 _0895_ (.B(net150),
    .C(\top_level.uart.bit_index_reg[1] ),
    .Y(_0362_),
    .A_N(net152));
 sg13g2_or2_1 _0896_ (.X(_0363_),
    .B(_0362_),
    .A(net148));
 sg13g2_o21ai_1 _0897_ (.B1(net71),
    .Y(_0364_),
    .A1(_0329_),
    .A2(_0363_));
 sg13g2_or3_1 _0898_ (.A(net147),
    .B(_0340_),
    .C(_0362_),
    .X(_0365_));
 sg13g2_o21ai_1 _0899_ (.B1(_0364_),
    .Y(_0018_),
    .A1(net136),
    .A2(_0365_));
 sg13g2_and2_2 _0900_ (.A(net150),
    .B(_0347_),
    .X(_0366_));
 sg13g2_nand2_1 _0901_ (.Y(_0367_),
    .A(net150),
    .B(_0347_));
 sg13g2_nand2b_1 _0902_ (.Y(_0368_),
    .B(_0366_),
    .A_N(net148));
 sg13g2_o21ai_1 _0903_ (.B1(net64),
    .Y(_0369_),
    .A1(_0329_),
    .A2(_0368_));
 sg13g2_nand2_1 _0904_ (.Y(_0370_),
    .A(_0341_),
    .B(_0366_));
 sg13g2_o21ai_1 _0905_ (.B1(_0369_),
    .Y(_0019_),
    .A1(net136),
    .A2(_0370_));
 sg13g2_nand2b_1 _0906_ (.Y(_0371_),
    .B(net153),
    .A_N(_0005_));
 sg13g2_nand2_1 _0907_ (.Y(_0372_),
    .A(net73),
    .B(_0337_));
 sg13g2_nand3_1 _0908_ (.B(net148),
    .C(_0336_),
    .A(net156),
    .Y(_0373_));
 sg13g2_a21oi_1 _0909_ (.A1(_0372_),
    .A2(_0373_),
    .Y(_0374_),
    .B1(net154));
 sg13g2_nand2_2 _0910_ (.Y(_0375_),
    .A(_0005_),
    .B(_0336_));
 sg13g2_nand2_1 _0911_ (.Y(_0376_),
    .A(net73),
    .B(_0375_));
 sg13g2_o21ai_1 _0912_ (.B1(_0376_),
    .Y(_0377_),
    .A1(net147),
    .A2(_0375_));
 sg13g2_a21oi_1 _0913_ (.A1(net154),
    .A2(_0377_),
    .Y(_0378_),
    .B1(_0374_));
 sg13g2_nand2_1 _0914_ (.Y(_0379_),
    .A(net73),
    .B(net136));
 sg13g2_o21ai_1 _0915_ (.B1(_0379_),
    .Y(_0020_),
    .A1(net136),
    .A2(_0378_));
 sg13g2_and2_1 _0916_ (.A(net156),
    .B(_0340_),
    .X(_0380_));
 sg13g2_nand2_1 _0917_ (.Y(_0381_),
    .A(_0371_),
    .B(_0380_));
 sg13g2_nor2_1 _0918_ (.A(_0332_),
    .B(_0381_),
    .Y(_0382_));
 sg13g2_a21oi_1 _0919_ (.A1(net138),
    .A2(_0382_),
    .Y(_0383_),
    .B1(net44));
 sg13g2_o21ai_1 _0920_ (.B1(_0371_),
    .Y(_0384_),
    .A1(net149),
    .A2(net153));
 sg13g2_inv_1 _0921_ (.Y(_0385_),
    .A(_0384_));
 sg13g2_nand2_1 _0922_ (.Y(_0386_),
    .A(net147),
    .B(_0385_));
 sg13g2_nor2_1 _0923_ (.A(_0332_),
    .B(_0386_),
    .Y(_0387_));
 sg13g2_a21oi_1 _0924_ (.A1(net138),
    .A2(_0387_),
    .Y(_0021_),
    .B1(_0383_));
 sg13g2_nand3_1 _0925_ (.B(_0371_),
    .C(_0380_),
    .A(_0343_),
    .Y(_0388_));
 sg13g2_nand2_1 _0926_ (.Y(_0389_),
    .A(_0343_),
    .B(_0385_));
 sg13g2_o21ai_1 _0927_ (.B1(net60),
    .Y(_0390_),
    .A1(net136),
    .A2(_0389_));
 sg13g2_o21ai_1 _0928_ (.B1(_0390_),
    .Y(_0022_),
    .A1(net136),
    .A2(_0388_));
 sg13g2_nor3_1 _0929_ (.A(net150),
    .B(_0348_),
    .C(_0381_),
    .Y(_0391_));
 sg13g2_a21oi_1 _0930_ (.A1(net138),
    .A2(_0391_),
    .Y(_0392_),
    .B1(net48));
 sg13g2_o21ai_1 _0931_ (.B1(_0386_),
    .Y(_0393_),
    .A1(net154),
    .A2(_0337_));
 sg13g2_and2_1 _0932_ (.A(_0349_),
    .B(_0393_),
    .X(_0394_));
 sg13g2_a21oi_1 _0933_ (.A1(net138),
    .A2(_0394_),
    .Y(_0023_),
    .B1(_0392_));
 sg13g2_nor3_1 _0934_ (.A(net136),
    .B(_0353_),
    .C(_0384_),
    .Y(_0395_));
 sg13g2_nor3_1 _0935_ (.A(net147),
    .B(_0353_),
    .C(_0384_),
    .Y(_0396_));
 sg13g2_mux2_1 _0936_ (.A0(net65),
    .A1(net156),
    .S(_0395_),
    .X(_0024_));
 sg13g2_nand3_1 _0937_ (.B(_0005_),
    .C(_0357_),
    .A(net156),
    .Y(_0397_));
 sg13g2_a21oi_1 _0938_ (.A1(_0357_),
    .A2(_0380_),
    .Y(_0398_),
    .B1(net153));
 sg13g2_a21oi_1 _0939_ (.A1(net153),
    .A2(_0397_),
    .Y(_0399_),
    .B1(_0398_));
 sg13g2_a21oi_1 _0940_ (.A1(net138),
    .A2(_0399_),
    .Y(_0400_),
    .B1(net45));
 sg13g2_nand3_1 _0941_ (.B(net153),
    .C(_0005_),
    .A(net147),
    .Y(_0401_));
 sg13g2_nand2_1 _0942_ (.Y(_0402_),
    .A(net149),
    .B(_0398_));
 sg13g2_a21oi_1 _0943_ (.A1(_0401_),
    .A2(_0402_),
    .Y(_0403_),
    .B1(_0358_));
 sg13g2_a21oi_1 _0944_ (.A1(net138),
    .A2(_0403_),
    .Y(_0025_),
    .B1(_0400_));
 sg13g2_nor3_1 _0945_ (.A(net136),
    .B(_0362_),
    .C(_0384_),
    .Y(_0404_));
 sg13g2_nor2_1 _0946_ (.A(net63),
    .B(_0404_),
    .Y(_0405_));
 sg13g2_a21oi_1 _0947_ (.A1(net147),
    .A2(_0404_),
    .Y(_0026_),
    .B1(_0405_));
 sg13g2_nand3_1 _0948_ (.B(_0005_),
    .C(_0366_),
    .A(net156),
    .Y(_0406_));
 sg13g2_a21oi_1 _0949_ (.A1(_0366_),
    .A2(_0380_),
    .Y(_0407_),
    .B1(net153));
 sg13g2_a21oi_1 _0950_ (.A1(net153),
    .A2(_0406_),
    .Y(_0408_),
    .B1(_0407_));
 sg13g2_a21oi_1 _0951_ (.A1(net138),
    .A2(_0408_),
    .Y(_0409_),
    .B1(net49));
 sg13g2_nand2_1 _0952_ (.Y(_0410_),
    .A(net149),
    .B(_0407_));
 sg13g2_a21oi_1 _0953_ (.A1(_0401_),
    .A2(_0410_),
    .Y(_0411_),
    .B1(_0367_));
 sg13g2_a21oi_1 _0954_ (.A1(net138),
    .A2(_0411_),
    .Y(_0027_),
    .B1(_0409_));
 sg13g2_nor3_1 _0955_ (.A(net2),
    .B(_0320_),
    .C(_0324_),
    .Y(_0412_));
 sg13g2_nand2b_2 _0956_ (.Y(_0413_),
    .B(_0325_),
    .A_N(net2));
 sg13g2_nor2_1 _0957_ (.A(net155),
    .B(_0413_),
    .Y(_0414_));
 sg13g2_nand2b_2 _0958_ (.Y(_0415_),
    .B(net140),
    .A_N(net153));
 sg13g2_o21ai_1 _0959_ (.B1(net41),
    .Y(_0416_),
    .A1(_0333_),
    .A2(_0415_));
 sg13g2_o21ai_1 _0960_ (.B1(_0416_),
    .Y(_0028_),
    .A1(_0342_),
    .A2(net135));
 sg13g2_o21ai_1 _0961_ (.B1(net31),
    .Y(_0417_),
    .A1(_0344_),
    .A2(_0415_));
 sg13g2_o21ai_1 _0962_ (.B1(net32),
    .Y(_0029_),
    .A1(_0346_),
    .A2(net135));
 sg13g2_o21ai_1 _0963_ (.B1(net33),
    .Y(_0418_),
    .A1(_0350_),
    .A2(_0415_));
 sg13g2_o21ai_1 _0964_ (.B1(_0418_),
    .Y(_0030_),
    .A1(_0352_),
    .A2(_0413_));
 sg13g2_o21ai_1 _0965_ (.B1(net29),
    .Y(_0419_),
    .A1(_0354_),
    .A2(_0415_));
 sg13g2_o21ai_1 _0966_ (.B1(_0419_),
    .Y(_0031_),
    .A1(_0356_),
    .A2(_0413_));
 sg13g2_o21ai_1 _0967_ (.B1(net51),
    .Y(_0420_),
    .A1(_0359_),
    .A2(_0415_));
 sg13g2_o21ai_1 _0968_ (.B1(_0420_),
    .Y(_0032_),
    .A1(_0361_),
    .A2(net135));
 sg13g2_o21ai_1 _0969_ (.B1(net36),
    .Y(_0421_),
    .A1(_0363_),
    .A2(_0415_));
 sg13g2_o21ai_1 _0970_ (.B1(_0421_),
    .Y(_0033_),
    .A1(_0365_),
    .A2(net135));
 sg13g2_o21ai_1 _0971_ (.B1(net52),
    .Y(_0422_),
    .A1(_0368_),
    .A2(_0415_));
 sg13g2_o21ai_1 _0972_ (.B1(_0422_),
    .Y(_0034_),
    .A1(_0370_),
    .A2(net135));
 sg13g2_nand2_1 _0973_ (.Y(_0423_),
    .A(net61),
    .B(_0337_));
 sg13g2_a21oi_1 _0974_ (.A1(_0373_),
    .A2(_0423_),
    .Y(_0424_),
    .B1(net154));
 sg13g2_nand2_1 _0975_ (.Y(_0425_),
    .A(net61),
    .B(_0375_));
 sg13g2_o21ai_1 _0976_ (.B1(_0425_),
    .Y(_0426_),
    .A1(net147),
    .A2(_0375_));
 sg13g2_a21oi_1 _0977_ (.A1(net154),
    .A2(_0426_),
    .Y(_0427_),
    .B1(_0424_));
 sg13g2_nor2_1 _0978_ (.A(net61),
    .B(net140),
    .Y(_0428_));
 sg13g2_a21oi_1 _0979_ (.A1(net140),
    .A2(_0427_),
    .Y(_0035_),
    .B1(_0428_));
 sg13g2_a21oi_1 _0980_ (.A1(_0382_),
    .A2(net139),
    .Y(_0429_),
    .B1(net21));
 sg13g2_a21oi_1 _0981_ (.A1(_0387_),
    .A2(net139),
    .Y(_0036_),
    .B1(_0429_));
 sg13g2_o21ai_1 _0982_ (.B1(net39),
    .Y(_0430_),
    .A1(_0389_),
    .A2(net135));
 sg13g2_o21ai_1 _0983_ (.B1(_0430_),
    .Y(_0037_),
    .A1(_0388_),
    .A2(net135));
 sg13g2_a21oi_1 _0984_ (.A1(_0391_),
    .A2(net140),
    .Y(_0431_),
    .B1(net22));
 sg13g2_a21oi_1 _0985_ (.A1(_0394_),
    .A2(net140),
    .Y(_0038_),
    .B1(_0431_));
 sg13g2_a21oi_1 _0986_ (.A1(_0396_),
    .A2(net139),
    .Y(_0432_),
    .B1(net27));
 sg13g2_nor2_1 _0987_ (.A(_0353_),
    .B(_0386_),
    .Y(_0433_));
 sg13g2_a21oi_1 _0988_ (.A1(net139),
    .A2(_0433_),
    .Y(_0039_),
    .B1(_0432_));
 sg13g2_a21oi_1 _0989_ (.A1(_0399_),
    .A2(net139),
    .Y(_0434_),
    .B1(net26));
 sg13g2_a21oi_1 _0990_ (.A1(_0403_),
    .A2(net139),
    .Y(_0040_),
    .B1(_0434_));
 sg13g2_nor3_1 _0991_ (.A(_0362_),
    .B(_0384_),
    .C(net135),
    .Y(_0435_));
 sg13g2_mux2_1 _0992_ (.A0(net40),
    .A1(net156),
    .S(_0435_),
    .X(_0041_));
 sg13g2_a21oi_1 _0993_ (.A1(_0408_),
    .A2(net139),
    .Y(_0436_),
    .B1(net28));
 sg13g2_a21oi_1 _0994_ (.A1(_0411_),
    .A2(net139),
    .Y(_0042_),
    .B1(_0436_));
 sg13g2_nand3_1 _0995_ (.B(\top_level.uart.clk_count_reg[0] ),
    .C(net69),
    .A(\top_level.uart.clk_count_reg[1] ),
    .Y(_0437_));
 sg13g2_and4_1 _0996_ (.A(\top_level.uart.clk_count_reg[1] ),
    .B(\top_level.uart.clk_count_reg[0] ),
    .C(\top_level.uart.clk_count_reg[3] ),
    .D(\top_level.uart.clk_count_reg[2] ),
    .X(_0438_));
 sg13g2_and2_1 _0997_ (.A(\top_level.uart.clk_count_reg[4] ),
    .B(_0438_),
    .X(_0439_));
 sg13g2_and2_1 _0998_ (.A(net46),
    .B(_0439_),
    .X(_0440_));
 sg13g2_and2_1 _0999_ (.A(net50),
    .B(_0440_),
    .X(_0441_));
 sg13g2_inv_1 _1000_ (.Y(_0442_),
    .A(_0441_));
 sg13g2_and3_1 _1001_ (.X(_0443_),
    .A(\top_level.uart.clk_count_reg[7] ),
    .B(\top_level.uart.clk_count_reg[8] ),
    .C(_0441_));
 sg13g2_a21oi_1 _1002_ (.A1(\top_level.uart.clk_count_reg[7] ),
    .A2(_0441_),
    .Y(_0444_),
    .B1(net58));
 sg13g2_or2_1 _1003_ (.X(_0445_),
    .B(_0444_),
    .A(_0443_));
 sg13g2_nor3_1 _1004_ (.A(\top_level.uart.clk_count_reg[1] ),
    .B(\top_level.uart.clk_count_reg[0] ),
    .C(\top_level.uart.clk_count_reg[3] ),
    .Y(_0446_));
 sg13g2_nand3_1 _1005_ (.B(_0317_),
    .C(_0446_),
    .A(net69),
    .Y(_0447_));
 sg13g2_nor3_2 _1006_ (.A(_0321_),
    .B(_0445_),
    .C(_0447_),
    .Y(_0448_));
 sg13g2_inv_1 _1007_ (.Y(_0449_),
    .A(_0448_));
 sg13g2_nor2b_1 _1008_ (.A(\top_level.uart.state_reg[0] ),
    .B_N(\top_level.uart.state_reg[1] ),
    .Y(_0450_));
 sg13g2_nand2_1 _1009_ (.Y(_0451_),
    .A(net84),
    .B(_0450_));
 sg13g2_nand3_1 _1010_ (.B(_0448_),
    .C(_0450_),
    .A(net84),
    .Y(_0452_));
 sg13g2_nand2_1 _1011_ (.Y(_0453_),
    .A(net155),
    .B(_0452_));
 sg13g2_o21ai_1 _1012_ (.B1(_0453_),
    .Y(_0043_),
    .A1(_0067_),
    .A2(net85));
 sg13g2_nor2_1 _1013_ (.A(\top_level.uart.state_reg[0] ),
    .B(\top_level.uart.state_reg[1] ),
    .Y(_0454_));
 sg13g2_nand2_1 _1014_ (.Y(_0455_),
    .A(net117),
    .B(_0323_));
 sg13g2_nor2_2 _1015_ (.A(_0454_),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_nand2_1 _1016_ (.Y(_0457_),
    .A(_0449_),
    .B(_0456_));
 sg13g2_nand2_1 _1017_ (.Y(_0458_),
    .A(net78),
    .B(_0454_));
 sg13g2_a21o_1 _1018_ (.A2(_0458_),
    .A1(_0324_),
    .B1(_0321_),
    .X(_0459_));
 sg13g2_nor3_1 _1019_ (.A(net149),
    .B(_0324_),
    .C(_0366_),
    .Y(_0460_));
 sg13g2_inv_1 _1020_ (.Y(_0461_),
    .A(_0460_));
 sg13g2_nand2_1 _1021_ (.Y(_0462_),
    .A(_0321_),
    .B(_0460_));
 sg13g2_nand3_1 _1022_ (.B(_0459_),
    .C(_0462_),
    .A(_0457_),
    .Y(_0463_));
 sg13g2_nand3_1 _1023_ (.B(_0067_),
    .C(_0454_),
    .A(net84),
    .Y(_0464_));
 sg13g2_nand3_1 _1024_ (.B(_0458_),
    .C(_0464_),
    .A(_0451_),
    .Y(_0465_));
 sg13g2_xor2_1 _1025_ (.B(_0465_),
    .A(_0463_),
    .X(_0044_));
 sg13g2_nor2_1 _1026_ (.A(\top_level.uart.state_reg[1] ),
    .B(_0322_),
    .Y(_0466_));
 sg13g2_inv_1 _1027_ (.Y(_0467_),
    .A(_0466_));
 sg13g2_o21ai_1 _1028_ (.B1(_0451_),
    .Y(_0468_),
    .A1(\top_level.uart.rx_data_reg ),
    .A2(_0467_));
 sg13g2_mux2_1 _1029_ (.A0(_0468_),
    .A1(net87),
    .S(_0463_),
    .X(_0045_));
 sg13g2_o21ai_1 _1030_ (.B1(_0458_),
    .Y(_0469_),
    .A1(net78),
    .A2(_0323_));
 sg13g2_mux2_1 _1031_ (.A0(_0469_),
    .A1(net78),
    .S(_0463_),
    .X(_0046_));
 sg13g2_a22oi_1 _1032_ (.Y(_0470_),
    .B1(_0469_),
    .B2(_0320_),
    .A2(_0456_),
    .A1(_0449_));
 sg13g2_nor2b_1 _1033_ (.A(_0469_),
    .B_N(_0455_),
    .Y(_0471_));
 sg13g2_nand3_1 _1034_ (.B(_0448_),
    .C(_0466_),
    .A(\top_level.uart.rx_data_reg ),
    .Y(_0472_));
 sg13g2_nor2b_2 _1035_ (.A(_0471_),
    .B_N(_0472_),
    .Y(_0473_));
 sg13g2_nand2b_1 _1036_ (.Y(_0474_),
    .B(_0472_),
    .A_N(_0471_));
 sg13g2_nand2_1 _1037_ (.Y(_0475_),
    .A(net91),
    .B(_0474_));
 sg13g2_o21ai_1 _1038_ (.B1(_0475_),
    .Y(_0047_),
    .A1(net91),
    .A2(_0470_));
 sg13g2_a21o_2 _1039_ (.A2(_0469_),
    .A1(_0320_),
    .B1(_0456_),
    .X(_0476_));
 sg13g2_o21ai_1 _1040_ (.B1(_0476_),
    .Y(_0477_),
    .A1(net82),
    .A2(\top_level.uart.clk_count_reg[0] ));
 sg13g2_a21oi_1 _1041_ (.A1(net82),
    .A2(\top_level.uart.clk_count_reg[0] ),
    .Y(_0478_),
    .B1(_0477_));
 sg13g2_a21o_1 _1042_ (.A2(net134),
    .A1(net82),
    .B1(_0478_),
    .X(_0048_));
 sg13g2_nand2_1 _1043_ (.Y(_0479_),
    .A(net69),
    .B(net134));
 sg13g2_a21o_1 _1044_ (.A2(\top_level.uart.clk_count_reg[0] ),
    .A1(\top_level.uart.clk_count_reg[1] ),
    .B1(net69),
    .X(_0480_));
 sg13g2_nand2_1 _1045_ (.Y(_0481_),
    .A(_0437_),
    .B(_0480_));
 sg13g2_o21ai_1 _1046_ (.B1(_0479_),
    .Y(_0049_),
    .A1(_0470_),
    .A2(_0481_));
 sg13g2_xnor2_1 _1047_ (.Y(_0482_),
    .A(net80),
    .B(_0437_));
 sg13g2_a22oi_1 _1048_ (.Y(_0483_),
    .B1(_0476_),
    .B2(_0482_),
    .A2(net134),
    .A1(net80));
 sg13g2_inv_1 _1049_ (.Y(_0050_),
    .A(net81));
 sg13g2_xor2_1 _1050_ (.B(_0438_),
    .A(net79),
    .X(_0484_));
 sg13g2_a22oi_1 _1051_ (.Y(_0485_),
    .B1(_0476_),
    .B2(_0484_),
    .A2(net134),
    .A1(net79));
 sg13g2_inv_1 _1052_ (.Y(_0051_),
    .A(_0485_));
 sg13g2_a21oi_1 _1053_ (.A1(_0439_),
    .A2(_0473_),
    .Y(_0486_),
    .B1(net46));
 sg13g2_nand2b_1 _1054_ (.Y(_0487_),
    .B(_0476_),
    .A_N(_0440_));
 sg13g2_a21oi_1 _1055_ (.A1(_0473_),
    .A2(_0487_),
    .Y(_0052_),
    .B1(net47));
 sg13g2_a21oi_1 _1056_ (.A1(_0442_),
    .A2(_0476_),
    .Y(_0488_),
    .B1(net134));
 sg13g2_a21oi_1 _1057_ (.A1(_0440_),
    .A2(_0473_),
    .Y(_0489_),
    .B1(net50));
 sg13g2_nor2_1 _1058_ (.A(_0488_),
    .B(_0489_),
    .Y(_0053_));
 sg13g2_a21oi_1 _1059_ (.A1(_0441_),
    .A2(_0476_),
    .Y(_0490_),
    .B1(net66));
 sg13g2_a21oi_1 _1060_ (.A1(net66),
    .A2(_0488_),
    .Y(_0054_),
    .B1(_0490_));
 sg13g2_nand2_1 _1061_ (.Y(_0491_),
    .A(net58),
    .B(net134));
 sg13g2_o21ai_1 _1062_ (.B1(_0491_),
    .Y(_0055_),
    .A1(_0445_),
    .A2(_0470_));
 sg13g2_a21oi_1 _1063_ (.A1(_0443_),
    .A2(_0473_),
    .Y(_0492_),
    .B1(net42));
 sg13g2_and2_1 _1064_ (.A(net42),
    .B(_0443_),
    .X(_0493_));
 sg13g2_inv_1 _1065_ (.Y(_0494_),
    .A(_0493_));
 sg13g2_a21oi_1 _1066_ (.A1(_0476_),
    .A2(_0494_),
    .Y(_0495_),
    .B1(net134));
 sg13g2_nor2_1 _1067_ (.A(net43),
    .B(_0495_),
    .Y(_0056_));
 sg13g2_nand2_1 _1068_ (.Y(_0496_),
    .A(net72),
    .B(_0493_));
 sg13g2_a21oi_1 _1069_ (.A1(_0456_),
    .A2(_0496_),
    .Y(_0497_),
    .B1(net134));
 sg13g2_a21oi_1 _1070_ (.A1(_0473_),
    .A2(_0493_),
    .Y(_0498_),
    .B1(net72));
 sg13g2_nor2_1 _1071_ (.A(_0497_),
    .B(_0498_),
    .Y(_0057_));
 sg13g2_nand4_1 _1072_ (.B(net72),
    .C(_0456_),
    .A(_0066_),
    .Y(_0499_),
    .D(_0493_));
 sg13g2_o21ai_1 _1073_ (.B1(_0499_),
    .Y(_0058_),
    .A1(_0066_),
    .A2(_0497_));
 sg13g2_nand2b_1 _1074_ (.Y(_0500_),
    .B(_0466_),
    .A_N(_0448_));
 sg13g2_a21oi_1 _1075_ (.A1(\top_level.uart.state_reg[2] ),
    .A2(\top_level.uart.state_reg[0] ),
    .Y(_0501_),
    .B1(_0450_));
 sg13g2_and4_2 _1076_ (.A(_0459_),
    .B(_0472_),
    .C(_0500_),
    .D(_0501_),
    .X(_0502_));
 sg13g2_nor2_1 _1077_ (.A(net152),
    .B(_0462_),
    .Y(_0503_));
 sg13g2_mux2_1 _1078_ (.A0(net152),
    .A1(_0503_),
    .S(_0502_),
    .X(_0059_));
 sg13g2_nor4_1 _1079_ (.A(net149),
    .B(_0324_),
    .C(_0335_),
    .D(_0347_),
    .Y(_0504_));
 sg13g2_nand2_1 _1080_ (.Y(_0505_),
    .A(_0502_),
    .B(_0504_));
 sg13g2_o21ai_1 _1081_ (.B1(_0505_),
    .Y(_0060_),
    .A1(_0068_),
    .A2(_0502_));
 sg13g2_a21oi_1 _1082_ (.A1(_0347_),
    .A2(_0502_),
    .Y(_0506_),
    .B1(net151));
 sg13g2_a21oi_1 _1083_ (.A1(_0461_),
    .A2(_0502_),
    .Y(_0061_),
    .B1(_0506_));
 sg13g2_nor2_1 _1084_ (.A(net111),
    .B(_0461_),
    .Y(_0507_));
 sg13g2_mux2_1 _1085_ (.A0(net149),
    .A1(_0507_),
    .S(_0502_),
    .X(_0062_));
 sg13g2_nor2_1 _1086_ (.A(net147),
    .B(_0338_),
    .Y(_0508_));
 sg13g2_a21oi_1 _1087_ (.A1(_0328_),
    .A2(_0508_),
    .Y(_0509_),
    .B1(\top_level.freq1_reg_out[0] ));
 sg13g2_o21ai_1 _1088_ (.B1(net37),
    .Y(_0510_),
    .A1(net156),
    .A2(_0338_));
 sg13g2_a21oi_1 _1089_ (.A1(_0328_),
    .A2(_0510_),
    .Y(_0063_),
    .B1(_0509_));
 sg13g2_a21oi_1 _1090_ (.A1(_0414_),
    .A2(_0508_),
    .Y(_0511_),
    .B1(net23));
 sg13g2_a21oi_1 _1091_ (.A1(_0414_),
    .A2(_0510_),
    .Y(_0064_),
    .B1(net24));
 sg13g2_dfrbp_1 _1092_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net174),
    .D(_0013_),
    .Q_N(_0560_),
    .Q(\top_level.freq1_reg_out[1] ));
 sg13g2_dfrbp_1 _1093_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net174),
    .D(_0014_),
    .Q_N(_0559_),
    .Q(\top_level.freq1_reg_out[2] ));
 sg13g2_dfrbp_1 _1094_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net175),
    .D(_0015_),
    .Q_N(_0558_),
    .Q(\top_level.freq1_reg_out[3] ));
 sg13g2_dfrbp_1 _1095_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net174),
    .D(net55),
    .Q_N(_0557_),
    .Q(\top_level.freq1_reg_out[4] ));
 sg13g2_dfrbp_1 _1096_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net176),
    .D(_0017_),
    .Q_N(_0556_),
    .Q(\top_level.freq1_reg_out[5] ));
 sg13g2_dfrbp_1 _1097_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net168),
    .D(_0018_),
    .Q_N(_0555_),
    .Q(\top_level.freq1_reg_out[6] ));
 sg13g2_dfrbp_1 _1098_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net168),
    .D(_0019_),
    .Q_N(_0554_),
    .Q(\top_level.freq1_reg_out[7] ));
 sg13g2_dfrbp_1 _1099_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net176),
    .D(_0020_),
    .Q_N(_0553_),
    .Q(\top_level.freq1_reg_out[8] ));
 sg13g2_dfrbp_1 _1100_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net167),
    .D(_0021_),
    .Q_N(_0552_),
    .Q(\top_level.freq1_reg_out[9] ));
 sg13g2_dfrbp_1 _1101_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net167),
    .D(_0022_),
    .Q_N(_0551_),
    .Q(\top_level.freq1_reg_out[10] ));
 sg13g2_dfrbp_1 _1102_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net167),
    .D(_0023_),
    .Q_N(_0550_),
    .Q(\top_level.freq1_reg_out[11] ));
 sg13g2_dfrbp_1 _1103_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net166),
    .D(_0024_),
    .Q_N(_0549_),
    .Q(\top_level.freq1_reg_out[12] ));
 sg13g2_dfrbp_1 _1104_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net166),
    .D(_0025_),
    .Q_N(_0548_),
    .Q(\top_level.freq1_reg_out[13] ));
 sg13g2_dfrbp_1 _1105_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net166),
    .D(_0026_),
    .Q_N(_0547_),
    .Q(\top_level.freq1_reg_out[14] ));
 sg13g2_dfrbp_1 _1106_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net170),
    .D(_0027_),
    .Q_N(_0561_),
    .Q(\top_level.freq1_reg_out[15] ));
 sg13g2_dfrbp_1 _1107_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net174),
    .D(net35),
    .Q_N(_0562_),
    .Q(\top_level.adder.b[0] ));
 sg13g2_dfrbp_1 _1108_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net174),
    .D(net77),
    .Q_N(_0563_),
    .Q(\top_level.adder.b[1] ));
 sg13g2_dfrbp_1 _1109_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net175),
    .D(\top_level.adder.sum[2] ),
    .Q_N(_0564_),
    .Q(\top_level.adder.b[2] ));
 sg13g2_dfrbp_1 _1110_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net175),
    .D(\top_level.adder.sum[3] ),
    .Q_N(_0000_),
    .Q(\top_level.adder.b[3] ));
 sg13g2_dfrbp_1 _1111_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net176),
    .D(net90),
    .Q_N(_0565_),
    .Q(\top_level.adder.b[4] ));
 sg13g2_dfrbp_1 _1112_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net176),
    .D(net101),
    .Q_N(_0001_),
    .Q(\top_level.adder.b[5] ));
 sg13g2_dfrbp_1 _1113_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net168),
    .D(\top_level.adder.sum[6] ),
    .Q_N(_0566_),
    .Q(\top_level.adder.b[6] ));
 sg13g2_dfrbp_1 _1114_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net167),
    .D(net96),
    .Q_N(_0002_),
    .Q(\top_level.adder.b[7] ));
 sg13g2_dfrbp_1 _1115_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net169),
    .D(\top_level.adder.sum[8] ),
    .Q_N(_0006_),
    .Q(\top_level.adder.b[8] ));
 sg13g2_dfrbp_1 _1116_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net169),
    .D(net110),
    .Q_N(_0008_),
    .Q(\top_level.adder.b[9] ));
 sg13g2_dfrbp_1 _1117_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net169),
    .D(\top_level.adder.sum[10] ),
    .Q_N(_0009_),
    .Q(\top_level.adder.b[10] ));
 sg13g2_dfrbp_1 _1118_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net169),
    .D(net99),
    .Q_N(_0010_),
    .Q(\top_level.adder.b[11] ));
 sg13g2_dfrbp_1 _1119_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net169),
    .D(net108),
    .Q_N(_0011_),
    .Q(\top_level.adder.b[12] ));
 sg13g2_dfrbp_1 _1120_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net166),
    .D(net104),
    .Q_N(_0012_),
    .Q(\top_level.adder.b[13] ));
 sg13g2_dfrbp_1 _1121_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net166),
    .D(\top_level.adder.sum[14] ),
    .Q_N(_0567_),
    .Q(\top_level.adder.b[14] ));
 sg13g2_dfrbp_1 _1122_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net166),
    .D(\top_level.adder.sum[15] ),
    .Q_N(_0007_),
    .Q(\top_level.adder.b[15] ));
 sg13g2_dfrbp_1 _1123_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net12),
    .D(net1),
    .Q_N(_0546_),
    .Q(\top_level.uart.rx_data_reg ));
 sg13g2_dfrbp_1 _1124_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net174),
    .D(_0028_),
    .Q_N(_0545_),
    .Q(\top_level.freq0_reg_out[1] ));
 sg13g2_dfrbp_1 _1125_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net175),
    .D(_0029_),
    .Q_N(_0544_),
    .Q(\top_level.freq0_reg_out[2] ));
 sg13g2_dfrbp_1 _1126_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net175),
    .D(_0030_),
    .Q_N(_0543_),
    .Q(\top_level.freq0_reg_out[3] ));
 sg13g2_dfrbp_1 _1127_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net176),
    .D(net30),
    .Q_N(_0542_),
    .Q(\top_level.freq0_reg_out[4] ));
 sg13g2_dfrbp_1 _1128_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net176),
    .D(_0032_),
    .Q_N(_0541_),
    .Q(\top_level.freq0_reg_out[5] ));
 sg13g2_dfrbp_1 _1129_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net168),
    .D(_0033_),
    .Q_N(_0540_),
    .Q(\top_level.freq0_reg_out[6] ));
 sg13g2_dfrbp_1 _1130_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net176),
    .D(_0034_),
    .Q_N(_0539_),
    .Q(\top_level.freq0_reg_out[7] ));
 sg13g2_dfrbp_1 _1131_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net176),
    .D(_0035_),
    .Q_N(_0538_),
    .Q(\top_level.freq0_reg_out[8] ));
 sg13g2_dfrbp_1 _1132_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net167),
    .D(_0036_),
    .Q_N(_0537_),
    .Q(\top_level.freq0_reg_out[9] ));
 sg13g2_dfrbp_1 _1133_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net167),
    .D(_0037_),
    .Q_N(_0536_),
    .Q(\top_level.freq0_reg_out[10] ));
 sg13g2_dfrbp_1 _1134_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net167),
    .D(_0038_),
    .Q_N(_0535_),
    .Q(\top_level.freq0_reg_out[11] ));
 sg13g2_dfrbp_1 _1135_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net167),
    .D(_0039_),
    .Q_N(_0534_),
    .Q(\top_level.freq0_reg_out[12] ));
 sg13g2_dfrbp_1 _1136_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net166),
    .D(_0040_),
    .Q_N(_0533_),
    .Q(\top_level.freq0_reg_out[13] ));
 sg13g2_dfrbp_1 _1137_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net166),
    .D(_0041_),
    .Q_N(_0532_),
    .Q(\top_level.freq0_reg_out[14] ));
 sg13g2_dfrbp_1 _1138_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net170),
    .D(_0042_),
    .Q_N(_0531_),
    .Q(\top_level.freq0_reg_out[15] ));
 sg13g2_dfrbp_1 _1139_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net172),
    .D(net86),
    .Q_N(_0004_),
    .Q(\top_level.uart.byte_number ));
 sg13g2_dfrbp_1 _1140_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net172),
    .D(_0044_),
    .Q_N(_0530_),
    .Q(\top_level.uart.state_reg[0] ));
 sg13g2_dfrbp_1 _1141_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net172),
    .D(net88),
    .Q_N(_0529_),
    .Q(\top_level.uart.state_reg[1] ));
 sg13g2_dfrbp_1 _1142_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net172),
    .D(_0046_),
    .Q_N(_0003_),
    .Q(\top_level.uart.state_reg[2] ));
 sg13g2_dfrbp_1 _1143_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net172),
    .D(net92),
    .Q_N(_0528_),
    .Q(\top_level.uart.clk_count_reg[0] ));
 sg13g2_dfrbp_1 _1144_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net172),
    .D(net83),
    .Q_N(_0527_),
    .Q(\top_level.uart.clk_count_reg[1] ));
 sg13g2_dfrbp_1 _1145_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net172),
    .D(net70),
    .Q_N(_0526_),
    .Q(\top_level.uart.clk_count_reg[2] ));
 sg13g2_dfrbp_1 _1146_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net172),
    .D(_0050_),
    .Q_N(_0525_),
    .Q(\top_level.uart.clk_count_reg[3] ));
 sg13g2_dfrbp_1 _1147_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net171),
    .D(_0051_),
    .Q_N(_0524_),
    .Q(\top_level.uart.clk_count_reg[4] ));
 sg13g2_dfrbp_1 _1148_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net171),
    .D(_0052_),
    .Q_N(_0523_),
    .Q(\top_level.uart.clk_count_reg[5] ));
 sg13g2_dfrbp_1 _1149_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net171),
    .D(_0053_),
    .Q_N(_0522_),
    .Q(\top_level.uart.clk_count_reg[6] ));
 sg13g2_dfrbp_1 _1150_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net171),
    .D(_0054_),
    .Q_N(_0521_),
    .Q(\top_level.uart.clk_count_reg[7] ));
 sg13g2_dfrbp_1 _1151_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net171),
    .D(net59),
    .Q_N(_0520_),
    .Q(\top_level.uart.clk_count_reg[8] ));
 sg13g2_dfrbp_1 _1152_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net171),
    .D(_0056_),
    .Q_N(_0519_),
    .Q(\top_level.uart.clk_count_reg[9] ));
 sg13g2_dfrbp_1 _1153_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net171),
    .D(_0057_),
    .Q_N(_0518_),
    .Q(\top_level.uart.clk_count_reg[10] ));
 sg13g2_dfrbp_1 _1154_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net173),
    .D(net75),
    .Q_N(_0517_),
    .Q(\top_level.uart.clk_count_reg[11] ));
 sg13g2_dfrbp_1 _1155_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net173),
    .D(_0059_),
    .Q_N(_0516_),
    .Q(\top_level.uart.bit_index_reg[0] ));
 sg13g2_dfrbp_1 _1156_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net173),
    .D(net106),
    .Q_N(_0515_),
    .Q(\top_level.uart.bit_index_reg[1] ));
 sg13g2_dfrbp_1 _1157_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net173),
    .D(_0061_),
    .Q_N(_0514_),
    .Q(\top_level.uart.bit_index_reg[2] ));
 sg13g2_dfrbp_1 _1158_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net171),
    .D(net112),
    .Q_N(_0005_),
    .Q(\top_level.uart.bit_index_reg[3] ));
 sg13g2_dfrbp_1 _1159_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net174),
    .D(net38),
    .Q_N(_0513_),
    .Q(\top_level.freq1_reg_out[0] ));
 sg13g2_dfrbp_1 _1160_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net174),
    .D(net25),
    .Q_N(_0512_),
    .Q(\top_level.freq0_reg_out[0] ));
 sg13g2_tiehi tt_um_DaDDS_13 (.L_HI(net13));
 sg13g2_tiehi tt_um_DaDDS_14 (.L_HI(net14));
 sg13g2_tiehi tt_um_DaDDS_15 (.L_HI(net15));
 sg13g2_tiehi tt_um_DaDDS_16 (.L_HI(net16));
 sg13g2_tiehi tt_um_DaDDS_17 (.L_HI(net17));
 sg13g2_tiehi tt_um_DaDDS_18 (.L_HI(net18));
 sg13g2_tiehi tt_um_DaDDS_19 (.L_HI(net19));
 sg13g2_tiehi tt_um_DaDDS_20 (.L_HI(net20));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_DaDDS_5 (.L_LO(net5));
 sg13g2_tielo tt_um_DaDDS_6 (.L_LO(net6));
 sg13g2_tielo tt_um_DaDDS_7 (.L_LO(net7));
 sg13g2_tielo tt_um_DaDDS_8 (.L_LO(net8));
 sg13g2_tielo tt_um_DaDDS_9 (.L_LO(net9));
 sg13g2_tielo tt_um_DaDDS_10 (.L_LO(net10));
 sg13g2_tielo tt_um_DaDDS_11 (.L_LO(net11));
 sg13g2_tiehi _1123__12 (.L_HI(net12));
 sg13g2_buf_2 fanout134 (.A(_0474_),
    .X(net134));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(_0413_));
 sg13g2_buf_2 fanout136 (.A(_0327_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_0327_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_0326_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_0412_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_0119_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_0114_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_0097_),
    .X(net143));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(_0088_));
 sg13g2_buf_2 fanout145 (.A(_0087_),
    .X(net145));
 sg13g2_buf_1 fanout146 (.A(_0087_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_0067_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(\top_level.uart.bit_index_reg[3] ),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(\top_level.uart.bit_index_reg[3] ),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(net118),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(net102),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(net114),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(net155),
    .X(net153));
 sg13g2_buf_1 fanout154 (.A(net155),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(\top_level.uart.byte_number ),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(\top_level.uart.rx_data_reg ),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(net158),
    .X(net157));
 sg13g2_buf_1 fanout158 (.A(net160),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(net160),
    .X(net159));
 sg13g2_buf_1 fanout160 (.A(\top_level.adder.b[15] ),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(\top_level.adder.b[14] ),
    .X(net162));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(net165));
 sg13g2_buf_2 fanout164 (.A(net165),
    .X(net164));
 sg13g2_buf_4 fanout165 (.X(net165),
    .A(net3));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(net170));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(net169));
 sg13g2_buf_2 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_4 fanout169 (.X(net169),
    .A(net170));
 sg13g2_buf_2 fanout170 (.A(rst_n),
    .X(net170));
 sg13g2_buf_4 fanout171 (.X(net171),
    .A(net173));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(net173));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(net177));
 sg13g2_buf_4 fanout174 (.X(net174),
    .A(net177));
 sg13g2_buf_2 fanout175 (.A(net177),
    .X(net175));
 sg13g2_buf_4 fanout176 (.X(net176),
    .A(net177));
 sg13g2_buf_2 fanout177 (.A(rst_n),
    .X(net177));
 sg13g2_buf_1 input1 (.A(ui_in[3]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[4]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[5]),
    .X(net3));
 sg13g2_tielo tt_um_DaDDS_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\top_level.freq0_reg_out[9] ),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold2 (.A(\top_level.freq0_reg_out[11] ),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold3 (.A(\top_level.freq0_reg_out[0] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0511_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0064_),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold6 (.A(\top_level.freq0_reg_out[13] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold7 (.A(\top_level.freq0_reg_out[12] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold8 (.A(\top_level.freq0_reg_out[15] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold9 (.A(\top_level.freq0_reg_out[4] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0031_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold11 (.A(\top_level.freq0_reg_out[2] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0417_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold13 (.A(\top_level.freq0_reg_out[3] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold14 (.A(\top_level.adder.b[0] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold15 (.A(\top_level.adder.sum[0] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold16 (.A(\top_level.freq0_reg_out[6] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0004_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0063_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold19 (.A(\top_level.freq0_reg_out[10] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold20 (.A(\top_level.freq0_reg_out[14] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold21 (.A(\top_level.freq0_reg_out[1] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold22 (.A(\top_level.uart.clk_count_reg[9] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0492_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold24 (.A(\top_level.freq1_reg_out[9] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold25 (.A(\top_level.freq1_reg_out[13] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold26 (.A(\top_level.uart.clk_count_reg[5] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0486_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold28 (.A(\top_level.freq1_reg_out[11] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold29 (.A(\top_level.freq1_reg_out[15] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold30 (.A(\top_level.uart.clk_count_reg[6] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold31 (.A(\top_level.freq0_reg_out[5] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold32 (.A(\top_level.freq0_reg_out[7] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold33 (.A(\top_level.freq1_reg_out[5] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold34 (.A(\top_level.freq1_reg_out[4] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0016_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold36 (.A(\top_level.freq1_reg_out[2] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0345_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold38 (.A(\top_level.uart.clk_count_reg[8] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0055_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold40 (.A(\top_level.freq1_reg_out[10] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold41 (.A(\top_level.freq0_reg_out[8] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold42 (.A(\top_level.freq1_reg_out[1] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold43 (.A(\top_level.freq1_reg_out[14] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold44 (.A(\top_level.freq1_reg_out[7] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold45 (.A(\top_level.freq1_reg_out[12] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold46 (.A(\top_level.uart.clk_count_reg[7] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold47 (.A(\top_level.freq1_reg_out[3] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0007_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold49 (.A(\top_level.uart.clk_count_reg[2] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0049_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold51 (.A(\top_level.freq1_reg_out[6] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold52 (.A(\top_level.uart.clk_count_reg[10] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold53 (.A(\top_level.freq1_reg_out[8] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold54 (.A(\top_level.uart.clk_count_reg[11] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0058_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold56 (.A(\top_level.adder.b[1] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold57 (.A(\top_level.adder.sum[1] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold58 (.A(\top_level.uart.state_reg[2] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold59 (.A(\top_level.uart.clk_count_reg[4] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold60 (.A(\top_level.uart.clk_count_reg[3] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0483_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold62 (.A(\top_level.uart.clk_count_reg[1] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0048_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0003_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0452_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0043_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold67 (.A(\top_level.uart.state_reg[1] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0045_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0000_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold70 (.A(\top_level.adder.sum[4] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold71 (.A(\top_level.uart.clk_count_reg[0] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0047_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold73 (.A(\top_level.adder.b[2] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0006_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0002_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold76 (.A(\top_level.adder.sum[7] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold77 (.A(\top_level.adder.b[10] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0293_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold79 (.A(\top_level.adder.sum[11] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0001_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold81 (.A(\top_level.adder.sum[5] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold82 (.A(\top_level.uart.bit_index_reg[2] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold83 (.A(\top_level.adder.b[12] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold84 (.A(\top_level.adder.sum[13] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold85 (.A(\top_level.uart.bit_index_reg[1] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0060_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0011_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold88 (.A(\top_level.adder.sum[12] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold89 (.A(\top_level.adder.b[8] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold90 (.A(\top_level.adder.sum[9] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0005_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0062_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold93 (.A(\top_level.adder.b[13] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold94 (.A(\top_level.uart.bit_index_reg[0] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold95 (.A(\top_level.adder.b[6] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0009_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0003_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold98 (.A(\top_level.uart.bit_index_reg[2] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0003_),
    .X(net119));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_fill_2 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_4 FILLER_16_301 ();
 sg13g2_fill_1 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_4 FILLER_16_352 ();
 sg13g2_fill_2 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_4 FILLER_17_273 ();
 sg13g2_fill_2 FILLER_17_277 ();
 sg13g2_fill_1 FILLER_17_323 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_4 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_fill_1 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_294 ();
 sg13g2_fill_1 FILLER_19_323 ();
 sg13g2_fill_2 FILLER_19_329 ();
 sg13g2_fill_1 FILLER_19_331 ();
 sg13g2_fill_2 FILLER_19_354 ();
 sg13g2_fill_1 FILLER_19_356 ();
 sg13g2_fill_2 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_4 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_270 ();
 sg13g2_fill_2 FILLER_20_328 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_fill_2 FILLER_21_325 ();
 sg13g2_fill_2 FILLER_21_359 ();
 sg13g2_fill_1 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_4 FILLER_22_147 ();
 sg13g2_fill_1 FILLER_22_151 ();
 sg13g2_decap_8 FILLER_22_160 ();
 sg13g2_decap_8 FILLER_22_167 ();
 sg13g2_decap_8 FILLER_22_174 ();
 sg13g2_decap_8 FILLER_22_181 ();
 sg13g2_decap_8 FILLER_22_188 ();
 sg13g2_decap_8 FILLER_22_195 ();
 sg13g2_decap_8 FILLER_22_202 ();
 sg13g2_decap_8 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_216 ();
 sg13g2_decap_8 FILLER_22_223 ();
 sg13g2_decap_8 FILLER_22_230 ();
 sg13g2_decap_8 FILLER_22_237 ();
 sg13g2_decap_8 FILLER_22_244 ();
 sg13g2_decap_8 FILLER_22_251 ();
 sg13g2_decap_8 FILLER_22_258 ();
 sg13g2_decap_4 FILLER_22_265 ();
 sg13g2_fill_2 FILLER_22_269 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_4 FILLER_23_91 ();
 sg13g2_fill_1 FILLER_23_95 ();
 sg13g2_decap_8 FILLER_23_104 ();
 sg13g2_decap_8 FILLER_23_111 ();
 sg13g2_fill_2 FILLER_23_118 ();
 sg13g2_decap_8 FILLER_23_137 ();
 sg13g2_decap_4 FILLER_23_144 ();
 sg13g2_fill_1 FILLER_23_148 ();
 sg13g2_fill_1 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_fill_2 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_263 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_decap_8 FILLER_23_281 ();
 sg13g2_fill_1 FILLER_23_288 ();
 sg13g2_decap_4 FILLER_23_297 ();
 sg13g2_fill_1 FILLER_23_336 ();
 sg13g2_decap_4 FILLER_23_344 ();
 sg13g2_fill_1 FILLER_23_348 ();
 sg13g2_fill_1 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_4 FILLER_24_49 ();
 sg13g2_fill_2 FILLER_24_53 ();
 sg13g2_fill_1 FILLER_24_72 ();
 sg13g2_fill_2 FILLER_24_82 ();
 sg13g2_fill_1 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_98 ();
 sg13g2_fill_2 FILLER_24_163 ();
 sg13g2_fill_2 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_227 ();
 sg13g2_fill_1 FILLER_24_229 ();
 sg13g2_decap_8 FILLER_24_240 ();
 sg13g2_fill_1 FILLER_24_247 ();
 sg13g2_decap_4 FILLER_24_262 ();
 sg13g2_fill_2 FILLER_24_266 ();
 sg13g2_fill_2 FILLER_24_298 ();
 sg13g2_fill_1 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_306 ();
 sg13g2_decap_8 FILLER_24_313 ();
 sg13g2_decap_8 FILLER_24_320 ();
 sg13g2_decap_4 FILLER_24_335 ();
 sg13g2_fill_2 FILLER_24_339 ();
 sg13g2_fill_2 FILLER_24_353 ();
 sg13g2_fill_1 FILLER_24_355 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_4 FILLER_25_35 ();
 sg13g2_fill_1 FILLER_25_39 ();
 sg13g2_fill_1 FILLER_25_66 ();
 sg13g2_decap_8 FILLER_25_127 ();
 sg13g2_fill_2 FILLER_25_134 ();
 sg13g2_fill_1 FILLER_25_136 ();
 sg13g2_fill_2 FILLER_25_163 ();
 sg13g2_decap_8 FILLER_25_208 ();
 sg13g2_fill_2 FILLER_25_215 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_269 ();
 sg13g2_fill_1 FILLER_25_271 ();
 sg13g2_fill_2 FILLER_25_290 ();
 sg13g2_fill_1 FILLER_25_292 ();
 sg13g2_fill_1 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_92 ();
 sg13g2_fill_2 FILLER_26_99 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_fill_2 FILLER_26_107 ();
 sg13g2_decap_4 FILLER_26_143 ();
 sg13g2_decap_4 FILLER_26_160 ();
 sg13g2_fill_2 FILLER_26_194 ();
 sg13g2_fill_1 FILLER_26_196 ();
 sg13g2_decap_4 FILLER_26_241 ();
 sg13g2_fill_1 FILLER_26_245 ();
 sg13g2_decap_4 FILLER_26_265 ();
 sg13g2_fill_1 FILLER_26_269 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_fill_2 FILLER_26_339 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_35 ();
 sg13g2_fill_2 FILLER_27_88 ();
 sg13g2_fill_1 FILLER_27_90 ();
 sg13g2_fill_2 FILLER_27_96 ();
 sg13g2_fill_1 FILLER_27_116 ();
 sg13g2_fill_2 FILLER_27_126 ();
 sg13g2_fill_2 FILLER_27_150 ();
 sg13g2_decap_4 FILLER_27_188 ();
 sg13g2_fill_1 FILLER_27_256 ();
 sg13g2_decap_4 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_266 ();
 sg13g2_fill_2 FILLER_27_319 ();
 sg13g2_fill_1 FILLER_27_392 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_4 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_46 ();
 sg13g2_fill_1 FILLER_28_61 ();
 sg13g2_fill_2 FILLER_28_91 ();
 sg13g2_fill_1 FILLER_28_93 ();
 sg13g2_fill_2 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_165 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_fill_2 FILLER_28_207 ();
 sg13g2_fill_2 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_321 ();
 sg13g2_fill_1 FILLER_28_323 ();
 sg13g2_fill_2 FILLER_28_352 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_4 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_46 ();
 sg13g2_decap_4 FILLER_29_53 ();
 sg13g2_fill_1 FILLER_29_57 ();
 sg13g2_fill_2 FILLER_29_63 ();
 sg13g2_decap_4 FILLER_29_90 ();
 sg13g2_fill_2 FILLER_29_94 ();
 sg13g2_decap_8 FILLER_29_106 ();
 sg13g2_fill_2 FILLER_29_113 ();
 sg13g2_fill_1 FILLER_29_115 ();
 sg13g2_decap_4 FILLER_29_125 ();
 sg13g2_fill_2 FILLER_29_129 ();
 sg13g2_fill_2 FILLER_29_176 ();
 sg13g2_fill_2 FILLER_29_192 ();
 sg13g2_fill_1 FILLER_29_194 ();
 sg13g2_fill_1 FILLER_29_230 ();
 sg13g2_fill_1 FILLER_29_235 ();
 sg13g2_fill_2 FILLER_29_240 ();
 sg13g2_fill_2 FILLER_29_271 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_329 ();
 sg13g2_fill_1 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_14 ();
 sg13g2_decap_4 FILLER_30_23 ();
 sg13g2_fill_1 FILLER_30_27 ();
 sg13g2_fill_1 FILLER_30_36 ();
 sg13g2_fill_1 FILLER_30_53 ();
 sg13g2_fill_1 FILLER_30_60 ();
 sg13g2_decap_4 FILLER_30_66 ();
 sg13g2_fill_2 FILLER_30_74 ();
 sg13g2_decap_8 FILLER_30_94 ();
 sg13g2_fill_2 FILLER_30_101 ();
 sg13g2_decap_4 FILLER_30_117 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_fill_1 FILLER_30_149 ();
 sg13g2_fill_2 FILLER_30_190 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_fill_2 FILLER_30_221 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_fill_2 FILLER_30_249 ();
 sg13g2_fill_1 FILLER_30_279 ();
 sg13g2_decap_4 FILLER_30_293 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_fill_2 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_383 ();
 sg13g2_fill_2 FILLER_30_396 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_24 ();
 sg13g2_decap_8 FILLER_31_36 ();
 sg13g2_decap_8 FILLER_31_61 ();
 sg13g2_fill_2 FILLER_31_68 ();
 sg13g2_fill_1 FILLER_31_70 ();
 sg13g2_decap_4 FILLER_31_86 ();
 sg13g2_fill_1 FILLER_31_110 ();
 sg13g2_fill_2 FILLER_31_150 ();
 sg13g2_decap_8 FILLER_31_218 ();
 sg13g2_fill_2 FILLER_31_225 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_decap_4 FILLER_31_292 ();
 sg13g2_fill_2 FILLER_31_319 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_fill_1 FILLER_31_332 ();
 sg13g2_fill_1 FILLER_31_338 ();
 sg13g2_fill_2 FILLER_31_370 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_22 ();
 sg13g2_fill_2 FILLER_32_29 ();
 sg13g2_fill_1 FILLER_32_31 ();
 sg13g2_decap_4 FILLER_32_63 ();
 sg13g2_fill_1 FILLER_32_67 ();
 sg13g2_fill_1 FILLER_32_79 ();
 sg13g2_decap_8 FILLER_32_85 ();
 sg13g2_fill_2 FILLER_32_92 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_decap_8 FILLER_32_107 ();
 sg13g2_fill_1 FILLER_32_114 ();
 sg13g2_fill_2 FILLER_32_119 ();
 sg13g2_fill_2 FILLER_32_130 ();
 sg13g2_fill_1 FILLER_32_132 ();
 sg13g2_fill_2 FILLER_32_148 ();
 sg13g2_fill_2 FILLER_32_186 ();
 sg13g2_decap_8 FILLER_32_204 ();
 sg13g2_decap_4 FILLER_32_211 ();
 sg13g2_decap_4 FILLER_32_224 ();
 sg13g2_fill_1 FILLER_32_228 ();
 sg13g2_decap_8 FILLER_32_255 ();
 sg13g2_decap_8 FILLER_32_262 ();
 sg13g2_decap_8 FILLER_32_269 ();
 sg13g2_decap_4 FILLER_32_276 ();
 sg13g2_fill_1 FILLER_32_280 ();
 sg13g2_fill_2 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_319 ();
 sg13g2_fill_2 FILLER_32_358 ();
 sg13g2_fill_1 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_14 ();
 sg13g2_decap_4 FILLER_33_19 ();
 sg13g2_fill_2 FILLER_33_23 ();
 sg13g2_fill_2 FILLER_33_39 ();
 sg13g2_fill_1 FILLER_33_41 ();
 sg13g2_fill_2 FILLER_33_47 ();
 sg13g2_decap_4 FILLER_33_62 ();
 sg13g2_fill_1 FILLER_33_66 ();
 sg13g2_fill_1 FILLER_33_77 ();
 sg13g2_fill_2 FILLER_33_83 ();
 sg13g2_fill_2 FILLER_33_101 ();
 sg13g2_fill_1 FILLER_33_128 ();
 sg13g2_fill_2 FILLER_33_133 ();
 sg13g2_fill_1 FILLER_33_143 ();
 sg13g2_fill_1 FILLER_33_157 ();
 sg13g2_decap_4 FILLER_33_174 ();
 sg13g2_fill_2 FILLER_33_208 ();
 sg13g2_fill_1 FILLER_33_210 ();
 sg13g2_fill_2 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_370 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_23 ();
 sg13g2_decap_4 FILLER_34_29 ();
 sg13g2_decap_4 FILLER_34_58 ();
 sg13g2_fill_2 FILLER_34_67 ();
 sg13g2_fill_2 FILLER_34_92 ();
 sg13g2_fill_1 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_103 ();
 sg13g2_fill_2 FILLER_34_110 ();
 sg13g2_fill_2 FILLER_34_133 ();
 sg13g2_fill_2 FILLER_34_195 ();
 sg13g2_fill_1 FILLER_34_197 ();
 sg13g2_decap_4 FILLER_34_271 ();
 sg13g2_fill_2 FILLER_34_284 ();
 sg13g2_fill_1 FILLER_34_286 ();
 sg13g2_fill_2 FILLER_34_327 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_decap_4 FILLER_34_373 ();
 sg13g2_fill_2 FILLER_34_377 ();
 sg13g2_fill_1 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_fill_2 FILLER_35_20 ();
 sg13g2_fill_1 FILLER_35_22 ();
 sg13g2_fill_2 FILLER_35_38 ();
 sg13g2_decap_4 FILLER_35_55 ();
 sg13g2_fill_2 FILLER_35_59 ();
 sg13g2_decap_8 FILLER_35_71 ();
 sg13g2_fill_1 FILLER_35_78 ();
 sg13g2_fill_1 FILLER_35_90 ();
 sg13g2_fill_2 FILLER_35_102 ();
 sg13g2_fill_2 FILLER_35_136 ();
 sg13g2_decap_8 FILLER_35_174 ();
 sg13g2_decap_4 FILLER_35_181 ();
 sg13g2_fill_1 FILLER_35_185 ();
 sg13g2_decap_4 FILLER_35_206 ();
 sg13g2_fill_2 FILLER_35_222 ();
 sg13g2_fill_2 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_305 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_fill_1 FILLER_35_313 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_11 ();
 sg13g2_fill_1 FILLER_36_29 ();
 sg13g2_fill_2 FILLER_36_35 ();
 sg13g2_fill_1 FILLER_36_53 ();
 sg13g2_fill_1 FILLER_36_64 ();
 sg13g2_fill_1 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_79 ();
 sg13g2_fill_1 FILLER_36_81 ();
 sg13g2_fill_1 FILLER_36_94 ();
 sg13g2_decap_4 FILLER_36_110 ();
 sg13g2_fill_1 FILLER_36_124 ();
 sg13g2_decap_8 FILLER_36_141 ();
 sg13g2_fill_2 FILLER_36_153 ();
 sg13g2_fill_1 FILLER_36_155 ();
 sg13g2_decap_4 FILLER_36_188 ();
 sg13g2_decap_4 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_308 ();
 sg13g2_fill_2 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_316 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_39 ();
 sg13g2_fill_1 FILLER_37_52 ();
 sg13g2_fill_1 FILLER_37_80 ();
 sg13g2_fill_2 FILLER_37_92 ();
 sg13g2_decap_8 FILLER_37_106 ();
 sg13g2_fill_2 FILLER_37_113 ();
 sg13g2_fill_2 FILLER_37_125 ();
 sg13g2_decap_8 FILLER_37_136 ();
 sg13g2_fill_2 FILLER_37_143 ();
 sg13g2_fill_2 FILLER_37_152 ();
 sg13g2_fill_2 FILLER_37_167 ();
 sg13g2_fill_2 FILLER_37_178 ();
 sg13g2_decap_4 FILLER_37_189 ();
 sg13g2_fill_1 FILLER_37_193 ();
 sg13g2_decap_8 FILLER_37_204 ();
 sg13g2_decap_4 FILLER_37_211 ();
 sg13g2_fill_1 FILLER_37_284 ();
 sg13g2_fill_1 FILLER_37_347 ();
 sg13g2_fill_2 FILLER_37_357 ();
 sg13g2_fill_2 FILLER_37_372 ();
 sg13g2_fill_1 FILLER_37_374 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_4 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_25 ();
 sg13g2_decap_8 FILLER_38_31 ();
 sg13g2_fill_2 FILLER_38_38 ();
 sg13g2_fill_2 FILLER_38_48 ();
 sg13g2_fill_2 FILLER_38_54 ();
 sg13g2_fill_1 FILLER_38_60 ();
 sg13g2_fill_2 FILLER_38_94 ();
 sg13g2_fill_1 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_135 ();
 sg13g2_fill_2 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_167 ();
 sg13g2_decap_4 FILLER_38_221 ();
 sg13g2_fill_1 FILLER_38_225 ();
 sg13g2_decap_8 FILLER_38_240 ();
 sg13g2_fill_2 FILLER_38_282 ();
 sg13g2_fill_1 FILLER_38_284 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_fill_1 FILLER_38_369 ();
 sg13g2_fill_1 FILLER_38_382 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net13;
 assign uio_oe[1] = net14;
 assign uio_oe[2] = net15;
 assign uio_oe[3] = net16;
 assign uio_oe[4] = net17;
 assign uio_oe[5] = net18;
 assign uio_oe[6] = net19;
 assign uio_oe[7] = net20;
 assign uio_out[0] = net4;
 assign uio_out[1] = net5;
 assign uio_out[2] = net6;
 assign uio_out[3] = net7;
 assign uio_out[4] = net8;
 assign uio_out[5] = net9;
 assign uio_out[6] = net10;
 assign uio_out[7] = net11;
endmodule

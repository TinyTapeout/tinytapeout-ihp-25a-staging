module tt_um_samuelm_pwm_generator (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire \pwm_generator_inst.counter[0] ;
 wire \pwm_generator_inst.counter[10] ;
 wire \pwm_generator_inst.counter[11] ;
 wire \pwm_generator_inst.counter[12] ;
 wire \pwm_generator_inst.counter[1] ;
 wire \pwm_generator_inst.counter[2] ;
 wire \pwm_generator_inst.counter[3] ;
 wire \pwm_generator_inst.counter[4] ;
 wire \pwm_generator_inst.counter[5] ;
 wire \pwm_generator_inst.counter[6] ;
 wire \pwm_generator_inst.counter[7] ;
 wire \pwm_generator_inst.counter[8] ;
 wire \pwm_generator_inst.counter[9] ;
 wire \pwm_generator_inst.duty_reg[0] ;
 wire \pwm_generator_inst.duty_reg[1] ;
 wire \pwm_generator_inst.duty_reg[2] ;
 wire \pwm_generator_inst.duty_reg[3] ;
 wire \pwm_generator_inst.duty_reg[4] ;
 wire \pwm_generator_inst.duty_reg[5] ;
 wire \pwm_generator_inst.duty_reg[6] ;
 wire \pwm_generator_inst.period_reg[0] ;
 wire \pwm_generator_inst.period_reg[10] ;
 wire \pwm_generator_inst.period_reg[11] ;
 wire \pwm_generator_inst.period_reg[1] ;
 wire \pwm_generator_inst.period_reg[2] ;
 wire \pwm_generator_inst.period_reg[3] ;
 wire \pwm_generator_inst.period_reg[4] ;
 wire \pwm_generator_inst.period_reg[5] ;
 wire \pwm_generator_inst.period_reg[6] ;
 wire \pwm_generator_inst.period_reg[7] ;
 wire \pwm_generator_inst.period_reg[8] ;
 wire \pwm_generator_inst.period_reg[9] ;
 wire \pwm_generator_inst.pwm_out ;
 wire \pwm_generator_inst.pwm_out_s ;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;

 sg13g2_inv_1 _0929_ (.Y(_0865_),
    .A(net12));
 sg13g2_inv_1 _0930_ (.Y(_0870_),
    .A(net11));
 sg13g2_inv_1 _0931_ (.Y(_0871_),
    .A(net10));
 sg13g2_inv_1 _0932_ (.Y(_0872_),
    .A(net9));
 sg13g2_inv_1 _0933_ (.Y(_0873_),
    .A(net8));
 sg13g2_inv_1 _0934_ (.Y(_0044_),
    .A(net7));
 sg13g2_inv_1 _0935_ (.Y(_0045_),
    .A(net6));
 sg13g2_inv_1 _0936_ (.Y(_0046_),
    .A(net5));
 sg13g2_inv_1 _0937_ (.Y(_0047_),
    .A(net4));
 sg13g2_inv_1 _0938_ (.Y(_0048_),
    .A(net3));
 sg13g2_inv_1 _0939_ (.Y(_0049_),
    .A(net2));
 sg13g2_inv_1 _0940_ (.Y(_0050_),
    .A(net1));
 sg13g2_inv_1 _0941_ (.Y(_0051_),
    .A(net204));
 sg13g2_inv_1 _0942_ (.Y(_0052_),
    .A(_0008_));
 sg13g2_inv_1 _0943_ (.Y(_0053_),
    .A(_0002_));
 sg13g2_nand2_1 _0944_ (.Y(_0054_),
    .A(net200),
    .B(net223));
 sg13g2_nand4_1 _0945_ (.B(net203),
    .C(net223),
    .A(net201),
    .Y(_0055_),
    .D(net225));
 sg13g2_nand2_1 _0946_ (.Y(_0056_),
    .A(net198),
    .B(net225));
 sg13g2_nand2_1 _0947_ (.Y(_0057_),
    .A(\pwm_generator_inst.period_reg[0] ),
    .B(net219));
 sg13g2_nor2_1 _0948_ (.A(_0054_),
    .B(_0057_),
    .Y(_0058_));
 sg13g2_xor2_1 _0949_ (.B(_0057_),
    .A(_0054_),
    .X(_0059_));
 sg13g2_nor2b_1 _0950_ (.A(_0056_),
    .B_N(_0059_),
    .Y(_0060_));
 sg13g2_xnor2_1 _0951_ (.Y(_0061_),
    .A(_0056_),
    .B(_0059_));
 sg13g2_nand2b_1 _0952_ (.Y(_0062_),
    .B(_0061_),
    .A_N(_0055_));
 sg13g2_nand2_1 _0953_ (.Y(_0063_),
    .A(net196),
    .B(net225));
 sg13g2_nand2_1 _0954_ (.Y(_0064_),
    .A(net198),
    .B(net223));
 sg13g2_and4_1 _0955_ (.A(net201),
    .B(net203),
    .C(\pwm_generator_inst.duty_reg[3] ),
    .D(net219),
    .X(_0065_));
 sg13g2_nand4_1 _0956_ (.B(net203),
    .C(net215),
    .A(net201),
    .Y(_0066_),
    .D(net219));
 sg13g2_a22oi_1 _0957_ (.Y(_0067_),
    .B1(net219),
    .B2(net201),
    .A2(net214),
    .A1(net203));
 sg13g2_nor2_1 _0958_ (.A(_0065_),
    .B(_0067_),
    .Y(_0068_));
 sg13g2_xnor2_1 _0959_ (.Y(_0069_),
    .A(_0064_),
    .B(_0068_));
 sg13g2_nand2_1 _0960_ (.Y(_0070_),
    .A(_0058_),
    .B(_0069_));
 sg13g2_nor2_1 _0961_ (.A(_0058_),
    .B(_0069_),
    .Y(_0071_));
 sg13g2_xor2_1 _0962_ (.B(_0069_),
    .A(_0058_),
    .X(_0072_));
 sg13g2_xnor2_1 _0963_ (.Y(_0073_),
    .A(_0063_),
    .B(_0072_));
 sg13g2_nand2_1 _0964_ (.Y(_0074_),
    .A(_0060_),
    .B(_0073_));
 sg13g2_xnor2_1 _0965_ (.Y(_0075_),
    .A(_0060_),
    .B(_0073_));
 sg13g2_nor2_1 _0966_ (.A(_0062_),
    .B(_0075_),
    .Y(_0076_));
 sg13g2_o21ai_1 _0967_ (.B1(_0070_),
    .Y(_0077_),
    .A1(_0063_),
    .A2(_0071_));
 sg13g2_nand2_1 _0968_ (.Y(_0078_),
    .A(net203),
    .B(net210));
 sg13g2_nand2_1 _0969_ (.Y(_0079_),
    .A(net195),
    .B(net225));
 sg13g2_nand2_1 _0970_ (.Y(_0080_),
    .A(net194),
    .B(net210));
 sg13g2_or2_1 _0971_ (.X(_0081_),
    .B(_0079_),
    .A(_0078_));
 sg13g2_xor2_1 _0972_ (.B(_0079_),
    .A(_0078_),
    .X(_0082_));
 sg13g2_inv_1 _0973_ (.Y(_0083_),
    .A(_0082_));
 sg13g2_o21ai_1 _0974_ (.B1(_0066_),
    .Y(_0084_),
    .A1(_0064_),
    .A2(_0067_));
 sg13g2_nand2_1 _0975_ (.Y(_0085_),
    .A(net197),
    .B(net223));
 sg13g2_and4_1 _0976_ (.A(net199),
    .B(\pwm_generator_inst.period_reg[1] ),
    .C(net214),
    .D(net220),
    .X(_0086_));
 sg13g2_nand4_1 _0977_ (.B(net201),
    .C(net214),
    .A(net199),
    .Y(_0087_),
    .D(net220));
 sg13g2_a22oi_1 _0978_ (.Y(_0088_),
    .B1(net219),
    .B2(net198),
    .A2(net214),
    .A1(net201));
 sg13g2_or3_1 _0979_ (.A(_0085_),
    .B(_0086_),
    .C(_0088_),
    .X(_0089_));
 sg13g2_o21ai_1 _0980_ (.B1(_0085_),
    .Y(_0090_),
    .A1(_0086_),
    .A2(_0088_));
 sg13g2_and3_1 _0981_ (.X(_0091_),
    .A(_0084_),
    .B(_0089_),
    .C(_0090_));
 sg13g2_nand3_1 _0982_ (.B(_0089_),
    .C(_0090_),
    .A(_0084_),
    .Y(_0092_));
 sg13g2_a21oi_1 _0983_ (.A1(_0089_),
    .A2(_0090_),
    .Y(_0093_),
    .B1(_0084_));
 sg13g2_nor2_1 _0984_ (.A(_0091_),
    .B(_0093_),
    .Y(_0094_));
 sg13g2_xnor2_1 _0985_ (.Y(_0095_),
    .A(_0082_),
    .B(_0094_));
 sg13g2_nand2b_1 _0986_ (.Y(_0096_),
    .B(_0077_),
    .A_N(_0095_));
 sg13g2_nor2b_1 _0987_ (.A(_0077_),
    .B_N(_0095_),
    .Y(_0097_));
 sg13g2_xnor2_1 _0988_ (.Y(_0098_),
    .A(_0077_),
    .B(_0095_));
 sg13g2_xor2_1 _0989_ (.B(_0098_),
    .A(_0074_),
    .X(_0099_));
 sg13g2_nand2_2 _0990_ (.Y(_0100_),
    .A(_0076_),
    .B(_0098_));
 sg13g2_o21ai_1 _0991_ (.B1(_0092_),
    .Y(_0101_),
    .A1(_0083_),
    .A2(_0093_));
 sg13g2_o21ai_1 _0992_ (.B1(_0087_),
    .Y(_0102_),
    .A1(_0085_),
    .A2(_0088_));
 sg13g2_nand2_1 _0993_ (.Y(_0103_),
    .A(net195),
    .B(net223));
 sg13g2_and4_1 _0994_ (.A(net197),
    .B(net198),
    .C(net214),
    .D(net219),
    .X(_0104_));
 sg13g2_nand4_1 _0995_ (.B(net198),
    .C(net214),
    .A(net196),
    .Y(_0105_),
    .D(net219));
 sg13g2_a22oi_1 _0996_ (.Y(_0106_),
    .B1(net219),
    .B2(net196),
    .A2(net214),
    .A1(net198));
 sg13g2_or3_1 _0997_ (.A(_0103_),
    .B(_0104_),
    .C(_0106_),
    .X(_0107_));
 sg13g2_o21ai_1 _0998_ (.B1(_0103_),
    .Y(_0108_),
    .A1(_0104_),
    .A2(_0106_));
 sg13g2_and3_1 _0999_ (.X(_0109_),
    .A(_0102_),
    .B(_0107_),
    .C(_0108_));
 sg13g2_nand3_1 _1000_ (.B(_0107_),
    .C(_0108_),
    .A(_0102_),
    .Y(_0110_));
 sg13g2_a21o_1 _1001_ (.A2(_0108_),
    .A1(_0107_),
    .B1(_0102_),
    .X(_0111_));
 sg13g2_nand2_1 _1002_ (.Y(_0112_),
    .A(net203),
    .B(\pwm_generator_inst.duty_reg[5] ));
 sg13g2_nand2_2 _1003_ (.Y(_0113_),
    .A(net192),
    .B(net224));
 sg13g2_nand2_1 _1004_ (.Y(_0114_),
    .A(net200),
    .B(net210));
 sg13g2_nor2_1 _1005_ (.A(_0113_),
    .B(_0114_),
    .Y(_0115_));
 sg13g2_xor2_1 _1006_ (.B(_0114_),
    .A(_0113_),
    .X(_0116_));
 sg13g2_nor2b_1 _1007_ (.A(_0112_),
    .B_N(_0116_),
    .Y(_0117_));
 sg13g2_xnor2_1 _1008_ (.Y(_0118_),
    .A(_0112_),
    .B(_0116_));
 sg13g2_nand3_1 _1009_ (.B(_0111_),
    .C(_0118_),
    .A(_0110_),
    .Y(_0119_));
 sg13g2_a21o_1 _1010_ (.A2(_0111_),
    .A1(_0110_),
    .B1(_0118_),
    .X(_0120_));
 sg13g2_and3_1 _1011_ (.X(_0121_),
    .A(_0101_),
    .B(_0119_),
    .C(_0120_));
 sg13g2_nand3_1 _1012_ (.B(_0119_),
    .C(_0120_),
    .A(_0101_),
    .Y(_0122_));
 sg13g2_a21oi_1 _1013_ (.A1(_0119_),
    .A2(_0120_),
    .Y(_0123_),
    .B1(_0101_));
 sg13g2_nor2_1 _1014_ (.A(_0121_),
    .B(_0123_),
    .Y(_0124_));
 sg13g2_xnor2_1 _1015_ (.Y(_0125_),
    .A(_0081_),
    .B(_0124_));
 sg13g2_o21ai_1 _1016_ (.B1(_0096_),
    .Y(_0126_),
    .A1(_0074_),
    .A2(_0097_));
 sg13g2_xnor2_1 _1017_ (.Y(_0127_),
    .A(_0125_),
    .B(_0126_));
 sg13g2_xnor2_1 _1018_ (.Y(_0128_),
    .A(_0100_),
    .B(_0127_));
 sg13g2_a21o_1 _1019_ (.A2(_0118_),
    .A1(_0111_),
    .B1(_0109_),
    .X(_0129_));
 sg13g2_o21ai_1 _1020_ (.B1(_0105_),
    .Y(_0130_),
    .A1(_0103_),
    .A2(_0106_));
 sg13g2_nand2_1 _1021_ (.Y(_0131_),
    .A(net193),
    .B(net222));
 sg13g2_and4_1 _1022_ (.A(net194),
    .B(net196),
    .C(net215),
    .D(net221),
    .X(_0132_));
 sg13g2_nand4_1 _1023_ (.B(net197),
    .C(net215),
    .A(net195),
    .Y(_0133_),
    .D(net221));
 sg13g2_a22oi_1 _1024_ (.Y(_0134_),
    .B1(net221),
    .B2(net195),
    .A2(net215),
    .A1(net196));
 sg13g2_or3_1 _1025_ (.A(_0131_),
    .B(_0132_),
    .C(_0134_),
    .X(_0135_));
 sg13g2_o21ai_1 _1026_ (.B1(_0131_),
    .Y(_0136_),
    .A1(_0132_),
    .A2(_0134_));
 sg13g2_and3_1 _1027_ (.X(_0137_),
    .A(_0130_),
    .B(_0135_),
    .C(_0136_));
 sg13g2_nand3_1 _1028_ (.B(_0135_),
    .C(_0136_),
    .A(_0130_),
    .Y(_0138_));
 sg13g2_a21oi_1 _1029_ (.A1(_0135_),
    .A2(_0136_),
    .Y(_0139_),
    .B1(_0130_));
 sg13g2_nand2_1 _1030_ (.Y(_0140_),
    .A(net200),
    .B(net208));
 sg13g2_nand2_1 _1031_ (.Y(_0141_),
    .A(net190),
    .B(net209));
 sg13g2_nand2_2 _1032_ (.Y(_0142_),
    .A(net190),
    .B(net224));
 sg13g2_nand2_1 _1033_ (.Y(_0143_),
    .A(net199),
    .B(net210));
 sg13g2_or2_1 _1034_ (.X(_0144_),
    .B(_0143_),
    .A(_0142_));
 sg13g2_xnor2_1 _1035_ (.Y(_0145_),
    .A(_0142_),
    .B(_0143_));
 sg13g2_xnor2_1 _1036_ (.Y(_0146_),
    .A(_0140_),
    .B(_0145_));
 sg13g2_or3_1 _1037_ (.A(_0137_),
    .B(_0139_),
    .C(_0146_),
    .X(_0147_));
 sg13g2_o21ai_1 _1038_ (.B1(_0146_),
    .Y(_0148_),
    .A1(_0137_),
    .A2(_0139_));
 sg13g2_and3_1 _1039_ (.X(_0149_),
    .A(_0129_),
    .B(_0147_),
    .C(_0148_));
 sg13g2_nand3_1 _1040_ (.B(_0147_),
    .C(_0148_),
    .A(_0129_),
    .Y(_0150_));
 sg13g2_nor2_1 _1041_ (.A(_0115_),
    .B(_0117_),
    .Y(_0151_));
 sg13g2_a21oi_1 _1042_ (.A1(_0147_),
    .A2(_0148_),
    .Y(_0152_),
    .B1(_0129_));
 sg13g2_or3_1 _1043_ (.A(_0149_),
    .B(_0151_),
    .C(_0152_),
    .X(_0153_));
 sg13g2_o21ai_1 _1044_ (.B1(_0150_),
    .Y(_0154_),
    .A1(_0151_),
    .A2(_0152_));
 sg13g2_o21ai_1 _1045_ (.B1(_0144_),
    .Y(_0155_),
    .A1(_0140_),
    .A2(_0145_));
 sg13g2_inv_1 _1046_ (.Y(_0156_),
    .A(_0155_));
 sg13g2_o21ai_1 _1047_ (.B1(_0138_),
    .Y(_0157_),
    .A1(_0139_),
    .A2(_0146_));
 sg13g2_o21ai_1 _1048_ (.B1(_0133_),
    .Y(_0158_),
    .A1(_0131_),
    .A2(_0134_));
 sg13g2_nand2_1 _1049_ (.Y(_0159_),
    .A(net191),
    .B(net223));
 sg13g2_and4_1 _1050_ (.A(net193),
    .B(net194),
    .C(net215),
    .D(net221),
    .X(_0160_));
 sg13g2_nand4_1 _1051_ (.B(net194),
    .C(net215),
    .A(net193),
    .Y(_0161_),
    .D(net221));
 sg13g2_a22oi_1 _1052_ (.Y(_0162_),
    .B1(net221),
    .B2(net193),
    .A2(net215),
    .A1(net194));
 sg13g2_or3_1 _1053_ (.A(_0159_),
    .B(_0160_),
    .C(_0162_),
    .X(_0163_));
 sg13g2_o21ai_1 _1054_ (.B1(_0159_),
    .Y(_0164_),
    .A1(_0160_),
    .A2(_0162_));
 sg13g2_and3_1 _1055_ (.X(_0165_),
    .A(_0158_),
    .B(_0163_),
    .C(_0164_));
 sg13g2_nand3_1 _1056_ (.B(_0163_),
    .C(_0164_),
    .A(_0158_),
    .Y(_0166_));
 sg13g2_a21oi_1 _1057_ (.A1(_0163_),
    .A2(_0164_),
    .Y(_0167_),
    .B1(_0158_));
 sg13g2_nand2_1 _1058_ (.Y(_0168_),
    .A(net199),
    .B(net208));
 sg13g2_nand2_1 _1059_ (.Y(_0169_),
    .A(net188),
    .B(net209));
 sg13g2_nand2_1 _1060_ (.Y(_0170_),
    .A(net189),
    .B(net224));
 sg13g2_nand2_1 _1061_ (.Y(_0171_),
    .A(net197),
    .B(net210));
 sg13g2_xor2_1 _1062_ (.B(_0171_),
    .A(_0170_),
    .X(_0172_));
 sg13g2_nand2b_1 _1063_ (.Y(_0173_),
    .B(_0172_),
    .A_N(_0168_));
 sg13g2_xor2_1 _1064_ (.B(_0172_),
    .A(_0168_),
    .X(_0174_));
 sg13g2_or3_1 _1065_ (.A(_0165_),
    .B(_0167_),
    .C(_0174_),
    .X(_0175_));
 sg13g2_o21ai_1 _1066_ (.B1(_0174_),
    .Y(_0176_),
    .A1(_0165_),
    .A2(_0167_));
 sg13g2_nand3_1 _1067_ (.B(_0175_),
    .C(_0176_),
    .A(_0157_),
    .Y(_0177_));
 sg13g2_a21oi_1 _1068_ (.A1(_0175_),
    .A2(_0176_),
    .Y(_0178_),
    .B1(_0157_));
 sg13g2_a21o_1 _1069_ (.A2(_0176_),
    .A1(_0175_),
    .B1(_0157_),
    .X(_0179_));
 sg13g2_nand3_1 _1070_ (.B(_0177_),
    .C(_0179_),
    .A(_0155_),
    .Y(_0180_));
 sg13g2_a21o_1 _1071_ (.A2(_0179_),
    .A1(_0177_),
    .B1(_0155_),
    .X(_0181_));
 sg13g2_nand3_1 _1072_ (.B(_0180_),
    .C(_0181_),
    .A(_0154_),
    .Y(_0182_));
 sg13g2_and2_1 _1073_ (.A(net200),
    .B(net206),
    .X(_0183_));
 sg13g2_nand2_1 _1074_ (.Y(_0184_),
    .A(net200),
    .B(net205));
 sg13g2_a21oi_1 _1075_ (.A1(_0180_),
    .A2(_0181_),
    .Y(_0185_),
    .B1(_0154_));
 sg13g2_a21o_1 _1076_ (.A2(_0181_),
    .A1(_0180_),
    .B1(_0154_),
    .X(_0186_));
 sg13g2_and3_1 _1077_ (.X(_0187_),
    .A(_0182_),
    .B(_0183_),
    .C(_0186_));
 sg13g2_o21ai_1 _1078_ (.B1(_0182_),
    .Y(_0188_),
    .A1(_0184_),
    .A2(_0185_));
 sg13g2_nand2_1 _1079_ (.Y(_0189_),
    .A(net199),
    .B(net205));
 sg13g2_o21ai_1 _1080_ (.B1(_0177_),
    .Y(_0190_),
    .A1(_0156_),
    .A2(_0178_));
 sg13g2_o21ai_1 _1081_ (.B1(_0173_),
    .Y(_0191_),
    .A1(_0170_),
    .A2(_0171_));
 sg13g2_inv_1 _1082_ (.Y(_0192_),
    .A(_0191_));
 sg13g2_o21ai_1 _1083_ (.B1(_0166_),
    .Y(_0193_),
    .A1(_0167_),
    .A2(_0174_));
 sg13g2_o21ai_1 _1084_ (.B1(_0161_),
    .Y(_0194_),
    .A1(_0159_),
    .A2(_0162_));
 sg13g2_nand2_1 _1085_ (.Y(_0195_),
    .A(net189),
    .B(net222));
 sg13g2_and4_1 _1086_ (.A(net190),
    .B(net192),
    .C(net213),
    .D(net218),
    .X(_0196_));
 sg13g2_nand4_1 _1087_ (.B(net192),
    .C(net213),
    .A(net191),
    .Y(_0197_),
    .D(net218));
 sg13g2_a22oi_1 _1088_ (.Y(_0198_),
    .B1(net218),
    .B2(net191),
    .A2(net213),
    .A1(net192));
 sg13g2_or3_1 _1089_ (.A(_0195_),
    .B(_0196_),
    .C(_0198_),
    .X(_0199_));
 sg13g2_o21ai_1 _1090_ (.B1(_0195_),
    .Y(_0200_),
    .A1(_0196_),
    .A2(_0198_));
 sg13g2_and3_1 _1091_ (.X(_0201_),
    .A(_0194_),
    .B(_0199_),
    .C(_0200_));
 sg13g2_nand3_1 _1092_ (.B(_0199_),
    .C(_0200_),
    .A(_0194_),
    .Y(_0202_));
 sg13g2_a21oi_1 _1093_ (.A1(_0199_),
    .A2(_0200_),
    .Y(_0203_),
    .B1(_0194_));
 sg13g2_nand2_1 _1094_ (.Y(_0204_),
    .A(net197),
    .B(net208));
 sg13g2_nand2_1 _1095_ (.Y(_0205_),
    .A(\pwm_generator_inst.period_reg[8] ),
    .B(net224));
 sg13g2_or2_1 _1096_ (.X(_0206_),
    .B(_0205_),
    .A(_0080_));
 sg13g2_xnor2_1 _1097_ (.Y(_0207_),
    .A(_0080_),
    .B(_0205_));
 sg13g2_xnor2_1 _1098_ (.Y(_0208_),
    .A(_0204_),
    .B(_0207_));
 sg13g2_or3_1 _1099_ (.A(_0201_),
    .B(_0203_),
    .C(_0208_),
    .X(_0209_));
 sg13g2_o21ai_1 _1100_ (.B1(_0208_),
    .Y(_0210_),
    .A1(_0201_),
    .A2(_0203_));
 sg13g2_nand3_1 _1101_ (.B(_0209_),
    .C(_0210_),
    .A(_0193_),
    .Y(_0211_));
 sg13g2_a21oi_1 _1102_ (.A1(_0209_),
    .A2(_0210_),
    .Y(_0212_),
    .B1(_0193_));
 sg13g2_a21o_1 _1103_ (.A2(_0210_),
    .A1(_0209_),
    .B1(_0193_),
    .X(_0213_));
 sg13g2_nand3_1 _1104_ (.B(_0211_),
    .C(_0213_),
    .A(_0191_),
    .Y(_0214_));
 sg13g2_a21o_1 _1105_ (.A2(_0213_),
    .A1(_0211_),
    .B1(_0191_),
    .X(_0215_));
 sg13g2_and3_1 _1106_ (.X(_0216_),
    .A(_0190_),
    .B(_0214_),
    .C(_0215_));
 sg13g2_nand3_1 _1107_ (.B(_0214_),
    .C(_0215_),
    .A(_0190_),
    .Y(_0217_));
 sg13g2_a21oi_1 _1108_ (.A1(_0214_),
    .A2(_0215_),
    .Y(_0218_),
    .B1(_0190_));
 sg13g2_or3_1 _1109_ (.A(_0189_),
    .B(_0216_),
    .C(_0218_),
    .X(_0219_));
 sg13g2_o21ai_1 _1110_ (.B1(_0189_),
    .Y(_0220_),
    .A1(_0216_),
    .A2(_0218_));
 sg13g2_nand3_1 _1111_ (.B(_0219_),
    .C(_0220_),
    .A(_0188_),
    .Y(_0221_));
 sg13g2_a21o_1 _1112_ (.A2(_0220_),
    .A1(_0219_),
    .B1(_0188_),
    .X(_0222_));
 sg13g2_and2_1 _1113_ (.A(_0221_),
    .B(_0222_),
    .X(_0223_));
 sg13g2_o21ai_1 _1114_ (.B1(_0122_),
    .Y(_0224_),
    .A1(_0081_),
    .A2(_0123_));
 sg13g2_o21ai_1 _1115_ (.B1(_0151_),
    .Y(_0225_),
    .A1(_0149_),
    .A2(_0152_));
 sg13g2_nand3_1 _1116_ (.B(_0224_),
    .C(_0225_),
    .A(_0153_),
    .Y(_0226_));
 sg13g2_a21o_1 _1117_ (.A2(_0225_),
    .A1(_0153_),
    .B1(_0224_),
    .X(_0227_));
 sg13g2_and4_1 _1118_ (.A(net202),
    .B(net205),
    .C(_0226_),
    .D(_0227_),
    .X(_0228_));
 sg13g2_nand4_1 _1119_ (.B(net205),
    .C(_0226_),
    .A(net202),
    .Y(_0229_),
    .D(_0227_));
 sg13g2_nand2_1 _1120_ (.Y(_0230_),
    .A(_0226_),
    .B(_0229_));
 sg13g2_a21oi_1 _1121_ (.A1(_0182_),
    .A2(_0186_),
    .Y(_0231_),
    .B1(_0183_));
 sg13g2_nor2_2 _1122_ (.A(_0187_),
    .B(_0231_),
    .Y(_0232_));
 sg13g2_nor2_1 _1123_ (.A(_0230_),
    .B(_0232_),
    .Y(_0233_));
 sg13g2_nand2b_1 _1124_ (.Y(_0234_),
    .B(_0125_),
    .A_N(_0096_));
 sg13g2_a22oi_1 _1125_ (.Y(_0235_),
    .B1(_0226_),
    .B2(_0227_),
    .A2(net205),
    .A1(net202));
 sg13g2_nor3_1 _1126_ (.A(_0228_),
    .B(_0234_),
    .C(_0235_),
    .Y(_0236_));
 sg13g2_nand4_1 _1127_ (.B(_0073_),
    .C(_0098_),
    .A(_0060_),
    .Y(_0237_),
    .D(_0125_));
 sg13g2_o21ai_1 _1128_ (.B1(_0237_),
    .Y(_0238_),
    .A1(_0100_),
    .A2(_0127_));
 sg13g2_o21ai_1 _1129_ (.B1(_0234_),
    .Y(_0239_),
    .A1(_0228_),
    .A2(_0235_));
 sg13g2_nor2b_1 _1130_ (.A(_0236_),
    .B_N(_0239_),
    .Y(_0240_));
 sg13g2_a21oi_1 _1131_ (.A1(_0238_),
    .A2(_0239_),
    .Y(_0241_),
    .B1(_0236_));
 sg13g2_a221oi_1 _1132_ (.B2(_0239_),
    .C1(_0236_),
    .B1(_0238_),
    .A1(_0230_),
    .Y(_0242_),
    .A2(_0232_));
 sg13g2_xnor2_1 _1133_ (.Y(_0243_),
    .A(_0230_),
    .B(_0232_));
 sg13g2_nor2_1 _1134_ (.A(_0233_),
    .B(_0242_),
    .Y(_0244_));
 sg13g2_nand2_1 _1135_ (.Y(_0245_),
    .A(_0223_),
    .B(_0244_));
 sg13g2_xnor2_1 _1136_ (.Y(_0246_),
    .A(_0223_),
    .B(_0244_));
 sg13g2_inv_1 _1137_ (.Y(_0247_),
    .A(_0246_));
 sg13g2_o21ai_1 _1138_ (.B1(_0211_),
    .Y(_0248_),
    .A1(_0192_),
    .A2(_0212_));
 sg13g2_o21ai_1 _1139_ (.B1(_0206_),
    .Y(_0249_),
    .A1(_0204_),
    .A2(_0207_));
 sg13g2_inv_1 _1140_ (.Y(_0250_),
    .A(_0249_));
 sg13g2_o21ai_1 _1141_ (.B1(_0202_),
    .Y(_0251_),
    .A1(_0203_),
    .A2(_0208_));
 sg13g2_o21ai_1 _1142_ (.B1(_0197_),
    .Y(_0252_),
    .A1(_0195_),
    .A2(_0198_));
 sg13g2_nand2_1 _1143_ (.Y(_0253_),
    .A(net187),
    .B(net222));
 sg13g2_and4_1 _1144_ (.A(net189),
    .B(net190),
    .C(net212),
    .D(net217),
    .X(_0254_));
 sg13g2_nand4_1 _1145_ (.B(net190),
    .C(net212),
    .A(net188),
    .Y(_0255_),
    .D(net216));
 sg13g2_a22oi_1 _1146_ (.Y(_0256_),
    .B1(net216),
    .B2(net188),
    .A2(net213),
    .A1(net190));
 sg13g2_or3_1 _1147_ (.A(_0253_),
    .B(_0254_),
    .C(_0256_),
    .X(_0257_));
 sg13g2_o21ai_1 _1148_ (.B1(_0253_),
    .Y(_0258_),
    .A1(_0254_),
    .A2(_0256_));
 sg13g2_and3_1 _1149_ (.X(_0259_),
    .A(_0252_),
    .B(_0257_),
    .C(_0258_));
 sg13g2_nand3_1 _1150_ (.B(_0257_),
    .C(_0258_),
    .A(_0252_),
    .Y(_0260_));
 sg13g2_a21o_1 _1151_ (.A2(_0258_),
    .A1(_0257_),
    .B1(_0252_),
    .X(_0261_));
 sg13g2_nand2_1 _1152_ (.Y(_0262_),
    .A(net194),
    .B(net208));
 sg13g2_nand2_2 _1153_ (.Y(_0263_),
    .A(net184),
    .B(net209));
 sg13g2_nand2_1 _1154_ (.Y(_0264_),
    .A(net192),
    .B(net210));
 sg13g2_nand2_1 _1155_ (.Y(_0265_),
    .A(net185),
    .B(net224));
 sg13g2_nor2_1 _1156_ (.A(_0113_),
    .B(_0263_),
    .Y(_0266_));
 sg13g2_xor2_1 _1157_ (.B(_0265_),
    .A(_0264_),
    .X(_0267_));
 sg13g2_nand2b_1 _1158_ (.Y(_0268_),
    .B(_0267_),
    .A_N(_0262_));
 sg13g2_xnor2_1 _1159_ (.Y(_0269_),
    .A(_0262_),
    .B(_0267_));
 sg13g2_nand3_1 _1160_ (.B(_0261_),
    .C(_0269_),
    .A(_0260_),
    .Y(_0270_));
 sg13g2_a21o_1 _1161_ (.A2(_0261_),
    .A1(_0260_),
    .B1(_0269_),
    .X(_0271_));
 sg13g2_nand3_1 _1162_ (.B(_0270_),
    .C(_0271_),
    .A(_0251_),
    .Y(_0272_));
 sg13g2_a21oi_1 _1163_ (.A1(_0270_),
    .A2(_0271_),
    .Y(_0273_),
    .B1(_0251_));
 sg13g2_a21o_1 _1164_ (.A2(_0271_),
    .A1(_0270_),
    .B1(_0251_),
    .X(_0274_));
 sg13g2_nand3_1 _1165_ (.B(_0272_),
    .C(_0274_),
    .A(_0249_),
    .Y(_0275_));
 sg13g2_a21o_1 _1166_ (.A2(_0274_),
    .A1(_0272_),
    .B1(_0249_),
    .X(_0276_));
 sg13g2_and3_1 _1167_ (.X(_0277_),
    .A(_0248_),
    .B(_0275_),
    .C(_0276_));
 sg13g2_nand3_1 _1168_ (.B(_0275_),
    .C(_0276_),
    .A(_0248_),
    .Y(_0278_));
 sg13g2_nand2_1 _1169_ (.Y(_0279_),
    .A(net197),
    .B(net205));
 sg13g2_a21oi_1 _1170_ (.A1(_0275_),
    .A2(_0276_),
    .Y(_0280_),
    .B1(_0248_));
 sg13g2_or3_1 _1171_ (.A(_0277_),
    .B(_0279_),
    .C(_0280_),
    .X(_0281_));
 sg13g2_o21ai_1 _1172_ (.B1(_0278_),
    .Y(_0282_),
    .A1(_0279_),
    .A2(_0280_));
 sg13g2_nand2_1 _1173_ (.Y(_0283_),
    .A(net194),
    .B(net206));
 sg13g2_o21ai_1 _1174_ (.B1(_0272_),
    .Y(_0284_),
    .A1(_0250_),
    .A2(_0273_));
 sg13g2_nor2b_1 _1175_ (.A(_0266_),
    .B_N(_0268_),
    .Y(_0285_));
 sg13g2_nand2b_1 _1176_ (.Y(_0286_),
    .B(_0268_),
    .A_N(_0266_));
 sg13g2_a21o_1 _1177_ (.A2(_0269_),
    .A1(_0261_),
    .B1(_0259_),
    .X(_0287_));
 sg13g2_o21ai_1 _1178_ (.B1(_0255_),
    .Y(_0288_),
    .A1(_0253_),
    .A2(_0256_));
 sg13g2_nand2_1 _1179_ (.Y(_0289_),
    .A(net184),
    .B(net222));
 sg13g2_and4_1 _1180_ (.A(net187),
    .B(net189),
    .C(net212),
    .D(net217),
    .X(_0290_));
 sg13g2_nand4_1 _1181_ (.B(net188),
    .C(net211),
    .A(net187),
    .Y(_0291_),
    .D(net216));
 sg13g2_a22oi_1 _1182_ (.Y(_0292_),
    .B1(net217),
    .B2(net186),
    .A2(net212),
    .A1(net188));
 sg13g2_or3_1 _1183_ (.A(_0289_),
    .B(_0290_),
    .C(_0292_),
    .X(_0293_));
 sg13g2_o21ai_1 _1184_ (.B1(_0289_),
    .Y(_0294_),
    .A1(_0290_),
    .A2(_0292_));
 sg13g2_and3_1 _1185_ (.X(_0295_),
    .A(_0288_),
    .B(_0293_),
    .C(_0294_));
 sg13g2_nand3_1 _1186_ (.B(_0293_),
    .C(_0294_),
    .A(_0288_),
    .Y(_0296_));
 sg13g2_a21oi_1 _1187_ (.A1(_0293_),
    .A2(_0294_),
    .Y(_0297_),
    .B1(_0288_));
 sg13g2_nand2_1 _1188_ (.Y(_0298_),
    .A(net192),
    .B(net208));
 sg13g2_nand2_2 _1189_ (.Y(_0299_),
    .A(net182),
    .B(net209));
 sg13g2_nand2_1 _1190_ (.Y(_0300_),
    .A(net182),
    .B(net224));
 sg13g2_nor2_1 _1191_ (.A(_0142_),
    .B(_0299_),
    .Y(_0301_));
 sg13g2_xnor2_1 _1192_ (.Y(_0302_),
    .A(_0141_),
    .B(_0300_));
 sg13g2_nor2_1 _1193_ (.A(_0298_),
    .B(_0302_),
    .Y(_0303_));
 sg13g2_xnor2_1 _1194_ (.Y(_0304_),
    .A(_0298_),
    .B(_0302_));
 sg13g2_or3_1 _1195_ (.A(_0295_),
    .B(_0297_),
    .C(_0304_),
    .X(_0305_));
 sg13g2_o21ai_1 _1196_ (.B1(_0304_),
    .Y(_0306_),
    .A1(_0295_),
    .A2(_0297_));
 sg13g2_nand3_1 _1197_ (.B(_0305_),
    .C(_0306_),
    .A(_0287_),
    .Y(_0307_));
 sg13g2_a21oi_1 _1198_ (.A1(_0305_),
    .A2(_0306_),
    .Y(_0308_),
    .B1(_0287_));
 sg13g2_a21o_1 _1199_ (.A2(_0306_),
    .A1(_0305_),
    .B1(_0287_),
    .X(_0309_));
 sg13g2_nand3_1 _1200_ (.B(_0307_),
    .C(_0309_),
    .A(_0286_),
    .Y(_0310_));
 sg13g2_a21o_1 _1201_ (.A2(_0309_),
    .A1(_0307_),
    .B1(_0286_),
    .X(_0311_));
 sg13g2_and3_1 _1202_ (.X(_0312_),
    .A(_0284_),
    .B(_0310_),
    .C(_0311_));
 sg13g2_nand3_1 _1203_ (.B(_0310_),
    .C(_0311_),
    .A(_0284_),
    .Y(_0313_));
 sg13g2_a21oi_1 _1204_ (.A1(_0310_),
    .A2(_0311_),
    .Y(_0314_),
    .B1(_0284_));
 sg13g2_or3_1 _1205_ (.A(_0283_),
    .B(_0312_),
    .C(_0314_),
    .X(_0315_));
 sg13g2_o21ai_1 _1206_ (.B1(_0283_),
    .Y(_0316_),
    .A1(_0312_),
    .A2(_0314_));
 sg13g2_nand3_1 _1207_ (.B(_0315_),
    .C(_0316_),
    .A(_0282_),
    .Y(_0317_));
 sg13g2_a21o_1 _1208_ (.A2(_0316_),
    .A1(_0315_),
    .B1(_0282_),
    .X(_0318_));
 sg13g2_and2_1 _1209_ (.A(_0317_),
    .B(_0318_),
    .X(_0319_));
 sg13g2_o21ai_1 _1210_ (.B1(_0217_),
    .Y(_0320_),
    .A1(_0189_),
    .A2(_0218_));
 sg13g2_o21ai_1 _1211_ (.B1(_0279_),
    .Y(_0321_),
    .A1(_0277_),
    .A2(_0280_));
 sg13g2_nand3_1 _1212_ (.B(_0320_),
    .C(_0321_),
    .A(_0281_),
    .Y(_0322_));
 sg13g2_a21oi_1 _1213_ (.A1(_0281_),
    .A2(_0321_),
    .Y(_0323_),
    .B1(_0320_));
 sg13g2_a21o_1 _1214_ (.A2(_0321_),
    .A1(_0281_),
    .B1(_0320_),
    .X(_0324_));
 sg13g2_nand2_1 _1215_ (.Y(_0325_),
    .A(_0322_),
    .B(_0324_));
 sg13g2_and2_1 _1216_ (.A(_0221_),
    .B(_0245_),
    .X(_0326_));
 sg13g2_or2_2 _1217_ (.X(_0327_),
    .B(_0326_),
    .A(_0325_));
 sg13g2_nand2_1 _1218_ (.Y(_0328_),
    .A(_0322_),
    .B(_0327_));
 sg13g2_nand2_1 _1219_ (.Y(_0329_),
    .A(_0319_),
    .B(_0328_));
 sg13g2_xor2_1 _1220_ (.B(_0328_),
    .A(_0319_),
    .X(_0330_));
 sg13g2_inv_1 _1221_ (.Y(_0331_),
    .A(_0330_));
 sg13g2_o21ai_1 _1222_ (.B1(_0296_),
    .Y(_0332_),
    .A1(_0297_),
    .A2(_0304_));
 sg13g2_o21ai_1 _1223_ (.B1(_0291_),
    .Y(_0333_),
    .A1(_0289_),
    .A2(_0292_));
 sg13g2_nand2_1 _1224_ (.Y(_0334_),
    .A(net182),
    .B(net222));
 sg13g2_and4_1 _1225_ (.A(net185),
    .B(net187),
    .C(net211),
    .D(net216),
    .X(_0335_));
 sg13g2_nand4_1 _1226_ (.B(net186),
    .C(net211),
    .A(net184),
    .Y(_0336_),
    .D(net216));
 sg13g2_a22oi_1 _1227_ (.Y(_0337_),
    .B1(net216),
    .B2(net184),
    .A2(net211),
    .A1(net186));
 sg13g2_or3_1 _1228_ (.A(_0334_),
    .B(_0335_),
    .C(_0337_),
    .X(_0338_));
 sg13g2_o21ai_1 _1229_ (.B1(_0334_),
    .Y(_0339_),
    .A1(_0335_),
    .A2(_0337_));
 sg13g2_and3_1 _1230_ (.X(_0340_),
    .A(_0333_),
    .B(_0338_),
    .C(_0339_));
 sg13g2_nand3_1 _1231_ (.B(_0338_),
    .C(_0339_),
    .A(_0333_),
    .Y(_0341_));
 sg13g2_a21oi_1 _1232_ (.A1(_0338_),
    .A2(_0339_),
    .Y(_0342_),
    .B1(_0333_));
 sg13g2_nand2_1 _1233_ (.Y(_0343_),
    .A(net190),
    .B(net207));
 sg13g2_nand2_1 _1234_ (.Y(_0344_),
    .A(net181),
    .B(net209));
 sg13g2_nand2_1 _1235_ (.Y(_0345_),
    .A(net181),
    .B(net224));
 sg13g2_or2_1 _1236_ (.X(_0346_),
    .B(_0345_),
    .A(_0169_));
 sg13g2_xnor2_1 _1237_ (.Y(_0347_),
    .A(_0169_),
    .B(_0345_));
 sg13g2_xnor2_1 _1238_ (.Y(_0348_),
    .A(_0343_),
    .B(_0347_));
 sg13g2_or3_1 _1239_ (.A(_0340_),
    .B(_0342_),
    .C(_0348_),
    .X(_0349_));
 sg13g2_o21ai_1 _1240_ (.B1(_0348_),
    .Y(_0350_),
    .A1(_0340_),
    .A2(_0342_));
 sg13g2_and3_1 _1241_ (.X(_0351_),
    .A(_0332_),
    .B(_0349_),
    .C(_0350_));
 sg13g2_nor2_1 _1242_ (.A(_0301_),
    .B(_0303_),
    .Y(_0352_));
 sg13g2_a21oi_1 _1243_ (.A1(_0349_),
    .A2(_0350_),
    .Y(_0353_),
    .B1(_0332_));
 sg13g2_or3_1 _1244_ (.A(_0351_),
    .B(_0352_),
    .C(_0353_),
    .X(_0354_));
 sg13g2_nand2b_1 _1245_ (.Y(_0355_),
    .B(_0354_),
    .A_N(_0351_));
 sg13g2_o21ai_1 _1246_ (.B1(_0346_),
    .Y(_0356_),
    .A1(_0343_),
    .A2(_0347_));
 sg13g2_o21ai_1 _1247_ (.B1(_0341_),
    .Y(_0357_),
    .A1(_0342_),
    .A2(_0348_));
 sg13g2_nand2_1 _1248_ (.Y(_0358_),
    .A(net186),
    .B(net207));
 sg13g2_nand4_1 _1249_ (.B(net188),
    .C(net207),
    .A(net186),
    .Y(_0359_),
    .D(net209));
 sg13g2_inv_1 _1250_ (.Y(_0360_),
    .A(_0359_));
 sg13g2_a22oi_1 _1251_ (.Y(_0361_),
    .B1(net209),
    .B2(net186),
    .A2(net207),
    .A1(net188));
 sg13g2_nor2_1 _1252_ (.A(_0360_),
    .B(_0361_),
    .Y(_0362_));
 sg13g2_o21ai_1 _1253_ (.B1(_0336_),
    .Y(_0363_),
    .A1(_0334_),
    .A2(_0337_));
 sg13g2_nand2_1 _1254_ (.Y(_0364_),
    .A(net181),
    .B(net222));
 sg13g2_nand2_1 _1255_ (.Y(_0365_),
    .A(net183),
    .B(net211));
 sg13g2_nand2_1 _1256_ (.Y(_0366_),
    .A(net182),
    .B(net217));
 sg13g2_and4_1 _1257_ (.A(net182),
    .B(net185),
    .C(net211),
    .D(net216),
    .X(_0367_));
 sg13g2_a22oi_1 _1258_ (.Y(_0368_),
    .B1(net216),
    .B2(net182),
    .A2(net211),
    .A1(net184));
 sg13g2_or3_1 _1259_ (.A(_0364_),
    .B(_0367_),
    .C(_0368_),
    .X(_0369_));
 sg13g2_o21ai_1 _1260_ (.B1(_0364_),
    .Y(_0370_),
    .A1(_0367_),
    .A2(_0368_));
 sg13g2_nand3_1 _1261_ (.B(_0369_),
    .C(_0370_),
    .A(_0363_),
    .Y(_0371_));
 sg13g2_a21o_1 _1262_ (.A2(_0370_),
    .A1(_0369_),
    .B1(_0363_),
    .X(_0372_));
 sg13g2_nand3_1 _1263_ (.B(_0371_),
    .C(_0372_),
    .A(_0362_),
    .Y(_0373_));
 sg13g2_a21o_1 _1264_ (.A2(_0372_),
    .A1(_0371_),
    .B1(_0362_),
    .X(_0374_));
 sg13g2_nand3_1 _1265_ (.B(_0373_),
    .C(_0374_),
    .A(_0357_),
    .Y(_0375_));
 sg13g2_a21o_1 _1266_ (.A2(_0374_),
    .A1(_0373_),
    .B1(_0357_),
    .X(_0376_));
 sg13g2_nand2_1 _1267_ (.Y(_0377_),
    .A(_0375_),
    .B(_0376_));
 sg13g2_nand3_1 _1268_ (.B(_0375_),
    .C(_0376_),
    .A(_0356_),
    .Y(_0378_));
 sg13g2_xnor2_1 _1269_ (.Y(_0379_),
    .A(_0356_),
    .B(_0377_));
 sg13g2_nand2_1 _1270_ (.Y(_0380_),
    .A(_0355_),
    .B(_0379_));
 sg13g2_nand2_1 _1271_ (.Y(_0381_),
    .A(net190),
    .B(net204));
 sg13g2_xnor2_1 _1272_ (.Y(_0382_),
    .A(_0355_),
    .B(_0379_));
 sg13g2_o21ai_1 _1273_ (.B1(_0380_),
    .Y(_0383_),
    .A1(_0381_),
    .A2(_0382_));
 sg13g2_nand2_1 _1274_ (.Y(_0384_),
    .A(net188),
    .B(net204));
 sg13g2_nand2_1 _1275_ (.Y(_0385_),
    .A(_0375_),
    .B(_0378_));
 sg13g2_nand2_1 _1276_ (.Y(_0386_),
    .A(_0371_),
    .B(_0373_));
 sg13g2_nand2_1 _1277_ (.Y(_0387_),
    .A(net184),
    .B(net207));
 sg13g2_nand4_1 _1278_ (.B(net186),
    .C(net207),
    .A(net184),
    .Y(_0388_),
    .D(net209));
 sg13g2_inv_1 _1279_ (.Y(_0389_),
    .A(_0388_));
 sg13g2_a21oi_1 _1280_ (.A1(_0263_),
    .A2(_0358_),
    .Y(_0390_),
    .B1(_0389_));
 sg13g2_inv_1 _1281_ (.Y(_0391_),
    .A(_0390_));
 sg13g2_nand2b_1 _1282_ (.Y(_0392_),
    .B(_0369_),
    .A_N(_0367_));
 sg13g2_nand2_1 _1283_ (.Y(_0393_),
    .A(net181),
    .B(net217));
 sg13g2_nand2_1 _1284_ (.Y(_0394_),
    .A(net181),
    .B(net211));
 sg13g2_xor2_1 _1285_ (.B(_0393_),
    .A(_0365_),
    .X(_0395_));
 sg13g2_nand2_1 _1286_ (.Y(_0396_),
    .A(_0392_),
    .B(_0395_));
 sg13g2_xnor2_1 _1287_ (.Y(_0397_),
    .A(_0392_),
    .B(_0395_));
 sg13g2_xnor2_1 _1288_ (.Y(_0398_),
    .A(_0390_),
    .B(_0397_));
 sg13g2_nand2_1 _1289_ (.Y(_0399_),
    .A(_0386_),
    .B(_0398_));
 sg13g2_xnor2_1 _1290_ (.Y(_0400_),
    .A(_0386_),
    .B(_0398_));
 sg13g2_xnor2_1 _1291_ (.Y(_0401_),
    .A(_0360_),
    .B(_0400_));
 sg13g2_nand2_1 _1292_ (.Y(_0402_),
    .A(_0385_),
    .B(_0401_));
 sg13g2_xnor2_1 _1293_ (.Y(_0403_),
    .A(_0385_),
    .B(_0401_));
 sg13g2_xor2_1 _1294_ (.B(_0403_),
    .A(_0384_),
    .X(_0404_));
 sg13g2_nand2_1 _1295_ (.Y(_0405_),
    .A(_0383_),
    .B(_0404_));
 sg13g2_nor2_1 _1296_ (.A(_0383_),
    .B(_0404_),
    .Y(_0406_));
 sg13g2_xnor2_1 _1297_ (.Y(_0407_),
    .A(_0383_),
    .B(_0404_));
 sg13g2_o21ai_1 _1298_ (.B1(_0307_),
    .Y(_0408_),
    .A1(_0285_),
    .A2(_0308_));
 sg13g2_o21ai_1 _1299_ (.B1(_0352_),
    .Y(_0409_),
    .A1(_0351_),
    .A2(_0353_));
 sg13g2_nand3_1 _1300_ (.B(_0408_),
    .C(_0409_),
    .A(_0354_),
    .Y(_0410_));
 sg13g2_and2_1 _1301_ (.A(net192),
    .B(net204),
    .X(_0411_));
 sg13g2_a21o_1 _1302_ (.A2(_0409_),
    .A1(_0354_),
    .B1(_0408_),
    .X(_0412_));
 sg13g2_nand3_1 _1303_ (.B(_0411_),
    .C(_0412_),
    .A(_0410_),
    .Y(_0413_));
 sg13g2_nand2_1 _1304_ (.Y(_0414_),
    .A(_0410_),
    .B(_0413_));
 sg13g2_xor2_1 _1305_ (.B(_0382_),
    .A(_0381_),
    .X(_0415_));
 sg13g2_nand2_1 _1306_ (.Y(_0416_),
    .A(_0414_),
    .B(_0415_));
 sg13g2_o21ai_1 _1307_ (.B1(_0313_),
    .Y(_0417_),
    .A1(_0283_),
    .A2(_0314_));
 sg13g2_a21o_1 _1308_ (.A2(_0412_),
    .A1(_0410_),
    .B1(_0411_),
    .X(_0418_));
 sg13g2_nand3_1 _1309_ (.B(_0417_),
    .C(_0418_),
    .A(_0413_),
    .Y(_0419_));
 sg13g2_a21o_1 _1310_ (.A2(_0418_),
    .A1(_0413_),
    .B1(_0417_),
    .X(_0420_));
 sg13g2_and2_1 _1311_ (.A(_0419_),
    .B(_0420_),
    .X(_0421_));
 sg13g2_and4_1 _1312_ (.A(_0317_),
    .B(_0318_),
    .C(_0419_),
    .D(_0420_),
    .X(_0422_));
 sg13g2_nand4_1 _1313_ (.B(_0318_),
    .C(_0419_),
    .A(_0317_),
    .Y(_0423_),
    .D(_0420_));
 sg13g2_nand4_1 _1314_ (.B(_0222_),
    .C(_0322_),
    .A(_0221_),
    .Y(_0424_),
    .D(_0324_));
 sg13g2_or4_1 _1315_ (.A(_0233_),
    .B(_0242_),
    .C(_0423_),
    .D(_0424_),
    .X(_0425_));
 sg13g2_o21ai_1 _1316_ (.B1(_0322_),
    .Y(_0426_),
    .A1(_0221_),
    .A2(_0323_));
 sg13g2_nand2_1 _1317_ (.Y(_0427_),
    .A(_0317_),
    .B(_0419_));
 sg13g2_a22oi_1 _1318_ (.Y(_0428_),
    .B1(_0427_),
    .B2(_0420_),
    .A2(_0426_),
    .A1(_0422_));
 sg13g2_nand2_1 _1319_ (.Y(_0429_),
    .A(_0425_),
    .B(_0428_));
 sg13g2_xor2_1 _1320_ (.B(_0415_),
    .A(_0414_),
    .X(_0430_));
 sg13g2_nand2_1 _1321_ (.Y(_0431_),
    .A(_0429_),
    .B(_0430_));
 sg13g2_and2_1 _1322_ (.A(_0416_),
    .B(_0431_),
    .X(_0432_));
 sg13g2_nand2_1 _1323_ (.Y(_0433_),
    .A(_0407_),
    .B(_0432_));
 sg13g2_or2_1 _1324_ (.X(_0434_),
    .B(_0432_),
    .A(_0407_));
 sg13g2_xnor2_1 _1325_ (.Y(_0435_),
    .A(_0407_),
    .B(_0432_));
 sg13g2_inv_1 _1326_ (.Y(_0436_),
    .A(_0435_));
 sg13g2_nand2b_1 _1327_ (.Y(_0437_),
    .B(_0430_),
    .A_N(_0407_));
 sg13g2_a21oi_1 _1328_ (.A1(_0425_),
    .A2(_0428_),
    .Y(_0438_),
    .B1(_0437_));
 sg13g2_o21ai_1 _1329_ (.B1(_0405_),
    .Y(_0439_),
    .A1(_0406_),
    .A2(_0416_));
 sg13g2_nor2_1 _1330_ (.A(_0438_),
    .B(_0439_),
    .Y(_0440_));
 sg13g2_o21ai_1 _1331_ (.B1(_0402_),
    .Y(_0441_),
    .A1(_0384_),
    .A2(_0403_));
 sg13g2_nand2_1 _1332_ (.Y(_0442_),
    .A(net186),
    .B(net204));
 sg13g2_o21ai_1 _1333_ (.B1(_0399_),
    .Y(_0443_),
    .A1(_0359_),
    .A2(_0400_));
 sg13g2_o21ai_1 _1334_ (.B1(_0396_),
    .Y(_0444_),
    .A1(_0391_),
    .A2(_0397_));
 sg13g2_nor2b_1 _1335_ (.A(_0394_),
    .B_N(_0366_),
    .Y(_0445_));
 sg13g2_nand2_1 _1336_ (.Y(_0446_),
    .A(net182),
    .B(net207));
 sg13g2_or2_1 _1337_ (.X(_0447_),
    .B(_0446_),
    .A(_0263_));
 sg13g2_inv_1 _1338_ (.Y(_0448_),
    .A(_0447_));
 sg13g2_a21oi_1 _1339_ (.A1(_0299_),
    .A2(_0387_),
    .Y(_0449_),
    .B1(_0448_));
 sg13g2_inv_1 _1340_ (.Y(_0450_),
    .A(_0449_));
 sg13g2_xnor2_1 _1341_ (.Y(_0451_),
    .A(_0445_),
    .B(_0449_));
 sg13g2_nand2b_1 _1342_ (.Y(_0452_),
    .B(_0444_),
    .A_N(_0451_));
 sg13g2_xor2_1 _1343_ (.B(_0451_),
    .A(_0444_),
    .X(_0453_));
 sg13g2_xnor2_1 _1344_ (.Y(_0454_),
    .A(_0389_),
    .B(_0453_));
 sg13g2_nand2_1 _1345_ (.Y(_0455_),
    .A(_0443_),
    .B(_0454_));
 sg13g2_xor2_1 _1346_ (.B(_0454_),
    .A(_0443_),
    .X(_0456_));
 sg13g2_nand2b_1 _1347_ (.Y(_0457_),
    .B(_0456_),
    .A_N(_0442_));
 sg13g2_xnor2_1 _1348_ (.Y(_0458_),
    .A(_0442_),
    .B(_0456_));
 sg13g2_nand2_1 _1349_ (.Y(_0459_),
    .A(_0441_),
    .B(_0458_));
 sg13g2_xnor2_1 _1350_ (.Y(_0460_),
    .A(_0441_),
    .B(_0458_));
 sg13g2_inv_1 _1351_ (.Y(_0461_),
    .A(_0460_));
 sg13g2_o21ai_1 _1352_ (.B1(_0461_),
    .Y(_0462_),
    .A1(_0438_),
    .A2(_0439_));
 sg13g2_xnor2_1 _1353_ (.Y(_0463_),
    .A(_0440_),
    .B(_0461_));
 sg13g2_and2_1 _1354_ (.A(_0455_),
    .B(_0457_),
    .X(_0464_));
 sg13g2_nand2_1 _1355_ (.Y(_0465_),
    .A(net184),
    .B(net204));
 sg13g2_o21ai_1 _1356_ (.B1(_0452_),
    .Y(_0466_),
    .A1(_0388_),
    .A2(_0453_));
 sg13g2_a21oi_1 _1357_ (.A1(_0366_),
    .A2(_0450_),
    .Y(_0467_),
    .B1(_0394_));
 sg13g2_or2_1 _1358_ (.X(_0468_),
    .B(_0446_),
    .A(_0344_));
 sg13g2_xor2_1 _1359_ (.B(_0446_),
    .A(_0344_),
    .X(_0469_));
 sg13g2_nand2_1 _1360_ (.Y(_0470_),
    .A(_0467_),
    .B(_0469_));
 sg13g2_xnor2_1 _1361_ (.Y(_0471_),
    .A(_0467_),
    .B(_0469_));
 sg13g2_xnor2_1 _1362_ (.Y(_0472_),
    .A(_0448_),
    .B(_0471_));
 sg13g2_nand2_1 _1363_ (.Y(_0473_),
    .A(_0466_),
    .B(_0472_));
 sg13g2_xnor2_1 _1364_ (.Y(_0474_),
    .A(_0466_),
    .B(_0472_));
 sg13g2_xnor2_1 _1365_ (.Y(_0475_),
    .A(_0465_),
    .B(_0474_));
 sg13g2_and2_1 _1366_ (.A(_0464_),
    .B(_0475_),
    .X(_0476_));
 sg13g2_or2_1 _1367_ (.X(_0477_),
    .B(_0475_),
    .A(_0464_));
 sg13g2_and2_1 _1368_ (.A(_0459_),
    .B(_0477_),
    .X(_0478_));
 sg13g2_a21oi_1 _1369_ (.A1(_0462_),
    .A2(_0478_),
    .Y(_0479_),
    .B1(_0476_));
 sg13g2_o21ai_1 _1370_ (.B1(_0473_),
    .Y(_0480_),
    .A1(_0465_),
    .A2(_0474_));
 sg13g2_nand2_1 _1371_ (.Y(_0481_),
    .A(net182),
    .B(net204));
 sg13g2_o21ai_1 _1372_ (.B1(_0470_),
    .Y(_0482_),
    .A1(_0447_),
    .A2(_0471_));
 sg13g2_nand3_1 _1373_ (.B(net207),
    .C(_0299_),
    .A(net181),
    .Y(_0483_));
 sg13g2_nand2b_1 _1374_ (.Y(_0484_),
    .B(_0482_),
    .A_N(_0483_));
 sg13g2_xor2_1 _1375_ (.B(_0483_),
    .A(_0482_),
    .X(_0485_));
 sg13g2_or2_1 _1376_ (.X(_0486_),
    .B(_0485_),
    .A(_0481_));
 sg13g2_xor2_1 _1377_ (.B(_0485_),
    .A(_0481_),
    .X(_0487_));
 sg13g2_and2_1 _1378_ (.A(_0480_),
    .B(_0487_),
    .X(_0488_));
 sg13g2_xnor2_1 _1379_ (.Y(_0489_),
    .A(_0480_),
    .B(_0487_));
 sg13g2_a221oi_1 _1380_ (.B2(_0462_),
    .C1(_0489_),
    .B1(_0478_),
    .A1(_0464_),
    .Y(_0490_),
    .A2(_0475_));
 sg13g2_xor2_1 _1381_ (.B(_0489_),
    .A(_0479_),
    .X(_0491_));
 sg13g2_nand2b_1 _1382_ (.Y(_0492_),
    .B(_0477_),
    .A_N(_0476_));
 sg13g2_inv_1 _1383_ (.Y(_0493_),
    .A(_0492_));
 sg13g2_a21oi_1 _1384_ (.A1(_0459_),
    .A2(_0462_),
    .Y(_0494_),
    .B1(_0493_));
 sg13g2_and3_1 _1385_ (.X(_0495_),
    .A(_0459_),
    .B(_0462_),
    .C(_0493_));
 sg13g2_nor2_1 _1386_ (.A(_0494_),
    .B(_0495_),
    .Y(_0496_));
 sg13g2_inv_1 _1387_ (.Y(_0497_),
    .A(_0496_));
 sg13g2_nor3_2 _1388_ (.A(_0463_),
    .B(_0494_),
    .C(_0495_),
    .Y(_0498_));
 sg13g2_nand2_1 _1389_ (.Y(_0499_),
    .A(_0491_),
    .B(_0498_));
 sg13g2_nand2_1 _1390_ (.Y(_0500_),
    .A(net181),
    .B(net204));
 sg13g2_nor2_1 _1391_ (.A(_0051_),
    .B(_0468_),
    .Y(_0501_));
 sg13g2_a21o_1 _1392_ (.A2(_0500_),
    .A1(_0468_),
    .B1(_0501_),
    .X(_0502_));
 sg13g2_and3_1 _1393_ (.X(_0503_),
    .A(_0484_),
    .B(_0486_),
    .C(_0502_));
 sg13g2_a21oi_1 _1394_ (.A1(_0484_),
    .A2(_0486_),
    .Y(_0504_),
    .B1(_0502_));
 sg13g2_or2_1 _1395_ (.X(_0505_),
    .B(_0504_),
    .A(_0503_));
 sg13g2_nor2_1 _1396_ (.A(_0488_),
    .B(_0490_),
    .Y(_0506_));
 sg13g2_o21ai_1 _1397_ (.B1(_0505_),
    .Y(_0507_),
    .A1(_0488_),
    .A2(_0490_));
 sg13g2_or3_1 _1398_ (.A(_0488_),
    .B(_0490_),
    .C(_0505_),
    .X(_0508_));
 sg13g2_nand2_1 _1399_ (.Y(_0509_),
    .A(_0507_),
    .B(_0508_));
 sg13g2_nand2_1 _1400_ (.Y(_0510_),
    .A(_0499_),
    .B(_0509_));
 sg13g2_nor2_1 _1401_ (.A(_0501_),
    .B(_0504_),
    .Y(_0511_));
 sg13g2_a221oi_1 _1402_ (.B2(_0508_),
    .C1(_0511_),
    .B1(_0507_),
    .A1(_0491_),
    .Y(_0512_),
    .A2(_0498_));
 sg13g2_nor2b_1 _1403_ (.A(_0463_),
    .B_N(_0512_),
    .Y(_0513_));
 sg13g2_xnor2_1 _1404_ (.Y(_0514_),
    .A(_0463_),
    .B(_0512_));
 sg13g2_inv_1 _1405_ (.Y(_0515_),
    .A(_0514_));
 sg13g2_nor2_1 _1406_ (.A(_0436_),
    .B(_0497_),
    .Y(_0516_));
 sg13g2_nand2_1 _1407_ (.Y(_0517_),
    .A(_0514_),
    .B(_0516_));
 sg13g2_nand2b_1 _1408_ (.Y(_0518_),
    .B(_0509_),
    .A_N(_0512_));
 sg13g2_a21o_1 _1409_ (.A2(_0512_),
    .A1(_0498_),
    .B1(_0491_),
    .X(_0519_));
 sg13g2_nand3b_1 _1410_ (.B(_0509_),
    .C(_0511_),
    .Y(_0520_),
    .A_N(_0491_));
 sg13g2_a21oi_1 _1411_ (.A1(_0514_),
    .A2(_0516_),
    .Y(_0521_),
    .B1(_0520_));
 sg13g2_a21o_2 _1412_ (.A2(_0516_),
    .A1(_0514_),
    .B1(_0520_),
    .X(_0522_));
 sg13g2_o21ai_1 _1413_ (.B1(_0511_),
    .Y(_0523_),
    .A1(_0505_),
    .A2(_0506_));
 sg13g2_and2_1 _1414_ (.A(_0510_),
    .B(_0523_),
    .X(_0524_));
 sg13g2_nand2_2 _1415_ (.Y(_0525_),
    .A(_0510_),
    .B(_0523_));
 sg13g2_nor2_1 _1416_ (.A(_0521_),
    .B(_0524_),
    .Y(_0526_));
 sg13g2_a21oi_2 _1417_ (.B1(_0436_),
    .Y(_0527_),
    .A2(_0525_),
    .A1(_0522_));
 sg13g2_nand3_1 _1418_ (.B(_0522_),
    .C(_0525_),
    .A(_0436_),
    .Y(_0528_));
 sg13g2_nor2b_1 _1419_ (.A(_0527_),
    .B_N(_0528_),
    .Y(_0529_));
 sg13g2_inv_1 _1420_ (.Y(_0530_),
    .A(_0529_));
 sg13g2_or2_1 _1421_ (.X(_0531_),
    .B(_0430_),
    .A(_0429_));
 sg13g2_nand2_1 _1422_ (.Y(_0532_),
    .A(_0431_),
    .B(_0531_));
 sg13g2_inv_1 _1423_ (.Y(_0533_),
    .A(_0532_));
 sg13g2_a221oi_1 _1424_ (.B2(_0525_),
    .C1(_0515_),
    .B1(_0522_),
    .A1(_0433_),
    .Y(_0534_),
    .A2(_0434_));
 sg13g2_o21ai_1 _1425_ (.B1(_0497_),
    .Y(_0535_),
    .A1(_0513_),
    .A2(_0534_));
 sg13g2_or3_1 _1426_ (.A(_0497_),
    .B(_0513_),
    .C(_0534_),
    .X(_0536_));
 sg13g2_nand2_1 _1427_ (.Y(_0537_),
    .A(_0535_),
    .B(_0536_));
 sg13g2_nor2_1 _1428_ (.A(_0515_),
    .B(_0533_),
    .Y(_0538_));
 sg13g2_nand3b_1 _1429_ (.B(_0528_),
    .C(_0538_),
    .Y(_0539_),
    .A_N(_0527_));
 sg13g2_o21ai_1 _1430_ (.B1(_0517_),
    .Y(_0540_),
    .A1(_0521_),
    .A2(_0524_));
 sg13g2_xor2_1 _1431_ (.B(_0540_),
    .A(_0519_),
    .X(_0541_));
 sg13g2_nand4_1 _1432_ (.B(_0536_),
    .C(_0539_),
    .A(_0535_),
    .Y(_0542_),
    .D(_0541_));
 sg13g2_o21ai_1 _1433_ (.B1(_0518_),
    .Y(_0543_),
    .A1(_0519_),
    .A2(_0540_));
 sg13g2_nand2_2 _1434_ (.Y(_0544_),
    .A(_0522_),
    .B(_0543_));
 sg13g2_nand2_1 _1435_ (.Y(_0545_),
    .A(_0542_),
    .B(_0544_));
 sg13g2_a21oi_2 _1436_ (.B1(_0533_),
    .Y(_0546_),
    .A2(_0544_),
    .A1(_0542_));
 sg13g2_a221oi_1 _1437_ (.B2(_0544_),
    .C1(_0530_),
    .B1(_0542_),
    .A1(_0431_),
    .Y(_0547_),
    .A2(_0531_));
 sg13g2_xnor2_1 _1438_ (.Y(_0548_),
    .A(_0515_),
    .B(_0527_));
 sg13g2_or2_1 _1439_ (.X(_0549_),
    .B(_0544_),
    .A(_0539_));
 sg13g2_mux2_1 _1440_ (.A0(_0548_),
    .A1(_0515_),
    .S(_0547_),
    .X(_0550_));
 sg13g2_o21ai_1 _1441_ (.B1(_0549_),
    .Y(_0551_),
    .A1(_0547_),
    .A2(_0548_));
 sg13g2_nand3_1 _1442_ (.B(_0542_),
    .C(_0544_),
    .A(_0533_),
    .Y(_0552_));
 sg13g2_nor2b_2 _1443_ (.A(_0546_),
    .B_N(_0552_),
    .Y(_0553_));
 sg13g2_inv_1 _1444_ (.Y(_0554_),
    .A(_0553_));
 sg13g2_nand2_1 _1445_ (.Y(_0555_),
    .A(_0317_),
    .B(_0329_));
 sg13g2_or2_1 _1446_ (.X(_0556_),
    .B(_0555_),
    .A(_0421_));
 sg13g2_nand2_1 _1447_ (.Y(_0557_),
    .A(_0421_),
    .B(_0555_));
 sg13g2_and2_1 _1448_ (.A(_0556_),
    .B(_0557_),
    .X(_0558_));
 sg13g2_nor2_1 _1449_ (.A(_0530_),
    .B(_0558_),
    .Y(_0559_));
 sg13g2_nand3b_1 _1450_ (.B(_0552_),
    .C(_0559_),
    .Y(_0560_),
    .A_N(_0546_));
 sg13g2_a22oi_1 _1451_ (.Y(_0561_),
    .B1(_0542_),
    .B2(_0544_),
    .A2(_0538_),
    .A1(_0529_));
 sg13g2_a221oi_1 _1452_ (.B2(_0544_),
    .C1(_0537_),
    .B1(_0542_),
    .A1(_0529_),
    .Y(_0562_),
    .A2(_0538_));
 sg13g2_xnor2_1 _1453_ (.Y(_0563_),
    .A(_0537_),
    .B(_0561_));
 sg13g2_and3_1 _1454_ (.X(_0564_),
    .A(_0551_),
    .B(_0560_),
    .C(_0563_));
 sg13g2_nand3b_1 _1455_ (.B(_0560_),
    .C(_0563_),
    .Y(_0565_),
    .A_N(_0550_));
 sg13g2_o21ai_1 _1456_ (.B1(_0542_),
    .Y(_0566_),
    .A1(_0541_),
    .A2(_0562_));
 sg13g2_inv_1 _1457_ (.Y(_0567_),
    .A(_0566_));
 sg13g2_nor2_1 _1458_ (.A(_0564_),
    .B(_0567_),
    .Y(_0568_));
 sg13g2_a221oi_1 _1459_ (.B2(_0566_),
    .C1(_0550_),
    .B1(_0565_),
    .A1(_0553_),
    .Y(_0569_),
    .A2(_0559_));
 sg13g2_nor2_1 _1460_ (.A(_0563_),
    .B(_0569_),
    .Y(_0570_));
 sg13g2_nor2_2 _1461_ (.A(_0564_),
    .B(_0570_),
    .Y(_0571_));
 sg13g2_o21ai_1 _1462_ (.B1(_0565_),
    .Y(_0572_),
    .A1(_0563_),
    .A2(_0569_));
 sg13g2_a21o_1 _1463_ (.A2(_0566_),
    .A1(_0565_),
    .B1(_0558_),
    .X(_0573_));
 sg13g2_a221oi_1 _1464_ (.B2(_0566_),
    .C1(_0554_),
    .B1(_0565_),
    .A1(_0556_),
    .Y(_0574_),
    .A2(_0557_));
 sg13g2_or3_1 _1465_ (.A(_0530_),
    .B(_0546_),
    .C(_0574_),
    .X(_0575_));
 sg13g2_o21ai_1 _1466_ (.B1(_0530_),
    .Y(_0576_),
    .A1(_0546_),
    .A2(_0574_));
 sg13g2_nand2_1 _1467_ (.Y(_0577_),
    .A(_0575_),
    .B(_0576_));
 sg13g2_a21oi_1 _1468_ (.A1(_0560_),
    .A2(_0567_),
    .Y(_0578_),
    .B1(_0551_));
 sg13g2_or2_1 _1469_ (.X(_0579_),
    .B(_0578_),
    .A(_0569_));
 sg13g2_nor3_1 _1470_ (.A(_0563_),
    .B(_0569_),
    .C(_0578_),
    .Y(_0580_));
 sg13g2_xnor2_1 _1471_ (.Y(_0581_),
    .A(_0553_),
    .B(_0573_));
 sg13g2_nand3_1 _1472_ (.B(_0565_),
    .C(_0566_),
    .A(_0558_),
    .Y(_0582_));
 sg13g2_and2_1 _1473_ (.A(_0573_),
    .B(_0582_),
    .X(_0583_));
 sg13g2_and2_1 _1474_ (.A(_0331_),
    .B(_0583_),
    .X(_0584_));
 sg13g2_nand4_1 _1475_ (.B(_0553_),
    .C(_0573_),
    .A(_0331_),
    .Y(_0585_),
    .D(_0582_));
 sg13g2_and4_1 _1476_ (.A(_0575_),
    .B(_0576_),
    .C(_0580_),
    .D(_0585_),
    .X(_0586_));
 sg13g2_nand4_1 _1477_ (.B(_0576_),
    .C(_0580_),
    .A(_0575_),
    .Y(_0587_),
    .D(_0585_));
 sg13g2_a21oi_2 _1478_ (.B1(_0330_),
    .Y(_0588_),
    .A2(_0587_),
    .A1(_0572_));
 sg13g2_nor3_1 _1479_ (.A(_0331_),
    .B(_0571_),
    .C(_0586_),
    .Y(_0589_));
 sg13g2_or2_1 _1480_ (.X(_0590_),
    .B(_0589_),
    .A(_0588_));
 sg13g2_nand2_2 _1481_ (.Y(_0591_),
    .A(_0325_),
    .B(_0326_));
 sg13g2_nand2_1 _1482_ (.Y(_0592_),
    .A(_0327_),
    .B(_0591_));
 sg13g2_o21ai_1 _1483_ (.B1(_0584_),
    .Y(_0593_),
    .A1(_0571_),
    .A2(_0586_));
 sg13g2_xnor2_1 _1484_ (.Y(_0594_),
    .A(_0581_),
    .B(_0593_));
 sg13g2_nand2_1 _1485_ (.Y(_0595_),
    .A(_0583_),
    .B(_0592_));
 sg13g2_nor3_2 _1486_ (.A(_0588_),
    .B(_0589_),
    .C(_0595_),
    .Y(_0596_));
 sg13g2_o21ai_1 _1487_ (.B1(_0585_),
    .Y(_0597_),
    .A1(_0571_),
    .A2(_0586_));
 sg13g2_nor2_1 _1488_ (.A(_0577_),
    .B(_0597_),
    .Y(_0598_));
 sg13g2_xnor2_1 _1489_ (.Y(_0599_),
    .A(_0577_),
    .B(_0597_));
 sg13g2_nor3_2 _1490_ (.A(_0594_),
    .B(_0596_),
    .C(_0599_),
    .Y(_0600_));
 sg13g2_or3_1 _1491_ (.A(_0594_),
    .B(_0596_),
    .C(_0599_),
    .X(_0601_));
 sg13g2_xnor2_1 _1492_ (.Y(_0602_),
    .A(_0579_),
    .B(_0598_));
 sg13g2_xor2_1 _1493_ (.B(_0598_),
    .A(_0579_),
    .X(_0603_));
 sg13g2_nor2_2 _1494_ (.A(_0600_),
    .B(_0602_),
    .Y(_0604_));
 sg13g2_a22oi_1 _1495_ (.Y(_0605_),
    .B1(_0601_),
    .B2(_0603_),
    .A2(_0591_),
    .A1(_0327_));
 sg13g2_nor3_1 _1496_ (.A(_0592_),
    .B(_0600_),
    .C(_0602_),
    .Y(_0606_));
 sg13g2_nor2_1 _1497_ (.A(_0605_),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_inv_1 _1498_ (.Y(_0608_),
    .A(_0607_));
 sg13g2_nor3_1 _1499_ (.A(_0590_),
    .B(_0605_),
    .C(_0606_),
    .Y(_0609_));
 sg13g2_or2_1 _1500_ (.X(_0610_),
    .B(_0588_),
    .A(_0583_));
 sg13g2_and2_1 _1501_ (.A(_0593_),
    .B(_0610_),
    .X(_0611_));
 sg13g2_a221oi_1 _1502_ (.B2(_0603_),
    .C1(_0590_),
    .B1(_0601_),
    .A1(_0327_),
    .Y(_0612_),
    .A2(_0591_));
 sg13g2_xnor2_1 _1503_ (.Y(_0613_),
    .A(_0611_),
    .B(_0612_));
 sg13g2_nor2_1 _1504_ (.A(_0246_),
    .B(_0611_),
    .Y(_0614_));
 sg13g2_mux2_1 _1505_ (.A0(_0613_),
    .A1(_0614_),
    .S(_0609_),
    .X(_0615_));
 sg13g2_or3_1 _1506_ (.A(_0594_),
    .B(_0596_),
    .C(_0604_),
    .X(_0616_));
 sg13g2_o21ai_1 _1507_ (.B1(_0594_),
    .Y(_0617_),
    .A1(_0596_),
    .A2(_0603_));
 sg13g2_and2_1 _1508_ (.A(_0616_),
    .B(_0617_),
    .X(_0618_));
 sg13g2_a21oi_1 _1509_ (.A1(_0599_),
    .A2(_0616_),
    .Y(_0619_),
    .B1(_0600_));
 sg13g2_a21oi_2 _1510_ (.B1(_0619_),
    .Y(_0620_),
    .A2(_0618_),
    .A1(_0615_));
 sg13g2_xnor2_1 _1511_ (.Y(_0621_),
    .A(_0246_),
    .B(_0620_));
 sg13g2_xnor2_1 _1512_ (.Y(_0622_),
    .A(_0241_),
    .B(_0243_));
 sg13g2_nor3_1 _1513_ (.A(_0247_),
    .B(_0608_),
    .C(_0620_),
    .Y(_0623_));
 sg13g2_or3_1 _1514_ (.A(_0590_),
    .B(_0605_),
    .C(_0623_),
    .X(_0624_));
 sg13g2_o21ai_1 _1515_ (.B1(_0590_),
    .Y(_0625_),
    .A1(_0605_),
    .A2(_0623_));
 sg13g2_nand2_1 _1516_ (.Y(_0626_),
    .A(_0624_),
    .B(_0625_));
 sg13g2_and2_1 _1517_ (.A(_0246_),
    .B(_0609_),
    .X(_0627_));
 sg13g2_or3_1 _1518_ (.A(_0613_),
    .B(_0620_),
    .C(_0627_),
    .X(_0628_));
 sg13g2_o21ai_1 _1519_ (.B1(_0613_),
    .Y(_0629_),
    .A1(_0620_),
    .A2(_0627_));
 sg13g2_nand2_1 _1520_ (.Y(_0630_),
    .A(_0628_),
    .B(_0629_));
 sg13g2_and2_1 _1521_ (.A(_0621_),
    .B(_0622_),
    .X(_0631_));
 sg13g2_and2_1 _1522_ (.A(_0607_),
    .B(_0622_),
    .X(_0632_));
 sg13g2_nand2_1 _1523_ (.Y(_0633_),
    .A(_0621_),
    .B(_0632_));
 sg13g2_inv_1 _1524_ (.Y(_0634_),
    .A(_0633_));
 sg13g2_a22oi_1 _1525_ (.Y(_0635_),
    .B1(_0632_),
    .B2(_0621_),
    .A2(_0629_),
    .A1(_0628_));
 sg13g2_and3_1 _1526_ (.X(_0636_),
    .A(_0624_),
    .B(_0625_),
    .C(_0633_));
 sg13g2_and3_1 _1527_ (.X(_0637_),
    .A(_0624_),
    .B(_0625_),
    .C(_0635_));
 sg13g2_nand3_1 _1528_ (.B(_0625_),
    .C(_0635_),
    .A(_0624_),
    .Y(_0638_));
 sg13g2_a21oi_1 _1529_ (.A1(_0615_),
    .A2(_0619_),
    .Y(_0639_),
    .B1(_0618_));
 sg13g2_a21oi_2 _1530_ (.B1(_0639_),
    .Y(_0640_),
    .A2(_0618_),
    .A1(_0615_));
 sg13g2_inv_1 _1531_ (.Y(_0641_),
    .A(_0640_));
 sg13g2_nor2_1 _1532_ (.A(_0637_),
    .B(_0640_),
    .Y(_0642_));
 sg13g2_o21ai_1 _1533_ (.B1(_0622_),
    .Y(_0643_),
    .A1(_0637_),
    .A2(_0640_));
 sg13g2_nand3b_1 _1534_ (.B(_0638_),
    .C(_0641_),
    .Y(_0644_),
    .A_N(_0622_));
 sg13g2_and2_1 _1535_ (.A(_0643_),
    .B(_0644_),
    .X(_0645_));
 sg13g2_xor2_1 _1536_ (.B(_0240_),
    .A(_0238_),
    .X(_0646_));
 sg13g2_inv_1 _1537_ (.Y(_0647_),
    .A(_0646_));
 sg13g2_nand3_1 _1538_ (.B(_0644_),
    .C(_0647_),
    .A(_0643_),
    .Y(_0648_));
 sg13g2_o21ai_1 _1539_ (.B1(_0636_),
    .Y(_0649_),
    .A1(_0630_),
    .A2(_0640_));
 sg13g2_a21o_1 _1540_ (.A2(_0640_),
    .A1(_0636_),
    .B1(_0630_),
    .X(_0650_));
 sg13g2_nand2_1 _1541_ (.Y(_0651_),
    .A(_0638_),
    .B(_0650_));
 sg13g2_o21ai_1 _1542_ (.B1(_0631_),
    .Y(_0652_),
    .A1(_0637_),
    .A2(_0640_));
 sg13g2_xnor2_1 _1543_ (.Y(_0653_),
    .A(_0621_),
    .B(_0643_));
 sg13g2_xor2_1 _1544_ (.B(_0643_),
    .A(_0621_),
    .X(_0654_));
 sg13g2_o21ai_1 _1545_ (.B1(_0608_),
    .Y(_0655_),
    .A1(_0247_),
    .A2(_0620_));
 sg13g2_nand2b_1 _1546_ (.Y(_0656_),
    .B(_0655_),
    .A_N(_0623_));
 sg13g2_o21ai_1 _1547_ (.B1(_0626_),
    .Y(_0657_),
    .A1(_0634_),
    .A2(_0641_));
 sg13g2_nand2_1 _1548_ (.Y(_0658_),
    .A(_0649_),
    .B(_0657_));
 sg13g2_nor2b_1 _1549_ (.A(_0650_),
    .B_N(_0657_),
    .Y(_0659_));
 sg13g2_a22oi_1 _1550_ (.Y(_0660_),
    .B1(_0652_),
    .B2(_0656_),
    .A2(_0640_),
    .A1(_0634_));
 sg13g2_nand4_1 _1551_ (.B(_0653_),
    .C(_0656_),
    .A(_0648_),
    .Y(_0661_),
    .D(_0659_));
 sg13g2_or4_1 _1552_ (.A(_0630_),
    .B(_0653_),
    .C(_0658_),
    .D(_0660_),
    .X(_0662_));
 sg13g2_nand2_1 _1553_ (.Y(_0663_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_and3_2 _1554_ (.X(_0664_),
    .A(_0651_),
    .B(_0661_),
    .C(_0662_));
 sg13g2_nand3_1 _1555_ (.B(_0661_),
    .C(_0662_),
    .A(_0651_),
    .Y(_0665_));
 sg13g2_nor2_1 _1556_ (.A(_0646_),
    .B(_0664_),
    .Y(_0666_));
 sg13g2_inv_1 _1557_ (.Y(_0667_),
    .A(_0666_));
 sg13g2_o21ai_1 _1558_ (.B1(_0653_),
    .Y(_0668_),
    .A1(_0648_),
    .A2(_0651_));
 sg13g2_nand4_1 _1559_ (.B(_0647_),
    .C(_0654_),
    .A(_0645_),
    .Y(_0669_),
    .D(_0665_));
 sg13g2_and2_1 _1560_ (.A(_0668_),
    .B(_0669_),
    .X(_0670_));
 sg13g2_xnor2_1 _1561_ (.Y(_0671_),
    .A(_0647_),
    .B(_0664_));
 sg13g2_inv_1 _1562_ (.Y(_0672_),
    .A(_0671_));
 sg13g2_and3_1 _1563_ (.X(_0673_),
    .A(_0128_),
    .B(_0645_),
    .C(_0671_));
 sg13g2_nand3_1 _1564_ (.B(_0645_),
    .C(_0671_),
    .A(_0128_),
    .Y(_0674_));
 sg13g2_nor2_1 _1565_ (.A(_0648_),
    .B(_0654_),
    .Y(_0675_));
 sg13g2_or3_1 _1566_ (.A(_0660_),
    .B(_0664_),
    .C(_0675_),
    .X(_0676_));
 sg13g2_o21ai_1 _1567_ (.B1(_0660_),
    .Y(_0677_),
    .A1(_0664_),
    .A2(_0675_));
 sg13g2_nand2_1 _1568_ (.Y(_0678_),
    .A(_0676_),
    .B(_0677_));
 sg13g2_nand4_1 _1569_ (.B(_0669_),
    .C(_0676_),
    .A(_0668_),
    .Y(_0679_),
    .D(_0677_));
 sg13g2_nor2_1 _1570_ (.A(_0673_),
    .B(_0679_),
    .Y(_0680_));
 sg13g2_a21o_1 _1571_ (.A2(_0676_),
    .A1(_0658_),
    .B1(_0663_),
    .X(_0681_));
 sg13g2_o21ai_1 _1572_ (.B1(_0681_),
    .Y(_0682_),
    .A1(_0673_),
    .A2(_0679_));
 sg13g2_inv_1 _1573_ (.Y(_0683_),
    .A(_0682_));
 sg13g2_xnor2_1 _1574_ (.Y(_0684_),
    .A(_0128_),
    .B(_0682_));
 sg13g2_nand2b_1 _1575_ (.Y(_0685_),
    .B(_0099_),
    .A_N(_0076_));
 sg13g2_and2_1 _1576_ (.A(_0100_),
    .B(_0685_),
    .X(_0686_));
 sg13g2_nand3_1 _1577_ (.B(_0671_),
    .C(_0682_),
    .A(_0128_),
    .Y(_0687_));
 sg13g2_nand3_1 _1578_ (.B(_0667_),
    .C(_0687_),
    .A(_0645_),
    .Y(_0688_));
 sg13g2_a21o_1 _1579_ (.A2(_0687_),
    .A1(_0667_),
    .B1(_0645_),
    .X(_0689_));
 sg13g2_and2_1 _1580_ (.A(_0688_),
    .B(_0689_),
    .X(_0690_));
 sg13g2_nand3_1 _1581_ (.B(_0674_),
    .C(_0682_),
    .A(_0670_),
    .Y(_0691_));
 sg13g2_a21o_1 _1582_ (.A2(_0682_),
    .A1(_0674_),
    .B1(_0670_),
    .X(_0692_));
 sg13g2_and2_1 _1583_ (.A(_0691_),
    .B(_0692_),
    .X(_0693_));
 sg13g2_or3_1 _1584_ (.A(_0672_),
    .B(_0684_),
    .C(_0686_),
    .X(_0694_));
 sg13g2_and2_1 _1585_ (.A(_0690_),
    .B(_0694_),
    .X(_0695_));
 sg13g2_and2_1 _1586_ (.A(_0693_),
    .B(_0695_),
    .X(_0696_));
 sg13g2_nand4_1 _1587_ (.B(_0689_),
    .C(_0693_),
    .A(_0688_),
    .Y(_0697_),
    .D(_0694_));
 sg13g2_a21o_2 _1588_ (.A2(_0691_),
    .A1(_0678_),
    .B1(_0680_),
    .X(_0698_));
 sg13g2_inv_1 _1589_ (.Y(_0699_),
    .A(_0698_));
 sg13g2_nand2_2 _1590_ (.Y(_0700_),
    .A(_0697_),
    .B(_0698_));
 sg13g2_a21oi_2 _1591_ (.B1(_0686_),
    .Y(_0701_),
    .A2(_0698_),
    .A1(_0697_));
 sg13g2_a221oi_1 _1592_ (.B2(_0698_),
    .C1(_0684_),
    .B1(_0697_),
    .A1(_0100_),
    .Y(_0702_),
    .A2(_0685_));
 sg13g2_xnor2_1 _1593_ (.Y(_0703_),
    .A(_0684_),
    .B(_0701_));
 sg13g2_and3_1 _1594_ (.X(_0704_),
    .A(_0686_),
    .B(_0697_),
    .C(_0698_));
 sg13g2_nor2_1 _1595_ (.A(_0701_),
    .B(_0704_),
    .Y(_0705_));
 sg13g2_xnor2_1 _1596_ (.Y(_0706_),
    .A(_0062_),
    .B(_0075_));
 sg13g2_inv_1 _1597_ (.Y(_0707_),
    .A(_0706_));
 sg13g2_a21oi_1 _1598_ (.A1(_0695_),
    .A2(_0700_),
    .Y(_0708_),
    .B1(_0693_));
 sg13g2_or2_1 _1599_ (.X(_0709_),
    .B(_0708_),
    .A(_0696_));
 sg13g2_a21o_1 _1600_ (.A2(_0682_),
    .A1(_0128_),
    .B1(_0671_),
    .X(_0710_));
 sg13g2_and2_1 _1601_ (.A(_0687_),
    .B(_0710_),
    .X(_0711_));
 sg13g2_mux2_1 _1602_ (.A0(_0711_),
    .A1(_0672_),
    .S(_0702_),
    .X(_0712_));
 sg13g2_nor2_1 _1603_ (.A(_0684_),
    .B(_0707_),
    .Y(_0713_));
 sg13g2_nor4_2 _1604_ (.A(_0684_),
    .B(_0701_),
    .C(_0704_),
    .Y(_0714_),
    .D(_0707_));
 sg13g2_a21oi_1 _1605_ (.A1(_0694_),
    .A2(_0699_),
    .Y(_0715_),
    .B1(_0690_));
 sg13g2_a21oi_1 _1606_ (.A1(_0695_),
    .A2(_0700_),
    .Y(_0716_),
    .B1(_0715_));
 sg13g2_a21o_1 _1607_ (.A2(_0700_),
    .A1(_0695_),
    .B1(_0715_),
    .X(_0717_));
 sg13g2_or3_1 _1608_ (.A(_0712_),
    .B(_0714_),
    .C(_0717_),
    .X(_0718_));
 sg13g2_nand2_1 _1609_ (.Y(_0719_),
    .A(_0709_),
    .B(_0718_));
 sg13g2_a21oi_1 _1610_ (.A1(_0709_),
    .A2(_0718_),
    .Y(_0720_),
    .B1(_0707_));
 sg13g2_a21o_1 _1611_ (.A2(_0720_),
    .A1(_0705_),
    .B1(_0703_),
    .X(_0721_));
 sg13g2_nand2_1 _1612_ (.Y(_0722_),
    .A(_0714_),
    .B(_0719_));
 sg13g2_a221oi_1 _1613_ (.B2(_0709_),
    .C1(_0712_),
    .B1(_0718_),
    .A1(_0705_),
    .Y(_0723_),
    .A2(_0713_));
 sg13g2_o21ai_1 _1614_ (.B1(_0712_),
    .Y(_0724_),
    .A1(_0709_),
    .A2(_0714_));
 sg13g2_nand2b_1 _1615_ (.Y(_0725_),
    .B(_0724_),
    .A_N(_0723_));
 sg13g2_nand3_1 _1616_ (.B(_0709_),
    .C(_0718_),
    .A(_0707_),
    .Y(_0726_));
 sg13g2_xnor2_1 _1617_ (.Y(_0727_),
    .A(_0055_),
    .B(_0061_));
 sg13g2_nor4_1 _1618_ (.A(_0701_),
    .B(_0704_),
    .C(_0720_),
    .D(_0727_),
    .Y(_0728_));
 sg13g2_a221oi_1 _1619_ (.B2(_0728_),
    .C1(_0725_),
    .B1(_0726_),
    .A1(_0721_),
    .Y(_0729_),
    .A2(_0722_));
 sg13g2_o21ai_1 _1620_ (.B1(_0718_),
    .Y(_0730_),
    .A1(_0716_),
    .A2(_0723_));
 sg13g2_inv_1 _1621_ (.Y(_0731_),
    .A(_0730_));
 sg13g2_nor2_1 _1622_ (.A(_0729_),
    .B(_0731_),
    .Y(_0732_));
 sg13g2_nor3_1 _1623_ (.A(_0011_),
    .B(_0729_),
    .C(_0731_),
    .Y(_0733_));
 sg13g2_xnor2_1 _1624_ (.Y(_0734_),
    .A(_0006_),
    .B(_0719_));
 sg13g2_nand2b_1 _1625_ (.Y(_0735_),
    .B(_0719_),
    .A_N(\pwm_generator_inst.counter[1] ));
 sg13g2_o21ai_1 _1626_ (.B1(_0735_),
    .Y(_0736_),
    .A1(_0733_),
    .A2(_0734_));
 sg13g2_xor2_1 _1627_ (.B(_0700_),
    .A(_0007_),
    .X(_0737_));
 sg13g2_nand2_1 _1628_ (.Y(_0738_),
    .A(_0008_),
    .B(_0665_));
 sg13g2_xnor2_1 _1629_ (.Y(_0739_),
    .A(_0010_),
    .B(_0642_));
 sg13g2_nor3_1 _1630_ (.A(_0002_),
    .B(_0571_),
    .C(_0586_),
    .Y(_0740_));
 sg13g2_a21oi_1 _1631_ (.A1(_0572_),
    .A2(_0587_),
    .Y(_0741_),
    .B1(_0053_));
 sg13g2_nor2_1 _1632_ (.A(\pwm_generator_inst.counter[11] ),
    .B(_0526_),
    .Y(_0742_));
 sg13g2_xnor2_1 _1633_ (.Y(_0743_),
    .A(\pwm_generator_inst.counter[11] ),
    .B(_0526_));
 sg13g2_xnor2_1 _1634_ (.Y(_0744_),
    .A(_0004_),
    .B(_0545_));
 sg13g2_nor2_1 _1635_ (.A(_0743_),
    .B(_0744_),
    .Y(_0745_));
 sg13g2_xnor2_1 _1636_ (.Y(_0746_),
    .A(_0003_),
    .B(_0568_));
 sg13g2_nand2_1 _1637_ (.Y(_0747_),
    .A(_0745_),
    .B(_0746_));
 sg13g2_nor3_2 _1638_ (.A(_0740_),
    .B(_0741_),
    .C(_0747_),
    .Y(_0748_));
 sg13g2_xnor2_1 _1639_ (.Y(_0749_),
    .A(\pwm_generator_inst.counter[7] ),
    .B(_0604_));
 sg13g2_xor2_1 _1640_ (.B(_0620_),
    .A(_0001_),
    .X(_0750_));
 sg13g2_nor2_1 _1641_ (.A(_0749_),
    .B(_0750_),
    .Y(_0751_));
 sg13g2_nand4_1 _1642_ (.B(_0739_),
    .C(_0748_),
    .A(_0738_),
    .Y(_0752_),
    .D(_0751_));
 sg13g2_a21oi_1 _1643_ (.A1(_0052_),
    .A2(_0664_),
    .Y(_0753_),
    .B1(_0752_));
 sg13g2_xnor2_1 _1644_ (.Y(_0754_),
    .A(\pwm_generator_inst.counter[3] ),
    .B(_0682_));
 sg13g2_and3_1 _1645_ (.X(_0755_),
    .A(_0737_),
    .B(_0753_),
    .C(_0754_));
 sg13g2_nand3b_1 _1646_ (.B(_0700_),
    .C(_0754_),
    .Y(_0756_),
    .A_N(\pwm_generator_inst.counter[2] ));
 sg13g2_o21ai_1 _1647_ (.B1(_0756_),
    .Y(_0757_),
    .A1(\pwm_generator_inst.counter[3] ),
    .A2(_0683_));
 sg13g2_nand3_1 _1648_ (.B(_0665_),
    .C(_0739_),
    .A(_0008_),
    .Y(_0758_));
 sg13g2_o21ai_1 _1649_ (.B1(_0758_),
    .Y(_0759_),
    .A1(\pwm_generator_inst.counter[5] ),
    .A2(_0642_));
 sg13g2_or3_1 _1650_ (.A(\pwm_generator_inst.counter[6] ),
    .B(_0620_),
    .C(_0749_),
    .X(_0760_));
 sg13g2_o21ai_1 _1651_ (.B1(_0760_),
    .Y(_0761_),
    .A1(\pwm_generator_inst.counter[7] ),
    .A2(_0604_));
 sg13g2_a21oi_1 _1652_ (.A1(_0751_),
    .A2(_0759_),
    .Y(_0762_),
    .B1(_0761_));
 sg13g2_nand2b_1 _1653_ (.Y(_0763_),
    .B(_0748_),
    .A_N(_0762_));
 sg13g2_nand2_1 _1654_ (.Y(_0764_),
    .A(_0741_),
    .B(_0746_));
 sg13g2_o21ai_1 _1655_ (.B1(_0764_),
    .Y(_0765_),
    .A1(\pwm_generator_inst.counter[9] ),
    .A2(_0568_));
 sg13g2_nor2_1 _1656_ (.A(\pwm_generator_inst.counter[10] ),
    .B(_0743_),
    .Y(_0766_));
 sg13g2_a221oi_1 _1657_ (.B2(_0545_),
    .C1(_0742_),
    .B1(_0766_),
    .A1(_0745_),
    .Y(_0767_),
    .A2(_0765_));
 sg13g2_nand2_1 _1658_ (.Y(_0768_),
    .A(_0763_),
    .B(_0767_));
 sg13g2_a221oi_1 _1659_ (.B2(_0753_),
    .C1(_0768_),
    .B1(_0757_),
    .A1(_0736_),
    .Y(_0769_),
    .A2(_0755_));
 sg13g2_nor2_1 _1660_ (.A(net74),
    .B(_0512_),
    .Y(_0770_));
 sg13g2_nor2b_1 _1661_ (.A(_0734_),
    .B_N(_0755_),
    .Y(_0771_));
 sg13g2_xor2_1 _1662_ (.B(_0732_),
    .A(\pwm_generator_inst.counter[0] ),
    .X(_0772_));
 sg13g2_a21o_1 _1663_ (.A2(_0772_),
    .A1(_0771_),
    .B1(_0770_),
    .X(_0773_));
 sg13g2_nand2_1 _1664_ (.Y(_0774_),
    .A(net74),
    .B(_0512_));
 sg13g2_o21ai_1 _1665_ (.B1(_0774_),
    .Y(_0000_),
    .A1(_0769_),
    .A2(_0773_));
 sg13g2_and2_1 _1666_ (.A(\pwm_generator_inst.pwm_out_s ),
    .B(net13),
    .X(\pwm_generator_inst.pwm_out ));
 sg13g2_nor2b_1 _1667_ (.A(net14),
    .B_N(net15),
    .Y(_0775_));
 sg13g2_o21ai_1 _1668_ (.B1(net233),
    .Y(_0776_),
    .A1(net225),
    .A2(net231));
 sg13g2_a21oi_1 _1669_ (.A1(_0050_),
    .A2(net231),
    .Y(_0012_),
    .B1(_0776_));
 sg13g2_o21ai_1 _1670_ (.B1(net233),
    .Y(_0777_),
    .A1(net222),
    .A2(net231));
 sg13g2_a21oi_1 _1671_ (.A1(_0049_),
    .A2(net231),
    .Y(_0013_),
    .B1(_0777_));
 sg13g2_o21ai_1 _1672_ (.B1(net233),
    .Y(_0778_),
    .A1(net220),
    .A2(net231));
 sg13g2_a21oi_1 _1673_ (.A1(_0048_),
    .A2(net231),
    .Y(_0014_),
    .B1(_0778_));
 sg13g2_o21ai_1 _1674_ (.B1(net232),
    .Y(_0779_),
    .A1(net214),
    .A2(net230));
 sg13g2_a21oi_1 _1675_ (.A1(_0047_),
    .A2(net230),
    .Y(_0015_),
    .B1(_0779_));
 sg13g2_o21ai_1 _1676_ (.B1(net232),
    .Y(_0780_),
    .A1(net210),
    .A2(net230));
 sg13g2_a21oi_1 _1677_ (.A1(_0046_),
    .A2(net230),
    .Y(_0016_),
    .B1(_0780_));
 sg13g2_o21ai_1 _1678_ (.B1(net232),
    .Y(_0781_),
    .A1(net208),
    .A2(net230));
 sg13g2_a21oi_1 _1679_ (.A1(_0045_),
    .A2(net230),
    .Y(_0017_),
    .B1(_0781_));
 sg13g2_o21ai_1 _1680_ (.B1(net234),
    .Y(_0782_),
    .A1(net205),
    .A2(net230));
 sg13g2_a21oi_1 _1681_ (.A1(_0044_),
    .A2(net230),
    .Y(_0018_),
    .B1(_0782_));
 sg13g2_nor3_1 _1682_ (.A(net199),
    .B(net200),
    .C(net202),
    .Y(_0783_));
 sg13g2_nor2b_1 _1683_ (.A(net196),
    .B_N(_0783_),
    .Y(_0784_));
 sg13g2_nor2_1 _1684_ (.A(net193),
    .B(net194),
    .Y(_0785_));
 sg13g2_and2_1 _1685_ (.A(_0784_),
    .B(_0785_),
    .X(_0786_));
 sg13g2_nor2b_1 _1686_ (.A(net191),
    .B_N(_0786_),
    .Y(_0787_));
 sg13g2_nor2b_1 _1687_ (.A(net189),
    .B_N(_0787_),
    .Y(_0788_));
 sg13g2_nand2b_1 _1688_ (.Y(_0789_),
    .B(_0788_),
    .A_N(net187));
 sg13g2_nor3_1 _1689_ (.A(net183),
    .B(net185),
    .C(_0789_),
    .Y(_0790_));
 sg13g2_o21ai_1 _1690_ (.B1(net183),
    .Y(_0791_),
    .A1(net185),
    .A2(_0789_));
 sg13g2_nand2b_1 _1691_ (.Y(_0792_),
    .B(_0791_),
    .A_N(_0790_));
 sg13g2_nand2b_1 _1692_ (.Y(_0793_),
    .B(\pwm_generator_inst.period_reg[11] ),
    .A_N(_0790_));
 sg13g2_or2_1 _1693_ (.X(_0794_),
    .B(_0793_),
    .A(\pwm_generator_inst.counter[11] ));
 sg13g2_nor2b_1 _1694_ (.A(\pwm_generator_inst.period_reg[11] ),
    .B_N(_0790_),
    .Y(_0795_));
 sg13g2_xnor2_1 _1695_ (.Y(_0796_),
    .A(net185),
    .B(_0789_));
 sg13g2_xnor2_1 _1696_ (.Y(_0797_),
    .A(_0003_),
    .B(_0796_));
 sg13g2_nor2_1 _1697_ (.A(_0795_),
    .B(_0797_),
    .Y(_0798_));
 sg13g2_xnor2_1 _1698_ (.Y(_0799_),
    .A(net187),
    .B(_0788_));
 sg13g2_xnor2_1 _1699_ (.Y(_0800_),
    .A(net191),
    .B(_0786_));
 sg13g2_xnor2_1 _1700_ (.Y(_0801_),
    .A(_0001_),
    .B(_0800_));
 sg13g2_o21ai_1 _1701_ (.B1(net198),
    .Y(_0802_),
    .A1(net200),
    .A2(net202));
 sg13g2_nand2b_1 _1702_ (.Y(_0803_),
    .B(_0802_),
    .A_N(_0783_));
 sg13g2_xor2_1 _1703_ (.B(_0010_),
    .A(net192),
    .X(_0804_));
 sg13g2_o21ai_1 _1704_ (.B1(_0804_),
    .Y(_0805_),
    .A1(_0009_),
    .A2(_0052_));
 sg13g2_xnor2_1 _1705_ (.Y(_0806_),
    .A(net200),
    .B(net202));
 sg13g2_a21oi_1 _1706_ (.A1(net202),
    .A2(\pwm_generator_inst.counter[0] ),
    .Y(_0807_),
    .B1(\pwm_generator_inst.counter[12] ));
 sg13g2_o21ai_1 _1707_ (.B1(_0807_),
    .Y(_0808_),
    .A1(net202),
    .A2(\pwm_generator_inst.counter[0] ));
 sg13g2_a22oi_1 _1708_ (.Y(_0809_),
    .B1(_0784_),
    .B2(_0804_),
    .A2(_0052_),
    .A1(_0009_));
 sg13g2_nand2_1 _1709_ (.Y(_0810_),
    .A(_0784_),
    .B(_0805_));
 sg13g2_mux2_1 _1710_ (.A0(_0810_),
    .A1(_0805_),
    .S(_0809_),
    .X(_0811_));
 sg13g2_inv_1 _1711_ (.Y(_0812_),
    .A(_0811_));
 sg13g2_xnor2_1 _1712_ (.Y(_0813_),
    .A(net196),
    .B(_0783_));
 sg13g2_xnor2_1 _1713_ (.Y(_0814_),
    .A(\pwm_generator_inst.counter[3] ),
    .B(_0813_));
 sg13g2_xnor2_1 _1714_ (.Y(_0815_),
    .A(_0006_),
    .B(_0806_));
 sg13g2_xnor2_1 _1715_ (.Y(_0816_),
    .A(_0007_),
    .B(_0803_));
 sg13g2_nor4_1 _1716_ (.A(_0808_),
    .B(_0814_),
    .C(_0815_),
    .D(_0816_),
    .Y(_0817_));
 sg13g2_xor2_1 _1717_ (.B(_0787_),
    .A(net189),
    .X(_0818_));
 sg13g2_xnor2_1 _1718_ (.Y(_0819_),
    .A(\pwm_generator_inst.counter[7] ),
    .B(_0818_));
 sg13g2_xnor2_1 _1719_ (.Y(_0820_),
    .A(_0004_),
    .B(_0792_));
 sg13g2_nand4_1 _1720_ (.B(_0812_),
    .C(_0817_),
    .A(_0801_),
    .Y(_0821_),
    .D(_0819_));
 sg13g2_a21oi_1 _1721_ (.A1(\pwm_generator_inst.counter[11] ),
    .A2(_0793_),
    .Y(_0822_),
    .B1(_0821_));
 sg13g2_xnor2_1 _1722_ (.Y(_0823_),
    .A(_0002_),
    .B(_0799_));
 sg13g2_nand4_1 _1723_ (.B(_0798_),
    .C(_0822_),
    .A(_0794_),
    .Y(_0824_),
    .D(_0823_));
 sg13g2_o21ai_1 _1724_ (.B1(net234),
    .Y(_0825_),
    .A1(_0820_),
    .A2(_0824_));
 sg13g2_nor3_1 _1725_ (.A(net218),
    .B(net222),
    .C(net224),
    .Y(_0826_));
 sg13g2_nor4_2 _1726_ (.A(net205),
    .B(net208),
    .C(\pwm_generator_inst.duty_reg[4] ),
    .Y(_0827_),
    .D(net213));
 sg13g2_a21oi_2 _1727_ (.B1(_0795_),
    .Y(_0828_),
    .A2(_0827_),
    .A1(_0826_));
 sg13g2_nand2b_1 _1728_ (.Y(_0829_),
    .B(\pwm_generator_inst.counter[0] ),
    .A_N(_0828_));
 sg13g2_nand2_1 _1729_ (.Y(_0830_),
    .A(net72),
    .B(_0828_));
 sg13g2_a21oi_1 _1730_ (.A1(_0829_),
    .A2(_0830_),
    .Y(_0019_),
    .B1(net180));
 sg13g2_and3_1 _1731_ (.X(_0831_),
    .A(net83),
    .B(\pwm_generator_inst.counter[0] ),
    .C(_0828_));
 sg13g2_a21oi_1 _1732_ (.A1(\pwm_generator_inst.counter[0] ),
    .A2(_0828_),
    .Y(_0832_),
    .B1(net83));
 sg13g2_nor3_1 _1733_ (.A(net180),
    .B(_0831_),
    .C(net84),
    .Y(_0020_));
 sg13g2_and2_1 _1734_ (.A(net90),
    .B(_0831_),
    .X(_0833_));
 sg13g2_nor2_1 _1735_ (.A(net90),
    .B(_0831_),
    .Y(_0834_));
 sg13g2_nor3_1 _1736_ (.A(net180),
    .B(_0833_),
    .C(net91),
    .Y(_0021_));
 sg13g2_nor2b_1 _1737_ (.A(net94),
    .B_N(_0831_),
    .Y(_0835_));
 sg13g2_xnor2_1 _1738_ (.Y(_0836_),
    .A(\pwm_generator_inst.counter[3] ),
    .B(_0835_));
 sg13g2_nor2_1 _1739_ (.A(net180),
    .B(net95),
    .Y(_0022_));
 sg13g2_a21oi_1 _1740_ (.A1(\pwm_generator_inst.counter[3] ),
    .A2(_0833_),
    .Y(_0837_),
    .B1(net75));
 sg13g2_and3_1 _1741_ (.X(_0838_),
    .A(net75),
    .B(\pwm_generator_inst.counter[3] ),
    .C(_0833_));
 sg13g2_nor3_1 _1742_ (.A(net180),
    .B(net76),
    .C(_0838_),
    .Y(_0023_));
 sg13g2_nand3_1 _1743_ (.B(_0052_),
    .C(_0833_),
    .A(\pwm_generator_inst.counter[3] ),
    .Y(_0839_));
 sg13g2_xor2_1 _1744_ (.B(_0839_),
    .A(net96),
    .X(_0840_));
 sg13g2_nor2_1 _1745_ (.A(net179),
    .B(net97),
    .Y(_0024_));
 sg13g2_a21oi_1 _1746_ (.A1(\pwm_generator_inst.counter[5] ),
    .A2(_0838_),
    .Y(_0841_),
    .B1(net80));
 sg13g2_and3_1 _1747_ (.X(_0842_),
    .A(net80),
    .B(\pwm_generator_inst.counter[5] ),
    .C(_0838_));
 sg13g2_nor3_1 _1748_ (.A(net179),
    .B(net81),
    .C(_0842_),
    .Y(_0025_));
 sg13g2_nand3b_1 _1749_ (.B(_0838_),
    .C(net96),
    .Y(_0843_),
    .A_N(_0001_));
 sg13g2_xor2_1 _1750_ (.B(_0843_),
    .A(net98),
    .X(_0844_));
 sg13g2_nor2_1 _1751_ (.A(net179),
    .B(net99),
    .Y(_0026_));
 sg13g2_and2_1 _1752_ (.A(\pwm_generator_inst.counter[7] ),
    .B(_0842_),
    .X(_0845_));
 sg13g2_nor2_1 _1753_ (.A(net88),
    .B(_0845_),
    .Y(_0846_));
 sg13g2_and2_1 _1754_ (.A(net88),
    .B(_0845_),
    .X(_0847_));
 sg13g2_nor3_1 _1755_ (.A(net179),
    .B(net89),
    .C(_0847_),
    .Y(_0027_));
 sg13g2_nor2b_1 _1756_ (.A(_0002_),
    .B_N(_0845_),
    .Y(_0848_));
 sg13g2_xnor2_1 _1757_ (.Y(_0849_),
    .A(net92),
    .B(_0848_));
 sg13g2_nor2_1 _1758_ (.A(net179),
    .B(net93),
    .Y(_0028_));
 sg13g2_a21oi_1 _1759_ (.A1(\pwm_generator_inst.counter[9] ),
    .A2(_0847_),
    .Y(_0850_),
    .B1(net85));
 sg13g2_and3_1 _1760_ (.X(_0851_),
    .A(net85),
    .B(\pwm_generator_inst.counter[9] ),
    .C(_0847_));
 sg13g2_nor3_1 _1761_ (.A(net179),
    .B(net86),
    .C(_0851_),
    .Y(_0029_));
 sg13g2_nand3b_1 _1762_ (.B(_0847_),
    .C(net92),
    .Y(_0852_),
    .A_N(_0004_));
 sg13g2_xor2_1 _1763_ (.B(_0852_),
    .A(net100),
    .X(_0853_));
 sg13g2_nor2_1 _1764_ (.A(net179),
    .B(net101),
    .Y(_0030_));
 sg13g2_and3_1 _1765_ (.X(_0854_),
    .A(net77),
    .B(\pwm_generator_inst.counter[11] ),
    .C(_0851_));
 sg13g2_a21oi_1 _1766_ (.A1(\pwm_generator_inst.counter[11] ),
    .A2(_0851_),
    .Y(_0855_),
    .B1(net77));
 sg13g2_nor3_1 _1767_ (.A(net179),
    .B(_0854_),
    .C(net78),
    .Y(_0031_));
 sg13g2_and2_1 _1768_ (.A(net15),
    .B(net14),
    .X(_0856_));
 sg13g2_o21ai_1 _1769_ (.B1(net233),
    .Y(_0857_),
    .A1(net203),
    .A2(net229));
 sg13g2_a21oi_1 _1770_ (.A1(_0050_),
    .A2(net228),
    .Y(_0032_),
    .B1(_0857_));
 sg13g2_o21ai_1 _1771_ (.B1(net232),
    .Y(_0858_),
    .A1(net201),
    .A2(net228));
 sg13g2_a21oi_1 _1772_ (.A1(_0049_),
    .A2(net228),
    .Y(_0033_),
    .B1(_0858_));
 sg13g2_o21ai_1 _1773_ (.B1(net232),
    .Y(_0859_),
    .A1(net198),
    .A2(net228));
 sg13g2_a21oi_1 _1774_ (.A1(_0048_),
    .A2(net229),
    .Y(_0034_),
    .B1(_0859_));
 sg13g2_o21ai_1 _1775_ (.B1(net232),
    .Y(_0860_),
    .A1(net196),
    .A2(net228));
 sg13g2_a21oi_1 _1776_ (.A1(_0047_),
    .A2(net229),
    .Y(_0035_),
    .B1(_0860_));
 sg13g2_o21ai_1 _1777_ (.B1(net232),
    .Y(_0861_),
    .A1(net195),
    .A2(net227));
 sg13g2_a21oi_1 _1778_ (.A1(_0046_),
    .A2(net228),
    .Y(_0036_),
    .B1(_0861_));
 sg13g2_o21ai_1 _1779_ (.B1(net232),
    .Y(_0862_),
    .A1(net193),
    .A2(net228));
 sg13g2_a21oi_1 _1780_ (.A1(_0045_),
    .A2(net228),
    .Y(_0037_),
    .B1(_0862_));
 sg13g2_o21ai_1 _1781_ (.B1(net234),
    .Y(_0863_),
    .A1(net191),
    .A2(net226));
 sg13g2_a21oi_1 _1782_ (.A1(_0044_),
    .A2(net227),
    .Y(_0038_),
    .B1(_0863_));
 sg13g2_o21ai_1 _1783_ (.B1(net234),
    .Y(_0864_),
    .A1(net189),
    .A2(net227));
 sg13g2_a21oi_1 _1784_ (.A1(_0873_),
    .A2(net227),
    .Y(_0039_),
    .B1(_0864_));
 sg13g2_o21ai_1 _1785_ (.B1(net234),
    .Y(_0866_),
    .A1(net187),
    .A2(net227));
 sg13g2_a21oi_1 _1786_ (.A1(_0872_),
    .A2(net226),
    .Y(_0040_),
    .B1(_0866_));
 sg13g2_o21ai_1 _1787_ (.B1(net234),
    .Y(_0867_),
    .A1(net185),
    .A2(net226));
 sg13g2_a21oi_1 _1788_ (.A1(_0871_),
    .A2(net226),
    .Y(_0041_),
    .B1(_0867_));
 sg13g2_o21ai_1 _1789_ (.B1(net234),
    .Y(_0868_),
    .A1(net183),
    .A2(net226));
 sg13g2_a21oi_1 _1790_ (.A1(_0870_),
    .A2(net226),
    .Y(_0042_),
    .B1(_0868_));
 sg13g2_o21ai_1 _1791_ (.B1(net234),
    .Y(_0869_),
    .A1(net181),
    .A2(net226));
 sg13g2_a21oi_1 _1792_ (.A1(_0865_),
    .A2(net226),
    .Y(_0043_),
    .B1(_0869_));
 sg13g2_dfrbp_1 _1793_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net45),
    .D(_0012_),
    .Q_N(_0894_),
    .Q(\pwm_generator_inst.duty_reg[0] ));
 sg13g2_dfrbp_1 _1794_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net59),
    .D(_0013_),
    .Q_N(_0893_),
    .Q(\pwm_generator_inst.duty_reg[1] ));
 sg13g2_dfrbp_1 _1795_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net57),
    .D(_0014_),
    .Q_N(_0892_),
    .Q(\pwm_generator_inst.duty_reg[2] ));
 sg13g2_dfrbp_1 _1796_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net55),
    .D(_0015_),
    .Q_N(_0891_),
    .Q(\pwm_generator_inst.duty_reg[3] ));
 sg13g2_dfrbp_1 _1797_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net53),
    .D(_0016_),
    .Q_N(_0890_),
    .Q(\pwm_generator_inst.duty_reg[4] ));
 sg13g2_dfrbp_1 _1798_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net51),
    .D(_0017_),
    .Q_N(_0889_),
    .Q(\pwm_generator_inst.duty_reg[5] ));
 sg13g2_dfrbp_1 _1799_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net60),
    .D(_0018_),
    .Q_N(_0895_),
    .Q(\pwm_generator_inst.duty_reg[6] ));
 sg13g2_dfrbp_1 _1800_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net49),
    .D(_0000_),
    .Q_N(_0888_),
    .Q(\pwm_generator_inst.pwm_out_s ));
 sg13g2_dfrbp_1 _1801_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net47),
    .D(net73),
    .Q_N(_0011_),
    .Q(\pwm_generator_inst.counter[0] ));
 sg13g2_dfrbp_1 _1802_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net44),
    .D(_0020_),
    .Q_N(_0006_),
    .Q(\pwm_generator_inst.counter[1] ));
 sg13g2_dfrbp_1 _1803_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net42),
    .D(_0021_),
    .Q_N(_0007_),
    .Q(\pwm_generator_inst.counter[2] ));
 sg13g2_dfrbp_1 _1804_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net40),
    .D(_0022_),
    .Q_N(_0887_),
    .Q(\pwm_generator_inst.counter[3] ));
 sg13g2_dfrbp_1 _1805_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net38),
    .D(_0023_),
    .Q_N(_0008_),
    .Q(\pwm_generator_inst.counter[4] ));
 sg13g2_dfrbp_1 _1806_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net69),
    .D(_0024_),
    .Q_N(_0010_),
    .Q(\pwm_generator_inst.counter[5] ));
 sg13g2_dfrbp_1 _1807_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net67),
    .D(net82),
    .Q_N(_0001_),
    .Q(\pwm_generator_inst.counter[6] ));
 sg13g2_dfrbp_1 _1808_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net65),
    .D(_0026_),
    .Q_N(_0886_),
    .Q(\pwm_generator_inst.counter[7] ));
 sg13g2_dfrbp_1 _1809_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net63),
    .D(_0027_),
    .Q_N(_0002_),
    .Q(\pwm_generator_inst.counter[8] ));
 sg13g2_dfrbp_1 _1810_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net61),
    .D(_0028_),
    .Q_N(_0003_),
    .Q(\pwm_generator_inst.counter[9] ));
 sg13g2_dfrbp_1 _1811_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net58),
    .D(net87),
    .Q_N(_0004_),
    .Q(\pwm_generator_inst.counter[10] ));
 sg13g2_dfrbp_1 _1812_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net54),
    .D(_0030_),
    .Q_N(_0885_),
    .Q(\pwm_generator_inst.counter[11] ));
 sg13g2_dfrbp_1 _1813_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net50),
    .D(net79),
    .Q_N(_0005_),
    .Q(\pwm_generator_inst.counter[12] ));
 sg13g2_dfrbp_1 _1814_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net46),
    .D(_0032_),
    .Q_N(_0884_),
    .Q(\pwm_generator_inst.period_reg[0] ));
 sg13g2_dfrbp_1 _1815_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net41),
    .D(_0033_),
    .Q_N(_0883_),
    .Q(\pwm_generator_inst.period_reg[1] ));
 sg13g2_dfrbp_1 _1816_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net70),
    .D(_0034_),
    .Q_N(_0882_),
    .Q(\pwm_generator_inst.period_reg[2] ));
 sg13g2_dfrbp_1 _1817_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net66),
    .D(_0035_),
    .Q_N(_0881_),
    .Q(\pwm_generator_inst.period_reg[3] ));
 sg13g2_dfrbp_1 _1818_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net62),
    .D(_0036_),
    .Q_N(_0009_),
    .Q(\pwm_generator_inst.period_reg[4] ));
 sg13g2_dfrbp_1 _1819_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net56),
    .D(_0037_),
    .Q_N(_0880_),
    .Q(\pwm_generator_inst.period_reg[5] ));
 sg13g2_dfrbp_1 _1820_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net48),
    .D(_0038_),
    .Q_N(_0879_),
    .Q(\pwm_generator_inst.period_reg[6] ));
 sg13g2_dfrbp_1 _1821_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net39),
    .D(_0039_),
    .Q_N(_0878_),
    .Q(\pwm_generator_inst.period_reg[7] ));
 sg13g2_dfrbp_1 _1822_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net64),
    .D(_0040_),
    .Q_N(_0877_),
    .Q(\pwm_generator_inst.period_reg[8] ));
 sg13g2_dfrbp_1 _1823_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net52),
    .D(_0041_),
    .Q_N(_0876_),
    .Q(\pwm_generator_inst.period_reg[9] ));
 sg13g2_dfrbp_1 _1824_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net68),
    .D(_0042_),
    .Q_N(_0875_),
    .Q(\pwm_generator_inst.period_reg[10] ));
 sg13g2_dfrbp_1 _1825_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net43),
    .D(_0043_),
    .Q_N(_0874_),
    .Q(\pwm_generator_inst.period_reg[11] ));
 sg13g2_tiehi _1821__39 (.L_HI(net39));
 sg13g2_tiehi _1804__40 (.L_HI(net40));
 sg13g2_tiehi _1815__41 (.L_HI(net41));
 sg13g2_tiehi _1803__42 (.L_HI(net42));
 sg13g2_tiehi _1825__43 (.L_HI(net43));
 sg13g2_tiehi _1802__44 (.L_HI(net44));
 sg13g2_tiehi _1793__45 (.L_HI(net45));
 sg13g2_tiehi _1814__46 (.L_HI(net46));
 sg13g2_tiehi _1801__47 (.L_HI(net47));
 sg13g2_tiehi _1820__48 (.L_HI(net48));
 sg13g2_tiehi _1800__49 (.L_HI(net49));
 sg13g2_tiehi _1813__50 (.L_HI(net50));
 sg13g2_tiehi _1798__51 (.L_HI(net51));
 sg13g2_tiehi _1823__52 (.L_HI(net52));
 sg13g2_tiehi _1797__53 (.L_HI(net53));
 sg13g2_tiehi _1812__54 (.L_HI(net54));
 sg13g2_tiehi _1796__55 (.L_HI(net55));
 sg13g2_tiehi _1819__56 (.L_HI(net56));
 sg13g2_tiehi _1795__57 (.L_HI(net57));
 sg13g2_tiehi _1811__58 (.L_HI(net58));
 sg13g2_tiehi _1794__59 (.L_HI(net59));
 sg13g2_tiehi _1799__60 (.L_HI(net60));
 sg13g2_tiehi _1810__61 (.L_HI(net61));
 sg13g2_tiehi _1818__62 (.L_HI(net62));
 sg13g2_tiehi _1809__63 (.L_HI(net63));
 sg13g2_tiehi _1822__64 (.L_HI(net64));
 sg13g2_tiehi _1808__65 (.L_HI(net65));
 sg13g2_tiehi _1817__66 (.L_HI(net66));
 sg13g2_tiehi _1807__67 (.L_HI(net67));
 sg13g2_tiehi _1824__68 (.L_HI(net68));
 sg13g2_tiehi _1806__69 (.L_HI(net69));
 sg13g2_tiehi _1816__70 (.L_HI(net70));
 sg13g2_tiehi tt_um_samuelm_pwm_generator_71 (.L_HI(net71));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_samuelm_pwm_generator_17 (.L_LO(net17));
 sg13g2_tielo tt_um_samuelm_pwm_generator_18 (.L_LO(net18));
 sg13g2_tielo tt_um_samuelm_pwm_generator_19 (.L_LO(net19));
 sg13g2_tielo tt_um_samuelm_pwm_generator_20 (.L_LO(net20));
 sg13g2_tielo tt_um_samuelm_pwm_generator_21 (.L_LO(net21));
 sg13g2_tielo tt_um_samuelm_pwm_generator_22 (.L_LO(net22));
 sg13g2_tielo tt_um_samuelm_pwm_generator_23 (.L_LO(net23));
 sg13g2_tielo tt_um_samuelm_pwm_generator_24 (.L_LO(net24));
 sg13g2_tielo tt_um_samuelm_pwm_generator_25 (.L_LO(net25));
 sg13g2_tielo tt_um_samuelm_pwm_generator_26 (.L_LO(net26));
 sg13g2_tielo tt_um_samuelm_pwm_generator_27 (.L_LO(net27));
 sg13g2_tielo tt_um_samuelm_pwm_generator_28 (.L_LO(net28));
 sg13g2_tielo tt_um_samuelm_pwm_generator_29 (.L_LO(net29));
 sg13g2_tielo tt_um_samuelm_pwm_generator_30 (.L_LO(net30));
 sg13g2_tielo tt_um_samuelm_pwm_generator_31 (.L_LO(net31));
 sg13g2_tielo tt_um_samuelm_pwm_generator_32 (.L_LO(net32));
 sg13g2_tielo tt_um_samuelm_pwm_generator_33 (.L_LO(net33));
 sg13g2_tielo tt_um_samuelm_pwm_generator_34 (.L_LO(net34));
 sg13g2_tielo tt_um_samuelm_pwm_generator_35 (.L_LO(net35));
 sg13g2_tielo tt_um_samuelm_pwm_generator_36 (.L_LO(net36));
 sg13g2_tielo tt_um_samuelm_pwm_generator_37 (.L_LO(net37));
 sg13g2_tiehi _1805__38 (.L_HI(net38));
 sg13g2_buf_2 _1882_ (.A(\pwm_generator_inst.pwm_out ),
    .X(uo_out[0]));
 sg13g2_buf_2 fanout179 (.A(_0825_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_0825_),
    .X(net180));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(net115));
 sg13g2_buf_2 fanout182 (.A(net183),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(net105),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(net185),
    .X(net184));
 sg13g2_buf_4 fanout185 (.X(net185),
    .A(net102));
 sg13g2_buf_2 fanout186 (.A(net187),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(net114),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(net189),
    .X(net188));
 sg13g2_buf_4 fanout189 (.X(net189),
    .A(net103));
 sg13g2_buf_4 fanout190 (.X(net190),
    .A(\pwm_generator_inst.period_reg[6] ));
 sg13g2_buf_2 fanout191 (.A(net113),
    .X(net191));
 sg13g2_buf_4 fanout192 (.X(net192),
    .A(\pwm_generator_inst.period_reg[5] ));
 sg13g2_buf_2 fanout193 (.A(net108),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(\pwm_generator_inst.period_reg[4] ),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(net107),
    .X(net195));
 sg13g2_buf_4 fanout196 (.X(net196),
    .A(net197));
 sg13g2_buf_2 fanout197 (.A(\pwm_generator_inst.period_reg[3] ),
    .X(net197));
 sg13g2_buf_4 fanout198 (.X(net198),
    .A(net199));
 sg13g2_buf_2 fanout199 (.A(\pwm_generator_inst.period_reg[2] ),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(net109),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(net203),
    .X(net202));
 sg13g2_buf_4 fanout203 (.X(net203),
    .A(net110));
 sg13g2_buf_2 fanout204 (.A(net206),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(net206),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(\pwm_generator_inst.duty_reg[6] ),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(net208),
    .X(net207));
 sg13g2_buf_4 fanout208 (.X(net208),
    .A(net111));
 sg13g2_buf_2 fanout209 (.A(net210),
    .X(net209));
 sg13g2_buf_4 fanout210 (.X(net210),
    .A(net112));
 sg13g2_buf_2 fanout211 (.A(net213),
    .X(net211));
 sg13g2_buf_1 fanout212 (.A(net213),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(\pwm_generator_inst.duty_reg[3] ),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(net215),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(\pwm_generator_inst.duty_reg[3] ),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(net217),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(net218),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(\pwm_generator_inst.duty_reg[2] ),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(net220),
    .X(net219));
 sg13g2_buf_1 fanout220 (.A(net221),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(\pwm_generator_inst.duty_reg[2] ),
    .X(net221));
 sg13g2_buf_4 fanout222 (.X(net222),
    .A(net106));
 sg13g2_buf_2 fanout223 (.A(\pwm_generator_inst.duty_reg[1] ),
    .X(net223));
 sg13g2_buf_4 fanout224 (.X(net224),
    .A(\pwm_generator_inst.duty_reg[0] ));
 sg13g2_buf_2 fanout225 (.A(net104),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(net227),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(net229),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(net229),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_0856_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_0775_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_0775_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(rst_n),
    .X(net232));
 sg13g2_buf_1 fanout233 (.A(rst_n),
    .X(net233));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[6]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[7]),
    .X(net15));
 sg13g2_tielo tt_um_samuelm_pwm_generator_16 (.L_LO(net16));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0011_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0019_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0005_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold4 (.A(\pwm_generator_inst.counter[4] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0837_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold6 (.A(\pwm_generator_inst.counter[12] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0855_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0031_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold9 (.A(\pwm_generator_inst.counter[6] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0841_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0025_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold12 (.A(\pwm_generator_inst.counter[1] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0832_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold14 (.A(\pwm_generator_inst.counter[10] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0850_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0029_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold17 (.A(\pwm_generator_inst.counter[8] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0846_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold19 (.A(\pwm_generator_inst.counter[2] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0834_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold21 (.A(\pwm_generator_inst.counter[9] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0849_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0007_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0836_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold25 (.A(\pwm_generator_inst.counter[5] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0840_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold27 (.A(\pwm_generator_inst.counter[7] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0844_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold29 (.A(\pwm_generator_inst.counter[11] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0853_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold31 (.A(\pwm_generator_inst.period_reg[9] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold32 (.A(\pwm_generator_inst.period_reg[7] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold33 (.A(\pwm_generator_inst.duty_reg[0] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold34 (.A(\pwm_generator_inst.period_reg[10] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold35 (.A(\pwm_generator_inst.duty_reg[1] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold36 (.A(\pwm_generator_inst.period_reg[4] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold37 (.A(\pwm_generator_inst.period_reg[5] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold38 (.A(\pwm_generator_inst.period_reg[1] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold39 (.A(\pwm_generator_inst.period_reg[0] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold40 (.A(\pwm_generator_inst.duty_reg[5] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold41 (.A(\pwm_generator_inst.duty_reg[4] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold42 (.A(\pwm_generator_inst.period_reg[6] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold43 (.A(\pwm_generator_inst.period_reg[8] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold44 (.A(\pwm_generator_inst.period_reg[11] ),
    .X(net115));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_fill_2 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_215 ();
 sg13g2_decap_8 FILLER_12_222 ();
 sg13g2_decap_4 FILLER_12_229 ();
 sg13g2_fill_2 FILLER_12_233 ();
 sg13g2_decap_8 FILLER_12_240 ();
 sg13g2_decap_8 FILLER_12_247 ();
 sg13g2_decap_8 FILLER_12_254 ();
 sg13g2_decap_8 FILLER_12_261 ();
 sg13g2_decap_8 FILLER_12_268 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_282 ();
 sg13g2_decap_8 FILLER_12_289 ();
 sg13g2_decap_8 FILLER_12_296 ();
 sg13g2_decap_4 FILLER_12_303 ();
 sg13g2_fill_1 FILLER_12_307 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_4 FILLER_13_140 ();
 sg13g2_fill_2 FILLER_13_144 ();
 sg13g2_decap_8 FILLER_13_151 ();
 sg13g2_decap_8 FILLER_13_158 ();
 sg13g2_fill_1 FILLER_13_165 ();
 sg13g2_decap_8 FILLER_13_174 ();
 sg13g2_decap_4 FILLER_13_181 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_4 FILLER_13_223 ();
 sg13g2_fill_1 FILLER_13_227 ();
 sg13g2_decap_4 FILLER_13_233 ();
 sg13g2_fill_2 FILLER_13_253 ();
 sg13g2_decap_8 FILLER_13_268 ();
 sg13g2_fill_2 FILLER_13_275 ();
 sg13g2_fill_2 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_319 ();
 sg13g2_fill_2 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_332 ();
 sg13g2_decap_8 FILLER_13_339 ();
 sg13g2_decap_8 FILLER_13_346 ();
 sg13g2_decap_8 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_367 ();
 sg13g2_decap_8 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_4 FILLER_14_138 ();
 sg13g2_fill_1 FILLER_14_142 ();
 sg13g2_fill_1 FILLER_14_172 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_decap_4 FILLER_14_198 ();
 sg13g2_fill_1 FILLER_14_202 ();
 sg13g2_fill_1 FILLER_14_218 ();
 sg13g2_fill_2 FILLER_14_227 ();
 sg13g2_fill_2 FILLER_14_239 ();
 sg13g2_fill_2 FILLER_14_274 ();
 sg13g2_fill_1 FILLER_14_276 ();
 sg13g2_fill_1 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_fill_1 FILLER_14_308 ();
 sg13g2_fill_1 FILLER_14_339 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_4 FILLER_15_112 ();
 sg13g2_fill_1 FILLER_15_116 ();
 sg13g2_decap_4 FILLER_15_145 ();
 sg13g2_fill_1 FILLER_15_167 ();
 sg13g2_decap_8 FILLER_15_176 ();
 sg13g2_fill_1 FILLER_15_195 ();
 sg13g2_decap_4 FILLER_15_222 ();
 sg13g2_fill_2 FILLER_15_226 ();
 sg13g2_fill_1 FILLER_15_237 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_4 FILLER_15_252 ();
 sg13g2_fill_1 FILLER_15_256 ();
 sg13g2_decap_4 FILLER_15_268 ();
 sg13g2_fill_2 FILLER_15_272 ();
 sg13g2_fill_1 FILLER_15_291 ();
 sg13g2_fill_2 FILLER_15_297 ();
 sg13g2_decap_8 FILLER_15_314 ();
 sg13g2_fill_1 FILLER_15_321 ();
 sg13g2_fill_1 FILLER_15_331 ();
 sg13g2_fill_2 FILLER_15_344 ();
 sg13g2_fill_1 FILLER_15_346 ();
 sg13g2_decap_4 FILLER_15_357 ();
 sg13g2_fill_1 FILLER_15_361 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_fill_1 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_143 ();
 sg13g2_fill_2 FILLER_16_150 ();
 sg13g2_fill_2 FILLER_16_162 ();
 sg13g2_fill_1 FILLER_16_164 ();
 sg13g2_decap_8 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_16_193 ();
 sg13g2_decap_4 FILLER_16_200 ();
 sg13g2_fill_2 FILLER_16_204 ();
 sg13g2_decap_4 FILLER_16_211 ();
 sg13g2_decap_4 FILLER_16_219 ();
 sg13g2_decap_4 FILLER_16_227 ();
 sg13g2_fill_1 FILLER_16_231 ();
 sg13g2_fill_2 FILLER_16_270 ();
 sg13g2_fill_1 FILLER_16_289 ();
 sg13g2_fill_2 FILLER_16_295 ();
 sg13g2_fill_2 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_4 FILLER_16_342 ();
 sg13g2_fill_1 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_fill_2 FILLER_17_98 ();
 sg13g2_fill_1 FILLER_17_100 ();
 sg13g2_decap_8 FILLER_17_114 ();
 sg13g2_fill_1 FILLER_17_121 ();
 sg13g2_decap_4 FILLER_17_137 ();
 sg13g2_fill_1 FILLER_17_141 ();
 sg13g2_fill_2 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_169 ();
 sg13g2_fill_2 FILLER_17_183 ();
 sg13g2_fill_1 FILLER_17_211 ();
 sg13g2_fill_2 FILLER_17_238 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_decap_4 FILLER_17_319 ();
 sg13g2_fill_2 FILLER_17_323 ();
 sg13g2_fill_1 FILLER_17_330 ();
 sg13g2_fill_2 FILLER_17_346 ();
 sg13g2_fill_1 FILLER_17_348 ();
 sg13g2_decap_4 FILLER_17_361 ();
 sg13g2_fill_2 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_fill_2 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_101 ();
 sg13g2_decap_8 FILLER_18_135 ();
 sg13g2_decap_4 FILLER_18_142 ();
 sg13g2_fill_2 FILLER_18_149 ();
 sg13g2_decap_4 FILLER_18_159 ();
 sg13g2_fill_2 FILLER_18_163 ();
 sg13g2_fill_1 FILLER_18_173 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_1 FILLER_18_207 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_fill_1 FILLER_18_279 ();
 sg13g2_fill_2 FILLER_18_324 ();
 sg13g2_fill_1 FILLER_18_326 ();
 sg13g2_decap_4 FILLER_18_339 ();
 sg13g2_fill_2 FILLER_18_343 ();
 sg13g2_fill_2 FILLER_18_362 ();
 sg13g2_fill_1 FILLER_18_364 ();
 sg13g2_fill_2 FILLER_18_389 ();
 sg13g2_fill_1 FILLER_18_391 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_4 FILLER_19_63 ();
 sg13g2_fill_2 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_81 ();
 sg13g2_fill_2 FILLER_19_88 ();
 sg13g2_fill_2 FILLER_19_167 ();
 sg13g2_fill_2 FILLER_19_198 ();
 sg13g2_fill_2 FILLER_19_208 ();
 sg13g2_fill_1 FILLER_19_210 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_fill_2 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_fill_2 FILLER_19_385 ();
 sg13g2_fill_1 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_4 FILLER_20_42 ();
 sg13g2_fill_2 FILLER_20_46 ();
 sg13g2_decap_4 FILLER_20_57 ();
 sg13g2_decap_4 FILLER_20_89 ();
 sg13g2_fill_2 FILLER_20_93 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_fill_1 FILLER_20_119 ();
 sg13g2_decap_4 FILLER_20_123 ();
 sg13g2_fill_2 FILLER_20_127 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_4 FILLER_20_147 ();
 sg13g2_fill_1 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_194 ();
 sg13g2_fill_1 FILLER_20_196 ();
 sg13g2_fill_1 FILLER_20_288 ();
 sg13g2_fill_2 FILLER_20_306 ();
 sg13g2_fill_2 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_341 ();
 sg13g2_fill_2 FILLER_20_348 ();
 sg13g2_decap_4 FILLER_20_355 ();
 sg13g2_fill_1 FILLER_20_362 ();
 sg13g2_decap_4 FILLER_20_373 ();
 sg13g2_fill_1 FILLER_20_377 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_2 FILLER_21_39 ();
 sg13g2_fill_2 FILLER_21_58 ();
 sg13g2_fill_1 FILLER_21_60 ();
 sg13g2_decap_4 FILLER_21_68 ();
 sg13g2_fill_2 FILLER_21_72 ();
 sg13g2_fill_2 FILLER_21_114 ();
 sg13g2_fill_1 FILLER_21_116 ();
 sg13g2_decap_4 FILLER_21_129 ();
 sg13g2_fill_1 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_fill_1 FILLER_21_150 ();
 sg13g2_decap_8 FILLER_21_155 ();
 sg13g2_fill_1 FILLER_21_183 ();
 sg13g2_fill_2 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_289 ();
 sg13g2_fill_1 FILLER_21_291 ();
 sg13g2_fill_2 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_303 ();
 sg13g2_decap_4 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_fill_1 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_48 ();
 sg13g2_decap_8 FILLER_22_71 ();
 sg13g2_fill_2 FILLER_22_87 ();
 sg13g2_decap_4 FILLER_22_92 ();
 sg13g2_fill_2 FILLER_22_96 ();
 sg13g2_decap_8 FILLER_22_103 ();
 sg13g2_decap_4 FILLER_22_110 ();
 sg13g2_fill_2 FILLER_22_114 ();
 sg13g2_fill_1 FILLER_22_129 ();
 sg13g2_fill_1 FILLER_22_139 ();
 sg13g2_fill_1 FILLER_22_214 ();
 sg13g2_fill_2 FILLER_22_266 ();
 sg13g2_fill_2 FILLER_22_278 ();
 sg13g2_fill_1 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_fill_2 FILLER_22_377 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_14 ();
 sg13g2_decap_4 FILLER_23_37 ();
 sg13g2_fill_2 FILLER_23_45 ();
 sg13g2_decap_4 FILLER_23_68 ();
 sg13g2_fill_2 FILLER_23_72 ();
 sg13g2_fill_2 FILLER_23_93 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_decap_4 FILLER_23_123 ();
 sg13g2_fill_2 FILLER_23_141 ();
 sg13g2_decap_4 FILLER_23_148 ();
 sg13g2_fill_1 FILLER_23_152 ();
 sg13g2_fill_2 FILLER_23_207 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_239 ();
 sg13g2_fill_2 FILLER_23_281 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_fill_1 FILLER_23_303 ();
 sg13g2_decap_4 FILLER_23_331 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_fill_2 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_11 ();
 sg13g2_decap_8 FILLER_24_31 ();
 sg13g2_fill_2 FILLER_24_38 ();
 sg13g2_fill_1 FILLER_24_40 ();
 sg13g2_fill_2 FILLER_24_64 ();
 sg13g2_fill_1 FILLER_24_66 ();
 sg13g2_decap_4 FILLER_24_77 ();
 sg13g2_fill_1 FILLER_24_93 ();
 sg13g2_fill_2 FILLER_24_97 ();
 sg13g2_fill_1 FILLER_24_99 ();
 sg13g2_decap_8 FILLER_24_104 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_1 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_172 ();
 sg13g2_fill_2 FILLER_24_187 ();
 sg13g2_fill_1 FILLER_24_194 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_decap_4 FILLER_24_207 ();
 sg13g2_fill_2 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_217 ();
 sg13g2_fill_2 FILLER_24_226 ();
 sg13g2_decap_4 FILLER_24_240 ();
 sg13g2_fill_2 FILLER_24_244 ();
 sg13g2_decap_4 FILLER_24_251 ();
 sg13g2_fill_1 FILLER_24_255 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_fill_2 FILLER_24_266 ();
 sg13g2_fill_1 FILLER_24_268 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_decap_4 FILLER_24_285 ();
 sg13g2_decap_4 FILLER_24_340 ();
 sg13g2_fill_2 FILLER_24_344 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_fill_2 FILLER_24_357 ();
 sg13g2_decap_4 FILLER_24_364 ();
 sg13g2_fill_1 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_fill_2 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_39 ();
 sg13g2_fill_1 FILLER_25_46 ();
 sg13g2_decap_8 FILLER_25_60 ();
 sg13g2_fill_1 FILLER_25_71 ();
 sg13g2_decap_8 FILLER_25_80 ();
 sg13g2_decap_4 FILLER_25_87 ();
 sg13g2_decap_4 FILLER_25_104 ();
 sg13g2_fill_2 FILLER_25_108 ();
 sg13g2_decap_4 FILLER_25_131 ();
 sg13g2_fill_1 FILLER_25_135 ();
 sg13g2_decap_8 FILLER_25_153 ();
 sg13g2_decap_4 FILLER_25_160 ();
 sg13g2_fill_2 FILLER_25_164 ();
 sg13g2_fill_2 FILLER_25_174 ();
 sg13g2_decap_4 FILLER_25_184 ();
 sg13g2_fill_1 FILLER_25_196 ();
 sg13g2_fill_2 FILLER_25_207 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_fill_2 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_264 ();
 sg13g2_fill_2 FILLER_25_271 ();
 sg13g2_fill_1 FILLER_25_273 ();
 sg13g2_fill_2 FILLER_25_285 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_4 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_decap_4 FILLER_25_340 ();
 sg13g2_fill_1 FILLER_25_344 ();
 sg13g2_fill_2 FILLER_25_350 ();
 sg13g2_fill_1 FILLER_25_352 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_decap_4 FILLER_25_385 ();
 sg13g2_fill_1 FILLER_25_389 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_34 ();
 sg13g2_fill_2 FILLER_26_38 ();
 sg13g2_decap_4 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_60 ();
 sg13g2_fill_2 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_106 ();
 sg13g2_decap_4 FILLER_26_113 ();
 sg13g2_fill_1 FILLER_26_117 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_fill_1 FILLER_26_133 ();
 sg13g2_fill_2 FILLER_26_139 ();
 sg13g2_decap_8 FILLER_26_153 ();
 sg13g2_decap_4 FILLER_26_177 ();
 sg13g2_fill_1 FILLER_26_181 ();
 sg13g2_decap_4 FILLER_26_197 ();
 sg13g2_fill_2 FILLER_26_201 ();
 sg13g2_decap_8 FILLER_26_220 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_246 ();
 sg13g2_fill_2 FILLER_26_253 ();
 sg13g2_decap_8 FILLER_26_281 ();
 sg13g2_decap_4 FILLER_26_288 ();
 sg13g2_fill_1 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_332 ();
 sg13g2_fill_2 FILLER_26_339 ();
 sg13g2_fill_1 FILLER_26_341 ();
 sg13g2_decap_4 FILLER_26_358 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_381 ();
 sg13g2_fill_2 FILLER_26_388 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_37 ();
 sg13g2_fill_2 FILLER_27_41 ();
 sg13g2_decap_4 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_67 ();
 sg13g2_decap_4 FILLER_27_74 ();
 sg13g2_fill_1 FILLER_27_78 ();
 sg13g2_decap_8 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_89 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_decap_4 FILLER_27_131 ();
 sg13g2_fill_1 FILLER_27_135 ();
 sg13g2_decap_4 FILLER_27_156 ();
 sg13g2_fill_2 FILLER_27_160 ();
 sg13g2_decap_8 FILLER_27_179 ();
 sg13g2_decap_8 FILLER_27_186 ();
 sg13g2_fill_2 FILLER_27_193 ();
 sg13g2_fill_1 FILLER_27_195 ();
 sg13g2_fill_2 FILLER_27_213 ();
 sg13g2_decap_4 FILLER_27_253 ();
 sg13g2_fill_1 FILLER_27_257 ();
 sg13g2_decap_4 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_284 ();
 sg13g2_fill_1 FILLER_27_291 ();
 sg13g2_fill_2 FILLER_27_296 ();
 sg13g2_decap_8 FILLER_27_303 ();
 sg13g2_decap_4 FILLER_27_310 ();
 sg13g2_fill_2 FILLER_27_314 ();
 sg13g2_decap_8 FILLER_27_328 ();
 sg13g2_fill_1 FILLER_27_335 ();
 sg13g2_decap_4 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_367 ();
 sg13g2_decap_4 FILLER_27_376 ();
 sg13g2_fill_1 FILLER_27_380 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_39 ();
 sg13g2_fill_1 FILLER_28_41 ();
 sg13g2_fill_2 FILLER_28_65 ();
 sg13g2_fill_2 FILLER_28_96 ();
 sg13g2_decap_8 FILLER_28_103 ();
 sg13g2_fill_2 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_125 ();
 sg13g2_fill_2 FILLER_28_131 ();
 sg13g2_fill_1 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_146 ();
 sg13g2_fill_1 FILLER_28_148 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_fill_2 FILLER_28_181 ();
 sg13g2_fill_1 FILLER_28_183 ();
 sg13g2_decap_8 FILLER_28_208 ();
 sg13g2_decap_4 FILLER_28_215 ();
 sg13g2_fill_2 FILLER_28_227 ();
 sg13g2_fill_2 FILLER_28_234 ();
 sg13g2_fill_1 FILLER_28_236 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_287 ();
 sg13g2_fill_1 FILLER_28_289 ();
 sg13g2_decap_4 FILLER_28_306 ();
 sg13g2_decap_8 FILLER_28_334 ();
 sg13g2_fill_1 FILLER_28_341 ();
 sg13g2_fill_2 FILLER_28_357 ();
 sg13g2_fill_1 FILLER_28_359 ();
 sg13g2_decap_4 FILLER_28_384 ();
 sg13g2_fill_1 FILLER_28_388 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_fill_2 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_31 ();
 sg13g2_fill_1 FILLER_29_33 ();
 sg13g2_fill_1 FILLER_29_39 ();
 sg13g2_fill_2 FILLER_29_44 ();
 sg13g2_decap_4 FILLER_29_51 ();
 sg13g2_fill_2 FILLER_29_55 ();
 sg13g2_fill_2 FILLER_29_65 ();
 sg13g2_fill_1 FILLER_29_67 ();
 sg13g2_fill_2 FILLER_29_80 ();
 sg13g2_fill_1 FILLER_29_94 ();
 sg13g2_fill_2 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_109 ();
 sg13g2_decap_4 FILLER_29_115 ();
 sg13g2_fill_1 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_125 ();
 sg13g2_fill_1 FILLER_29_127 ();
 sg13g2_decap_4 FILLER_29_140 ();
 sg13g2_fill_2 FILLER_29_156 ();
 sg13g2_fill_1 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_186 ();
 sg13g2_decap_4 FILLER_29_193 ();
 sg13g2_decap_8 FILLER_29_202 ();
 sg13g2_decap_4 FILLER_29_209 ();
 sg13g2_fill_1 FILLER_29_213 ();
 sg13g2_decap_8 FILLER_29_233 ();
 sg13g2_decap_8 FILLER_29_249 ();
 sg13g2_decap_4 FILLER_29_256 ();
 sg13g2_fill_1 FILLER_29_260 ();
 sg13g2_fill_2 FILLER_29_271 ();
 sg13g2_decap_8 FILLER_29_285 ();
 sg13g2_fill_2 FILLER_29_292 ();
 sg13g2_decap_4 FILLER_29_329 ();
 sg13g2_fill_2 FILLER_29_333 ();
 sg13g2_decap_4 FILLER_29_361 ();
 sg13g2_fill_1 FILLER_29_365 ();
 sg13g2_fill_2 FILLER_29_383 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_4 FILLER_30_52 ();
 sg13g2_decap_8 FILLER_30_64 ();
 sg13g2_fill_2 FILLER_30_71 ();
 sg13g2_fill_1 FILLER_30_73 ();
 sg13g2_fill_1 FILLER_30_78 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_fill_1 FILLER_30_117 ();
 sg13g2_decap_8 FILLER_30_130 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_fill_2 FILLER_30_161 ();
 sg13g2_fill_1 FILLER_30_163 ();
 sg13g2_fill_2 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_178 ();
 sg13g2_fill_1 FILLER_30_188 ();
 sg13g2_decap_8 FILLER_30_211 ();
 sg13g2_fill_2 FILLER_30_218 ();
 sg13g2_decap_4 FILLER_30_230 ();
 sg13g2_fill_1 FILLER_30_234 ();
 sg13g2_decap_4 FILLER_30_256 ();
 sg13g2_fill_2 FILLER_30_260 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_fill_2 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_325 ();
 sg13g2_decap_4 FILLER_30_332 ();
 sg13g2_fill_2 FILLER_30_336 ();
 sg13g2_fill_2 FILLER_30_354 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_fill_2 FILLER_30_402 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_4 FILLER_31_28 ();
 sg13g2_fill_1 FILLER_31_37 ();
 sg13g2_decap_8 FILLER_31_46 ();
 sg13g2_fill_2 FILLER_31_53 ();
 sg13g2_fill_2 FILLER_31_67 ();
 sg13g2_fill_2 FILLER_31_86 ();
 sg13g2_fill_1 FILLER_31_88 ();
 sg13g2_fill_2 FILLER_31_106 ();
 sg13g2_fill_1 FILLER_31_108 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_fill_1 FILLER_31_126 ();
 sg13g2_decap_4 FILLER_31_139 ();
 sg13g2_decap_8 FILLER_31_155 ();
 sg13g2_decap_4 FILLER_31_162 ();
 sg13g2_fill_1 FILLER_31_166 ();
 sg13g2_fill_2 FILLER_31_181 ();
 sg13g2_fill_1 FILLER_31_183 ();
 sg13g2_fill_2 FILLER_31_204 ();
 sg13g2_fill_1 FILLER_31_206 ();
 sg13g2_fill_2 FILLER_31_236 ();
 sg13g2_decap_8 FILLER_31_251 ();
 sg13g2_decap_4 FILLER_31_258 ();
 sg13g2_decap_4 FILLER_31_292 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_decap_4 FILLER_31_323 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_353 ();
 sg13g2_decap_4 FILLER_31_360 ();
 sg13g2_fill_2 FILLER_31_370 ();
 sg13g2_fill_1 FILLER_31_380 ();
 sg13g2_fill_1 FILLER_31_397 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_4 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_46 ();
 sg13g2_fill_1 FILLER_32_64 ();
 sg13g2_fill_2 FILLER_32_88 ();
 sg13g2_fill_2 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_108 ();
 sg13g2_decap_4 FILLER_32_121 ();
 sg13g2_fill_2 FILLER_32_125 ();
 sg13g2_decap_8 FILLER_32_135 ();
 sg13g2_fill_1 FILLER_32_142 ();
 sg13g2_fill_2 FILLER_32_148 ();
 sg13g2_fill_1 FILLER_32_150 ();
 sg13g2_fill_2 FILLER_32_198 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_fill_1 FILLER_32_218 ();
 sg13g2_decap_4 FILLER_32_224 ();
 sg13g2_fill_1 FILLER_32_228 ();
 sg13g2_fill_1 FILLER_32_254 ();
 sg13g2_decap_8 FILLER_32_260 ();
 sg13g2_fill_1 FILLER_32_267 ();
 sg13g2_decap_4 FILLER_32_273 ();
 sg13g2_fill_2 FILLER_32_296 ();
 sg13g2_fill_1 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_318 ();
 sg13g2_decap_8 FILLER_32_325 ();
 sg13g2_decap_4 FILLER_32_332 ();
 sg13g2_fill_2 FILLER_32_336 ();
 sg13g2_fill_2 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_346 ();
 sg13g2_decap_4 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_decap_4 FILLER_32_372 ();
 sg13g2_fill_2 FILLER_32_376 ();
 sg13g2_decap_4 FILLER_32_383 ();
 sg13g2_fill_1 FILLER_32_387 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_fill_2 FILLER_33_49 ();
 sg13g2_fill_1 FILLER_33_51 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_4 FILLER_33_70 ();
 sg13g2_fill_1 FILLER_33_74 ();
 sg13g2_decap_8 FILLER_33_80 ();
 sg13g2_decap_8 FILLER_33_87 ();
 sg13g2_fill_1 FILLER_33_94 ();
 sg13g2_decap_4 FILLER_33_107 ();
 sg13g2_fill_1 FILLER_33_141 ();
 sg13g2_fill_1 FILLER_33_154 ();
 sg13g2_decap_4 FILLER_33_160 ();
 sg13g2_decap_8 FILLER_33_169 ();
 sg13g2_decap_8 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_183 ();
 sg13g2_fill_1 FILLER_33_198 ();
 sg13g2_decap_8 FILLER_33_227 ();
 sg13g2_decap_8 FILLER_33_251 ();
 sg13g2_fill_2 FILLER_33_258 ();
 sg13g2_decap_4 FILLER_33_280 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_fill_2 FILLER_33_308 ();
 sg13g2_fill_2 FILLER_33_351 ();
 sg13g2_fill_2 FILLER_33_358 ();
 sg13g2_fill_1 FILLER_33_360 ();
 sg13g2_fill_2 FILLER_33_374 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_124 ();
 sg13g2_decap_8 FILLER_34_131 ();
 sg13g2_fill_2 FILLER_34_138 ();
 sg13g2_decap_8 FILLER_34_149 ();
 sg13g2_fill_1 FILLER_34_156 ();
 sg13g2_decap_8 FILLER_34_186 ();
 sg13g2_fill_2 FILLER_34_193 ();
 sg13g2_fill_1 FILLER_34_195 ();
 sg13g2_fill_2 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_272 ();
 sg13g2_fill_2 FILLER_34_299 ();
 sg13g2_fill_1 FILLER_34_316 ();
 sg13g2_fill_2 FILLER_34_320 ();
 sg13g2_fill_1 FILLER_34_322 ();
 sg13g2_fill_2 FILLER_34_350 ();
 sg13g2_fill_1 FILLER_34_352 ();
 sg13g2_fill_2 FILLER_34_358 ();
 sg13g2_fill_1 FILLER_34_368 ();
 sg13g2_fill_1 FILLER_34_374 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_fill_2 FILLER_35_161 ();
 sg13g2_fill_2 FILLER_35_168 ();
 sg13g2_fill_1 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_4 FILLER_35_182 ();
 sg13g2_fill_2 FILLER_35_186 ();
 sg13g2_fill_2 FILLER_35_257 ();
 sg13g2_fill_1 FILLER_35_259 ();
 sg13g2_fill_2 FILLER_35_274 ();
 sg13g2_decap_4 FILLER_35_284 ();
 sg13g2_fill_1 FILLER_35_288 ();
 sg13g2_fill_1 FILLER_35_294 ();
 sg13g2_decap_4 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_154 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_decap_4 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_205 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_4 FILLER_36_217 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_231 ();
 sg13g2_decap_4 FILLER_36_237 ();
 sg13g2_fill_2 FILLER_36_241 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_decap_4 FILLER_36_273 ();
 sg13g2_fill_2 FILLER_36_325 ();
 sg13g2_fill_2 FILLER_36_336 ();
 sg13g2_fill_1 FILLER_36_338 ();
 sg13g2_fill_2 FILLER_36_343 ();
 sg13g2_fill_1 FILLER_36_345 ();
 sg13g2_fill_2 FILLER_36_360 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_fill_1 FILLER_37_211 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_fill_2 FILLER_37_224 ();
 sg13g2_fill_2 FILLER_37_366 ();
 sg13g2_fill_1 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_decap_4 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_240 ();
 sg13g2_fill_1 FILLER_38_249 ();
 sg13g2_fill_2 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_344 ();
 sg13g2_fill_1 FILLER_38_346 ();
 sg13g2_fill_2 FILLER_38_352 ();
 sg13g2_fill_2 FILLER_38_380 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net16;
 assign uio_oe[1] = net17;
 assign uio_oe[2] = net18;
 assign uio_oe[3] = net19;
 assign uio_oe[4] = net71;
 assign uio_oe[5] = net20;
 assign uio_oe[6] = net21;
 assign uio_oe[7] = net22;
 assign uio_out[0] = net23;
 assign uio_out[1] = net24;
 assign uio_out[2] = net25;
 assign uio_out[3] = net26;
 assign uio_out[4] = net27;
 assign uio_out[5] = net28;
 assign uio_out[6] = net29;
 assign uio_out[7] = net30;
 assign uo_out[1] = net31;
 assign uo_out[2] = net32;
 assign uo_out[3] = net33;
 assign uo_out[4] = net34;
 assign uo_out[5] = net35;
 assign uo_out[6] = net36;
 assign uo_out[7] = net37;
endmodule

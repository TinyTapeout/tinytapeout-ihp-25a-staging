module tt_um_gfcwfzkm_scope_bfh_mht1_3 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire \champlitude[0] ;
 wire \champlitude[1] ;
 wire \champlitude[2] ;
 wire \choffset[0] ;
 wire \choffset[1] ;
 wire \choffset[2] ;
 wire \choffset[3] ;
 wire \choffset[4] ;
 wire \display_x[0] ;
 wire \display_x[1] ;
 wire \display_x[2] ;
 wire \display_x[3] ;
 wire \display_x[4] ;
 wire \display_x[5] ;
 wire \display_x[6] ;
 wire \display_x[7] ;
 wire \display_x[8] ;
 wire \display_x[9] ;
 wire \dsgfreqshift[0] ;
 wire \dsgfreqshift[1] ;
 wire \lastsample[0] ;
 wire \lastsample[1] ;
 wire \lastsample[2] ;
 wire \lastsample[3] ;
 wire \lastsample[4] ;
 wire \lastsample[5] ;
 wire \lastsample[6] ;
 wire \lastsample[7] ;
 wire \measurements.adc_cs ;
 wire \measurements.adc_sclk ;
 wire \measurements.address_counter_reg[0] ;
 wire \measurements.address_counter_reg[10] ;
 wire \measurements.address_counter_reg[11] ;
 wire \measurements.address_counter_reg[12] ;
 wire \measurements.address_counter_reg[13] ;
 wire \measurements.address_counter_reg[14] ;
 wire \measurements.address_counter_reg[1] ;
 wire \measurements.address_counter_reg[2] ;
 wire \measurements.address_counter_reg[3] ;
 wire \measurements.address_counter_reg[4] ;
 wire \measurements.address_counter_reg[5] ;
 wire \measurements.address_counter_reg[6] ;
 wire \measurements.address_counter_reg[7] ;
 wire \measurements.address_counter_reg[8] ;
 wire \measurements.address_counter_reg[9] ;
 wire \measurements.alreadytriggered_reg ;
 wire \measurements.enough_samples_in_fram_reg ;
 wire \measurements.fram_cs ;
 wire \measurements.fram_mosi ;
 wire \measurements.fram_sclk ;
 wire \measurements.memoryShift[0] ;
 wire \measurements.memoryShift[1] ;
 wire \measurements.memoryShift[2] ;
 wire \measurements.memoryShift[3] ;
 wire \measurements.memoryShift[4] ;
 wire \measurements.memoryShift[5] ;
 wire \measurements.memoryShift[6] ;
 wire \measurements.memoryShift[7] ;
 wire \measurements.memoryShift[8] ;
 wire \measurements.n163_o[0] ;
 wire \measurements.n163_o[1] ;
 wire \measurements.n163_o[2] ;
 wire \measurements.n175_o[0] ;
 wire \measurements.n175_o[1] ;
 wire \measurements.n175_o[2] ;
 wire \measurements.n175_o[3] ;
 wire \measurements.n175_o[4] ;
 wire \measurements.n175_o[5] ;
 wire \measurements.n182_o ;
 wire \measurements.n200_o[0] ;
 wire \measurements.n200_o[1] ;
 wire \measurements.n200_o[2] ;
 wire \measurements.n244_o[0] ;
 wire \measurements.n244_o[1] ;
 wire \measurements.n244_o[2] ;
 wire \measurements.n244_o[3] ;
 wire \measurements.n246_q[0] ;
 wire \measurements.n246_q[10] ;
 wire \measurements.n246_q[11] ;
 wire \measurements.n246_q[12] ;
 wire \measurements.n246_q[13] ;
 wire \measurements.n246_q[14] ;
 wire \measurements.n246_q[1] ;
 wire \measurements.n246_q[2] ;
 wire \measurements.n246_q[3] ;
 wire \measurements.n246_q[4] ;
 wire \measurements.n246_q[5] ;
 wire \measurements.n246_q[6] ;
 wire \measurements.n246_q[7] ;
 wire \measurements.n246_q[8] ;
 wire \measurements.n246_q[9] ;
 wire \measurements.n249_q[0] ;
 wire \measurements.n249_q[1] ;
 wire \measurements.n249_q[2] ;
 wire \measurements.n249_q[3] ;
 wire \measurements.n249_q[4] ;
 wire \measurements.n249_q[5] ;
 wire \measurements.n250_q[0] ;
 wire \measurements.n250_q[1] ;
 wire \measurements.n250_q[2] ;
 wire \measurements.n250_q[3] ;
 wire \measurements.n253_q ;
 wire \measurements.n98_o[0] ;
 wire \measurements.n98_o[1] ;
 wire \measurements.n98_o[2] ;
 wire \measurements.n98_o[3] ;
 wire \measurements.samples_adc.cnt_reg[0] ;
 wire \measurements.samples_adc.cnt_reg[1] ;
 wire \measurements.samples_adc.cnt_reg[2] ;
 wire \measurements.samples_adc.cnt_reg[3] ;
 wire \measurements.samples_adc.n84_q[0] ;
 wire \measurements.samples_adc.n84_q[1] ;
 wire \measurements.samples_storage.n101_o ;
 wire \measurements.samples_storage.n170_o ;
 wire \measurements.samples_storage.n230_q[0] ;
 wire \measurements.samples_storage.n230_q[1] ;
 wire \measurements.samples_storage.n230_q[2] ;
 wire \measurements.samples_storage.n230_q[3] ;
 wire \measurements.samples_storage.n232_q ;
 wire \measurements.samples_storage.spi_master_inst.n100_q[0] ;
 wire \measurements.samples_storage.spi_master_inst.n100_q[1] ;
 wire \measurements.samples_storage.spi_master_inst.n103_q[1] ;
 wire \measurements.samples_storage.spi_master_inst.n103_q[2] ;
 wire \measurements.samples_storage.spi_master_inst.n103_q[3] ;
 wire \measurements.samples_storage.spi_master_inst.n18_o ;
 wire \measurements.samples_storage.spi_master_inst.n20_o ;
 wire \measurements.samples_storage.spi_master_inst.n22_o ;
 wire \measurements.samples_storage.spi_master_inst.n24_o ;
 wire \measurements.samples_storage.spi_master_inst.n26_o ;
 wire \measurements.samples_storage.spi_master_inst.n28_o ;
 wire \measurements.samples_storage.spi_master_inst.n30_o ;
 wire \measurements.samples_storage.spi_master_inst.n96_o ;
 wire \measurements.trigger.sample_on_rising_edge ;
 wire \measurements.trigger.trigger_threshold[0] ;
 wire \measurements.trigger.trigger_threshold[1] ;
 wire \measurements.trigger.trigger_threshold[2] ;
 wire \measurements.trigger.trigger_threshold[3] ;
 wire \oscilloscope_control.button_debouncer_n1_debounce_buttons.counter_next[0] ;
 wire \oscilloscope_control.button_debouncer_n1_debounce_buttons.counter_reg[0] ;
 wire \oscilloscope_control.button_debouncer_n1_debounce_buttons.counter_reg[1] ;
 wire \oscilloscope_control.button_debouncer_n1_debounce_buttons.counter_reg[2] ;
 wire \oscilloscope_control.button_debouncer_n1_debounce_buttons.debounced ;
 wire \oscilloscope_control.button_debouncer_n1_debounce_buttons.in_raw ;
 wire \oscilloscope_control.button_debouncer_n2_debounce_buttons.counter_next[0] ;
 wire \oscilloscope_control.button_debouncer_n2_debounce_buttons.counter_reg[0] ;
 wire \oscilloscope_control.button_debouncer_n2_debounce_buttons.counter_reg[1] ;
 wire \oscilloscope_control.button_debouncer_n2_debounce_buttons.counter_reg[2] ;
 wire \oscilloscope_control.button_debouncer_n2_debounce_buttons.debounced ;
 wire \oscilloscope_control.button_debouncer_n2_debounce_buttons.in_raw ;
 wire \oscilloscope_control.button_debouncer_n3_debounce_buttons.counter_next[0] ;
 wire \oscilloscope_control.button_debouncer_n3_debounce_buttons.counter_reg[0] ;
 wire \oscilloscope_control.button_debouncer_n3_debounce_buttons.counter_reg[1] ;
 wire \oscilloscope_control.button_debouncer_n3_debounce_buttons.counter_reg[2] ;
 wire \oscilloscope_control.button_debouncer_n3_debounce_buttons.debounced ;
 wire \oscilloscope_control.button_debouncer_n3_debounce_buttons.in_raw ;
 wire \oscilloscope_control.button_debouncer_n4_debounce_buttons.counter_next[0] ;
 wire \oscilloscope_control.button_debouncer_n4_debounce_buttons.counter_reg[0] ;
 wire \oscilloscope_control.button_debouncer_n4_debounce_buttons.counter_reg[1] ;
 wire \oscilloscope_control.button_debouncer_n4_debounce_buttons.counter_reg[2] ;
 wire \oscilloscope_control.button_debouncer_n4_debounce_buttons.debounced ;
 wire \oscilloscope_control.button_debouncer_n4_debounce_buttons.in_raw ;
 wire \oscilloscope_control.button_ff_stage_1_reg[0] ;
 wire \oscilloscope_control.button_ff_stage_1_reg[1] ;
 wire \oscilloscope_control.button_ff_stage_1_reg[2] ;
 wire \oscilloscope_control.button_ff_stage_1_reg[3] ;
 wire \oscilloscope_control.n111_o[0] ;
 wire \oscilloscope_control.n114_o[0] ;
 wire \oscilloscope_control.n146_o[0] ;
 wire \oscilloscope_control.n171_o[0] ;
 wire \oscilloscope_control.n206_o ;
 wire \oscilloscope_control.n208_o ;
 wire \oscilloscope_control.n220_q[0] ;
 wire \oscilloscope_control.n220_q[1] ;
 wire \oscilloscope_control.n223_q[0] ;
 wire \oscilloscope_control.n223_q[1] ;
 wire \oscilloscope_control.switch_debouncer_n1_debounce_switches.counter_next[0] ;
 wire \oscilloscope_control.switch_debouncer_n1_debounce_switches.counter_reg[0] ;
 wire \oscilloscope_control.switch_debouncer_n1_debounce_switches.counter_reg[1] ;
 wire \oscilloscope_control.switch_debouncer_n1_debounce_switches.counter_reg[2] ;
 wire \oscilloscope_control.switch_debouncer_n1_debounce_switches.debounced ;
 wire \oscilloscope_control.switch_debouncer_n2_debounce_switches.counter_next[0] ;
 wire \oscilloscope_control.switch_debouncer_n2_debounce_switches.counter_reg[0] ;
 wire \oscilloscope_control.switch_debouncer_n2_debounce_switches.counter_reg[1] ;
 wire \oscilloscope_control.switch_debouncer_n2_debounce_switches.counter_reg[2] ;
 wire \oscilloscope_control.switch_debouncer_n2_debounce_switches.debounced ;
 wire \settings_uart_printer.n103_q[0] ;
 wire \settings_uart_printer.n103_q[1] ;
 wire \settings_uart_printer.n103_q[2] ;
 wire \settings_uart_printer.n103_q[3] ;
 wire \settings_uart_printer.n103_q[4] ;
 wire \settings_uart_printer.n103_q[5] ;
 wire \settings_uart_printer.n104_q[0] ;
 wire \settings_uart_printer.n104_q[1] ;
 wire \settings_uart_printer.tx ;
 wire \settings_uart_printer.uart_tx_module.counter_reg[0] ;
 wire \settings_uart_printer.uart_tx_module.counter_reg[10] ;
 wire \settings_uart_printer.uart_tx_module.counter_reg[11] ;
 wire \settings_uart_printer.uart_tx_module.counter_reg[1] ;
 wire \settings_uart_printer.uart_tx_module.counter_reg[2] ;
 wire \settings_uart_printer.uart_tx_module.counter_reg[3] ;
 wire \settings_uart_printer.uart_tx_module.counter_reg[4] ;
 wire \settings_uart_printer.uart_tx_module.counter_reg[5] ;
 wire \settings_uart_printer.uart_tx_module.counter_reg[6] ;
 wire \settings_uart_printer.uart_tx_module.counter_reg[7] ;
 wire \settings_uart_printer.uart_tx_module.counter_reg[8] ;
 wire \settings_uart_printer.uart_tx_module.counter_reg[9] ;
 wire \settings_uart_printer.uart_tx_module.data_reg[0] ;
 wire \settings_uart_printer.uart_tx_module.data_reg[1] ;
 wire \settings_uart_printer.uart_tx_module.data_reg[2] ;
 wire \settings_uart_printer.uart_tx_module.data_reg[3] ;
 wire \settings_uart_printer.uart_tx_module.data_reg[4] ;
 wire \settings_uart_printer.uart_tx_module.data_reg[5] ;
 wire \settings_uart_printer.uart_tx_module.data_reg[6] ;
 wire \settings_uart_printer.uart_tx_module.datacnt_reg[0] ;
 wire \settings_uart_printer.uart_tx_module.datacnt_reg[1] ;
 wire \settings_uart_printer.uart_tx_module.datacnt_reg[2] ;
 wire \settings_uart_printer.uart_tx_module.n88_q[0] ;
 wire \settings_uart_printer.uart_tx_module.n88_q[1] ;
 wire \siggen.da_cs ;
 wire \siggen.da_mosi ;
 wire \siggen.da_sclk ;
 wire \siggen.dac_pmod.cnt_reg[0] ;
 wire \siggen.dac_pmod.cnt_reg[1] ;
 wire \siggen.dac_pmod.cnt_reg[2] ;
 wire \siggen.dac_pmod.cnt_reg[3] ;
 wire \siggen.dac_pmod.n50_o[0] ;
 wire \siggen.dac_pmod.n50_o[1] ;
 wire \siggen.dac_pmod.n50_o[2] ;
 wire \siggen.dac_pmod.n50_o[3] ;
 wire \siggen.dac_pmod.n50_o[4] ;
 wire \siggen.dac_pmod.n50_o[5] ;
 wire \siggen.dac_pmod.n50_o[6] ;
 wire \siggen.dac_pmod.n66_o ;
 wire \siggen.dac_pmod.n85_q[0] ;
 wire \siggen.dac_pmod.n85_q[1] ;
 wire \siggen.dac_pmod.n88_q ;
 wire \siggen.n20_o ;
 wire \siggen.n22_o ;
 wire \siggen.n49_o[3] ;
 wire \siggen.n49_o[4] ;
 wire \siggen.n49_o[5] ;
 wire \siggen.n49_o[6] ;
 wire \siggen.n49_o[7] ;
 wire \siggen.n66_q[0] ;
 wire \siggen.n66_q[1] ;
 wire \siggen.n66_q[2] ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire \videogen.b ;
 wire \videogen.de ;
 wire \videogen.draw_y[0] ;
 wire \videogen.draw_y[1] ;
 wire \videogen.draw_y[2] ;
 wire \videogen.draw_y[3] ;
 wire \videogen.draw_y[4] ;
 wire \videogen.draw_y[5] ;
 wire \videogen.draw_y[6] ;
 wire \videogen.draw_y[7] ;
 wire \videogen.draw_y[8] ;
 wire \videogen.draw_y[9] ;
 wire \videogen.g ;
 wire \videogen.hsync ;
 wire \videogen.r ;
 wire \videogen.video_timing_generator.hdmi_vsync ;
 wire \videogen.video_timing_generator.n21_o[0] ;
 wire \videogen.video_timing_generator.n21_o[1] ;
 wire \videogen.video_timing_generator.n21_o[2] ;
 wire \videogen.video_timing_generator.n21_o[3] ;
 wire \videogen.video_timing_generator.n21_o[4] ;
 wire \videogen.video_timing_generator.n21_o[5] ;
 wire \videogen.video_timing_generator.n21_o[6] ;
 wire \videogen.video_timing_generator.n21_o[7] ;
 wire \videogen.video_timing_generator.n21_o[8] ;
 wire \videogen.video_timing_generator.n21_o[9] ;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;

 sg13g2_inv_1 _2514_ (.Y(_1974_),
    .A(net128));
 sg13g2_inv_1 _2515_ (.Y(_1975_),
    .A(net95));
 sg13g2_inv_1 _2516_ (.Y(_1976_),
    .A(net140));
 sg13g2_inv_1 _2517_ (.Y(_1977_),
    .A(net730));
 sg13g2_inv_2 _2518_ (.Y(_1978_),
    .A(net975));
 sg13g2_inv_1 _2519_ (.Y(_1979_),
    .A(net620));
 sg13g2_inv_2 _2520_ (.Y(_1980_),
    .A(net576));
 sg13g2_inv_1 _2521_ (.Y(_1981_),
    .A(net579));
 sg13g2_inv_1 _2522_ (.Y(_1982_),
    .A(net497));
 sg13g2_inv_1 _2523_ (.Y(_1983_),
    .A(net347));
 sg13g2_inv_1 _2524_ (.Y(_1984_),
    .A(net117));
 sg13g2_inv_2 _2525_ (.Y(_1985_),
    .A(net479));
 sg13g2_inv_2 _2526_ (.Y(_1986_),
    .A(net991));
 sg13g2_inv_2 _2527_ (.Y(_1987_),
    .A(net534));
 sg13g2_inv_1 _2528_ (.Y(_1988_),
    .A(net894));
 sg13g2_inv_2 _2529_ (.Y(_1989_),
    .A(net410));
 sg13g2_inv_1 _2530_ (.Y(_1990_),
    .A(net378));
 sg13g2_inv_1 _2531_ (.Y(_1991_),
    .A(net328));
 sg13g2_inv_1 _2532_ (.Y(_1992_),
    .A(net588));
 sg13g2_inv_4 _2533_ (.A(net397),
    .Y(_1993_));
 sg13g2_inv_1 _2534_ (.Y(\videogen.video_timing_generator.n21_o[0] ),
    .A(net560));
 sg13g2_inv_2 _2535_ (.Y(_1994_),
    .A(\videogen.draw_y[5] ));
 sg13g2_inv_1 _2536_ (.Y(_1995_),
    .A(\videogen.draw_y[6] ));
 sg13g2_inv_1 _2537_ (.Y(_1996_),
    .A(net785));
 sg13g2_inv_2 _2538_ (.Y(_1997_),
    .A(net955));
 sg13g2_inv_1 _2539_ (.Y(_1998_),
    .A(net407));
 sg13g2_inv_1 _2540_ (.Y(_1999_),
    .A(net627));
 sg13g2_inv_1 _2541_ (.Y(_2000_),
    .A(\display_x[4] ));
 sg13g2_inv_1 _2542_ (.Y(_2001_),
    .A(net932));
 sg13g2_inv_1 _2543_ (.Y(_2002_),
    .A(net540));
 sg13g2_inv_1 _2544_ (.Y(_2003_),
    .A(net731));
 sg13g2_inv_1 _2545_ (.Y(_2004_),
    .A(\measurements.n246_q[4] ));
 sg13g2_inv_1 _2546_ (.Y(_2005_),
    .A(\measurements.n246_q[5] ));
 sg13g2_inv_1 _2547_ (.Y(_2006_),
    .A(net101));
 sg13g2_inv_1 _2548_ (.Y(_2007_),
    .A(net350));
 sg13g2_inv_1 _2549_ (.Y(_2008_),
    .A(net787));
 sg13g2_inv_2 _2550_ (.Y(_2009_),
    .A(net933));
 sg13g2_inv_1 _2551_ (.Y(_2010_),
    .A(net292));
 sg13g2_inv_1 _2552_ (.Y(_2011_),
    .A(net333));
 sg13g2_inv_1 _2553_ (.Y(_2012_),
    .A(net849));
 sg13g2_inv_1 _2554_ (.Y(_2013_),
    .A(net927));
 sg13g2_inv_1 _2555_ (.Y(_2014_),
    .A(net163));
 sg13g2_inv_1 _2556_ (.Y(_2015_),
    .A(net269));
 sg13g2_inv_1 _2557_ (.Y(_2016_),
    .A(net170));
 sg13g2_inv_1 _2558_ (.Y(_2017_),
    .A(net204));
 sg13g2_inv_1 _2559_ (.Y(_2018_),
    .A(net488));
 sg13g2_inv_2 _2560_ (.Y(_2019_),
    .A(net567));
 sg13g2_inv_1 _2561_ (.Y(_2020_),
    .A(\measurements.memoryShift[0] ));
 sg13g2_inv_1 _2562_ (.Y(_2021_),
    .A(net402));
 sg13g2_inv_1 _2563_ (.Y(_2022_),
    .A(net418));
 sg13g2_inv_1 _2564_ (.Y(_2023_),
    .A(net343));
 sg13g2_inv_1 _2565_ (.Y(_2024_),
    .A(net752));
 sg13g2_inv_1 _2566_ (.Y(_2025_),
    .A(net749));
 sg13g2_inv_2 _2567_ (.Y(_2026_),
    .A(net582));
 sg13g2_inv_1 _2568_ (.Y(_2027_),
    .A(net592));
 sg13g2_inv_1 _2569_ (.Y(_2028_),
    .A(net782));
 sg13g2_inv_2 _2570_ (.Y(_2029_),
    .A(net773));
 sg13g2_inv_1 _2571_ (.Y(_2030_),
    .A(net996));
 sg13g2_inv_1 _2572_ (.Y(_2031_),
    .A(net160));
 sg13g2_inv_2 _2573_ (.Y(_2032_),
    .A(net790));
 sg13g2_inv_1 _2574_ (.Y(_2033_),
    .A(net856));
 sg13g2_inv_1 _2575_ (.Y(_2034_),
    .A(_0004_));
 sg13g2_inv_1 _2576_ (.Y(_2035_),
    .A(\oscilloscope_control.n220_q[0] ));
 sg13g2_inv_1 _2577_ (.Y(_2036_),
    .A(net1005));
 sg13g2_inv_1 _2578_ (.Y(_2037_),
    .A(_0010_));
 sg13g2_inv_1 _2579_ (.Y(_2038_),
    .A(net114));
 sg13g2_inv_2 _2580_ (.Y(_2039_),
    .A(net442));
 sg13g2_inv_1 _2581_ (.Y(_2040_),
    .A(net892));
 sg13g2_inv_2 _2582_ (.Y(_2041_),
    .A(net26));
 sg13g2_inv_1 _2583_ (.Y(_2042_),
    .A(_0029_));
 sg13g2_inv_1 _2584_ (.Y(_2043_),
    .A(net525));
 sg13g2_inv_1 _2585_ (.Y(_2044_),
    .A(net528));
 sg13g2_inv_1 _2586_ (.Y(_2045_),
    .A(net456));
 sg13g2_inv_1 _2587_ (.Y(_2046_),
    .A(net316));
 sg13g2_inv_1 _2588_ (.Y(_2047_),
    .A(net375));
 sg13g2_inv_1 _2589_ (.Y(_2048_),
    .A(net467));
 sg13g2_inv_1 _2590_ (.Y(_2049_),
    .A(net244));
 sg13g2_inv_1 _2591_ (.Y(_2050_),
    .A(net617));
 sg13g2_inv_1 _2592_ (.Y(_2051_),
    .A(net709));
 sg13g2_inv_1 _2593_ (.Y(_2052_),
    .A(net624));
 sg13g2_inv_1 _2594_ (.Y(_2053_),
    .A(net714));
 sg13g2_inv_1 _2595_ (.Y(_2054_),
    .A(_0039_));
 sg13g2_inv_1 _2596_ (.Y(_2055_),
    .A(net319));
 sg13g2_inv_2 _2597_ (.Y(_2056_),
    .A(net708));
 sg13g2_inv_1 _2598_ (.Y(_2057_),
    .A(net137));
 sg13g2_inv_1 _2599_ (.Y(_2058_),
    .A(net98));
 sg13g2_inv_1 _2600_ (.Y(_2059_),
    .A(net104));
 sg13g2_inv_1 _2601_ (.Y(_2060_),
    .A(_0048_));
 sg13g2_inv_1 _2602_ (.Y(_2061_),
    .A(_0050_));
 sg13g2_inv_1 _2603_ (.Y(_2062_),
    .A(_0051_));
 sg13g2_inv_1 _2604_ (.Y(_2063_),
    .A(net1));
 sg13g2_inv_1 _2605_ (.Y(_2064_),
    .A(\siggen.dac_pmod.n66_o ));
 sg13g2_nor2_1 _2606_ (.A(_1979_),
    .B(net576),
    .Y(_2065_));
 sg13g2_nand2_2 _2607_ (.Y(_2066_),
    .A(net620),
    .B(_1980_));
 sg13g2_nor2_2 _2608_ (.A(net953),
    .B(net579),
    .Y(_2067_));
 sg13g2_nor2_1 _2609_ (.A(net953),
    .B(_2066_),
    .Y(_2068_));
 sg13g2_nand2_2 _2610_ (.Y(_2069_),
    .A(_2065_),
    .B(_2067_));
 sg13g2_nor2_1 _2611_ (.A(net413),
    .B(_2069_),
    .Y(_2070_));
 sg13g2_or2_2 _2612_ (.X(_2071_),
    .B(_2069_),
    .A(net413));
 sg13g2_nor2_2 _2613_ (.A(net588),
    .B(net603),
    .Y(_2072_));
 sg13g2_nor2_1 _2614_ (.A(net548),
    .B(net734),
    .Y(_2073_));
 sg13g2_or2_2 _2615_ (.X(_2074_),
    .B(net735),
    .A(net548));
 sg13g2_nor3_1 _2616_ (.A(net548),
    .B(net588),
    .C(net733),
    .Y(_2075_));
 sg13g2_nand2_2 _2617_ (.Y(_2076_),
    .A(_2072_),
    .B(_2073_));
 sg13g2_nor2_2 _2618_ (.A(net944),
    .B(_2069_),
    .Y(_2077_));
 sg13g2_nand2_1 _2619_ (.Y(_2078_),
    .A(net629),
    .B(net560));
 sg13g2_nand3_1 _2620_ (.B(net629),
    .C(net560),
    .A(net940),
    .Y(_2079_));
 sg13g2_nor2_1 _2621_ (.A(_1993_),
    .B(_2079_),
    .Y(_2080_));
 sg13g2_and2_2 _2622_ (.A(net613),
    .B(_2080_),
    .X(_2081_));
 sg13g2_nand2_1 _2623_ (.Y(_2082_),
    .A(net925),
    .B(_2081_));
 sg13g2_nor2_1 _2624_ (.A(\videogen.draw_y[7] ),
    .B(\videogen.draw_y[8] ),
    .Y(_2083_));
 sg13g2_nand3_1 _2625_ (.B(net785),
    .C(net956),
    .A(net943),
    .Y(_2084_));
 sg13g2_nor2_2 _2626_ (.A(_2082_),
    .B(_2084_),
    .Y(_2085_));
 sg13g2_and2_2 _2627_ (.A(net275),
    .B(net259),
    .X(_2086_));
 sg13g2_nand2_2 _2628_ (.Y(_2087_),
    .A(net275),
    .B(net259));
 sg13g2_and3_1 _2629_ (.X(_2088_),
    .A(net736),
    .B(net381),
    .C(_2086_));
 sg13g2_and2_2 _2630_ (.A(net405),
    .B(net738),
    .X(_2089_));
 sg13g2_nand3_1 _2631_ (.B(net900),
    .C(_2089_),
    .A(net407),
    .Y(_2090_));
 sg13g2_inv_1 _2632_ (.Y(_2091_),
    .A(_2090_));
 sg13g2_nand2_2 _2633_ (.Y(_2092_),
    .A(net381),
    .B(_2001_));
 sg13g2_nand2b_1 _2634_ (.Y(_2093_),
    .B(net518),
    .A_N(net736));
 sg13g2_nor4_1 _2635_ (.A(_2087_),
    .B(_2090_),
    .C(_2092_),
    .D(_2093_),
    .Y(_2094_));
 sg13g2_or4_1 _2636_ (.A(_2087_),
    .B(_2090_),
    .C(_2092_),
    .D(_2093_),
    .X(_2095_));
 sg13g2_nand2_1 _2637_ (.Y(_2096_),
    .A(net518),
    .B(_2086_));
 sg13g2_nor4_2 _2638_ (.A(net736),
    .B(_2090_),
    .C(_2092_),
    .Y(_2097_),
    .D(_2096_));
 sg13g2_o21ai_1 _2639_ (.B1(net656),
    .Y(_2098_),
    .A1(_2002_),
    .A2(_2088_));
 sg13g2_nand2_2 _2640_ (.Y(_2099_),
    .A(_2085_),
    .B(_2098_));
 sg13g2_nor3_1 _2641_ (.A(net944),
    .B(_2069_),
    .C(_2099_),
    .Y(_2100_));
 sg13g2_nor2_1 _2642_ (.A(_2076_),
    .B(_2100_),
    .Y(_2101_));
 sg13g2_nand2_1 _2643_ (.Y(_2102_),
    .A(_2071_),
    .B(_2101_));
 sg13g2_nor2_1 _2644_ (.A(net734),
    .B(net733),
    .Y(_2103_));
 sg13g2_nand2b_1 _2645_ (.Y(_2104_),
    .B(net548),
    .A_N(net734));
 sg13g2_nor2_1 _2646_ (.A(net733),
    .B(_2104_),
    .Y(_2105_));
 sg13g2_nand2_1 _2647_ (.Y(_2106_),
    .A(net588),
    .B(_2105_));
 sg13g2_nand2_1 _2648_ (.Y(_2107_),
    .A(_2076_),
    .B(_2106_));
 sg13g2_a21oi_1 _2649_ (.A1(_2102_),
    .A2(_2107_),
    .Y(_2108_),
    .B1(_2011_));
 sg13g2_nor2b_2 _2650_ (.A(_2076_),
    .B_N(_2100_),
    .Y(_2109_));
 sg13g2_nor2b_1 _2651_ (.A(net552),
    .B_N(net503),
    .Y(_2110_));
 sg13g2_nand2b_2 _2652_ (.Y(_2111_),
    .B(net503),
    .A_N(\measurements.samples_storage.spi_master_inst.n100_q[1] ));
 sg13g2_nor2_1 _2653_ (.A(net186),
    .B(net691),
    .Y(_2112_));
 sg13g2_nor2_1 _2654_ (.A(net333),
    .B(_2112_),
    .Y(_2113_));
 sg13g2_nor2_1 _2655_ (.A(_2106_),
    .B(net334),
    .Y(_2114_));
 sg13g2_nor3_1 _2656_ (.A(_2108_),
    .B(_2109_),
    .C(net335),
    .Y(_0092_));
 sg13g2_nor2_1 _2657_ (.A(\measurements.samples_storage.spi_master_inst.n100_q[0] ),
    .B(\measurements.samples_storage.spi_master_inst.n100_q[1] ),
    .Y(\measurements.fram_cs ));
 sg13g2_nand3_1 _2658_ (.B(_2065_),
    .C(_2067_),
    .A(net944),
    .Y(_2115_));
 sg13g2_nor2_2 _2659_ (.A(_2076_),
    .B(_2115_),
    .Y(_2116_));
 sg13g2_nor2b_1 _2660_ (.A(_2112_),
    .B_N(_2105_),
    .Y(_2117_));
 sg13g2_o21ai_1 _2661_ (.B1(_2107_),
    .Y(_2118_),
    .A1(_2106_),
    .A2(_2112_));
 sg13g2_o21ai_1 _2662_ (.B1(net225),
    .Y(_2119_),
    .A1(_2101_),
    .A2(_2118_));
 sg13g2_nand2b_1 _2663_ (.Y(_0000_),
    .B(net226),
    .A_N(_2116_));
 sg13g2_nand2b_1 _2664_ (.Y(\measurements.adc_cs ),
    .B(\measurements.samples_adc.n84_q[0] ),
    .A_N(\measurements.samples_adc.n84_q[1] ));
 sg13g2_nand2b_2 _2665_ (.Y(\siggen.da_cs ),
    .B(net292),
    .A_N(net569));
 sg13g2_nand3_1 _2666_ (.B(net880),
    .C(net368),
    .A(net295),
    .Y(_2120_));
 sg13g2_and3_1 _2667_ (.X(_2121_),
    .A(net921),
    .B(net295),
    .C(net880));
 sg13g2_nand2_1 _2668_ (.Y(_2122_),
    .A(net368),
    .B(_2121_));
 sg13g2_nor2_2 _2669_ (.A(net269),
    .B(_2122_),
    .Y(_2123_));
 sg13g2_nand3_1 _2670_ (.B(_2015_),
    .C(_2121_),
    .A(net368),
    .Y(_2124_));
 sg13g2_nand2_2 _2671_ (.Y(_2125_),
    .A(net849),
    .B(net927));
 sg13g2_inv_2 _2672_ (.Y(_2126_),
    .A(_2125_));
 sg13g2_nand2_1 _2673_ (.Y(_2127_),
    .A(net655),
    .B(_2126_));
 sg13g2_nand2_1 _2674_ (.Y(_2128_),
    .A(net345),
    .B(_1987_));
 sg13g2_nand2b_1 _2675_ (.Y(_2129_),
    .B(\measurements.trigger.trigger_threshold[3] ),
    .A_N(net345));
 sg13g2_o21ai_1 _2676_ (.B1(_2129_),
    .Y(_2130_),
    .A1(\measurements.n244_o[2] ),
    .A2(_1989_));
 sg13g2_o21ai_1 _2677_ (.B1(_2128_),
    .Y(_2131_),
    .A1(_1988_),
    .A2(net410));
 sg13g2_nor2_1 _2678_ (.A(_2130_),
    .B(_2131_),
    .Y(_2132_));
 sg13g2_xnor2_1 _2679_ (.Y(_2133_),
    .A(net357),
    .B(\measurements.trigger.trigger_threshold[1] ));
 sg13g2_o21ai_1 _2680_ (.B1(_2133_),
    .Y(_2134_),
    .A1(\measurements.trigger.trigger_threshold[0] ),
    .A2(_1985_));
 sg13g2_o21ai_1 _2681_ (.B1(_2134_),
    .Y(_2135_),
    .A1(net357),
    .A2(_1986_));
 sg13g2_a22oi_1 _2682_ (.Y(_2136_),
    .B1(_2132_),
    .B2(_2135_),
    .A2(_2130_),
    .A1(_2128_));
 sg13g2_o21ai_1 _2683_ (.B1(_2132_),
    .Y(_2137_),
    .A1(_1978_),
    .A2(net479));
 sg13g2_nor2_1 _2684_ (.A(_2134_),
    .B(_2137_),
    .Y(_2138_));
 sg13g2_nor2_1 _2685_ (.A(_2136_),
    .B(_2138_),
    .Y(_2139_));
 sg13g2_a22oi_1 _2686_ (.Y(_2140_),
    .B1(net378),
    .B2(_1989_),
    .A2(\lastsample[7] ),
    .A1(_1987_));
 sg13g2_nor2_1 _2687_ (.A(_1987_),
    .B(\lastsample[7] ),
    .Y(_2141_));
 sg13g2_o21ai_1 _2688_ (.B1(_2140_),
    .Y(_2142_),
    .A1(_1989_),
    .A2(net378));
 sg13g2_nor2_1 _2689_ (.A(_2141_),
    .B(_2142_),
    .Y(_2143_));
 sg13g2_nor2_1 _2690_ (.A(\measurements.trigger.trigger_threshold[1] ),
    .B(_1991_),
    .Y(_2144_));
 sg13g2_nor2_1 _2691_ (.A(_1986_),
    .B(net328),
    .Y(_2145_));
 sg13g2_nor2_1 _2692_ (.A(_1978_),
    .B(\lastsample[4] ),
    .Y(_2146_));
 sg13g2_nor3_1 _2693_ (.A(_2144_),
    .B(_2145_),
    .C(_2146_),
    .Y(_2147_));
 sg13g2_o21ai_1 _2694_ (.B1(_2143_),
    .Y(_2148_),
    .A1(_2144_),
    .A2(_2147_));
 sg13g2_o21ai_1 _2695_ (.B1(_2148_),
    .Y(_2149_),
    .A1(_2140_),
    .A2(_2141_));
 sg13g2_nor3_1 _2696_ (.A(\measurements.trigger.sample_on_rising_edge ),
    .B(_2139_),
    .C(_2149_),
    .Y(_2150_));
 sg13g2_nand2_1 _2697_ (.Y(_2151_),
    .A(_1978_),
    .B(\lastsample[4] ));
 sg13g2_nand3_1 _2698_ (.B(_2147_),
    .C(_2151_),
    .A(_2143_),
    .Y(_2152_));
 sg13g2_nand3_1 _2699_ (.B(_2149_),
    .C(_2152_),
    .A(\measurements.trigger.sample_on_rising_edge ),
    .Y(_2153_));
 sg13g2_o21ai_1 _2700_ (.B1(net413),
    .Y(_2154_),
    .A1(_2136_),
    .A2(_2153_));
 sg13g2_o21ai_1 _2701_ (.B1(net134),
    .Y(_2155_),
    .A1(_2150_),
    .A2(_2154_));
 sg13g2_o21ai_1 _2702_ (.B1(net576),
    .Y(_2156_),
    .A1(net347),
    .A2(_2155_));
 sg13g2_nand2b_2 _2703_ (.Y(_2157_),
    .B(net579),
    .A_N(net953));
 sg13g2_nor3_2 _2704_ (.A(net620),
    .B(net577),
    .C(_2157_),
    .Y(_2158_));
 sg13g2_nor2_2 _2705_ (.A(net197),
    .B(net497),
    .Y(_2159_));
 sg13g2_inv_4 _2706_ (.A(_2159_),
    .Y(_2160_));
 sg13g2_and2_1 _2707_ (.A(_2158_),
    .B(_2160_),
    .X(_2161_));
 sg13g2_nor2b_2 _2708_ (.A(net588),
    .B_N(net733),
    .Y(_2162_));
 sg13g2_nand2_2 _2709_ (.Y(_2163_),
    .A(_1992_),
    .B(net733));
 sg13g2_nand2_2 _2710_ (.Y(_2164_),
    .A(net548),
    .B(net734));
 sg13g2_nor2_2 _2711_ (.A(_2163_),
    .B(_2164_),
    .Y(_2165_));
 sg13g2_nand3_1 _2712_ (.B(net734),
    .C(_2162_),
    .A(net548),
    .Y(_2166_));
 sg13g2_nor2_1 _2713_ (.A(net620),
    .B(net576),
    .Y(_2167_));
 sg13g2_nand2b_2 _2714_ (.Y(_2168_),
    .B(_1980_),
    .A_N(_2157_));
 sg13g2_nor3_2 _2715_ (.A(net620),
    .B(_2165_),
    .C(_2168_),
    .Y(_2169_));
 sg13g2_nor4_1 _2716_ (.A(net620),
    .B(_2157_),
    .C(_2161_),
    .D(_2169_),
    .Y(_2170_));
 sg13g2_a22oi_1 _2717_ (.Y(\measurements.n182_o ),
    .B1(_2156_),
    .B2(_2170_),
    .A2(_2127_),
    .A1(net413));
 sg13g2_nor2_2 _2718_ (.A(net483),
    .B(net616),
    .Y(_2171_));
 sg13g2_or2_1 _2719_ (.X(_2172_),
    .B(net616),
    .A(net483));
 sg13g2_o21ai_1 _2720_ (.B1(\settings_uart_printer.uart_tx_module.n88_q[1] ),
    .Y(_2173_),
    .A1(\settings_uart_printer.uart_tx_module.n88_q[0] ),
    .A2(\settings_uart_printer.uart_tx_module.data_reg[0] ));
 sg13g2_nand2_1 _2721_ (.Y(\settings_uart_printer.tx ),
    .A(net689),
    .B(_2173_));
 sg13g2_nor2_2 _2722_ (.A(_2066_),
    .B(_2157_),
    .Y(_2174_));
 sg13g2_nor2_1 _2723_ (.A(_2169_),
    .B(_2174_),
    .Y(_2175_));
 sg13g2_nand2_1 _2724_ (.Y(_2176_),
    .A(net23),
    .B(_2168_));
 sg13g2_o21ai_1 _2725_ (.B1(net24),
    .Y(\measurements.n175_o[0] ),
    .A1(net878),
    .A2(_2175_));
 sg13g2_nand2b_1 _2726_ (.Y(_2177_),
    .B(net978),
    .A_N(net241));
 sg13g2_nand2_1 _2727_ (.Y(_2178_),
    .A(net280),
    .B(net272));
 sg13g2_nor4_1 _2728_ (.A(net216),
    .B(net131),
    .C(_2177_),
    .D(_2178_),
    .Y(_2179_));
 sg13g2_nor3_2 _2729_ (.A(_2066_),
    .B(_2157_),
    .C(_2179_),
    .Y(_2180_));
 sg13g2_nor3_2 _2730_ (.A(_2168_),
    .B(_2169_),
    .C(_2180_),
    .Y(_2181_));
 sg13g2_xnor2_1 _2731_ (.Y(_2182_),
    .A(\measurements.n249_q[0] ),
    .B(net241));
 sg13g2_nor2_1 _2732_ (.A(_2181_),
    .B(net242),
    .Y(\measurements.n175_o[1] ));
 sg13g2_nor3_1 _2733_ (.A(net620),
    .B(_2166_),
    .C(_2168_),
    .Y(_2183_));
 sg13g2_and3_1 _2734_ (.X(_2184_),
    .A(net878),
    .B(net241),
    .C(net131));
 sg13g2_a21oi_1 _2735_ (.A1(\measurements.n249_q[0] ),
    .A2(net954),
    .Y(_2185_),
    .B1(net131));
 sg13g2_nor3_1 _2736_ (.A(_2183_),
    .B(_2184_),
    .C(net132),
    .Y(\measurements.n175_o[2] ));
 sg13g2_and2_1 _2737_ (.A(net216),
    .B(_2184_),
    .X(_2186_));
 sg13g2_nor2_1 _2738_ (.A(net216),
    .B(_2184_),
    .Y(_2187_));
 sg13g2_nor3_1 _2739_ (.A(_2183_),
    .B(_2186_),
    .C(net217),
    .Y(\measurements.n175_o[3] ));
 sg13g2_nand2_1 _2740_ (.Y(_2188_),
    .A(\measurements.n249_q[4] ),
    .B(_2186_));
 sg13g2_xnor2_1 _2741_ (.Y(_2189_),
    .A(net280),
    .B(_2186_));
 sg13g2_nor2_1 _2742_ (.A(_2181_),
    .B(net281),
    .Y(\measurements.n175_o[4] ));
 sg13g2_xor2_1 _2743_ (.B(_2188_),
    .A(net272),
    .X(_2190_));
 sg13g2_nor2_1 _2744_ (.A(_2181_),
    .B(net273),
    .Y(\measurements.n175_o[5] ));
 sg13g2_or2_1 _2745_ (.X(_2191_),
    .B(net560),
    .A(net629));
 sg13g2_and2_1 _2746_ (.A(net630),
    .B(_2191_),
    .X(\videogen.video_timing_generator.n21_o[1] ));
 sg13g2_nand3_1 _2747_ (.B(_1995_),
    .C(net785),
    .A(_1994_),
    .Y(_2192_));
 sg13g2_nor3_2 _2748_ (.A(net906),
    .B(_1997_),
    .C(_2192_),
    .Y(_2193_));
 sg13g2_and2_2 _2749_ (.A(_2081_),
    .B(_2193_),
    .X(_2194_));
 sg13g2_nand2_2 _2750_ (.Y(_2195_),
    .A(_2081_),
    .B(_2193_));
 sg13g2_xnor2_1 _2751_ (.Y(_2196_),
    .A(net337),
    .B(_2078_));
 sg13g2_nor2_1 _2752_ (.A(_2194_),
    .B(net338),
    .Y(\videogen.video_timing_generator.n21_o[2] ));
 sg13g2_xnor2_1 _2753_ (.Y(\videogen.video_timing_generator.n21_o[3] ),
    .A(net397),
    .B(_2079_));
 sg13g2_or2_1 _2754_ (.X(_2197_),
    .B(_2080_),
    .A(net613));
 sg13g2_nor2b_1 _2755_ (.A(_2081_),
    .B_N(net614),
    .Y(\videogen.video_timing_generator.n21_o[4] ));
 sg13g2_nand3b_1 _2756_ (.B(_2081_),
    .C(net495),
    .Y(_2198_),
    .A_N(_2193_));
 sg13g2_o21ai_1 _2757_ (.B1(_2198_),
    .Y(\videogen.video_timing_generator.n21_o[5] ),
    .A1(net495),
    .A2(_2081_));
 sg13g2_or2_1 _2758_ (.X(_2199_),
    .B(_2082_),
    .A(net465));
 sg13g2_nand2_1 _2759_ (.Y(_2200_),
    .A(net653),
    .B(_2199_));
 sg13g2_a21oi_1 _2760_ (.A1(net465),
    .A2(_2082_),
    .Y(\videogen.video_timing_generator.n21_o[6] ),
    .B1(_2200_));
 sg13g2_o21ai_1 _2761_ (.B1(_2195_),
    .Y(_2201_),
    .A1(net574),
    .A2(_2199_));
 sg13g2_a21oi_1 _2762_ (.A1(net574),
    .A2(_2199_),
    .Y(\videogen.video_timing_generator.n21_o[7] ),
    .B1(_2201_));
 sg13g2_nand2_1 _2763_ (.Y(_2202_),
    .A(\videogen.draw_y[5] ),
    .B(\videogen.draw_y[6] ));
 sg13g2_nand4_1 _2764_ (.B(net906),
    .C(\videogen.draw_y[6] ),
    .A(\videogen.draw_y[5] ),
    .Y(_2203_),
    .D(_2081_));
 sg13g2_nand2b_1 _2765_ (.Y(_2204_),
    .B(_2041_),
    .A_N(net907));
 sg13g2_nand2_1 _2766_ (.Y(_2205_),
    .A(_2195_),
    .B(_2204_));
 sg13g2_a21oi_1 _2767_ (.A1(net26),
    .A2(net907),
    .Y(\videogen.video_timing_generator.n21_o[8] ),
    .B1(_2205_));
 sg13g2_a21oi_1 _2768_ (.A1(net537),
    .A2(_2204_),
    .Y(_2206_),
    .B1(_2194_));
 sg13g2_o21ai_1 _2769_ (.B1(_2206_),
    .Y(_2207_),
    .A1(net537),
    .A2(_2204_));
 sg13g2_inv_1 _2770_ (.Y(\videogen.video_timing_generator.n21_o[9] ),
    .A(net538));
 sg13g2_o21ai_1 _2771_ (.B1(_0026_),
    .Y(_2208_),
    .A1(\videogen.draw_y[4] ),
    .A2(_2192_));
 sg13g2_nand2b_1 _2772_ (.Y(_2209_),
    .B(_2197_),
    .A_N(_2202_));
 sg13g2_nor3_1 _2773_ (.A(\videogen.draw_y[5] ),
    .B(\videogen.draw_y[6] ),
    .C(_2197_),
    .Y(_2210_));
 sg13g2_nand3_1 _2774_ (.B(_1997_),
    .C(_2209_),
    .A(\videogen.draw_y[7] ),
    .Y(_2211_));
 sg13g2_o21ai_1 _2775_ (.B1(net785),
    .Y(_2212_),
    .A1(_2210_),
    .A2(_2211_));
 sg13g2_nand2_1 _2776_ (.Y(\videogen.hsync ),
    .A(_2208_),
    .B(_2212_));
 sg13g2_nor2_2 _2777_ (.A(net405),
    .B(net738),
    .Y(_2213_));
 sg13g2_nor3_1 _2778_ (.A(_2089_),
    .B(_2092_),
    .C(_2213_),
    .Y(_2214_));
 sg13g2_nor3_1 _2779_ (.A(_1998_),
    .B(\display_x[2] ),
    .C(net518),
    .Y(_2215_));
 sg13g2_nand4_1 _2780_ (.B(_2086_),
    .C(_2214_),
    .A(\display_x[5] ),
    .Y(\videogen.video_timing_generator.hdmi_vsync ),
    .D(_2215_));
 sg13g2_o21ai_1 _2781_ (.B1(_2098_),
    .Y(_2216_),
    .A1(_1996_),
    .A2(_2083_));
 sg13g2_inv_1 _2782_ (.Y(\videogen.de ),
    .A(_2216_));
 sg13g2_nand2b_1 _2783_ (.Y(_2217_),
    .B(\measurements.fram_mosi ),
    .A_N(net765));
 sg13g2_nor2_1 _2784_ (.A(net779),
    .B(_2217_),
    .Y(_2218_));
 sg13g2_nor2_1 _2785_ (.A(net763),
    .B(_2043_),
    .Y(_2219_));
 sg13g2_a21oi_1 _2786_ (.A1(net779),
    .A2(_2219_),
    .Y(_2220_),
    .B1(_2218_));
 sg13g2_or2_2 _2787_ (.X(_2221_),
    .B(net775),
    .A(net781));
 sg13g2_and2_1 _2788_ (.A(_0042_),
    .B(_2221_),
    .X(_2222_));
 sg13g2_o21ai_1 _2789_ (.B1(_0042_),
    .Y(_2223_),
    .A1(net781),
    .A2(net772));
 sg13g2_nor2_2 _2790_ (.A(_0009_),
    .B(net686),
    .Y(_2224_));
 sg13g2_nor2b_1 _2791_ (.A(_2220_),
    .B_N(_2224_),
    .Y(_2225_));
 sg13g2_nor2b_1 _2792_ (.A(net763),
    .B_N(\measurements.samples_storage.spi_master_inst.n28_o ),
    .Y(_2226_));
 sg13g2_nand2b_1 _2793_ (.Y(_2227_),
    .B(\measurements.samples_storage.spi_master_inst.n28_o ),
    .A_N(net764));
 sg13g2_nor2_1 _2794_ (.A(net699),
    .B(_2227_),
    .Y(_2228_));
 sg13g2_a21oi_1 _2795_ (.A1(net698),
    .A2(_2219_),
    .Y(_2229_),
    .B1(_2228_));
 sg13g2_nor2_1 _2796_ (.A(\oscilloscope_control.n114_o[0] ),
    .B(_2217_),
    .Y(_2230_));
 sg13g2_a21oi_1 _2797_ (.A1(net776),
    .A2(_2229_),
    .Y(_2231_),
    .B1(net687));
 sg13g2_o21ai_1 _2798_ (.B1(_2231_),
    .Y(_2232_),
    .A1(net771),
    .A2(_2230_));
 sg13g2_inv_1 _2799_ (.Y(_2233_),
    .A(_2232_));
 sg13g2_nand2_1 _2800_ (.Y(_2234_),
    .A(net740),
    .B(_2233_));
 sg13g2_nor2_1 _2801_ (.A(net766),
    .B(_2221_),
    .Y(_2235_));
 sg13g2_or3_1 _2802_ (.A(net779),
    .B(net771),
    .C(net763),
    .X(_2236_));
 sg13g2_nand2b_1 _2803_ (.Y(_2237_),
    .B(\measurements.samples_storage.spi_master_inst.n26_o ),
    .A_N(net764));
 sg13g2_nor2_1 _2804_ (.A(net699),
    .B(_2237_),
    .Y(_2238_));
 sg13g2_a21oi_1 _2805_ (.A1(net699),
    .A2(_2226_),
    .Y(_2239_),
    .B1(_2238_));
 sg13g2_nand2_1 _2806_ (.Y(_2240_),
    .A(net775),
    .B(_2239_));
 sg13g2_a21oi_1 _2807_ (.A1(_2029_),
    .A2(_2220_),
    .Y(_2241_),
    .B1(net687));
 sg13g2_a22oi_1 _2808_ (.Y(_2242_),
    .B1(_2240_),
    .B2(_2241_),
    .A2(_2235_),
    .A1(_2061_));
 sg13g2_nor2b_1 _2809_ (.A(_2242_),
    .B_N(net742),
    .Y(_2243_));
 sg13g2_and2_1 _2810_ (.A(net687),
    .B(net685),
    .X(_2244_));
 sg13g2_nand2_1 _2811_ (.Y(_2245_),
    .A(net687),
    .B(_2236_));
 sg13g2_o21ai_1 _2812_ (.B1(net763),
    .Y(_2246_),
    .A1(net779),
    .A2(net771));
 sg13g2_nand2_1 _2813_ (.Y(_2247_),
    .A(net685),
    .B(_2246_));
 sg13g2_a21o_1 _2814_ (.A2(_2246_),
    .A1(net685),
    .B1(_2050_),
    .X(_2248_));
 sg13g2_a21o_1 _2815_ (.A2(_2246_),
    .A1(net685),
    .B1(_2043_),
    .X(_2249_));
 sg13g2_mux2_1 _2816_ (.A0(_2248_),
    .A1(_2249_),
    .S(net698),
    .X(_2250_));
 sg13g2_nand2_2 _2817_ (.Y(_2251_),
    .A(net782),
    .B(net774));
 sg13g2_and2_2 _2818_ (.A(_2221_),
    .B(_2251_),
    .X(_2252_));
 sg13g2_xnor2_1 _2819_ (.Y(_2253_),
    .A(net783),
    .B(net773));
 sg13g2_nor2_2 _2820_ (.A(_0042_),
    .B(net684),
    .Y(_2254_));
 sg13g2_or2_2 _2821_ (.X(_2255_),
    .B(_2253_),
    .A(_0042_));
 sg13g2_nand2b_1 _2822_ (.Y(_2256_),
    .B(\measurements.samples_storage.spi_master_inst.n24_o ),
    .A_N(net766));
 sg13g2_mux2_1 _2823_ (.A0(_2237_),
    .A1(_2256_),
    .S(net781),
    .X(_2257_));
 sg13g2_a21oi_1 _2824_ (.A1(net780),
    .A2(_2226_),
    .Y(_2258_),
    .B1(net775));
 sg13g2_a21o_1 _2825_ (.A2(_2257_),
    .A1(net772),
    .B1(_2258_),
    .X(_2259_));
 sg13g2_a21oi_1 _2826_ (.A1(_2062_),
    .A2(net687),
    .Y(_2260_),
    .B1(net679));
 sg13g2_a221oi_1 _2827_ (.B2(_2260_),
    .C1(_2254_),
    .B1(_2259_),
    .A1(net679),
    .Y(_2261_),
    .A2(_2250_));
 sg13g2_nand2b_1 _2828_ (.Y(_2262_),
    .B(_2261_),
    .A_N(_0007_));
 sg13g2_a21o_1 _2829_ (.A2(_2246_),
    .A1(net685),
    .B1(_2044_),
    .X(_2263_));
 sg13g2_a21oi_1 _2830_ (.A1(net764),
    .A2(\measurements.samples_storage.spi_master_inst.n30_o ),
    .Y(_2264_),
    .B1(net699));
 sg13g2_a21oi_1 _2831_ (.A1(net699),
    .A2(_2263_),
    .Y(_2265_),
    .B1(_2264_));
 sg13g2_a221oi_1 _2832_ (.B2(net699),
    .C1(_2264_),
    .B1(_2263_),
    .A1(_2221_),
    .Y(_2266_),
    .A2(_2251_));
 sg13g2_nor2_2 _2833_ (.A(net783),
    .B(_2029_),
    .Y(_2267_));
 sg13g2_nand2_2 _2834_ (.Y(_2268_),
    .A(net697),
    .B(net771));
 sg13g2_o21ai_1 _2835_ (.B1(net679),
    .Y(_2269_),
    .A1(_2248_),
    .A2(_2268_));
 sg13g2_nand2b_1 _2836_ (.Y(_2270_),
    .B(\measurements.samples_storage.spi_master_inst.n22_o ),
    .A_N(net766));
 sg13g2_mux2_1 _2837_ (.A0(_2256_),
    .A1(_2270_),
    .S(net782),
    .X(_2271_));
 sg13g2_inv_1 _2838_ (.Y(_2272_),
    .A(_2271_));
 sg13g2_mux4_1 _2839_ (.S0(net781),
    .A0(_2227_),
    .A1(_2237_),
    .A2(_2256_),
    .A3(_2270_),
    .S1(net772),
    .X(_2273_));
 sg13g2_nor4_1 _2840_ (.A(net780),
    .B(net772),
    .C(net764),
    .D(_0052_),
    .Y(_2274_));
 sg13g2_a21oi_1 _2841_ (.A1(net687),
    .A2(net685),
    .Y(_2275_),
    .B1(_2274_));
 sg13g2_o21ai_1 _2842_ (.B1(_2275_),
    .Y(_2276_),
    .A1(net680),
    .A2(_2273_));
 sg13g2_o21ai_1 _2843_ (.B1(_2276_),
    .Y(_2277_),
    .A1(_2266_),
    .A2(_2269_));
 sg13g2_or2_1 _2844_ (.X(_2278_),
    .B(_2277_),
    .A(_2009_));
 sg13g2_xor2_1 _2845_ (.B(_2261_),
    .A(_0007_),
    .X(_2279_));
 sg13g2_or2_1 _2846_ (.X(_2280_),
    .B(_2279_),
    .A(_2278_));
 sg13g2_o21ai_1 _2847_ (.B1(_2262_),
    .Y(_2281_),
    .A1(_2278_),
    .A2(_2279_));
 sg13g2_nand2b_1 _2848_ (.Y(_2282_),
    .B(_2242_),
    .A_N(net742));
 sg13g2_nand2b_1 _2849_ (.Y(_2283_),
    .B(_2282_),
    .A_N(_2243_));
 sg13g2_nand2b_1 _2850_ (.Y(_2284_),
    .B(_2281_),
    .A_N(_2283_));
 sg13g2_a21oi_1 _2851_ (.A1(_2281_),
    .A2(_2282_),
    .Y(_2285_),
    .B1(_2243_));
 sg13g2_nor2_1 _2852_ (.A(net740),
    .B(_2233_),
    .Y(_2286_));
 sg13g2_xnor2_1 _2853_ (.Y(_2287_),
    .A(net740),
    .B(_2232_));
 sg13g2_o21ai_1 _2854_ (.B1(_2234_),
    .Y(_2288_),
    .A1(_2285_),
    .A2(_2286_));
 sg13g2_xnor2_1 _2855_ (.Y(_2289_),
    .A(_0043_),
    .B(_2225_));
 sg13g2_a22oi_1 _2856_ (.Y(_2290_),
    .B1(_2288_),
    .B2(_2289_),
    .A2(_2225_),
    .A1(\choffset[4] ));
 sg13g2_and2_1 _2857_ (.A(_2224_),
    .B(_2230_),
    .X(_2291_));
 sg13g2_xor2_1 _2858_ (.B(_2291_),
    .A(_2290_),
    .X(_2292_));
 sg13g2_inv_2 _2859_ (.Y(_2293_),
    .A(_2292_));
 sg13g2_xnor2_1 _2860_ (.Y(_2294_),
    .A(_2285_),
    .B(_2287_));
 sg13g2_nand2_1 _2861_ (.Y(_2295_),
    .A(_2292_),
    .B(_2294_));
 sg13g2_xor2_1 _2862_ (.B(_2289_),
    .A(_2288_),
    .X(_2296_));
 sg13g2_o21ai_1 _2863_ (.B1(_1996_),
    .Y(_2297_),
    .A1(_2293_),
    .A2(_2296_));
 sg13g2_xnor2_1 _2864_ (.Y(_2298_),
    .A(_1997_),
    .B(_2295_));
 sg13g2_nand2b_1 _2865_ (.Y(_2299_),
    .B(_2283_),
    .A_N(_2281_));
 sg13g2_and3_1 _2866_ (.X(_2300_),
    .A(_2284_),
    .B(_2292_),
    .C(_2299_));
 sg13g2_nor2_1 _2867_ (.A(_0024_),
    .B(_2300_),
    .Y(_2301_));
 sg13g2_nand3b_1 _2868_ (.B(net785),
    .C(_2292_),
    .Y(_2302_),
    .A_N(_2296_));
 sg13g2_nand3_1 _2869_ (.B(_2298_),
    .C(_2302_),
    .A(_2297_),
    .Y(_2303_));
 sg13g2_nor2_1 _2870_ (.A(_2301_),
    .B(_2303_),
    .Y(_2304_));
 sg13g2_nand2_1 _2871_ (.Y(_2305_),
    .A(_2278_),
    .B(_2279_));
 sg13g2_a21o_1 _2872_ (.A2(_2305_),
    .A1(_2280_),
    .B1(_2293_),
    .X(_2306_));
 sg13g2_xor2_1 _2873_ (.B(_2306_),
    .A(_0023_),
    .X(_2307_));
 sg13g2_xnor2_1 _2874_ (.Y(_2308_),
    .A(\oscilloscope_control.n111_o[0] ),
    .B(_2277_));
 sg13g2_nand2_1 _2875_ (.Y(_2309_),
    .A(_2292_),
    .B(_2308_));
 sg13g2_nor2_2 _2876_ (.A(net676),
    .B(_2252_),
    .Y(_2310_));
 sg13g2_nand2_1 _2877_ (.Y(_2311_),
    .A(net678),
    .B(net684));
 sg13g2_a21oi_1 _2878_ (.A1(\measurements.samples_storage.spi_master_inst.n26_o ),
    .A2(net675),
    .Y(_2312_),
    .B1(net780));
 sg13g2_a21o_1 _2879_ (.A2(_2263_),
    .A1(net780),
    .B1(_2312_),
    .X(_2313_));
 sg13g2_nor2_1 _2880_ (.A(_2250_),
    .B(_2255_),
    .Y(_2314_));
 sg13g2_nor2_1 _2881_ (.A(net767),
    .B(_2048_),
    .Y(_2315_));
 sg13g2_nand2_1 _2882_ (.Y(_2316_),
    .A(net782),
    .B(_2315_));
 sg13g2_o21ai_1 _2883_ (.B1(_2316_),
    .Y(_2317_),
    .A1(net782),
    .A2(_2270_));
 sg13g2_nand2_1 _2884_ (.Y(_2318_),
    .A(net774),
    .B(_2317_));
 sg13g2_o21ai_1 _2885_ (.B1(_2318_),
    .Y(_2319_),
    .A1(net774),
    .A2(_2257_));
 sg13g2_a21oi_1 _2886_ (.A1(net677),
    .A2(_2319_),
    .Y(_2320_),
    .B1(_2314_));
 sg13g2_o21ai_1 _2887_ (.B1(_2320_),
    .Y(_2321_),
    .A1(_2311_),
    .A2(_2313_));
 sg13g2_nor2_1 _2888_ (.A(_2293_),
    .B(_2321_),
    .Y(_2322_));
 sg13g2_xnor2_1 _2889_ (.Y(_2323_),
    .A(_0022_),
    .B(_2309_));
 sg13g2_a21oi_1 _2890_ (.A1(_2060_),
    .A2(_2322_),
    .Y(_2324_),
    .B1(_2323_));
 sg13g2_o21ai_1 _2891_ (.B1(_0048_),
    .Y(_2325_),
    .A1(_2293_),
    .A2(_2321_));
 sg13g2_nand3_1 _2892_ (.B(\measurements.samples_storage.spi_master_inst.n24_o ),
    .C(net675),
    .A(net700),
    .Y(_2326_));
 sg13g2_nand3_1 _2893_ (.B(net766),
    .C(\measurements.samples_storage.spi_master_inst.n26_o ),
    .A(net780),
    .Y(_2327_));
 sg13g2_and2_1 _2894_ (.A(_2326_),
    .B(_2327_),
    .X(_2328_));
 sg13g2_o21ai_1 _2895_ (.B1(_2255_),
    .Y(_2329_),
    .A1(net677),
    .A2(_2328_));
 sg13g2_o21ai_1 _2896_ (.B1(_2329_),
    .Y(_2330_),
    .A1(net684),
    .A2(_2265_));
 sg13g2_nand2b_1 _2897_ (.Y(_2331_),
    .B(\measurements.samples_storage.spi_master_inst.n18_o ),
    .A_N(net767));
 sg13g2_nor2_1 _2898_ (.A(net700),
    .B(_2331_),
    .Y(_2332_));
 sg13g2_a21oi_1 _2899_ (.A1(net700),
    .A2(_2315_),
    .Y(_2333_),
    .B1(_2332_));
 sg13g2_a21oi_1 _2900_ (.A1(net773),
    .A2(_2333_),
    .Y(_2334_),
    .B1(net678));
 sg13g2_o21ai_1 _2901_ (.B1(_2334_),
    .Y(_2335_),
    .A1(net773),
    .A2(_2272_));
 sg13g2_nand3_1 _2902_ (.B(_2330_),
    .C(_2335_),
    .A(_2292_),
    .Y(_2336_));
 sg13g2_nor2_1 _2903_ (.A(_1993_),
    .B(_2336_),
    .Y(_2337_));
 sg13g2_nand3_1 _2904_ (.B(\measurements.samples_storage.spi_master_inst.n22_o ),
    .C(net675),
    .A(net699),
    .Y(_2338_));
 sg13g2_nand3_1 _2905_ (.B(net766),
    .C(\measurements.samples_storage.spi_master_inst.n24_o ),
    .A(net782),
    .Y(_2339_));
 sg13g2_nand2_1 _2906_ (.Y(_2340_),
    .A(_2338_),
    .B(_2339_));
 sg13g2_nor2_1 _2907_ (.A(net684),
    .B(_2340_),
    .Y(_2341_));
 sg13g2_nor2_2 _2908_ (.A(_0042_),
    .B(_2246_),
    .Y(_2342_));
 sg13g2_a21oi_1 _2909_ (.A1(_2048_),
    .A2(net684),
    .Y(_2343_),
    .B1(_2341_));
 sg13g2_nor2_1 _2910_ (.A(_2029_),
    .B(_0009_),
    .Y(_2344_));
 sg13g2_nor3_1 _2911_ (.A(net783),
    .B(_2331_),
    .C(_2344_),
    .Y(_2345_));
 sg13g2_a22oi_1 _2912_ (.Y(_2346_),
    .B1(_2345_),
    .B2(net676),
    .A2(_2343_),
    .A1(_2342_));
 sg13g2_and2_1 _2913_ (.A(_2292_),
    .B(_2346_),
    .X(_2347_));
 sg13g2_nand2_1 _2914_ (.Y(_2348_),
    .A(\videogen.draw_y[0] ),
    .B(_2347_));
 sg13g2_o21ai_1 _2915_ (.B1(net774),
    .Y(_2349_),
    .A1(net782),
    .A2(_2331_));
 sg13g2_o21ai_1 _2916_ (.B1(_2349_),
    .Y(_2350_),
    .A1(net774),
    .A2(_2317_));
 sg13g2_nor2_1 _2917_ (.A(net678),
    .B(_2350_),
    .Y(_2351_));
 sg13g2_a21oi_1 _2918_ (.A1(_2310_),
    .A2(_2340_),
    .Y(_2352_),
    .B1(_2351_));
 sg13g2_o21ai_1 _2919_ (.B1(_2352_),
    .Y(_2353_),
    .A1(_2255_),
    .A2(_2313_));
 sg13g2_nor2_1 _2920_ (.A(_2293_),
    .B(_2353_),
    .Y(_2354_));
 sg13g2_xnor2_1 _2921_ (.Y(_2355_),
    .A(_0021_),
    .B(_2354_));
 sg13g2_a21oi_1 _2922_ (.A1(\measurements.samples_storage.spi_master_inst.n22_o ),
    .A2(net675),
    .Y(_2356_),
    .B1(_2251_));
 sg13g2_a21oi_1 _2923_ (.A1(_2252_),
    .A2(_2328_),
    .Y(_2357_),
    .B1(_2356_));
 sg13g2_nand3b_1 _2924_ (.B(_0009_),
    .C(net677),
    .Y(_2358_),
    .A_N(_2333_));
 sg13g2_a22oi_1 _2925_ (.Y(_2359_),
    .B1(_2342_),
    .B2(_2357_),
    .A2(net680),
    .A1(\measurements.samples_storage.spi_master_inst.n20_o ));
 sg13g2_nand3_1 _2926_ (.B(_2358_),
    .C(_2359_),
    .A(_2292_),
    .Y(_2360_));
 sg13g2_xor2_1 _2927_ (.B(_2360_),
    .A(_0047_),
    .X(_2361_));
 sg13g2_nand2_1 _2928_ (.Y(_2362_),
    .A(_1993_),
    .B(_2336_));
 sg13g2_o21ai_1 _2929_ (.B1(_2362_),
    .Y(_2363_),
    .A1(\videogen.draw_y[2] ),
    .A2(_2354_));
 sg13g2_nor2b_1 _2930_ (.A(\videogen.draw_y[1] ),
    .B_N(_2360_),
    .Y(_2364_));
 sg13g2_a21o_1 _2931_ (.A2(_2361_),
    .A1(_2348_),
    .B1(_2364_),
    .X(_2365_));
 sg13g2_a21oi_1 _2932_ (.A1(_2355_),
    .A2(_2365_),
    .Y(_2366_),
    .B1(_2363_));
 sg13g2_o21ai_1 _2933_ (.B1(_2325_),
    .Y(_2367_),
    .A1(_2337_),
    .A2(_2366_));
 sg13g2_a22oi_1 _2934_ (.Y(_2368_),
    .B1(_2324_),
    .B2(_2367_),
    .A2(_2309_),
    .A1(_1994_));
 sg13g2_nand2b_1 _2935_ (.Y(_2369_),
    .B(_2307_),
    .A_N(_2368_));
 sg13g2_nand2_1 _2936_ (.Y(_2370_),
    .A(_0024_),
    .B(_2300_));
 sg13g2_a22oi_1 _2937_ (.Y(_2371_),
    .B1(_2306_),
    .B2(_1995_),
    .A2(_2300_),
    .A1(net786));
 sg13g2_nand2_1 _2938_ (.Y(_2372_),
    .A(_2369_),
    .B(_2371_));
 sg13g2_o21ai_1 _2939_ (.B1(_2297_),
    .Y(_2373_),
    .A1(_2041_),
    .A2(_2295_));
 sg13g2_a22oi_1 _2940_ (.Y(_2374_),
    .B1(_2373_),
    .B2(_2302_),
    .A2(_2372_),
    .A1(_2304_));
 sg13g2_nand2b_1 _2941_ (.Y(_2375_),
    .B(\lastsample[7] ),
    .A_N(net762));
 sg13g2_nand2b_1 _2942_ (.Y(_2376_),
    .B(\lastsample[6] ),
    .A_N(net762));
 sg13g2_mux2_1 _2943_ (.A0(_2375_),
    .A1(_2376_),
    .S(net777),
    .X(_2377_));
 sg13g2_nor2b_1 _2944_ (.A(_2377_),
    .B_N(_2224_),
    .Y(_2378_));
 sg13g2_nand2b_1 _2945_ (.Y(_2379_),
    .B(\lastsample[5] ),
    .A_N(net762));
 sg13g2_mux2_1 _2946_ (.A0(_2376_),
    .A1(_2379_),
    .S(net777),
    .X(_2380_));
 sg13g2_nor2_1 _2947_ (.A(\oscilloscope_control.n114_o[0] ),
    .B(_2375_),
    .Y(_2381_));
 sg13g2_a21oi_1 _2948_ (.A1(net770),
    .A2(_2380_),
    .Y(_2382_),
    .B1(net686));
 sg13g2_o21ai_1 _2949_ (.B1(_2382_),
    .Y(_2383_),
    .A1(net770),
    .A2(_2381_));
 sg13g2_nor2_1 _2950_ (.A(_2027_),
    .B(_2383_),
    .Y(_2384_));
 sg13g2_nor2_1 _2951_ (.A(net777),
    .B(_2379_),
    .Y(_0294_));
 sg13g2_nor2b_1 _2952_ (.A(net764),
    .B_N(\lastsample[4] ),
    .Y(_0295_));
 sg13g2_nand2b_1 _2953_ (.Y(_0296_),
    .B(\lastsample[4] ),
    .A_N(net763));
 sg13g2_nor2_1 _2954_ (.A(net697),
    .B(_0296_),
    .Y(_0297_));
 sg13g2_o21ai_1 _2955_ (.B1(net771),
    .Y(_0298_),
    .A1(_0294_),
    .A2(_0297_));
 sg13g2_nor2_1 _2956_ (.A(net770),
    .B(_2377_),
    .Y(_0299_));
 sg13g2_nor2_1 _2957_ (.A(net680),
    .B(_0299_),
    .Y(_0300_));
 sg13g2_a221oi_1 _2958_ (.B2(_0300_),
    .C1(net678),
    .B1(_0298_),
    .A1(_0044_),
    .Y(_0301_),
    .A2(net686));
 sg13g2_nand2_1 _2959_ (.Y(_0302_),
    .A(net742),
    .B(_0301_));
 sg13g2_xnor2_1 _2960_ (.Y(_0303_),
    .A(net742),
    .B(_0301_));
 sg13g2_a21o_1 _2961_ (.A2(_2246_),
    .A1(net685),
    .B1(_1990_),
    .X(_0304_));
 sg13g2_and2_1 _2962_ (.A(\lastsample[7] ),
    .B(net674),
    .X(_0305_));
 sg13g2_a21oi_1 _2963_ (.A1(\lastsample[7] ),
    .A2(net763),
    .Y(_0306_),
    .B1(net697));
 sg13g2_a21o_1 _2964_ (.A2(_0304_),
    .A1(net697),
    .B1(_0306_),
    .X(_0307_));
 sg13g2_a21oi_1 _2965_ (.A1(net698),
    .A2(_0304_),
    .Y(_0308_),
    .B1(_0306_));
 sg13g2_or2_1 _2966_ (.X(_0309_),
    .B(_2380_),
    .A(net771));
 sg13g2_nand2b_1 _2967_ (.Y(_0310_),
    .B(\lastsample[3] ),
    .A_N(net767));
 sg13g2_nand3b_1 _2968_ (.B(\lastsample[3] ),
    .C(net780),
    .Y(_0311_),
    .A_N(net763));
 sg13g2_o21ai_1 _2969_ (.B1(_0311_),
    .Y(_0312_),
    .A1(net779),
    .A2(_0296_));
 sg13g2_a21oi_1 _2970_ (.A1(net771),
    .A2(_0312_),
    .Y(_0313_),
    .B1(net686));
 sg13g2_a21o_1 _2971_ (.A2(net680),
    .A1(_0045_),
    .B1(_2254_),
    .X(_0314_));
 sg13g2_a221oi_1 _2972_ (.B2(_0313_),
    .C1(_0314_),
    .B1(_0309_),
    .A1(net678),
    .Y(_0315_),
    .A2(_0307_));
 sg13g2_nor2b_1 _2973_ (.A(_0007_),
    .B_N(_0315_),
    .Y(_0316_));
 sg13g2_a21oi_1 _2974_ (.A1(net685),
    .A2(_2246_),
    .Y(_0317_),
    .B1(_1991_));
 sg13g2_and3_1 _2975_ (.X(_0318_),
    .A(\lastsample[6] ),
    .B(net779),
    .C(net763));
 sg13g2_a21o_1 _2976_ (.A2(_0317_),
    .A1(net698),
    .B1(_0318_),
    .X(_0319_));
 sg13g2_a221oi_1 _2977_ (.B2(net684),
    .C1(net676),
    .B1(_0319_),
    .A1(_2267_),
    .Y(_0320_),
    .A2(_0305_));
 sg13g2_nand2b_1 _2978_ (.Y(_0321_),
    .B(\lastsample[2] ),
    .A_N(net766));
 sg13g2_mux2_2 _2979_ (.A0(_0310_),
    .A1(_0321_),
    .S(net784),
    .X(_0322_));
 sg13g2_inv_1 _2980_ (.Y(_0323_),
    .A(_0322_));
 sg13g2_a21oi_1 _2981_ (.A1(net780),
    .A2(_0295_),
    .Y(_0324_),
    .B1(net772));
 sg13g2_a21oi_1 _2982_ (.A1(net772),
    .A2(_0322_),
    .Y(_0325_),
    .B1(_0324_));
 sg13g2_o21ai_1 _2983_ (.B1(net676),
    .Y(_0326_),
    .A1(_0046_),
    .A2(_2222_));
 sg13g2_nor2_1 _2984_ (.A(_0325_),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_nor2_1 _2985_ (.A(_0320_),
    .B(_0327_),
    .Y(_0328_));
 sg13g2_nor3_1 _2986_ (.A(_2009_),
    .B(_0320_),
    .C(_0327_),
    .Y(_0329_));
 sg13g2_xnor2_1 _2987_ (.Y(_0330_),
    .A(_0007_),
    .B(_0315_));
 sg13g2_a21oi_1 _2988_ (.A1(_0329_),
    .A2(_0330_),
    .Y(_0331_),
    .B1(_0316_));
 sg13g2_o21ai_1 _2989_ (.B1(_0302_),
    .Y(_0332_),
    .A1(_0303_),
    .A2(_0331_));
 sg13g2_xnor2_1 _2990_ (.Y(_0333_),
    .A(net739),
    .B(_2383_));
 sg13g2_a21oi_1 _2991_ (.A1(_0332_),
    .A2(_0333_),
    .Y(_0334_),
    .B1(_2384_));
 sg13g2_xor2_1 _2992_ (.B(_2378_),
    .A(_0043_),
    .X(_0335_));
 sg13g2_nor2_1 _2993_ (.A(_0334_),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_a21o_1 _2994_ (.A2(_2378_),
    .A1(\choffset[4] ),
    .B1(_0336_),
    .X(_0337_));
 sg13g2_and2_1 _2995_ (.A(_2224_),
    .B(_2381_),
    .X(_0338_));
 sg13g2_xnor2_1 _2996_ (.Y(_0339_),
    .A(_0337_),
    .B(_0338_));
 sg13g2_a21o_1 _2997_ (.A2(net674),
    .A1(\lastsample[4] ),
    .B1(net779),
    .X(_0340_));
 sg13g2_o21ai_1 _2998_ (.B1(_0340_),
    .Y(_0341_),
    .A1(net698),
    .A2(_0317_));
 sg13g2_o21ai_1 _2999_ (.B1(_2255_),
    .Y(_0342_),
    .A1(net676),
    .A2(_0341_));
 sg13g2_o21ai_1 _3000_ (.B1(_0342_),
    .Y(_0343_),
    .A1(net684),
    .A2(_0308_));
 sg13g2_nor2_1 _3001_ (.A(net784),
    .B(_0321_),
    .Y(_0344_));
 sg13g2_nor2b_1 _3002_ (.A(net766),
    .B_N(\lastsample[1] ),
    .Y(_0345_));
 sg13g2_a21oi_2 _3003_ (.B1(_0344_),
    .Y(_0346_),
    .A2(_0345_),
    .A1(net784));
 sg13g2_o21ai_1 _3004_ (.B1(net676),
    .Y(_0347_),
    .A1(net772),
    .A2(_0312_));
 sg13g2_a21o_1 _3005_ (.A2(_0346_),
    .A1(net772),
    .B1(_0347_),
    .X(_0348_));
 sg13g2_nand3_1 _3006_ (.B(_0343_),
    .C(_0348_),
    .A(net638),
    .Y(_0349_));
 sg13g2_and2_1 _3007_ (.A(_0048_),
    .B(_0349_),
    .X(_0350_));
 sg13g2_a21oi_1 _3008_ (.A1(\lastsample[4] ),
    .A2(net764),
    .Y(_0351_),
    .B1(net698));
 sg13g2_a21oi_1 _3009_ (.A1(\lastsample[3] ),
    .A2(net675),
    .Y(_0352_),
    .B1(net780));
 sg13g2_or2_1 _3010_ (.X(_0353_),
    .B(_0352_),
    .A(_0351_));
 sg13g2_o21ai_1 _3011_ (.B1(_2255_),
    .Y(_0354_),
    .A1(net676),
    .A2(_0353_));
 sg13g2_o21ai_1 _3012_ (.B1(_0354_),
    .Y(_0355_),
    .A1(net684),
    .A2(_0319_));
 sg13g2_nand2b_2 _3013_ (.Y(_0356_),
    .B(\lastsample[0] ),
    .A_N(net767));
 sg13g2_nor2_1 _3014_ (.A(net700),
    .B(_0356_),
    .Y(_0357_));
 sg13g2_a21oi_1 _3015_ (.A1(net700),
    .A2(_0345_),
    .Y(_0358_),
    .B1(_0357_));
 sg13g2_a21oi_1 _3016_ (.A1(net773),
    .A2(_0358_),
    .Y(_0359_),
    .B1(net679));
 sg13g2_o21ai_1 _3017_ (.B1(_0359_),
    .Y(_0360_),
    .A1(net773),
    .A2(_0323_));
 sg13g2_nand3_1 _3018_ (.B(_0355_),
    .C(_0360_),
    .A(_0339_),
    .Y(_0361_));
 sg13g2_or2_1 _3019_ (.X(_0362_),
    .B(_0361_),
    .A(_1993_));
 sg13g2_a21oi_1 _3020_ (.A1(\lastsample[2] ),
    .A2(net675),
    .Y(_0363_),
    .B1(_2251_));
 sg13g2_a21oi_1 _3021_ (.A1(_2252_),
    .A2(_0353_),
    .Y(_0364_),
    .B1(_0363_));
 sg13g2_nand3b_1 _3022_ (.B(_0009_),
    .C(net676),
    .Y(_0365_),
    .A_N(_0358_));
 sg13g2_a22oi_1 _3023_ (.Y(_0366_),
    .B1(_2342_),
    .B2(_0364_),
    .A2(net680),
    .A1(\lastsample[1] ));
 sg13g2_nand3_1 _3024_ (.B(_0365_),
    .C(_0366_),
    .A(net638),
    .Y(_0367_));
 sg13g2_nand2b_1 _3025_ (.Y(_0368_),
    .B(_0367_),
    .A_N(\videogen.draw_y[1] ));
 sg13g2_xnor2_1 _3026_ (.Y(_0369_),
    .A(_0047_),
    .B(_0367_));
 sg13g2_nor3_1 _3027_ (.A(net783),
    .B(_2036_),
    .C(_0356_),
    .Y(_0370_));
 sg13g2_o21ai_1 _3028_ (.B1(net686),
    .Y(_0371_),
    .A1(_2221_),
    .A2(_0356_));
 sg13g2_o21ai_1 _3029_ (.B1(_0371_),
    .Y(_0372_),
    .A1(net680),
    .A2(_0370_));
 sg13g2_a21oi_1 _3030_ (.A1(net766),
    .A2(\lastsample[3] ),
    .Y(_0373_),
    .B1(net699));
 sg13g2_a21oi_1 _3031_ (.A1(\lastsample[2] ),
    .A2(net674),
    .Y(_0374_),
    .B1(net782));
 sg13g2_or2_1 _3032_ (.X(_0375_),
    .B(_0374_),
    .A(_0373_));
 sg13g2_o21ai_1 _3033_ (.B1(_2342_),
    .Y(_0376_),
    .A1(\lastsample[1] ),
    .A2(_2252_));
 sg13g2_a21o_1 _3034_ (.A2(_0375_),
    .A1(_2252_),
    .B1(_0376_),
    .X(_0377_));
 sg13g2_nand3_1 _3035_ (.B(_0372_),
    .C(_0377_),
    .A(net638),
    .Y(_0378_));
 sg13g2_nor2_1 _3036_ (.A(_0049_),
    .B(_0378_),
    .Y(_0379_));
 sg13g2_o21ai_1 _3037_ (.B1(_0368_),
    .Y(_0380_),
    .A1(_0369_),
    .A2(_0379_));
 sg13g2_nor2_1 _3038_ (.A(_2255_),
    .B(_0341_),
    .Y(_0381_));
 sg13g2_nand2_1 _3039_ (.Y(_0382_),
    .A(_2029_),
    .B(_0346_));
 sg13g2_o21ai_1 _3040_ (.B1(net773),
    .Y(_0383_),
    .A1(net783),
    .A2(_0356_));
 sg13g2_nand3_1 _3041_ (.B(_0382_),
    .C(_0383_),
    .A(net677),
    .Y(_0384_));
 sg13g2_o21ai_1 _3042_ (.B1(_0384_),
    .Y(_0385_),
    .A1(_2311_),
    .A2(_0375_));
 sg13g2_nor2_1 _3043_ (.A(_0381_),
    .B(_0385_),
    .Y(_0386_));
 sg13g2_and2_1 _3044_ (.A(_0339_),
    .B(_0386_),
    .X(_0387_));
 sg13g2_xnor2_1 _3045_ (.Y(_0388_),
    .A(_0021_),
    .B(_0387_));
 sg13g2_nand2_1 _3046_ (.Y(_0389_),
    .A(_1993_),
    .B(_0361_));
 sg13g2_nor2_1 _3047_ (.A(\videogen.draw_y[2] ),
    .B(_0387_),
    .Y(_0390_));
 sg13g2_and3_1 _3048_ (.X(_0391_),
    .A(_0362_),
    .B(_0388_),
    .C(_0389_));
 sg13g2_a21o_1 _3049_ (.A2(_0361_),
    .A1(_1993_),
    .B1(_0350_),
    .X(_0392_));
 sg13g2_a221oi_1 _3050_ (.B2(_0380_),
    .C1(_0392_),
    .B1(_0391_),
    .A1(_0362_),
    .Y(_0393_),
    .A2(_0390_));
 sg13g2_xor2_1 _3051_ (.B(_0328_),
    .A(\oscilloscope_control.n111_o[0] ),
    .X(_0394_));
 sg13g2_nand2_1 _3052_ (.Y(_0395_),
    .A(_0339_),
    .B(_0394_));
 sg13g2_xnor2_1 _3053_ (.Y(_0396_),
    .A(_0329_),
    .B(_0330_));
 sg13g2_nand2_1 _3054_ (.Y(_0397_),
    .A(net638),
    .B(_0396_));
 sg13g2_xnor2_1 _3055_ (.Y(_0398_),
    .A(_0023_),
    .B(_0397_));
 sg13g2_nor2_1 _3056_ (.A(_0048_),
    .B(_0349_),
    .Y(_0399_));
 sg13g2_xnor2_1 _3057_ (.Y(_0400_),
    .A(_0303_),
    .B(_0331_));
 sg13g2_nor2b_1 _3058_ (.A(_0400_),
    .B_N(net638),
    .Y(_0401_));
 sg13g2_and2_1 _3059_ (.A(net786),
    .B(_0401_),
    .X(_0402_));
 sg13g2_nand2_1 _3060_ (.Y(_0403_),
    .A(_1994_),
    .B(_0395_));
 sg13g2_a21oi_1 _3061_ (.A1(_0022_),
    .A2(_0395_),
    .Y(_0404_),
    .B1(_0399_));
 sg13g2_o21ai_1 _3062_ (.B1(_0404_),
    .Y(_0405_),
    .A1(_0022_),
    .A2(_0395_));
 sg13g2_o21ai_1 _3063_ (.B1(_0403_),
    .Y(_0406_),
    .A1(_0393_),
    .A2(_0405_));
 sg13g2_nor2b_1 _3064_ (.A(_0398_),
    .B_N(_0406_),
    .Y(_0407_));
 sg13g2_a221oi_1 _3065_ (.B2(net786),
    .C1(_0407_),
    .B1(_0401_),
    .A1(_1995_),
    .Y(_0408_),
    .A2(_0397_));
 sg13g2_nor2_1 _3066_ (.A(net786),
    .B(_0401_),
    .Y(_0409_));
 sg13g2_xnor2_1 _3067_ (.Y(_0410_),
    .A(_0332_),
    .B(_0333_));
 sg13g2_nor2b_1 _3068_ (.A(_0410_),
    .B_N(net638),
    .Y(_0411_));
 sg13g2_xnor2_1 _3069_ (.Y(_0412_),
    .A(_1997_),
    .B(_0411_));
 sg13g2_xnor2_1 _3070_ (.Y(_0413_),
    .A(_0334_),
    .B(_0335_));
 sg13g2_nand3_1 _3071_ (.B(net638),
    .C(_0413_),
    .A(\videogen.draw_y[9] ),
    .Y(_0414_));
 sg13g2_inv_1 _3072_ (.Y(_0415_),
    .A(_0414_));
 sg13g2_a21oi_1 _3073_ (.A1(net638),
    .A2(_0413_),
    .Y(_0416_),
    .B1(net785));
 sg13g2_nor3_2 _3074_ (.A(_0412_),
    .B(_0415_),
    .C(_0416_),
    .Y(_0417_));
 sg13g2_nand2b_1 _3075_ (.Y(_0418_),
    .B(_0417_),
    .A_N(_0409_));
 sg13g2_a21oi_1 _3076_ (.A1(_0025_),
    .A2(_0411_),
    .Y(_0419_),
    .B1(_0416_));
 sg13g2_or2_1 _3077_ (.X(_0420_),
    .B(_0419_),
    .A(_0415_));
 sg13g2_o21ai_1 _3078_ (.B1(_0420_),
    .Y(_0421_),
    .A1(_0408_),
    .A2(_0418_));
 sg13g2_nor2_1 _3079_ (.A(_2374_),
    .B(_0421_),
    .Y(_0422_));
 sg13g2_and2_1 _3080_ (.A(_2374_),
    .B(_0421_),
    .X(_0423_));
 sg13g2_xnor2_1 _3081_ (.Y(_0424_),
    .A(_0049_),
    .B(_2347_));
 sg13g2_nor4_1 _3082_ (.A(_0350_),
    .B(_0369_),
    .C(_0398_),
    .D(_0402_),
    .Y(_0425_));
 sg13g2_xnor2_1 _3083_ (.Y(_0426_),
    .A(\videogen.video_timing_generator.n21_o[0] ),
    .B(_0378_));
 sg13g2_nor3_1 _3084_ (.A(_0405_),
    .B(_0409_),
    .C(_0426_),
    .Y(_0427_));
 sg13g2_nand4_1 _3085_ (.B(_0417_),
    .C(_0425_),
    .A(_0391_),
    .Y(_0428_),
    .D(_0427_));
 sg13g2_nand3b_1 _3086_ (.B(_2325_),
    .C(_2361_),
    .Y(_0429_),
    .A_N(_2301_));
 sg13g2_nand3b_1 _3087_ (.B(_2362_),
    .C(_2370_),
    .Y(_0430_),
    .A_N(_2337_));
 sg13g2_nand4_1 _3088_ (.B(_2324_),
    .C(_2355_),
    .A(_2307_),
    .Y(_0431_),
    .D(_0424_));
 sg13g2_nor4_1 _3089_ (.A(_2303_),
    .B(_0429_),
    .C(_0430_),
    .D(_0431_),
    .Y(_0432_));
 sg13g2_nor3_1 _3090_ (.A(_0422_),
    .B(_0423_),
    .C(_0432_),
    .Y(_0433_));
 sg13g2_a21oi_2 _3091_ (.B1(_2069_),
    .Y(_0434_),
    .A2(_0433_),
    .A1(_0428_));
 sg13g2_xnor2_1 _3092_ (.Y(_0435_),
    .A(net785),
    .B(\choffset[4] ));
 sg13g2_nor2_2 _3093_ (.A(net381),
    .B(\display_x[9] ),
    .Y(_0436_));
 sg13g2_nor2_2 _3094_ (.A(net275),
    .B(net259),
    .Y(_0437_));
 sg13g2_and2_1 _3095_ (.A(_0436_),
    .B(_0437_),
    .X(_0438_));
 sg13g2_xor2_1 _3096_ (.B(\choffset[0] ),
    .A(\videogen.draw_y[5] ),
    .X(_0439_));
 sg13g2_nor4_2 _3097_ (.A(\videogen.draw_y[3] ),
    .B(\videogen.draw_y[2] ),
    .C(\videogen.draw_y[4] ),
    .Y(_0440_),
    .D(_2191_));
 sg13g2_xor2_1 _3098_ (.B(net740),
    .A(\videogen.draw_y[8] ),
    .X(_0441_));
 sg13g2_xnor2_1 _3099_ (.Y(_0442_),
    .A(\videogen.draw_y[6] ),
    .B(\choffset[1] ));
 sg13g2_nor2b_2 _3100_ (.A(net736),
    .B_N(_0438_),
    .Y(_0443_));
 sg13g2_nand4_1 _3101_ (.B(_0440_),
    .C(_0442_),
    .A(_0435_),
    .Y(_0444_),
    .D(_0443_));
 sg13g2_xor2_1 _3102_ (.B(net741),
    .A(\videogen.draw_y[7] ),
    .X(_0445_));
 sg13g2_nor4_2 _3103_ (.A(_0439_),
    .B(_0441_),
    .C(_0444_),
    .Y(_0446_),
    .D(_0445_));
 sg13g2_xor2_1 _3104_ (.B(net550),
    .A(net743),
    .X(_0447_));
 sg13g2_xnor2_1 _3105_ (.Y(_0448_),
    .A(_0015_),
    .B(_0447_));
 sg13g2_nor2_1 _3106_ (.A(net550),
    .B(net929),
    .Y(_0449_));
 sg13g2_nand2b_2 _3107_ (.Y(_0450_),
    .B(_0449_),
    .A_N(net743));
 sg13g2_o21ai_1 _3108_ (.B1(net929),
    .Y(_0451_),
    .A1(net743),
    .A2(net550));
 sg13g2_inv_1 _3109_ (.Y(_0452_),
    .A(_0451_));
 sg13g2_and2_1 _3110_ (.A(_0450_),
    .B(_0451_),
    .X(_0453_));
 sg13g2_nor2_1 _3111_ (.A(net737),
    .B(_0453_),
    .Y(_0454_));
 sg13g2_nor2_2 _3112_ (.A(net743),
    .B(_0449_),
    .Y(_0455_));
 sg13g2_xnor2_1 _3113_ (.Y(_0456_),
    .A(_0018_),
    .B(_0455_));
 sg13g2_a21oi_1 _3114_ (.A1(net743),
    .A2(net550),
    .Y(_0457_),
    .B1(net929));
 sg13g2_nor2_2 _3115_ (.A(_0447_),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_and2_1 _3116_ (.A(_0019_),
    .B(_0458_),
    .X(_0459_));
 sg13g2_nor2_1 _3117_ (.A(_0017_),
    .B(_0450_),
    .Y(_0460_));
 sg13g2_xnor2_1 _3118_ (.Y(_0461_),
    .A(\display_x[2] ),
    .B(net743));
 sg13g2_nand4_1 _3119_ (.B(_2001_),
    .C(_2213_),
    .A(net785),
    .Y(_0462_),
    .D(_0461_));
 sg13g2_nand2_1 _3120_ (.Y(_0463_),
    .A(net737),
    .B(_0453_));
 sg13g2_o21ai_1 _3121_ (.B1(_0463_),
    .Y(_0464_),
    .A1(_0019_),
    .A2(_0458_));
 sg13g2_nor4_1 _3122_ (.A(_0459_),
    .B(_0460_),
    .C(_0462_),
    .D(_0464_),
    .Y(_0465_));
 sg13g2_o21ai_1 _3123_ (.B1(_2083_),
    .Y(_0466_),
    .A1(_2202_),
    .A2(_0440_));
 sg13g2_nand2_1 _3124_ (.Y(_0467_),
    .A(_0020_),
    .B(_0452_));
 sg13g2_a22oi_1 _3125_ (.Y(_0468_),
    .B1(_0451_),
    .B2(_2040_),
    .A2(_0450_),
    .A1(_0017_));
 sg13g2_nand4_1 _3126_ (.B(_0466_),
    .C(_0467_),
    .A(_0465_),
    .Y(_0469_),
    .D(_0468_));
 sg13g2_nor4_2 _3127_ (.A(_0448_),
    .B(_0454_),
    .C(_0456_),
    .Y(_0470_),
    .D(_0469_));
 sg13g2_nand2b_1 _3128_ (.Y(_0471_),
    .B(\measurements.trigger.trigger_threshold[3] ),
    .A_N(net762));
 sg13g2_nor2_1 _3129_ (.A(net777),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_nor2_1 _3130_ (.A(_1989_),
    .B(net762),
    .Y(_0473_));
 sg13g2_a21oi_1 _3131_ (.A1(net777),
    .A2(_0473_),
    .Y(_0474_),
    .B1(_0472_));
 sg13g2_nor2b_1 _3132_ (.A(_0474_),
    .B_N(_2224_),
    .Y(_0475_));
 sg13g2_nand2_1 _3133_ (.Y(_0476_),
    .A(\choffset[4] ),
    .B(_0475_));
 sg13g2_or2_1 _3134_ (.X(_0477_),
    .B(_0474_),
    .A(net770));
 sg13g2_nor2_1 _3135_ (.A(_1986_),
    .B(net762),
    .Y(_0478_));
 sg13g2_nand2_1 _3136_ (.Y(_0479_),
    .A(net697),
    .B(_0478_));
 sg13g2_nand2b_1 _3137_ (.Y(_0480_),
    .B(\measurements.trigger.trigger_threshold[0] ),
    .A_N(net762));
 sg13g2_o21ai_1 _3138_ (.B1(_0479_),
    .Y(_0481_),
    .A1(net697),
    .A2(_0480_));
 sg13g2_a21oi_1 _3139_ (.A1(net770),
    .A2(_0481_),
    .Y(_0482_),
    .B1(net680));
 sg13g2_a221oi_1 _3140_ (.B2(_0482_),
    .C1(net678),
    .B1(_0477_),
    .A1(_0011_),
    .Y(_0483_),
    .A2(net686));
 sg13g2_nand2_1 _3141_ (.Y(_0484_),
    .A(net741),
    .B(_0483_));
 sg13g2_nand2_1 _3142_ (.Y(_0485_),
    .A(\measurements.trigger.trigger_threshold[3] ),
    .B(net674));
 sg13g2_a21oi_1 _3143_ (.A1(\measurements.trigger.trigger_threshold[2] ),
    .A2(net674),
    .Y(_0486_),
    .B1(net778));
 sg13g2_a21o_1 _3144_ (.A2(_0485_),
    .A1(net777),
    .B1(_0486_),
    .X(_0487_));
 sg13g2_nand2_1 _3145_ (.Y(_0488_),
    .A(net678),
    .B(_0487_));
 sg13g2_nor3_1 _3146_ (.A(_1989_),
    .B(net777),
    .C(net769),
    .Y(_0489_));
 sg13g2_a21oi_1 _3147_ (.A1(net777),
    .A2(_0478_),
    .Y(_0490_),
    .B1(_0489_));
 sg13g2_nor2_1 _3148_ (.A(_2268_),
    .B(_0480_),
    .Y(_0491_));
 sg13g2_nor2_1 _3149_ (.A(net686),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_o21ai_1 _3150_ (.B1(_0492_),
    .Y(_0493_),
    .A1(net770),
    .A2(_0490_));
 sg13g2_a21oi_1 _3151_ (.A1(_0010_),
    .A2(net680),
    .Y(_0494_),
    .B1(_2254_));
 sg13g2_nand3_1 _3152_ (.B(_0493_),
    .C(_0494_),
    .A(_0488_),
    .Y(_0495_));
 sg13g2_nor2_1 _3153_ (.A(_2026_),
    .B(_0495_),
    .Y(_0496_));
 sg13g2_nand2_1 _3154_ (.Y(_0497_),
    .A(\measurements.trigger.trigger_threshold[1] ),
    .B(net674));
 sg13g2_nand3_1 _3155_ (.B(net778),
    .C(net769),
    .A(\measurements.trigger.trigger_threshold[2] ),
    .Y(_0498_));
 sg13g2_o21ai_1 _3156_ (.B1(_0498_),
    .Y(_0499_),
    .A1(net778),
    .A2(_0497_));
 sg13g2_nor3_1 _3157_ (.A(_0042_),
    .B(_2268_),
    .C(_0485_),
    .Y(_0500_));
 sg13g2_nor2_1 _3158_ (.A(net776),
    .B(net678),
    .Y(_0501_));
 sg13g2_a221oi_1 _3159_ (.B2(_0481_),
    .C1(_0500_),
    .B1(_0501_),
    .A1(_2310_),
    .Y(_0502_),
    .A2(_0499_));
 sg13g2_nor2_1 _3160_ (.A(_2009_),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_xnor2_1 _3161_ (.Y(_0504_),
    .A(_2026_),
    .B(_0495_));
 sg13g2_inv_1 _3162_ (.Y(_0505_),
    .A(_0504_));
 sg13g2_a21oi_1 _3163_ (.A1(_0503_),
    .A2(_0505_),
    .Y(_0506_),
    .B1(_0496_));
 sg13g2_xnor2_1 _3164_ (.Y(_0507_),
    .A(net741),
    .B(_0483_));
 sg13g2_or2_1 _3165_ (.X(_0508_),
    .B(_0507_),
    .A(_0506_));
 sg13g2_nor2_1 _3166_ (.A(\oscilloscope_control.n114_o[0] ),
    .B(_0471_),
    .Y(_0509_));
 sg13g2_a21oi_1 _3167_ (.A1(net770),
    .A2(_0490_),
    .Y(_0510_),
    .B1(net686));
 sg13g2_o21ai_1 _3168_ (.B1(_0510_),
    .Y(_0511_),
    .A1(net770),
    .A2(_0509_));
 sg13g2_inv_1 _3169_ (.Y(_0512_),
    .A(_0511_));
 sg13g2_xnor2_1 _3170_ (.Y(_0513_),
    .A(_0041_),
    .B(_0511_));
 sg13g2_a21oi_1 _3171_ (.A1(_0484_),
    .A2(_0508_),
    .Y(_0514_),
    .B1(_0513_));
 sg13g2_a21oi_1 _3172_ (.A1(net739),
    .A2(_0512_),
    .Y(_0515_),
    .B1(_0514_));
 sg13g2_xnor2_1 _3173_ (.Y(_0516_),
    .A(\choffset[4] ),
    .B(_0475_));
 sg13g2_o21ai_1 _3174_ (.B1(_0476_),
    .Y(_0517_),
    .A1(_0515_),
    .A2(_0516_));
 sg13g2_nand2_1 _3175_ (.Y(_0518_),
    .A(_2224_),
    .B(_0509_));
 sg13g2_and2_1 _3176_ (.A(_0517_),
    .B(_0518_),
    .X(_0519_));
 sg13g2_and3_1 _3177_ (.X(_0520_),
    .A(_0484_),
    .B(_0508_),
    .C(_0513_));
 sg13g2_nor3_1 _3178_ (.A(_2041_),
    .B(_0514_),
    .C(_0520_),
    .Y(_0521_));
 sg13g2_o21ai_1 _3179_ (.B1(_2041_),
    .Y(_0522_),
    .A1(_0514_),
    .A2(_0520_));
 sg13g2_xor2_1 _3180_ (.B(_0507_),
    .A(_0506_),
    .X(_0523_));
 sg13g2_xnor2_1 _3181_ (.Y(_0524_),
    .A(_0503_),
    .B(_0504_));
 sg13g2_xnor2_1 _3182_ (.Y(_0525_),
    .A(\choffset[0] ),
    .B(_0502_));
 sg13g2_xnor2_1 _3183_ (.Y(_0526_),
    .A(_0022_),
    .B(_0525_));
 sg13g2_nand2_1 _3184_ (.Y(_0527_),
    .A(\measurements.trigger.trigger_threshold[0] ),
    .B(net674));
 sg13g2_nor2_1 _3185_ (.A(\oscilloscope_control.n114_o[0] ),
    .B(_0527_),
    .Y(_0528_));
 sg13g2_nor3_1 _3186_ (.A(\oscilloscope_control.n114_o[0] ),
    .B(_2255_),
    .C(_0527_),
    .Y(_0529_));
 sg13g2_nand2b_1 _3187_ (.Y(_0530_),
    .B(\videogen.draw_y[1] ),
    .A_N(_0529_));
 sg13g2_nor2b_1 _3188_ (.A(\videogen.draw_y[1] ),
    .B_N(_0529_),
    .Y(_0531_));
 sg13g2_nor4_2 _3189_ (.A(net407),
    .B(\display_x[2] ),
    .C(net736),
    .Y(_0532_),
    .D(\display_x[4] ));
 sg13g2_a21oi_1 _3190_ (.A1(_2213_),
    .A2(_0532_),
    .Y(_0533_),
    .B1(_2087_));
 sg13g2_nor2_1 _3191_ (.A(_2092_),
    .B(_0533_),
    .Y(_0534_));
 sg13g2_nor4_1 _3192_ (.A(\videogen.draw_y[0] ),
    .B(_0436_),
    .C(_0531_),
    .D(_0534_),
    .Y(_0535_));
 sg13g2_nand3_1 _3193_ (.B(net697),
    .C(net674),
    .A(\measurements.trigger.trigger_threshold[0] ),
    .Y(_0536_));
 sg13g2_o21ai_1 _3194_ (.B1(_0536_),
    .Y(_0537_),
    .A1(net697),
    .A2(_0497_));
 sg13g2_nand2_1 _3195_ (.Y(_0538_),
    .A(_2254_),
    .B(_0537_));
 sg13g2_xor2_1 _3196_ (.B(_0538_),
    .A(\videogen.draw_y[2] ),
    .X(_0539_));
 sg13g2_a22oi_1 _3197_ (.Y(_0540_),
    .B1(_0528_),
    .B2(_2310_),
    .A2(_0499_),
    .A1(_2254_));
 sg13g2_xnor2_1 _3198_ (.Y(_0541_),
    .A(_1993_),
    .B(_0540_));
 sg13g2_nand4_1 _3199_ (.B(_0535_),
    .C(_0539_),
    .A(_0530_),
    .Y(_0542_),
    .D(_0541_));
 sg13g2_a22oi_1 _3200_ (.Y(_0543_),
    .B1(_2252_),
    .B2(_0487_),
    .A2(_2222_),
    .A1(net765));
 sg13g2_o21ai_1 _3201_ (.B1(_0543_),
    .Y(_0544_),
    .A1(_2252_),
    .A2(_0537_));
 sg13g2_xnor2_1 _3202_ (.Y(_0545_),
    .A(_2060_),
    .B(_0544_));
 sg13g2_xor2_1 _3203_ (.B(_0516_),
    .A(_0515_),
    .X(_0546_));
 sg13g2_nor2_1 _3204_ (.A(_0517_),
    .B(_0518_),
    .Y(_0547_));
 sg13g2_xnor2_1 _3205_ (.Y(_0548_),
    .A(_0026_),
    .B(_0546_));
 sg13g2_xnor2_1 _3206_ (.Y(_0549_),
    .A(_0023_),
    .B(_0524_));
 sg13g2_nor4_1 _3207_ (.A(_0526_),
    .B(_0542_),
    .C(_0545_),
    .D(_0549_),
    .Y(_0550_));
 sg13g2_o21ai_1 _3208_ (.B1(_0550_),
    .Y(_0551_),
    .A1(net786),
    .A2(_0523_));
 sg13g2_a21oi_1 _3209_ (.A1(net786),
    .A2(_0523_),
    .Y(_0552_),
    .B1(_0551_));
 sg13g2_nand3b_1 _3210_ (.B(_0522_),
    .C(_0552_),
    .Y(_0553_),
    .A_N(_0521_));
 sg13g2_nor4_1 _3211_ (.A(_0519_),
    .B(_0547_),
    .C(_0548_),
    .D(_0553_),
    .Y(_0554_));
 sg13g2_nor4_2 _3212_ (.A(_0434_),
    .B(_0446_),
    .C(_0470_),
    .Y(_0555_),
    .D(_0554_));
 sg13g2_nor2_1 _3213_ (.A(_2216_),
    .B(_0555_),
    .Y(\videogen.b ));
 sg13g2_nand3_1 _3214_ (.B(\display_x[9] ),
    .C(_2086_),
    .A(\display_x[8] ),
    .Y(_0556_));
 sg13g2_nor2b_1 _3215_ (.A(_0018_),
    .B_N(_0556_),
    .Y(_0557_));
 sg13g2_nand3_1 _3216_ (.B(net737),
    .C(_0556_),
    .A(\display_x[4] ),
    .Y(_0558_));
 sg13g2_nor2b_1 _3217_ (.A(_0019_),
    .B_N(_0557_),
    .Y(_0559_));
 sg13g2_nand3b_1 _3218_ (.B(_0558_),
    .C(_0559_),
    .Y(_0560_),
    .A_N(_0017_));
 sg13g2_nor2_1 _3219_ (.A(_2092_),
    .B(_0560_),
    .Y(_0561_));
 sg13g2_xnor2_1 _3220_ (.Y(_0562_),
    .A(_0055_),
    .B(_0556_));
 sg13g2_nor2b_1 _3221_ (.A(_0561_),
    .B_N(_0562_),
    .Y(_0563_));
 sg13g2_nor2_1 _3222_ (.A(_0017_),
    .B(_0563_),
    .Y(_0564_));
 sg13g2_nand2_1 _3223_ (.Y(_0565_),
    .A(_0558_),
    .B(_0564_));
 sg13g2_xor2_1 _3224_ (.B(_0565_),
    .A(_0557_),
    .X(_0566_));
 sg13g2_a21oi_2 _3225_ (.B1(_0564_),
    .Y(_0567_),
    .A2(_0562_),
    .A1(_0017_));
 sg13g2_nand3b_1 _3226_ (.B(_0559_),
    .C(_0567_),
    .Y(_0568_),
    .A_N(net737));
 sg13g2_and2_1 _3227_ (.A(_2040_),
    .B(_0556_),
    .X(_0569_));
 sg13g2_nor2_1 _3228_ (.A(_0560_),
    .B(_0563_),
    .Y(_0570_));
 sg13g2_nor2_1 _3229_ (.A(_0055_),
    .B(_0560_),
    .Y(_0571_));
 sg13g2_nor3_1 _3230_ (.A(_2092_),
    .B(_0560_),
    .C(_0569_),
    .Y(_0572_));
 sg13g2_a22oi_1 _3231_ (.Y(_0573_),
    .B1(_0572_),
    .B2(_0562_),
    .A2(_0571_),
    .A1(_0569_));
 sg13g2_xnor2_1 _3232_ (.Y(_0574_),
    .A(_0569_),
    .B(_0570_));
 sg13g2_and2_1 _3233_ (.A(_0573_),
    .B(_0574_),
    .X(_0575_));
 sg13g2_a21oi_1 _3234_ (.A1(_0568_),
    .A2(_0575_),
    .Y(_0576_),
    .B1(net737));
 sg13g2_nand2_1 _3235_ (.Y(_0577_),
    .A(_0567_),
    .B(_0576_));
 sg13g2_xnor2_1 _3236_ (.Y(_0578_),
    .A(_0566_),
    .B(_0577_));
 sg13g2_a21o_1 _3237_ (.A2(_0575_),
    .A1(_0016_),
    .B1(_0576_),
    .X(_0579_));
 sg13g2_a21oi_1 _3238_ (.A1(_0568_),
    .A2(_0575_),
    .Y(_0580_),
    .B1(_2000_));
 sg13g2_xnor2_1 _3239_ (.Y(_0581_),
    .A(_0567_),
    .B(_0580_));
 sg13g2_nor2_1 _3240_ (.A(_0579_),
    .B(_0581_),
    .Y(_0582_));
 sg13g2_a21oi_1 _3241_ (.A1(\display_x[3] ),
    .A2(_0582_),
    .Y(_0583_),
    .B1(_0578_));
 sg13g2_nand3_1 _3242_ (.B(_0579_),
    .C(_0581_),
    .A(_1998_),
    .Y(_0584_));
 sg13g2_nand2_1 _3243_ (.Y(_0585_),
    .A(_0578_),
    .B(_0584_));
 sg13g2_o21ai_1 _3244_ (.B1(_0556_),
    .Y(_0586_),
    .A1(_0018_),
    .A2(_0565_));
 sg13g2_xor2_1 _3245_ (.B(_0586_),
    .A(_0019_),
    .X(_0587_));
 sg13g2_o21ai_1 _3246_ (.B1(_0587_),
    .Y(_0588_),
    .A1(_0566_),
    .A2(_0577_));
 sg13g2_and2_1 _3247_ (.A(_0568_),
    .B(_0588_),
    .X(_0589_));
 sg13g2_nor3_1 _3248_ (.A(\display_x[2] ),
    .B(_0583_),
    .C(_0589_),
    .Y(_0590_));
 sg13g2_nand2_1 _3249_ (.Y(_0591_),
    .A(_0585_),
    .B(_0590_));
 sg13g2_nor2_1 _3250_ (.A(_2039_),
    .B(_0578_),
    .Y(_0592_));
 sg13g2_o21ai_1 _3251_ (.B1(\display_x[2] ),
    .Y(_0593_),
    .A1(_0582_),
    .A2(_0592_));
 sg13g2_a22oi_1 _3252_ (.Y(_0594_),
    .B1(_0579_),
    .B2(_0581_),
    .A2(_0578_),
    .A1(_2039_));
 sg13g2_a21oi_1 _3253_ (.A1(\display_x[3] ),
    .A2(_0589_),
    .Y(_0595_),
    .B1(_0594_));
 sg13g2_o21ai_1 _3254_ (.B1(_0595_),
    .Y(_0596_),
    .A1(\display_x[3] ),
    .A2(_0589_));
 sg13g2_or2_1 _3255_ (.X(_0597_),
    .B(_0596_),
    .A(_0593_));
 sg13g2_a21oi_1 _3256_ (.A1(_0568_),
    .A2(_0573_),
    .Y(_0598_),
    .B1(_0575_));
 sg13g2_nand2b_1 _3257_ (.Y(_0599_),
    .B(_2213_),
    .A_N(_0598_));
 sg13g2_a21oi_2 _3258_ (.B1(_0599_),
    .Y(_0600_),
    .A2(_0597_),
    .A1(_0591_));
 sg13g2_and2_1 _3259_ (.A(_1994_),
    .B(_0440_),
    .X(_0601_));
 sg13g2_nor4_2 _3260_ (.A(_2085_),
    .B(net660),
    .C(_0600_),
    .Y(_0602_),
    .D(_0601_));
 sg13g2_nor2_1 _3261_ (.A(_2216_),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_a21oi_1 _3262_ (.A1(_0555_),
    .A2(_0602_),
    .Y(\videogen.r ),
    .B1(_2216_));
 sg13g2_and2_1 _3263_ (.A(_0555_),
    .B(_0603_),
    .X(\videogen.g ));
 sg13g2_nor2_1 _3264_ (.A(net470),
    .B(net310),
    .Y(_0604_));
 sg13g2_xnor2_1 _3265_ (.Y(_0605_),
    .A(net470),
    .B(net310));
 sg13g2_nor3_1 _3266_ (.A(_2064_),
    .B(\siggen.da_cs ),
    .C(_0605_),
    .Y(\siggen.da_mosi ));
 sg13g2_nor2_1 _3267_ (.A(net233),
    .B(net107),
    .Y(_0606_));
 sg13g2_nand2b_1 _3268_ (.Y(_0607_),
    .B(_0606_),
    .A_N(net425));
 sg13g2_xnor2_1 _3269_ (.Y(_0608_),
    .A(net425),
    .B(_0606_));
 sg13g2_mux2_1 _3270_ (.A0(_0608_),
    .A1(net425),
    .S(net262),
    .X(_0609_));
 sg13g2_nand3b_1 _3271_ (.B(net497),
    .C(net562),
    .Y(_0610_),
    .A_N(net197));
 sg13g2_and3_1 _3272_ (.X(_0611_),
    .A(net953),
    .B(_1981_),
    .C(_2167_));
 sg13g2_nor2_1 _3273_ (.A(_2077_),
    .B(_2180_),
    .Y(_0612_));
 sg13g2_o21ai_1 _3274_ (.B1(_0612_),
    .Y(_0613_),
    .A1(_2068_),
    .A2(_0611_));
 sg13g2_inv_2 _3275_ (.Y(_0614_),
    .A(net649));
 sg13g2_nor2_2 _3276_ (.A(_1981_),
    .B(net649),
    .Y(_0615_));
 sg13g2_nand2_1 _3277_ (.Y(_0616_),
    .A(net579),
    .B(_0614_));
 sg13g2_a21oi_1 _3278_ (.A1(_1982_),
    .A2(net646),
    .Y(_0617_),
    .B1(net197));
 sg13g2_nand2b_1 _3279_ (.Y(_0618_),
    .B(net497),
    .A_N(net425));
 sg13g2_or4_1 _3280_ (.A(_1982_),
    .B(net562),
    .C(net262),
    .D(_0607_),
    .X(_0619_));
 sg13g2_and2_1 _3281_ (.A(_0617_),
    .B(net563),
    .X(_0213_));
 sg13g2_nand2_2 _3282_ (.Y(_0620_),
    .A(_0610_),
    .B(_0213_));
 sg13g2_nor2_1 _3283_ (.A(net197),
    .B(_0619_),
    .Y(_0214_));
 sg13g2_a21oi_1 _3284_ (.A1(net497),
    .A2(_0609_),
    .Y(_0621_),
    .B1(_0620_));
 sg13g2_nor2b_1 _3285_ (.A(_2159_),
    .B_N(net322),
    .Y(_0622_));
 sg13g2_mux2_1 _3286_ (.A0(net427),
    .A1(_0622_),
    .S(net635),
    .X(_0093_));
 sg13g2_nor2b_1 _3287_ (.A(_2159_),
    .B_N(net427),
    .Y(_0623_));
 sg13g2_mux2_1 _3288_ (.A0(net399),
    .A1(_0623_),
    .S(net498),
    .X(_0094_));
 sg13g2_nor2b_1 _3289_ (.A(_2159_),
    .B_N(net399),
    .Y(_0624_));
 sg13g2_mux2_1 _3290_ (.A0(net305),
    .A1(net400),
    .S(net635),
    .X(_0095_));
 sg13g2_nand3_1 _3291_ (.B(_2160_),
    .C(net635),
    .A(net305),
    .Y(_0625_));
 sg13g2_o21ai_1 _3292_ (.B1(net306),
    .Y(_0096_),
    .A1(_1985_),
    .A2(net635));
 sg13g2_nor2_1 _3293_ (.A(net480),
    .B(_2159_),
    .Y(_0626_));
 sg13g2_mux2_1 _3294_ (.A0(net357),
    .A1(net481),
    .S(net635),
    .X(_0097_));
 sg13g2_nand3_1 _3295_ (.B(_2160_),
    .C(net635),
    .A(net357),
    .Y(_0627_));
 sg13g2_o21ai_1 _3296_ (.B1(net358),
    .Y(_0098_),
    .A1(_1988_),
    .A2(net635));
 sg13g2_nor2_1 _3297_ (.A(_1988_),
    .B(_2159_),
    .Y(_0628_));
 sg13g2_mux2_1 _3298_ (.A0(net345),
    .A1(_0628_),
    .S(net635),
    .X(_0099_));
 sg13g2_or2_1 _3299_ (.X(_0629_),
    .B(net870),
    .A(\settings_uart_printer.uart_tx_module.counter_reg[0] ));
 sg13g2_nor2_1 _3300_ (.A(\settings_uart_printer.uart_tx_module.counter_reg[2] ),
    .B(_0629_),
    .Y(_0630_));
 sg13g2_nor3_1 _3301_ (.A(net942),
    .B(net886),
    .C(_0629_),
    .Y(_0631_));
 sg13g2_nor2b_1 _3302_ (.A(net181),
    .B_N(_0631_),
    .Y(_0632_));
 sg13g2_nor2b_1 _3303_ (.A(net882),
    .B_N(_0632_),
    .Y(_0633_));
 sg13g2_nor2b_1 _3304_ (.A(net222),
    .B_N(_0633_),
    .Y(_0634_));
 sg13g2_nand2b_2 _3305_ (.Y(_0635_),
    .B(_0634_),
    .A_N(net151));
 sg13g2_nor3_2 _3306_ (.A(net352),
    .B(net876),
    .C(_0635_),
    .Y(_0636_));
 sg13g2_nand2b_2 _3307_ (.Y(_0637_),
    .B(_0636_),
    .A_N(net157));
 sg13g2_nor2_1 _3308_ (.A(net901),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_nor3_2 _3309_ (.A(\settings_uart_printer.uart_tx_module.datacnt_reg[0] ),
    .B(\settings_uart_printer.uart_tx_module.datacnt_reg[1] ),
    .C(net421),
    .Y(_0639_));
 sg13g2_nand2b_1 _3310_ (.Y(_0640_),
    .B(\settings_uart_printer.uart_tx_module.n88_q[1] ),
    .A_N(\settings_uart_printer.uart_tx_module.n88_q[0] ));
 sg13g2_a21oi_1 _3311_ (.A1(_0638_),
    .A2(net422),
    .Y(_0641_),
    .B1(_0640_));
 sg13g2_and2_2 _3312_ (.A(net594),
    .B(_2171_),
    .X(_0642_));
 sg13g2_inv_2 _3313_ (.Y(_0121_),
    .A(net595));
 sg13g2_and2_1 _3314_ (.A(net616),
    .B(_0638_),
    .X(_0643_));
 sg13g2_nor3_1 _3315_ (.A(net423),
    .B(net595),
    .C(_0643_),
    .Y(_0100_));
 sg13g2_and2_2 _3316_ (.A(net483),
    .B(_0643_),
    .X(_0644_));
 sg13g2_or2_2 _3317_ (.X(_0645_),
    .B(_0644_),
    .A(_2171_));
 sg13g2_inv_1 _3318_ (.Y(_0646_),
    .A(_0645_));
 sg13g2_nor2_1 _3319_ (.A(net483),
    .B(_0638_),
    .Y(_0647_));
 sg13g2_nor2_1 _3320_ (.A(_0645_),
    .B(net484),
    .Y(_0101_));
 sg13g2_nor2_2 _3321_ (.A(net799),
    .B(net793),
    .Y(_0648_));
 sg13g2_or2_1 _3322_ (.X(_0649_),
    .B(net793),
    .A(net798));
 sg13g2_nand2_2 _3323_ (.Y(_0650_),
    .A(_2032_),
    .B(_0648_));
 sg13g2_or3_1 _3324_ (.A(net789),
    .B(net984),
    .C(_0650_),
    .X(_0651_));
 sg13g2_nor2_1 _3325_ (.A(net500),
    .B(_0651_),
    .Y(_0652_));
 sg13g2_nor2_1 _3326_ (.A(_0121_),
    .B(net501),
    .Y(_0653_));
 sg13g2_a22oi_1 _3327_ (.Y(_0654_),
    .B1(_0653_),
    .B2(net199),
    .A2(_0121_),
    .A1(net798));
 sg13g2_inv_1 _3328_ (.Y(_0102_),
    .A(net200));
 sg13g2_and2_1 _3329_ (.A(net800),
    .B(net796),
    .X(_0655_));
 sg13g2_nand2_2 _3330_ (.Y(_0656_),
    .A(net799),
    .B(net793));
 sg13g2_nand2_2 _3331_ (.Y(_0657_),
    .A(_0649_),
    .B(_0656_));
 sg13g2_mux2_1 _3332_ (.A0(net793),
    .A1(_0657_),
    .S(net595),
    .X(_0103_));
 sg13g2_nor2_1 _3333_ (.A(_0121_),
    .B(_0650_),
    .Y(_0658_));
 sg13g2_o21ai_1 _3334_ (.B1(net791),
    .Y(_0659_),
    .A1(_0121_),
    .A2(_0649_));
 sg13g2_nand2b_1 _3335_ (.Y(_0104_),
    .B(net847),
    .A_N(_0658_));
 sg13g2_xnor2_1 _3336_ (.Y(_0105_),
    .A(net696),
    .B(_0658_));
 sg13g2_o21ai_1 _3337_ (.B1(net984),
    .Y(_0660_),
    .A1(net789),
    .A2(_0650_));
 sg13g2_and2_2 _3338_ (.A(_0651_),
    .B(_0660_),
    .X(_0661_));
 sg13g2_nand2_1 _3339_ (.Y(_0662_),
    .A(_0651_),
    .B(_0660_));
 sg13g2_a22oi_1 _3340_ (.Y(_0106_),
    .B1(_0653_),
    .B2(net652),
    .A2(_0121_),
    .A1(net141));
 sg13g2_nand3_1 _3341_ (.B(_0642_),
    .C(_0651_),
    .A(\settings_uart_printer.n103_q[5] ),
    .Y(_0663_));
 sg13g2_o21ai_1 _3342_ (.B1(_0663_),
    .Y(_0664_),
    .A1(net178),
    .A2(_0642_));
 sg13g2_inv_1 _3343_ (.Y(_0107_),
    .A(net179));
 sg13g2_nor4_2 _3344_ (.A(net901),
    .B(net616),
    .C(_0637_),
    .Y(_0665_),
    .D(net422));
 sg13g2_nor2_2 _3345_ (.A(_2171_),
    .B(_0665_),
    .Y(_0666_));
 sg13g2_nand2_2 _3346_ (.Y(_0667_),
    .A(net483),
    .B(_0665_));
 sg13g2_inv_1 _3347_ (.Y(_0668_),
    .A(_0667_));
 sg13g2_a22oi_1 _3348_ (.Y(_0669_),
    .B1(_0668_),
    .B2(\settings_uart_printer.uart_tx_module.datacnt_reg[0] ),
    .A2(_0666_),
    .A1(net61));
 sg13g2_inv_1 _3349_ (.Y(_0108_),
    .A(net62));
 sg13g2_nand2_1 _3350_ (.Y(_0670_),
    .A(net49),
    .B(_0666_));
 sg13g2_xnor2_1 _3351_ (.Y(_0671_),
    .A(\settings_uart_printer.uart_tx_module.datacnt_reg[0] ),
    .B(net895));
 sg13g2_o21ai_1 _3352_ (.B1(net50),
    .Y(_0109_),
    .A1(_0667_),
    .A2(net896));
 sg13g2_o21ai_1 _3353_ (.B1(net421),
    .Y(_0672_),
    .A1(net937),
    .A2(net895));
 sg13g2_nor2b_1 _3354_ (.A(_0667_),
    .B_N(_0672_),
    .Y(_0673_));
 sg13g2_a21o_1 _3355_ (.A2(_0666_),
    .A1(net112),
    .B1(_0673_),
    .X(_0110_));
 sg13g2_o21ai_1 _3356_ (.B1(_0121_),
    .Y(_0674_),
    .A1(_2171_),
    .A2(_0665_));
 sg13g2_nand2_1 _3357_ (.Y(_0675_),
    .A(net791),
    .B(_0649_));
 sg13g2_and2_1 _3358_ (.A(_0650_),
    .B(_0675_),
    .X(_0676_));
 sg13g2_a21oi_1 _3359_ (.A1(_2032_),
    .A2(_0648_),
    .Y(_0677_),
    .B1(net695));
 sg13g2_xnor2_1 _3360_ (.Y(_0678_),
    .A(net696),
    .B(_0650_));
 sg13g2_xnor2_1 _3361_ (.Y(_0679_),
    .A(net789),
    .B(_0650_));
 sg13g2_nand2_1 _3362_ (.Y(_0680_),
    .A(_0004_),
    .B(_0678_));
 sg13g2_nand2_1 _3363_ (.Y(_0681_),
    .A(net793),
    .B(net789));
 sg13g2_a21oi_1 _3364_ (.A1(_0680_),
    .A2(_0681_),
    .Y(_0682_),
    .B1(_0676_));
 sg13g2_nand2b_2 _3365_ (.Y(_0683_),
    .B(_0661_),
    .A_N(net1003));
 sg13g2_inv_1 _3366_ (.Y(_0684_),
    .A(_0683_));
 sg13g2_nor2b_1 _3367_ (.A(net790),
    .B_N(net794),
    .Y(_0685_));
 sg13g2_nand2_2 _3368_ (.Y(_0686_),
    .A(net793),
    .B(_2032_));
 sg13g2_nor3_2 _3369_ (.A(net791),
    .B(\settings_uart_printer.n103_q[3] ),
    .C(_0656_),
    .Y(_0687_));
 sg13g2_nor2_1 _3370_ (.A(net790),
    .B(_0657_),
    .Y(_0688_));
 sg13g2_nor3_1 _3371_ (.A(net790),
    .B(net695),
    .C(_0657_),
    .Y(_0689_));
 sg13g2_nor4_1 _3372_ (.A(_0682_),
    .B(_0683_),
    .C(_0687_),
    .D(_0689_),
    .Y(_0690_));
 sg13g2_nand2_1 _3373_ (.Y(_0691_),
    .A(net798),
    .B(_0003_));
 sg13g2_o21ai_1 _3374_ (.B1(_0691_),
    .Y(_0692_),
    .A1(net798),
    .A2(_0676_));
 sg13g2_a221oi_1 _3375_ (.B2(_0692_),
    .C1(_0661_),
    .B1(_0678_),
    .A1(_0675_),
    .Y(_0693_),
    .A2(_0677_));
 sg13g2_xor2_1 _3376_ (.B(_0660_),
    .A(\settings_uart_printer.n103_q[5] ),
    .X(_0694_));
 sg13g2_nand2_1 _3377_ (.Y(_0695_),
    .A(net794),
    .B(net695));
 sg13g2_nand2_1 _3378_ (.Y(_0696_),
    .A(net790),
    .B(_0657_));
 sg13g2_a21oi_1 _3379_ (.A1(_0695_),
    .A2(_0696_),
    .Y(_0697_),
    .B1(_0662_));
 sg13g2_nor3_1 _3380_ (.A(_0693_),
    .B(_0694_),
    .C(_0697_),
    .Y(_0698_));
 sg13g2_nor3_2 _3381_ (.A(net788),
    .B(_0690_),
    .C(_0698_),
    .Y(_0699_));
 sg13g2_nor2b_2 _3382_ (.A(net800),
    .B_N(net796),
    .Y(_0700_));
 sg13g2_nand2_1 _3383_ (.Y(_0701_),
    .A(net796),
    .B(\oscilloscope_control.n114_o[0] ));
 sg13g2_a22oi_1 _3384_ (.Y(_0702_),
    .B1(_0701_),
    .B2(net801),
    .A2(_0700_),
    .A1(\measurements.trigger.trigger_threshold[0] ));
 sg13g2_xnor2_1 _3385_ (.Y(_0703_),
    .A(net792),
    .B(net683));
 sg13g2_nor2_1 _3386_ (.A(_0006_),
    .B(_0656_),
    .Y(_0704_));
 sg13g2_xnor2_1 _3387_ (.Y(_0705_),
    .A(\settings_uart_printer.n103_q[3] ),
    .B(_0704_));
 sg13g2_xnor2_1 _3388_ (.Y(_0706_),
    .A(net696),
    .B(_0704_));
 sg13g2_and2_1 _3389_ (.A(_0703_),
    .B(_0706_),
    .X(_0707_));
 sg13g2_nand2b_1 _3390_ (.Y(_0708_),
    .B(_0707_),
    .A_N(_0702_));
 sg13g2_nor2b_2 _3391_ (.A(net797),
    .B_N(net800),
    .Y(_0709_));
 sg13g2_nand2b_1 _3392_ (.Y(_0710_),
    .B(net799),
    .A_N(net796));
 sg13g2_a22oi_1 _3393_ (.Y(_0711_),
    .B1(_0709_),
    .B2(_2035_),
    .A2(_0700_),
    .A1(_2030_));
 sg13g2_nand3_1 _3394_ (.B(_0705_),
    .C(_0711_),
    .A(_0703_),
    .Y(_0712_));
 sg13g2_nor2_2 _3395_ (.A(_0703_),
    .B(_0705_),
    .Y(_0713_));
 sg13g2_nor2_1 _3396_ (.A(net46),
    .B(_0656_),
    .Y(_0714_));
 sg13g2_a21oi_1 _3397_ (.A1(_0713_),
    .A2(_0714_),
    .Y(_0715_),
    .B1(_2008_));
 sg13g2_nor2_2 _3398_ (.A(_0703_),
    .B(_0706_),
    .Y(_0716_));
 sg13g2_a21oi_1 _3399_ (.A1(net800),
    .A2(net331),
    .Y(_0717_),
    .B1(net796));
 sg13g2_nor2_1 _3400_ (.A(net800),
    .B(\oscilloscope_control.n111_o[0] ),
    .Y(_0718_));
 sg13g2_o21ai_1 _3401_ (.B1(_0716_),
    .Y(_0719_),
    .A1(_0717_),
    .A2(_0718_));
 sg13g2_nand4_1 _3402_ (.B(_0712_),
    .C(_0715_),
    .A(_0708_),
    .Y(_0720_),
    .D(_0719_));
 sg13g2_nor2_1 _3403_ (.A(net688),
    .B(_0699_),
    .Y(_0721_));
 sg13g2_a221oi_1 _3404_ (.B2(_0721_),
    .C1(net642),
    .B1(net997),
    .A1(net122),
    .Y(_0722_),
    .A2(net688));
 sg13g2_a21oi_1 _3405_ (.A1(net115),
    .A2(net642),
    .Y(_0111_),
    .B1(_0722_));
 sg13g2_nor2_1 _3406_ (.A(\settings_uart_printer.n103_q[3] ),
    .B(_0710_),
    .Y(_0723_));
 sg13g2_nand2_1 _3407_ (.Y(_0724_),
    .A(net793),
    .B(net790));
 sg13g2_o21ai_1 _3408_ (.B1(_0649_),
    .Y(_0725_),
    .A1(net791),
    .A2(_0656_));
 sg13g2_a21oi_1 _3409_ (.A1(_0678_),
    .A2(_0725_),
    .Y(_0726_),
    .B1(_0689_));
 sg13g2_a221oi_1 _3410_ (.B2(net790),
    .C1(net652),
    .B1(_0723_),
    .A1(net794),
    .Y(_0727_),
    .A2(net789));
 sg13g2_a21oi_1 _3411_ (.A1(net652),
    .A2(_0726_),
    .Y(_0728_),
    .B1(_0727_));
 sg13g2_and3_1 _3412_ (.X(_0729_),
    .A(_0657_),
    .B(_0676_),
    .C(_0679_));
 sg13g2_o21ai_1 _3413_ (.B1(_0686_),
    .Y(_0730_),
    .A1(net794),
    .A2(net987));
 sg13g2_nor2_1 _3414_ (.A(_0679_),
    .B(_0730_),
    .Y(_0731_));
 sg13g2_nor3_1 _3415_ (.A(_0683_),
    .B(_0729_),
    .C(_0731_),
    .Y(_0732_));
 sg13g2_nor2_1 _3416_ (.A(net787),
    .B(_0732_),
    .Y(_0733_));
 sg13g2_o21ai_1 _3417_ (.B1(_0733_),
    .Y(_0734_),
    .A1(_0694_),
    .A2(_0728_));
 sg13g2_nand2_1 _3418_ (.Y(_0735_),
    .A(net695),
    .B(_0688_));
 sg13g2_nor2b_1 _3419_ (.A(net801),
    .B_N(\dsgfreqshift[1] ),
    .Y(_0736_));
 sg13g2_a21oi_1 _3420_ (.A1(net801),
    .A2(\oscilloscope_control.n220_q[1] ),
    .Y(_0737_),
    .B1(_0736_));
 sg13g2_a221oi_1 _3421_ (.B2(_1986_),
    .C1(_0705_),
    .B1(_0700_),
    .A1(net792),
    .Y(_0738_),
    .A2(_0009_));
 sg13g2_a221oi_1 _3422_ (.B2(_0008_),
    .C1(_0703_),
    .B1(_0709_),
    .A1(_0007_),
    .Y(_0739_),
    .A2(_0700_));
 sg13g2_nor3_1 _3423_ (.A(_0713_),
    .B(_0738_),
    .C(_0739_),
    .Y(_0740_));
 sg13g2_o21ai_1 _3424_ (.B1(_0740_),
    .Y(_0741_),
    .A1(_0735_),
    .A2(_0737_));
 sg13g2_nand2_1 _3425_ (.Y(_0742_),
    .A(net799),
    .B(net993));
 sg13g2_nand3_1 _3426_ (.B(_0713_),
    .C(_0742_),
    .A(net795),
    .Y(_0743_));
 sg13g2_nand3_1 _3427_ (.B(_0741_),
    .C(_0743_),
    .A(net787),
    .Y(_0744_));
 sg13g2_a21oi_1 _3428_ (.A1(_0734_),
    .A2(net994),
    .Y(_0745_),
    .B1(net688));
 sg13g2_a21oi_1 _3429_ (.A1(net195),
    .A2(net689),
    .Y(_0746_),
    .B1(_0745_));
 sg13g2_nand2_1 _3430_ (.Y(_0747_),
    .A(net122),
    .B(net641));
 sg13g2_o21ai_1 _3431_ (.B1(net123),
    .Y(_0112_),
    .A1(net641),
    .A2(_0746_));
 sg13g2_nand2_1 _3432_ (.Y(_0748_),
    .A(_0656_),
    .B(_0724_));
 sg13g2_a21oi_1 _3433_ (.A1(net652),
    .A2(_0748_),
    .Y(_0749_),
    .B1(_0678_));
 sg13g2_o21ai_1 _3434_ (.B1(_0749_),
    .Y(_0750_),
    .A1(net683),
    .A2(net652));
 sg13g2_o21ai_1 _3435_ (.B1(_0696_),
    .Y(_0751_),
    .A1(net798),
    .A2(_0686_));
 sg13g2_a21oi_1 _3436_ (.A1(_0678_),
    .A2(_0751_),
    .Y(_0752_),
    .B1(_0694_));
 sg13g2_o21ai_1 _3437_ (.B1(net789),
    .Y(_0753_),
    .A1(net798),
    .A2(_0685_));
 sg13g2_and2_1 _3438_ (.A(_0680_),
    .B(_0753_),
    .X(_0754_));
 sg13g2_a221oi_1 _3439_ (.B2(_0684_),
    .C1(net788),
    .B1(_0754_),
    .A1(_0750_),
    .Y(_0755_),
    .A2(_0752_));
 sg13g2_nand3_1 _3440_ (.B(_0703_),
    .C(_0705_),
    .A(_0657_),
    .Y(_0756_));
 sg13g2_a21oi_1 _3441_ (.A1(_0002_),
    .A2(net800),
    .Y(_0757_),
    .B1(net796));
 sg13g2_nor2b_1 _3442_ (.A(net800),
    .B_N(net741),
    .Y(_0758_));
 sg13g2_o21ai_1 _3443_ (.B1(_0716_),
    .Y(_0759_),
    .A1(_0757_),
    .A2(_0758_));
 sg13g2_a22oi_1 _3444_ (.Y(_0760_),
    .B1(_0700_),
    .B2(_2037_),
    .A2(_0655_),
    .A1(net762));
 sg13g2_nand2b_1 _3445_ (.Y(_0761_),
    .B(_0707_),
    .A_N(_0760_));
 sg13g2_nand3_1 _3446_ (.B(net929),
    .C(_0713_),
    .A(net795),
    .Y(_0762_));
 sg13g2_nand2_1 _3447_ (.Y(_0763_),
    .A(net788),
    .B(_0762_));
 sg13g2_nor3_1 _3448_ (.A(net799),
    .B(_2032_),
    .C(net695),
    .Y(_0764_));
 sg13g2_o21ai_1 _3449_ (.B1(_0764_),
    .Y(_0765_),
    .A1(\measurements.trigger.sample_on_rising_edge ),
    .A2(net797));
 sg13g2_nand4_1 _3450_ (.B(_0759_),
    .C(_0761_),
    .A(_0756_),
    .Y(_0766_),
    .D(_0765_));
 sg13g2_o21ai_1 _3451_ (.B1(_2171_),
    .Y(_0767_),
    .A1(_0763_),
    .A2(_0766_));
 sg13g2_nand2_1 _3452_ (.Y(_0768_),
    .A(net84),
    .B(net689));
 sg13g2_o21ai_1 _3453_ (.B1(_0768_),
    .Y(_0769_),
    .A1(_0755_),
    .A2(_0767_));
 sg13g2_mux2_1 _3454_ (.A0(_0769_),
    .A1(net195),
    .S(net641),
    .X(_0113_));
 sg13g2_a22oi_1 _3455_ (.Y(_0770_),
    .B1(_0657_),
    .B2(_0679_),
    .A2(net695),
    .A1(net793));
 sg13g2_a21oi_1 _3456_ (.A1(_2032_),
    .A2(_0723_),
    .Y(_0771_),
    .B1(_0683_));
 sg13g2_o21ai_1 _3457_ (.B1(_0771_),
    .Y(_0772_),
    .A1(_0685_),
    .A2(_0770_));
 sg13g2_nand2b_1 _3458_ (.Y(_0773_),
    .B(_0006_),
    .A_N(net798));
 sg13g2_a21oi_1 _3459_ (.A1(_0691_),
    .A2(_0773_),
    .Y(_0774_),
    .B1(_0679_));
 sg13g2_o21ai_1 _3460_ (.B1(net652),
    .Y(_0775_),
    .A1(_0729_),
    .A2(_0774_));
 sg13g2_nand2_2 _3461_ (.Y(_0776_),
    .A(net792),
    .B(_0709_));
 sg13g2_o21ai_1 _3462_ (.B1(_0776_),
    .Y(_0777_),
    .A1(net798),
    .A2(_0686_));
 sg13g2_o21ai_1 _3463_ (.B1(_0696_),
    .Y(_0778_),
    .A1(net792),
    .A2(net683));
 sg13g2_a22oi_1 _3464_ (.Y(_0779_),
    .B1(_0778_),
    .B2(_0679_),
    .A2(_0777_),
    .A1(net696));
 sg13g2_o21ai_1 _3465_ (.B1(_0775_),
    .Y(_0780_),
    .A1(net652),
    .A2(_0779_));
 sg13g2_o21ai_1 _3466_ (.B1(_0772_),
    .Y(_0781_),
    .A1(_0694_),
    .A2(_0780_));
 sg13g2_nand2_1 _3467_ (.Y(_0782_),
    .A(_2008_),
    .B(_0781_));
 sg13g2_a21oi_1 _3468_ (.A1(net796),
    .A2(net989),
    .Y(_0783_),
    .B1(net800));
 sg13g2_a21o_1 _3469_ (.A2(net796),
    .A1(net739),
    .B1(net683),
    .X(_0784_));
 sg13g2_a22oi_1 _3470_ (.Y(_0785_),
    .B1(_0784_),
    .B2(_0716_),
    .A2(_0783_),
    .A1(_0707_));
 sg13g2_o21ai_1 _3471_ (.B1(net787),
    .Y(_0786_),
    .A1(_0705_),
    .A2(_0776_));
 sg13g2_nor2b_1 _3472_ (.A(_0786_),
    .B_N(_0756_),
    .Y(_0787_));
 sg13g2_a21oi_1 _3473_ (.A1(_0785_),
    .A2(_0787_),
    .Y(_0788_),
    .B1(net689));
 sg13g2_a22oi_1 _3474_ (.Y(_0789_),
    .B1(_0782_),
    .B2(_0788_),
    .A2(net689),
    .A1(net67));
 sg13g2_nand2_1 _3475_ (.Y(_0790_),
    .A(net84),
    .B(net642));
 sg13g2_o21ai_1 _3476_ (.B1(net85),
    .Y(_0114_),
    .A1(net642),
    .A2(_0789_));
 sg13g2_a21oi_1 _3477_ (.A1(net792),
    .A2(_0700_),
    .Y(_0791_),
    .B1(_0687_));
 sg13g2_nand2_1 _3478_ (.Y(_0792_),
    .A(_0661_),
    .B(_0791_));
 sg13g2_nand2_1 _3479_ (.Y(_0793_),
    .A(net790),
    .B(net683));
 sg13g2_a22oi_1 _3480_ (.Y(_0794_),
    .B1(_0793_),
    .B2(net695),
    .A2(_0675_),
    .A1(_2034_));
 sg13g2_nand2_1 _3481_ (.Y(_0795_),
    .A(_0650_),
    .B(_0794_));
 sg13g2_a21oi_1 _3482_ (.A1(net652),
    .A2(_0795_),
    .Y(_0796_),
    .B1(_0694_));
 sg13g2_a21oi_1 _3483_ (.A1(net789),
    .A2(_0686_),
    .Y(_0797_),
    .B1(net683));
 sg13g2_a21oi_1 _3484_ (.A1(net792),
    .A2(net683),
    .Y(_0798_),
    .B1(_0797_));
 sg13g2_a221oi_1 _3485_ (.B2(_0684_),
    .C1(net788),
    .B1(_0798_),
    .A1(_0792_),
    .Y(_0799_),
    .A2(_0796_));
 sg13g2_a21oi_1 _3486_ (.A1(_0707_),
    .A2(_0710_),
    .Y(_0800_),
    .B1(_2008_));
 sg13g2_nand2_1 _3487_ (.Y(_0801_),
    .A(_0735_),
    .B(_0800_));
 sg13g2_a21oi_1 _3488_ (.A1(net917),
    .A2(_0648_),
    .Y(_0802_),
    .B1(_0703_));
 sg13g2_nor3_1 _3489_ (.A(_0716_),
    .B(_0801_),
    .C(_0802_),
    .Y(_0803_));
 sg13g2_nor3_1 _3490_ (.A(net688),
    .B(_0799_),
    .C(_0803_),
    .Y(_0804_));
 sg13g2_a21oi_1 _3491_ (.A1(net64),
    .A2(net689),
    .Y(_0805_),
    .B1(_0804_));
 sg13g2_nand2_1 _3492_ (.Y(_0806_),
    .A(net67),
    .B(net641));
 sg13g2_o21ai_1 _3493_ (.B1(net68),
    .Y(_0115_),
    .A1(net641),
    .A2(_0805_));
 sg13g2_nor2b_1 _3494_ (.A(_0688_),
    .B_N(_0724_),
    .Y(_0807_));
 sg13g2_a21oi_1 _3495_ (.A1(_0679_),
    .A2(_0807_),
    .Y(_0808_),
    .B1(_0723_));
 sg13g2_nor2_1 _3496_ (.A(_0661_),
    .B(_0808_),
    .Y(_0809_));
 sg13g2_a21o_1 _3497_ (.A2(_0724_),
    .A1(_0650_),
    .B1(_0678_),
    .X(_0810_));
 sg13g2_a21oi_1 _3498_ (.A1(_0661_),
    .A2(_0810_),
    .Y(_0811_),
    .B1(_0809_));
 sg13g2_o21ai_1 _3499_ (.B1(_0771_),
    .Y(_0812_),
    .A1(_0678_),
    .A2(_0730_));
 sg13g2_o21ai_1 _3500_ (.B1(net988),
    .Y(_0813_),
    .A1(_0694_),
    .A2(_0811_));
 sg13g2_nor2_1 _3501_ (.A(net787),
    .B(_0813_),
    .Y(_0814_));
 sg13g2_a21oi_1 _3502_ (.A1(net801),
    .A2(_0713_),
    .Y(_0815_),
    .B1(_0801_));
 sg13g2_o21ai_1 _3503_ (.B1(_0815_),
    .Y(_0816_),
    .A1(_0713_),
    .A2(_0778_));
 sg13g2_nor2_1 _3504_ (.A(net688),
    .B(_0814_),
    .Y(_0817_));
 sg13g2_a22oi_1 _3505_ (.Y(_0818_),
    .B1(_0816_),
    .B2(_0817_),
    .A2(net688),
    .A1(net70));
 sg13g2_nand2_1 _3506_ (.Y(_0819_),
    .A(net64),
    .B(net641));
 sg13g2_o21ai_1 _3507_ (.B1(net65),
    .Y(_0116_),
    .A1(net641),
    .A2(_0818_));
 sg13g2_nand2_1 _3508_ (.Y(_0820_),
    .A(net70),
    .B(net641));
 sg13g2_a21o_1 _3509_ (.A2(_0776_),
    .A1(_0686_),
    .B1(_0678_),
    .X(_0821_));
 sg13g2_nand3_1 _3510_ (.B(_0735_),
    .C(_0821_),
    .A(_0661_),
    .Y(_0822_));
 sg13g2_a22oi_1 _3511_ (.Y(_0823_),
    .B1(net683),
    .B2(net792),
    .A2(_0648_),
    .A1(net695));
 sg13g2_nor2_1 _3512_ (.A(_0694_),
    .B(_0823_),
    .Y(_0824_));
 sg13g2_a221oi_1 _3513_ (.B2(_0661_),
    .C1(_0809_),
    .B1(_0824_),
    .A1(_0694_),
    .Y(_0825_),
    .A2(_0822_));
 sg13g2_a22oi_1 _3514_ (.Y(_0826_),
    .B1(_0713_),
    .B2(net799),
    .A2(_0710_),
    .A1(_0703_));
 sg13g2_o21ai_1 _3515_ (.B1(_0826_),
    .Y(_0827_),
    .A1(_0648_),
    .A2(_0706_));
 sg13g2_a21oi_1 _3516_ (.A1(net787),
    .A2(_0827_),
    .Y(_0828_),
    .B1(net594));
 sg13g2_o21ai_1 _3517_ (.B1(_0828_),
    .Y(_0829_),
    .A1(net787),
    .A2(_0825_));
 sg13g2_o21ai_1 _3518_ (.B1(net71),
    .Y(_0117_),
    .A1(net688),
    .A2(net970));
 sg13g2_or2_1 _3519_ (.X(_0830_),
    .B(net960),
    .A(net930));
 sg13g2_and2_2 _3520_ (.A(_2085_),
    .B(net660),
    .X(_0831_));
 sg13g2_nand2_2 _3521_ (.Y(_0832_),
    .A(_2085_),
    .B(net660));
 sg13g2_and3_1 _3522_ (.X(_0833_),
    .A(net930),
    .B(net184),
    .C(net249));
 sg13g2_nand2_1 _3523_ (.Y(_0834_),
    .A(net228),
    .B(_0833_));
 sg13g2_nor3_1 _3524_ (.A(\oscilloscope_control.n208_o ),
    .B(net184),
    .C(net249),
    .Y(_0835_));
 sg13g2_nor2b_1 _3525_ (.A(net228),
    .B_N(net250),
    .Y(_0836_));
 sg13g2_a221oi_1 _3526_ (.B2(net228),
    .C1(_0836_),
    .B1(_0833_),
    .A1(_0830_),
    .Y(_0837_),
    .A2(_0832_));
 sg13g2_mux2_1 _3527_ (.A0(net249),
    .A1(net168),
    .S(_0837_),
    .X(_0118_));
 sg13g2_xor2_1 _3528_ (.B(net168),
    .A(net930),
    .X(_0838_));
 sg13g2_nand2_1 _3529_ (.Y(_0839_),
    .A(_0837_),
    .B(_0838_));
 sg13g2_xnor2_1 _3530_ (.Y(_0119_),
    .A(net184),
    .B(net931));
 sg13g2_o21ai_1 _3531_ (.B1(_0837_),
    .Y(_0840_),
    .A1(_0833_),
    .A2(net250));
 sg13g2_xnor2_1 _3532_ (.Y(_0120_),
    .A(net228),
    .B(net251));
 sg13g2_a21o_1 _3533_ (.A2(net501),
    .A1(net595),
    .B1(net787),
    .X(_0122_));
 sg13g2_nor2_2 _3534_ (.A(net292),
    .B(net569),
    .Y(_0841_));
 sg13g2_inv_1 _3535_ (.Y(_0842_),
    .A(net682));
 sg13g2_and2_1 _3536_ (.A(net40),
    .B(net570),
    .X(_0843_));
 sg13g2_nor2_1 _3537_ (.A(net148),
    .B(net265),
    .Y(_0844_));
 sg13g2_or2_1 _3538_ (.X(_0845_),
    .B(net265),
    .A(net148));
 sg13g2_nand3_1 _3539_ (.B(_0604_),
    .C(_0844_),
    .A(net256),
    .Y(_0846_));
 sg13g2_nand2b_1 _3540_ (.Y(_0847_),
    .B(_0846_),
    .A_N(net293));
 sg13g2_nand2b_1 _3541_ (.Y(_0123_),
    .B(_0847_),
    .A_N(net571));
 sg13g2_nor2_1 _3542_ (.A(net293),
    .B(_0846_),
    .Y(_0124_));
 sg13g2_o21ai_1 _3543_ (.B1(net229),
    .Y(_0125_),
    .A1(_2013_),
    .A2(_0836_));
 sg13g2_nand3_1 _3544_ (.B(net355),
    .C(net190),
    .A(net890),
    .Y(_0848_));
 sg13g2_nor3_1 _3545_ (.A(net890),
    .B(net355),
    .C(net190),
    .Y(_0849_));
 sg13g2_o21ai_1 _3546_ (.B1(net946),
    .Y(_0850_),
    .A1(_0832_),
    .A2(_0849_));
 sg13g2_o21ai_1 _3547_ (.B1(_0850_),
    .Y(_0851_),
    .A1(net946),
    .A2(_0848_));
 sg13g2_a21o_1 _3548_ (.A2(_0832_),
    .A1(net488),
    .B1(_0851_),
    .X(_0852_));
 sg13g2_mux2_1 _3549_ (.A0(net82),
    .A1(net890),
    .S(_0852_),
    .X(_0126_));
 sg13g2_xnor2_1 _3550_ (.Y(_0853_),
    .A(net488),
    .B(net82));
 sg13g2_nor2_1 _3551_ (.A(_0852_),
    .B(_0853_),
    .Y(_0854_));
 sg13g2_xor2_1 _3552_ (.B(_0854_),
    .A(net355),
    .X(_0127_));
 sg13g2_nand3_1 _3553_ (.B(net488),
    .C(net355),
    .A(net890),
    .Y(_0855_));
 sg13g2_or3_1 _3554_ (.A(net890),
    .B(net488),
    .C(net355),
    .X(_0856_));
 sg13g2_a21oi_1 _3555_ (.A1(_0855_),
    .A2(_0856_),
    .Y(_0857_),
    .B1(_0852_));
 sg13g2_xor2_1 _3556_ (.B(_0857_),
    .A(net190),
    .X(_0128_));
 sg13g2_or2_1 _3557_ (.X(_0858_),
    .B(_0848_),
    .A(net489));
 sg13g2_a22oi_1 _3558_ (.Y(_0129_),
    .B1(_0858_),
    .B2(_2012_),
    .A2(_0849_),
    .A1(net489));
 sg13g2_nor3_1 _3559_ (.A(net300),
    .B(net874),
    .C(net247),
    .Y(_0859_));
 sg13g2_nand2b_1 _3560_ (.Y(_0860_),
    .B(_0831_),
    .A_N(_0859_));
 sg13g2_nand3_1 _3561_ (.B(net874),
    .C(net247),
    .A(net300),
    .Y(_0861_));
 sg13g2_nor2_1 _3562_ (.A(net919),
    .B(_0861_),
    .Y(_0862_));
 sg13g2_a221oi_1 _3563_ (.B2(net919),
    .C1(_0862_),
    .B1(_0860_),
    .A1(net893),
    .Y(_0863_),
    .A2(_0832_));
 sg13g2_mux2_1 _3564_ (.A0(net874),
    .A1(net188),
    .S(_0863_),
    .X(_0130_));
 sg13g2_xor2_1 _3565_ (.B(net188),
    .A(net893),
    .X(_0864_));
 sg13g2_nand2_1 _3566_ (.Y(_0865_),
    .A(_0863_),
    .B(_0864_));
 sg13g2_xnor2_1 _3567_ (.Y(_0131_),
    .A(net300),
    .B(_0865_));
 sg13g2_and3_1 _3568_ (.X(_0866_),
    .A(net893),
    .B(net300),
    .C(net874));
 sg13g2_nor3_1 _3569_ (.A(net893),
    .B(net300),
    .C(net874),
    .Y(_0867_));
 sg13g2_o21ai_1 _3570_ (.B1(_0863_),
    .Y(_0868_),
    .A1(_0866_),
    .A2(_0867_));
 sg13g2_xnor2_1 _3571_ (.Y(_0132_),
    .A(net247),
    .B(_0868_));
 sg13g2_nor2b_1 _3572_ (.A(net893),
    .B_N(_0859_),
    .Y(_0869_));
 sg13g2_nand2_1 _3573_ (.Y(_0870_),
    .A(net247),
    .B(_0866_));
 sg13g2_o21ai_1 _3574_ (.B1(_0870_),
    .Y(_0133_),
    .A1(net164),
    .A2(_0869_));
 sg13g2_nand2_1 _3575_ (.Y(_0871_),
    .A(net278),
    .B(\oscilloscope_control.button_debouncer_n3_debounce_buttons.counter_reg[0] ));
 sg13g2_nand3_1 _3576_ (.B(net888),
    .C(net905),
    .A(net278),
    .Y(_0872_));
 sg13g2_nand4_1 _3577_ (.B(net888),
    .C(net231),
    .A(net278),
    .Y(_0873_),
    .D(net905));
 sg13g2_or3_1 _3578_ (.A(net278),
    .B(net888),
    .C(net905),
    .X(_0874_));
 sg13g2_or2_1 _3579_ (.X(_0875_),
    .B(_0874_),
    .A(net231));
 sg13g2_nand4_1 _3580_ (.B(_2097_),
    .C(_0873_),
    .A(_2085_),
    .Y(_0876_),
    .D(_0875_));
 sg13g2_mux2_1 _3581_ (.A0(net93),
    .A1(net888),
    .S(_0876_),
    .X(_0134_));
 sg13g2_xnor2_1 _3582_ (.Y(_0877_),
    .A(net905),
    .B(net93));
 sg13g2_nor2_1 _3583_ (.A(_0876_),
    .B(_0877_),
    .Y(_0878_));
 sg13g2_xor2_1 _3584_ (.B(_0878_),
    .A(net278),
    .X(_0135_));
 sg13g2_a21oi_1 _3585_ (.A1(_0872_),
    .A2(_0874_),
    .Y(_0879_),
    .B1(_0876_));
 sg13g2_xor2_1 _3586_ (.B(_0879_),
    .A(net231),
    .X(_0136_));
 sg13g2_nand2_1 _3587_ (.Y(_0880_),
    .A(net170),
    .B(_0875_));
 sg13g2_nand2_1 _3588_ (.Y(_0137_),
    .A(_0873_),
    .B(net171));
 sg13g2_nor3_1 _3589_ (.A(net283),
    .B(net872),
    .C(net350),
    .Y(_0881_));
 sg13g2_nand2b_1 _3590_ (.Y(_0882_),
    .B(_0831_),
    .A_N(_0881_));
 sg13g2_nand3_1 _3591_ (.B(net872),
    .C(net350),
    .A(net283),
    .Y(_0883_));
 sg13g2_nor2_1 _3592_ (.A(net911),
    .B(_0883_),
    .Y(_0884_));
 sg13g2_a221oi_1 _3593_ (.B2(net911),
    .C1(_0884_),
    .B1(_0882_),
    .A1(\oscilloscope_control.button_debouncer_n2_debounce_buttons.in_raw ),
    .Y(_0885_),
    .A2(_0832_));
 sg13g2_mux2_1 _3594_ (.A0(net872),
    .A1(net166),
    .S(_0885_),
    .X(_0138_));
 sg13g2_xor2_1 _3595_ (.B(net166),
    .A(\oscilloscope_control.button_debouncer_n2_debounce_buttons.in_raw ),
    .X(_0886_));
 sg13g2_nand2_1 _3596_ (.Y(_0887_),
    .A(net912),
    .B(_0886_));
 sg13g2_xnor2_1 _3597_ (.Y(_0139_),
    .A(net283),
    .B(net913));
 sg13g2_and3_1 _3598_ (.X(_0888_),
    .A(net923),
    .B(net283),
    .C(net872));
 sg13g2_nor3_1 _3599_ (.A(net923),
    .B(net283),
    .C(net872),
    .Y(_0889_));
 sg13g2_o21ai_1 _3600_ (.B1(net912),
    .Y(_0890_),
    .A1(_0888_),
    .A2(_0889_));
 sg13g2_xnor2_1 _3601_ (.Y(_0140_),
    .A(net350),
    .B(_0890_));
 sg13g2_nand2_2 _3602_ (.Y(_0891_),
    .A(net350),
    .B(_0888_));
 sg13g2_a22oi_1 _3603_ (.Y(_0141_),
    .B1(_0891_),
    .B2(net205),
    .A2(_0889_),
    .A1(_2007_));
 sg13g2_nor3_1 _3604_ (.A(net295),
    .B(net880),
    .C(net368),
    .Y(_0892_));
 sg13g2_a21oi_1 _3605_ (.A1(net939),
    .A2(_0892_),
    .Y(_0893_),
    .B1(_0831_));
 sg13g2_nor3_1 _3606_ (.A(net921),
    .B(net295),
    .C(net880),
    .Y(_0894_));
 sg13g2_nor2b_1 _3607_ (.A(net368),
    .B_N(_0894_),
    .Y(_0895_));
 sg13g2_nor2_1 _3608_ (.A(net939),
    .B(_2120_),
    .Y(_0896_));
 sg13g2_nor3_2 _3609_ (.A(_0893_),
    .B(_0895_),
    .C(_0896_),
    .Y(_0897_));
 sg13g2_mux2_1 _3610_ (.A0(net880),
    .A1(net202),
    .S(_0897_),
    .X(_0142_));
 sg13g2_xor2_1 _3611_ (.B(net202),
    .A(net921),
    .X(_0898_));
 sg13g2_nand2_1 _3612_ (.Y(_0899_),
    .A(_0897_),
    .B(_0898_));
 sg13g2_xnor2_1 _3613_ (.Y(_0143_),
    .A(net295),
    .B(net922));
 sg13g2_o21ai_1 _3614_ (.B1(_0897_),
    .Y(_0900_),
    .A1(_2121_),
    .A2(_0894_));
 sg13g2_xnor2_1 _3615_ (.Y(_0144_),
    .A(net368),
    .B(_0900_));
 sg13g2_o21ai_1 _3616_ (.B1(_2122_),
    .Y(_0145_),
    .A1(net270),
    .A2(_0895_));
 sg13g2_o21ai_1 _3617_ (.B1(_2124_),
    .Y(_0901_),
    .A1(net204),
    .A2(_0891_));
 sg13g2_nand2_2 _3618_ (.Y(_0902_),
    .A(net849),
    .B(_2013_));
 sg13g2_nand2b_1 _3619_ (.Y(_0903_),
    .B(_0901_),
    .A_N(net850));
 sg13g2_xnor2_1 _3620_ (.Y(_0904_),
    .A(net768),
    .B(_2124_));
 sg13g2_a21oi_2 _3621_ (.B1(_0903_),
    .Y(_0905_),
    .A2(_0904_),
    .A1(_2267_));
 sg13g2_a22oi_1 _3622_ (.Y(_0906_),
    .B1(_0905_),
    .B2(net600),
    .A2(_0903_),
    .A1(net783));
 sg13g2_inv_1 _3623_ (.Y(_0146_),
    .A(net601));
 sg13g2_xnor2_1 _3624_ (.Y(_0907_),
    .A(net773),
    .B(_2123_));
 sg13g2_xor2_1 _3625_ (.B(_0907_),
    .A(net600),
    .X(_0908_));
 sg13g2_a22oi_1 _3626_ (.Y(_0147_),
    .B1(_0905_),
    .B2(_0908_),
    .A2(_0903_),
    .A1(_2029_));
 sg13g2_nor2_1 _3627_ (.A(net768),
    .B(_0905_),
    .Y(_0909_));
 sg13g2_a22oi_1 _3628_ (.Y(_0910_),
    .B1(_0907_),
    .B2(net783),
    .A2(_2124_),
    .A1(_2036_));
 sg13g2_xnor2_1 _3629_ (.Y(_0911_),
    .A(_0904_),
    .B(net1006));
 sg13g2_a21oi_1 _3630_ (.A1(_0905_),
    .A2(_0911_),
    .Y(_0148_),
    .B1(net843));
 sg13g2_nand2_2 _3631_ (.Y(_0912_),
    .A(_2012_),
    .B(net927));
 sg13g2_nand2_2 _3632_ (.Y(_0913_),
    .A(net758),
    .B(net510));
 sg13g2_inv_1 _3633_ (.Y(_0914_),
    .A(_0913_));
 sg13g2_nand2_1 _3634_ (.Y(_0915_),
    .A(net586),
    .B(_0914_));
 sg13g2_nor3_2 _3635_ (.A(net204),
    .B(_2123_),
    .C(_0891_),
    .Y(_0916_));
 sg13g2_nor2_2 _3636_ (.A(net760),
    .B(net753),
    .Y(_0917_));
 sg13g2_nand2_1 _3637_ (.Y(_0918_),
    .A(net990),
    .B(_0917_));
 sg13g2_a22oi_1 _3638_ (.Y(_0919_),
    .B1(_0916_),
    .B2(_0918_),
    .A2(_0915_),
    .A1(net655));
 sg13g2_nor2_2 _3639_ (.A(_0912_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_mux2_1 _3640_ (.A0(net758),
    .A1(net331),
    .S(_0920_),
    .X(_0149_));
 sg13g2_xnor2_1 _3641_ (.Y(_0921_),
    .A(net331),
    .B(_2124_));
 sg13g2_nand2_1 _3642_ (.Y(_0922_),
    .A(_0920_),
    .B(_0921_));
 sg13g2_xnor2_1 _3643_ (.Y(_0150_),
    .A(net510),
    .B(_0922_));
 sg13g2_nor2b_2 _3644_ (.A(net752),
    .B_N(net758),
    .Y(_0923_));
 sg13g2_nor2b_1 _3645_ (.A(_0923_),
    .B_N(net966),
    .Y(_0924_));
 sg13g2_nor2_1 _3646_ (.A(net655),
    .B(_0924_),
    .Y(_0925_));
 sg13g2_a21oi_1 _3647_ (.A1(net655),
    .A2(_0913_),
    .Y(_0926_),
    .B1(_0925_));
 sg13g2_nand2_1 _3648_ (.Y(_0927_),
    .A(_0920_),
    .B(net967));
 sg13g2_xnor2_1 _3649_ (.Y(_0151_),
    .A(net586),
    .B(net968));
 sg13g2_nand2_2 _3650_ (.Y(_0928_),
    .A(_2126_),
    .B(_0916_));
 sg13g2_xnor2_1 _3651_ (.Y(_0152_),
    .A(net558),
    .B(_0928_));
 sg13g2_o21ai_1 _3652_ (.B1(net515),
    .Y(_0929_),
    .A1(_2035_),
    .A2(_0928_));
 sg13g2_nand2b_2 _3653_ (.Y(_0930_),
    .B(net558),
    .A_N(net515));
 sg13g2_o21ai_1 _3654_ (.B1(net516),
    .Y(_0153_),
    .A1(_0928_),
    .A2(_0930_));
 sg13g2_nor2_2 _3655_ (.A(net849),
    .B(net927),
    .Y(_0931_));
 sg13g2_nor2b_1 _3656_ (.A(_0901_),
    .B_N(_0931_),
    .Y(_0932_));
 sg13g2_nor2_2 _3657_ (.A(net170),
    .B(_0873_),
    .Y(_0933_));
 sg13g2_nand2b_2 _3658_ (.Y(_0934_),
    .B(_2016_),
    .A_N(_0873_));
 sg13g2_nor2_2 _3659_ (.A(net163),
    .B(_0870_),
    .Y(_0935_));
 sg13g2_nand3_1 _3660_ (.B(net668),
    .C(_0935_),
    .A(_0932_),
    .Y(_0936_));
 sg13g2_mux2_1 _3661_ (.A0(net917),
    .A1(net146),
    .S(_0936_),
    .X(_0154_));
 sg13g2_nand3_1 _3662_ (.B(_2162_),
    .C(_2164_),
    .A(_2074_),
    .Y(_0937_));
 sg13g2_inv_1 _3663_ (.Y(_0938_),
    .A(_0937_));
 sg13g2_nor3_2 _3664_ (.A(net588),
    .B(net733),
    .C(_2164_),
    .Y(_0939_));
 sg13g2_nand3_1 _3665_ (.B(net734),
    .C(net604),
    .A(net548),
    .Y(_0940_));
 sg13g2_nor2_2 _3666_ (.A(_2074_),
    .B(_2163_),
    .Y(_0941_));
 sg13g2_nand2_1 _3667_ (.Y(_0942_),
    .A(net609),
    .B(_2162_));
 sg13g2_and2_1 _3668_ (.A(net735),
    .B(_2075_),
    .X(_0943_));
 sg13g2_a21oi_1 _3669_ (.A1(net734),
    .A2(_2072_),
    .Y(_0944_),
    .B1(_0941_));
 sg13g2_a21oi_1 _3670_ (.A1(_0937_),
    .A2(_0944_),
    .Y(_0945_),
    .B1(net690));
 sg13g2_or2_1 _3671_ (.X(_0946_),
    .B(_0945_),
    .A(_2109_));
 sg13g2_nand2_1 _3672_ (.Y(_0947_),
    .A(net503),
    .B(net552));
 sg13g2_nor3_1 _3673_ (.A(net552),
    .B(_2071_),
    .C(_2076_),
    .Y(_0948_));
 sg13g2_nor2b_1 _3674_ (.A(net503),
    .B_N(net552),
    .Y(_0949_));
 sg13g2_a21oi_2 _3675_ (.B1(_0948_),
    .Y(_0950_),
    .A2(_0947_),
    .A1(_0946_));
 sg13g2_nand2_1 _3676_ (.Y(_0951_),
    .A(net504),
    .B(_0950_));
 sg13g2_and3_1 _3677_ (.X(_0952_),
    .A(net506),
    .B(net238),
    .C(net160));
 sg13g2_and3_1 _3678_ (.X(_0953_),
    .A(net210),
    .B(net692),
    .C(_0952_));
 sg13g2_or2_2 _3679_ (.X(_0954_),
    .B(_0950_),
    .A(net691));
 sg13g2_a21oi_1 _3680_ (.A1(net504),
    .A2(_0950_),
    .Y(_0155_),
    .B1(_0953_));
 sg13g2_nor3_2 _3681_ (.A(_1992_),
    .B(net733),
    .C(_2074_),
    .Y(_0955_));
 sg13g2_and2_1 _3682_ (.A(net225),
    .B(_0955_),
    .X(_0956_));
 sg13g2_inv_1 _3683_ (.Y(_0957_),
    .A(_0956_));
 sg13g2_nand2_2 _3684_ (.Y(_0958_),
    .A(_2158_),
    .B(_2159_));
 sg13g2_nor3_2 _3685_ (.A(\measurements.n246_q[0] ),
    .B(\measurements.n246_q[1] ),
    .C(\measurements.n246_q[2] ),
    .Y(_0959_));
 sg13g2_nor2b_1 _3686_ (.A(\measurements.n246_q[3] ),
    .B_N(_0959_),
    .Y(_0960_));
 sg13g2_and2_1 _3687_ (.A(_2004_),
    .B(_0960_),
    .X(_0961_));
 sg13g2_and2_1 _3688_ (.A(_2005_),
    .B(_0961_),
    .X(_0962_));
 sg13g2_nor2b_2 _3689_ (.A(\measurements.n246_q[6] ),
    .B_N(_0962_),
    .Y(_0963_));
 sg13g2_nand2b_2 _3690_ (.Y(_0964_),
    .B(_0963_),
    .A_N(\measurements.n246_q[7] ));
 sg13g2_nor3_2 _3691_ (.A(\measurements.n246_q[8] ),
    .B(\measurements.n246_q[9] ),
    .C(_0964_),
    .Y(_0965_));
 sg13g2_nand2b_2 _3692_ (.Y(_0966_),
    .B(_0965_),
    .A_N(\measurements.n246_q[10] ));
 sg13g2_nor3_2 _3693_ (.A(\measurements.n246_q[11] ),
    .B(net308),
    .C(_0966_),
    .Y(_0967_));
 sg13g2_o21ai_1 _3694_ (.B1(net308),
    .Y(_0968_),
    .A1(\measurements.n246_q[11] ),
    .A2(_0966_));
 sg13g2_nor2b_1 _3695_ (.A(_0967_),
    .B_N(_0968_),
    .Y(_0969_));
 sg13g2_xnor2_1 _3696_ (.Y(_0970_),
    .A(net909),
    .B(_0969_));
 sg13g2_nor2b_1 _3697_ (.A(net373),
    .B_N(_0967_),
    .Y(_0971_));
 sg13g2_xor2_1 _3698_ (.B(net253),
    .A(net949),
    .X(_0972_));
 sg13g2_nand2_1 _3699_ (.Y(_0973_),
    .A(_0971_),
    .B(_0972_));
 sg13g2_xor2_1 _3700_ (.B(_0966_),
    .A(net958),
    .X(_0974_));
 sg13g2_xnor2_1 _3701_ (.Y(_0975_),
    .A(net390),
    .B(_0974_));
 sg13g2_xnor2_1 _3702_ (.Y(_0976_),
    .A(net373),
    .B(_0967_));
 sg13g2_nor2b_1 _3703_ (.A(_0976_),
    .B_N(net903),
    .Y(_0977_));
 sg13g2_nor2b_1 _3704_ (.A(net903),
    .B_N(_0976_),
    .Y(_0978_));
 sg13g2_nor2_1 _3705_ (.A(_0971_),
    .B(_0972_),
    .Y(_0979_));
 sg13g2_xnor2_1 _3706_ (.Y(_0980_),
    .A(\measurements.n246_q[10] ),
    .B(_0965_));
 sg13g2_xnor2_1 _3707_ (.Y(_0981_),
    .A(net285),
    .B(_0980_));
 sg13g2_xnor2_1 _3708_ (.Y(_0982_),
    .A(\measurements.n246_q[1] ),
    .B(_0056_));
 sg13g2_nand2_1 _3709_ (.Y(_0983_),
    .A(net731),
    .B(\measurements.n246_q[0] ));
 sg13g2_o21ai_1 _3710_ (.B1(_0983_),
    .Y(_0984_),
    .A1(\measurements.n246_q[0] ),
    .A2(_0982_));
 sg13g2_a21oi_1 _3711_ (.A1(_2003_),
    .A2(_0982_),
    .Y(_0985_),
    .B1(_0984_));
 sg13g2_o21ai_1 _3712_ (.B1(\measurements.n246_q[2] ),
    .Y(_0986_),
    .A1(\measurements.n246_q[0] ),
    .A2(\measurements.n246_q[1] ));
 sg13g2_nor2b_1 _3713_ (.A(_0959_),
    .B_N(_0986_),
    .Y(_0987_));
 sg13g2_xnor2_1 _3714_ (.Y(_0988_),
    .A(_0057_),
    .B(_0987_));
 sg13g2_xnor2_1 _3715_ (.Y(_0989_),
    .A(\measurements.n246_q[3] ),
    .B(_0959_));
 sg13g2_xnor2_1 _3716_ (.Y(_0990_),
    .A(net449),
    .B(_0989_));
 sg13g2_xnor2_1 _3717_ (.Y(_0991_),
    .A(net235),
    .B(_0960_));
 sg13g2_xnor2_1 _3718_ (.Y(_0992_),
    .A(net473),
    .B(_0991_));
 sg13g2_nand4_1 _3719_ (.B(_0988_),
    .C(_0990_),
    .A(_0985_),
    .Y(_0993_),
    .D(_0992_));
 sg13g2_xnor2_1 _3720_ (.Y(_0994_),
    .A(_2005_),
    .B(_0961_));
 sg13g2_xnor2_1 _3721_ (.Y(_0995_),
    .A(net476),
    .B(_0994_));
 sg13g2_xor2_1 _3722_ (.B(_0962_),
    .A(\measurements.n246_q[6] ),
    .X(_0996_));
 sg13g2_xnor2_1 _3723_ (.Y(_0997_),
    .A(net432),
    .B(_0996_));
 sg13g2_xor2_1 _3724_ (.B(_0963_),
    .A(\measurements.n246_q[7] ),
    .X(_0998_));
 sg13g2_xnor2_1 _3725_ (.Y(_0999_),
    .A(_0062_),
    .B(_0998_));
 sg13g2_nor4_2 _3726_ (.A(_0993_),
    .B(_0995_),
    .C(_0997_),
    .Y(_1000_),
    .D(_0999_));
 sg13g2_xor2_1 _3727_ (.B(_0964_),
    .A(\measurements.n246_q[8] ),
    .X(_1001_));
 sg13g2_xnor2_1 _3728_ (.Y(_1002_),
    .A(net289),
    .B(_1001_));
 sg13g2_o21ai_1 _3729_ (.B1(\measurements.n246_q[9] ),
    .Y(_1003_),
    .A1(\measurements.n246_q[8] ),
    .A2(_0964_));
 sg13g2_nor2b_1 _3730_ (.A(_0965_),
    .B_N(_1003_),
    .Y(_1004_));
 sg13g2_xnor2_1 _3731_ (.Y(_1005_),
    .A(net302),
    .B(_1004_));
 sg13g2_nand4_1 _3732_ (.B(_1000_),
    .C(_1002_),
    .A(_0981_),
    .Y(_1006_),
    .D(_1005_));
 sg13g2_nor4_1 _3733_ (.A(_0977_),
    .B(_0978_),
    .C(_0979_),
    .D(_1006_),
    .Y(_1007_));
 sg13g2_nand4_1 _3734_ (.B(_0973_),
    .C(_0975_),
    .A(_0970_),
    .Y(_1008_),
    .D(_1007_));
 sg13g2_nor3_2 _3735_ (.A(net117),
    .B(_0958_),
    .C(net959),
    .Y(_0234_));
 sg13g2_nand3b_1 _3736_ (.B(_0970_),
    .C(_0973_),
    .Y(_1009_),
    .A_N(_0979_));
 sg13g2_nand2b_1 _3737_ (.Y(_1010_),
    .B(_0975_),
    .A_N(_1006_));
 sg13g2_or4_1 _3738_ (.A(_0977_),
    .B(_0978_),
    .C(_1009_),
    .D(_1010_),
    .X(_1011_));
 sg13g2_nor3_2 _3739_ (.A(net117),
    .B(_0958_),
    .C(_1011_),
    .Y(_1012_));
 sg13g2_o21ai_1 _3740_ (.B1(_0957_),
    .Y(_1013_),
    .A1(_2166_),
    .A2(_1012_));
 sg13g2_a21o_1 _3741_ (.A2(_1013_),
    .A1(net553),
    .B1(_0953_),
    .X(_0156_));
 sg13g2_nand2_1 _3742_ (.Y(_1014_),
    .A(_1989_),
    .B(_2124_));
 sg13g2_or4_1 _3743_ (.A(\measurements.trigger.trigger_threshold[0] ),
    .B(net999),
    .C(net534),
    .D(_1014_),
    .X(_1015_));
 sg13g2_nand2_1 _3744_ (.Y(_1016_),
    .A(net410),
    .B(net655));
 sg13g2_or4_1 _3745_ (.A(_1978_),
    .B(_1986_),
    .C(_1987_),
    .D(_1016_),
    .X(_1017_));
 sg13g2_nand4_1 _3746_ (.B(_0931_),
    .C(_1015_),
    .A(_0901_),
    .Y(_1018_),
    .D(_1017_));
 sg13g2_nand2_1 _3747_ (.Y(_1019_),
    .A(net34),
    .B(_1018_));
 sg13g2_o21ai_1 _3748_ (.B1(net35),
    .Y(_0157_),
    .A1(_1978_),
    .A2(_1018_));
 sg13g2_xnor2_1 _3749_ (.Y(_1020_),
    .A(net991),
    .B(net655));
 sg13g2_nand2_1 _3750_ (.Y(_1021_),
    .A(net975),
    .B(_1020_));
 sg13g2_xnor2_1 _3751_ (.Y(_1022_),
    .A(_1978_),
    .B(_1020_));
 sg13g2_nand2_1 _3752_ (.Y(_1023_),
    .A(net28),
    .B(_1018_));
 sg13g2_o21ai_1 _3753_ (.B1(net29),
    .Y(_0158_),
    .A1(_1018_),
    .A2(_1022_));
 sg13g2_nand2_1 _3754_ (.Y(_1024_),
    .A(net410),
    .B(_1018_));
 sg13g2_o21ai_1 _3755_ (.B1(_1021_),
    .Y(_1025_),
    .A1(_1986_),
    .A2(net655));
 sg13g2_nand2_1 _3756_ (.Y(_1026_),
    .A(_1014_),
    .B(_1016_));
 sg13g2_xnor2_1 _3757_ (.Y(_1027_),
    .A(_1025_),
    .B(_1026_));
 sg13g2_o21ai_1 _3758_ (.B1(net411),
    .Y(_0159_),
    .A1(_1018_),
    .A2(_1027_));
 sg13g2_or2_1 _3759_ (.X(_1028_),
    .B(_1021_),
    .A(_1016_));
 sg13g2_nand2_1 _3760_ (.Y(_1029_),
    .A(net973),
    .B(_2124_));
 sg13g2_a21o_1 _3761_ (.A2(_1026_),
    .A1(_1025_),
    .B1(_1029_),
    .X(_1030_));
 sg13g2_a21oi_1 _3762_ (.A1(_1028_),
    .A2(_1030_),
    .Y(_1031_),
    .B1(_1018_));
 sg13g2_xnor2_1 _3763_ (.Y(_0160_),
    .A(net535),
    .B(net974));
 sg13g2_nor3_2 _3764_ (.A(net463),
    .B(net440),
    .C(_2023_),
    .Y(_1032_));
 sg13g2_nor4_1 _3765_ (.A(net402),
    .B(net454),
    .C(net418),
    .D(net486),
    .Y(_1033_));
 sg13g2_nand4_1 _3766_ (.B(net565),
    .C(_1032_),
    .A(_2019_),
    .Y(_1034_),
    .D(_1033_));
 sg13g2_a21oi_1 _3767_ (.A1(_0935_),
    .A2(_1034_),
    .Y(_1035_),
    .B1(net672));
 sg13g2_nand4_1 _3768_ (.B(\oscilloscope_control.button_debouncer_n3_debounce_buttons.in_raw ),
    .C(_2016_),
    .A(net231),
    .Y(_1036_),
    .D(net567));
 sg13g2_nand4_1 _3769_ (.B(net463),
    .C(net440),
    .A(net486),
    .Y(_1037_),
    .D(_2023_));
 sg13g2_nand4_1 _3770_ (.B(net402),
    .C(net454),
    .A(net565),
    .Y(_1038_),
    .D(net418));
 sg13g2_nor4_1 _3771_ (.A(_0871_),
    .B(_1036_),
    .C(_1037_),
    .D(_1038_),
    .Y(_1039_));
 sg13g2_nor4_2 _3772_ (.A(_0901_),
    .B(_0912_),
    .C(_1035_),
    .Y(_1040_),
    .D(_1039_));
 sg13g2_a21oi_1 _3773_ (.A1(net655),
    .A2(_2126_),
    .Y(_1041_),
    .B1(_1040_));
 sg13g2_mux2_1 _3774_ (.A0(net651),
    .A1(net647),
    .S(net565),
    .X(_0161_));
 sg13g2_xnor2_1 _3775_ (.Y(_1042_),
    .A(net567),
    .B(net670));
 sg13g2_nand2_1 _3776_ (.Y(_1043_),
    .A(net565),
    .B(_1042_));
 sg13g2_o21ai_1 _3777_ (.B1(net651),
    .Y(_1044_),
    .A1(net565),
    .A2(_1042_));
 sg13g2_nor2b_1 _3778_ (.A(_1044_),
    .B_N(_1043_),
    .Y(_1045_));
 sg13g2_a21o_1 _3779_ (.A2(net647),
    .A1(net567),
    .B1(_1045_),
    .X(_0162_));
 sg13g2_o21ai_1 _3780_ (.B1(_1043_),
    .Y(_1046_),
    .A1(_2019_),
    .A2(net670));
 sg13g2_xnor2_1 _3781_ (.Y(_1047_),
    .A(net454),
    .B(net670));
 sg13g2_nand2_1 _3782_ (.Y(_1048_),
    .A(_1046_),
    .B(_1047_));
 sg13g2_o21ai_1 _3783_ (.B1(net651),
    .Y(_1049_),
    .A1(_1046_),
    .A2(_1047_));
 sg13g2_nor2b_1 _3784_ (.A(_1049_),
    .B_N(_1048_),
    .Y(_1050_));
 sg13g2_a21o_1 _3785_ (.A2(net647),
    .A1(net454),
    .B1(_1050_),
    .X(_0163_));
 sg13g2_o21ai_1 _3786_ (.B1(_1048_),
    .Y(_1051_),
    .A1(net1000),
    .A2(net670));
 sg13g2_xnor2_1 _3787_ (.Y(_1052_),
    .A(_2021_),
    .B(net670));
 sg13g2_xnor2_1 _3788_ (.Y(_1053_),
    .A(_1051_),
    .B(_1052_));
 sg13g2_a22oi_1 _3789_ (.Y(_1054_),
    .B1(_1053_),
    .B2(net651),
    .A2(net647),
    .A1(net402));
 sg13g2_inv_1 _3790_ (.Y(_0164_),
    .A(net403));
 sg13g2_a21oi_1 _3791_ (.A1(net402),
    .A2(_0934_),
    .Y(_1055_),
    .B1(_1051_));
 sg13g2_a21oi_1 _3792_ (.A1(_2021_),
    .A2(net670),
    .Y(_1056_),
    .B1(_1055_));
 sg13g2_xnor2_1 _3793_ (.Y(_1057_),
    .A(net486),
    .B(net670));
 sg13g2_nand2_1 _3794_ (.Y(_1058_),
    .A(_1056_),
    .B(_1057_));
 sg13g2_o21ai_1 _3795_ (.B1(net651),
    .Y(_1059_),
    .A1(_1056_),
    .A2(_1057_));
 sg13g2_nor2b_1 _3796_ (.A(_1059_),
    .B_N(_1058_),
    .Y(_1060_));
 sg13g2_a21o_1 _3797_ (.A2(net647),
    .A1(net486),
    .B1(_1060_),
    .X(_0165_));
 sg13g2_o21ai_1 _3798_ (.B1(_1058_),
    .Y(_1061_),
    .A1(net1001),
    .A2(net671));
 sg13g2_xnor2_1 _3799_ (.Y(_1062_),
    .A(_2022_),
    .B(net671));
 sg13g2_xnor2_1 _3800_ (.Y(_1063_),
    .A(_1061_),
    .B(_1062_));
 sg13g2_a22oi_1 _3801_ (.Y(_1064_),
    .B1(_1063_),
    .B2(net651),
    .A2(net647),
    .A1(net418));
 sg13g2_inv_1 _3802_ (.Y(_0166_),
    .A(net419));
 sg13g2_a21oi_1 _3803_ (.A1(net418),
    .A2(net668),
    .Y(_1065_),
    .B1(_1061_));
 sg13g2_a21oi_1 _3804_ (.A1(_2022_),
    .A2(net671),
    .Y(_1066_),
    .B1(_1065_));
 sg13g2_xnor2_1 _3805_ (.Y(_1067_),
    .A(net440),
    .B(net670));
 sg13g2_nand2_1 _3806_ (.Y(_1068_),
    .A(_1066_),
    .B(_1067_));
 sg13g2_o21ai_1 _3807_ (.B1(_1040_),
    .Y(_1069_),
    .A1(_1066_),
    .A2(_1067_));
 sg13g2_nor2b_1 _3808_ (.A(_1069_),
    .B_N(_1068_),
    .Y(_1070_));
 sg13g2_a21o_1 _3809_ (.A2(_1041_),
    .A1(net440),
    .B1(_1070_),
    .X(_0167_));
 sg13g2_o21ai_1 _3810_ (.B1(_1068_),
    .Y(_1071_),
    .A1(net965),
    .A2(net672));
 sg13g2_xnor2_1 _3811_ (.Y(_1072_),
    .A(net463),
    .B(net672));
 sg13g2_nand2_1 _3812_ (.Y(_1073_),
    .A(_1071_),
    .B(_1072_));
 sg13g2_o21ai_1 _3813_ (.B1(net651),
    .Y(_1074_),
    .A1(_1071_),
    .A2(_1072_));
 sg13g2_nor2b_1 _3814_ (.A(_1074_),
    .B_N(_1073_),
    .Y(_1075_));
 sg13g2_a21o_1 _3815_ (.A2(net647),
    .A1(net463),
    .B1(_1075_),
    .X(_0168_));
 sg13g2_o21ai_1 _3816_ (.B1(_1073_),
    .Y(_1076_),
    .A1(_0031_),
    .A2(net672));
 sg13g2_xnor2_1 _3817_ (.Y(_1077_),
    .A(net935),
    .B(net668));
 sg13g2_o21ai_1 _3818_ (.B1(net651),
    .Y(_1078_),
    .A1(_1076_),
    .A2(_1077_));
 sg13g2_a21oi_1 _3819_ (.A1(_1076_),
    .A2(_1077_),
    .Y(_1079_),
    .B1(_1078_));
 sg13g2_a21o_1 _3820_ (.A2(net647),
    .A1(net343),
    .B1(net936),
    .X(_0169_));
 sg13g2_nand2_2 _3821_ (.Y(_1080_),
    .A(_0932_),
    .B(net669));
 sg13g2_nand3_1 _3822_ (.B(net550),
    .C(net929),
    .A(net743),
    .Y(_1081_));
 sg13g2_nand2_1 _3823_ (.Y(_1082_),
    .A(net46),
    .B(_1081_));
 sg13g2_nand2_1 _3824_ (.Y(_1083_),
    .A(net743),
    .B(_1080_));
 sg13g2_o21ai_1 _3825_ (.B1(_1083_),
    .Y(_0170_),
    .A1(_1080_),
    .A2(net47));
 sg13g2_mux2_1 _3826_ (.A0(_0447_),
    .A1(net550),
    .S(_1080_),
    .X(_0171_));
 sg13g2_nor2b_1 _3827_ (.A(_0457_),
    .B_N(_1081_),
    .Y(_1084_));
 sg13g2_nand2_1 _3828_ (.Y(_1085_),
    .A(net43),
    .B(_1080_));
 sg13g2_o21ai_1 _3829_ (.B1(net44),
    .Y(_0172_),
    .A1(_1080_),
    .A2(_1084_));
 sg13g2_or2_1 _3830_ (.X(_1086_),
    .B(net884),
    .A(net360));
 sg13g2_a21oi_1 _3831_ (.A1(_0935_),
    .A2(_1086_),
    .Y(_1087_),
    .B1(net669));
 sg13g2_and2_1 _3832_ (.A(net360),
    .B(net884),
    .X(_1088_));
 sg13g2_and2_1 _3833_ (.A(net669),
    .B(_1088_),
    .X(_1089_));
 sg13g2_nor4_2 _3834_ (.A(_2125_),
    .B(_0901_),
    .C(_1087_),
    .Y(_1090_),
    .D(_1089_));
 sg13g2_mux2_1 _3835_ (.A0(net884),
    .A1(net176),
    .S(_1090_),
    .X(_0173_));
 sg13g2_xnor2_1 _3836_ (.Y(_1091_),
    .A(net176),
    .B(net668));
 sg13g2_nand2_1 _3837_ (.Y(_1092_),
    .A(_1090_),
    .B(_1091_));
 sg13g2_xnor2_1 _3838_ (.Y(_0174_),
    .A(net360),
    .B(_1092_));
 sg13g2_nor4_1 _3839_ (.A(\choffset[0] ),
    .B(net739),
    .C(net741),
    .D(\choffset[4] ),
    .Y(_1093_));
 sg13g2_nand2_1 _3840_ (.Y(_1094_),
    .A(_2026_),
    .B(_1093_));
 sg13g2_a21oi_1 _3841_ (.A1(_0935_),
    .A2(_1094_),
    .Y(_1095_),
    .B1(net669));
 sg13g2_nand3_1 _3842_ (.B(net582),
    .C(\choffset[4] ),
    .A(net933),
    .Y(_1096_));
 sg13g2_nor4_1 _3843_ (.A(net739),
    .B(net741),
    .C(net668),
    .D(_1096_),
    .Y(_1097_));
 sg13g2_or4_1 _3844_ (.A(_0901_),
    .B(_0902_),
    .C(_1095_),
    .D(_1097_),
    .X(_1098_));
 sg13g2_nor2_1 _3845_ (.A(net555),
    .B(net650),
    .Y(_1099_));
 sg13g2_a21oi_1 _3846_ (.A1(_2009_),
    .A2(net650),
    .Y(_0175_),
    .B1(net556));
 sg13g2_xnor2_1 _3847_ (.Y(_1100_),
    .A(net582),
    .B(_0933_));
 sg13g2_xnor2_1 _3848_ (.Y(_1101_),
    .A(net555),
    .B(_1100_));
 sg13g2_nor2_1 _3849_ (.A(_1098_),
    .B(_1101_),
    .Y(_1102_));
 sg13g2_a21oi_1 _3850_ (.A1(net583),
    .A2(net650),
    .Y(_0176_),
    .B1(_1102_));
 sg13g2_and2_1 _3851_ (.A(net741),
    .B(net668),
    .X(_1103_));
 sg13g2_xnor2_1 _3852_ (.Y(_1104_),
    .A(net741),
    .B(net669));
 sg13g2_o21ai_1 _3853_ (.B1(net933),
    .Y(_1105_),
    .A1(net582),
    .A2(net668));
 sg13g2_o21ai_1 _3854_ (.B1(_1105_),
    .Y(_1106_),
    .A1(_2026_),
    .A2(net669));
 sg13g2_nor2_1 _3855_ (.A(_1104_),
    .B(_1106_),
    .Y(_1107_));
 sg13g2_and2_1 _3856_ (.A(_1104_),
    .B(_1106_),
    .X(_1108_));
 sg13g2_nor3_1 _3857_ (.A(net650),
    .B(_1107_),
    .C(_1108_),
    .Y(_1109_));
 sg13g2_a21oi_1 _3858_ (.A1(net96),
    .A2(net650),
    .Y(_0177_),
    .B1(_1109_));
 sg13g2_xnor2_1 _3859_ (.Y(_1110_),
    .A(net592),
    .B(net669));
 sg13g2_o21ai_1 _3860_ (.B1(_1110_),
    .Y(_1111_),
    .A1(_1103_),
    .A2(_1108_));
 sg13g2_or3_1 _3861_ (.A(_1103_),
    .B(_1108_),
    .C(_1110_),
    .X(_1112_));
 sg13g2_a21oi_1 _3862_ (.A1(_1111_),
    .A2(_1112_),
    .Y(_1113_),
    .B1(net650));
 sg13g2_a21oi_1 _3863_ (.A1(_2027_),
    .A2(net650),
    .Y(_0178_),
    .B1(_1113_));
 sg13g2_nand3_1 _3864_ (.B(net669),
    .C(_1108_),
    .A(net739),
    .Y(_1114_));
 sg13g2_nand3_1 _3865_ (.B(net668),
    .C(_1111_),
    .A(net544),
    .Y(_1115_));
 sg13g2_a21oi_1 _3866_ (.A1(_1114_),
    .A2(net545),
    .Y(_1116_),
    .B1(net650));
 sg13g2_xor2_1 _3867_ (.B(net546),
    .A(net928),
    .X(_0179_));
 sg13g2_nand2_2 _3868_ (.Y(_1117_),
    .A(net506),
    .B(net692));
 sg13g2_and2_1 _3869_ (.A(_0954_),
    .B(_1117_),
    .X(_1118_));
 sg13g2_o21ai_1 _3870_ (.B1(net634),
    .Y(_1119_),
    .A1(net340),
    .A2(_0951_));
 sg13g2_a21oi_1 _3871_ (.A1(_2063_),
    .A2(net692),
    .Y(_0180_),
    .B1(net341));
 sg13g2_nand2_1 _3872_ (.Y(_1120_),
    .A(net738),
    .B(_2194_));
 sg13g2_xnor2_1 _3873_ (.Y(_0181_),
    .A(_1999_),
    .B(_2194_));
 sg13g2_xnor2_1 _3874_ (.Y(_0182_),
    .A(net405),
    .B(_1120_));
 sg13g2_nand2_1 _3875_ (.Y(_1121_),
    .A(net900),
    .B(net653));
 sg13g2_nand2_1 _3876_ (.Y(_1122_),
    .A(_2039_),
    .B(_2089_));
 sg13g2_xnor2_1 _3877_ (.Y(_1123_),
    .A(net443),
    .B(_2089_));
 sg13g2_nor3_1 _3878_ (.A(net736),
    .B(net381),
    .C(_2001_),
    .Y(_1124_));
 sg13g2_and4_1 _3879_ (.A(_2089_),
    .B(_2215_),
    .C(_0437_),
    .D(_1124_),
    .X(_1125_));
 sg13g2_nand2b_2 _3880_ (.Y(_1126_),
    .B(_2194_),
    .A_N(_1125_));
 sg13g2_o21ai_1 _3881_ (.B1(_1121_),
    .Y(_0183_),
    .A1(net444),
    .A2(_1126_));
 sg13g2_nand2_1 _3882_ (.Y(_1127_),
    .A(net407),
    .B(net653));
 sg13g2_xnor2_1 _3883_ (.Y(_1128_),
    .A(net910),
    .B(_1122_));
 sg13g2_o21ai_1 _3884_ (.B1(net408),
    .Y(_0184_),
    .A1(_1126_),
    .A2(_1128_));
 sg13g2_nand2_1 _3885_ (.Y(_1129_),
    .A(net518),
    .B(net653));
 sg13g2_nor2_1 _3886_ (.A(net737),
    .B(_2090_),
    .Y(_1130_));
 sg13g2_xnor2_1 _3887_ (.Y(_1131_),
    .A(net737),
    .B(_2090_));
 sg13g2_o21ai_1 _3888_ (.B1(net519),
    .Y(_0185_),
    .A1(_1126_),
    .A2(_1131_));
 sg13g2_nand2_1 _3889_ (.Y(_1132_),
    .A(net522),
    .B(net653));
 sg13g2_xor2_1 _3890_ (.B(_1130_),
    .A(net947),
    .X(_1133_));
 sg13g2_o21ai_1 _3891_ (.B1(net523),
    .Y(_0186_),
    .A1(_1126_),
    .A2(net948));
 sg13g2_nand2_1 _3892_ (.Y(_1134_),
    .A(net275),
    .B(net653));
 sg13g2_nand3_1 _3893_ (.B(net518),
    .C(_2091_),
    .A(net522),
    .Y(_1135_));
 sg13g2_nor2_1 _3894_ (.A(net951),
    .B(_1135_),
    .Y(_1136_));
 sg13g2_xnor2_1 _3895_ (.Y(_1137_),
    .A(net951),
    .B(_1135_));
 sg13g2_o21ai_1 _3896_ (.B1(net276),
    .Y(_0187_),
    .A1(_1126_),
    .A2(_1137_));
 sg13g2_nand2_1 _3897_ (.Y(_1138_),
    .A(net259),
    .B(net653));
 sg13g2_xor2_1 _3898_ (.B(_1136_),
    .A(net952),
    .X(_1139_));
 sg13g2_o21ai_1 _3899_ (.B1(net260),
    .Y(_0188_),
    .A1(_1126_),
    .A2(_1139_));
 sg13g2_nand2_1 _3900_ (.Y(_1140_),
    .A(net381),
    .B(net653));
 sg13g2_o21ai_1 _3901_ (.B1(net892),
    .Y(_1141_),
    .A1(_2087_),
    .A2(_1135_));
 sg13g2_nand3b_1 _3902_ (.B(_2040_),
    .C(_2086_),
    .Y(_1142_),
    .A_N(_1135_));
 sg13g2_nand2_1 _3903_ (.Y(_1143_),
    .A(_1141_),
    .B(_1142_));
 sg13g2_o21ai_1 _3904_ (.B1(net382),
    .Y(_0189_),
    .A1(_1126_),
    .A2(_1143_));
 sg13g2_a21oi_1 _3905_ (.A1(net540),
    .A2(_1142_),
    .Y(_1144_),
    .B1(_1126_));
 sg13g2_o21ai_1 _3906_ (.B1(net541),
    .Y(_1145_),
    .A1(net540),
    .A2(_1142_));
 sg13g2_o21ai_1 _3907_ (.B1(net542),
    .Y(_0190_),
    .A1(_2001_),
    .A2(_2194_));
 sg13g2_o21ai_1 _3908_ (.B1(_0617_),
    .Y(_1146_),
    .A1(net262),
    .A2(_0618_));
 sg13g2_nand2_1 _3909_ (.Y(_1147_),
    .A(net5),
    .B(_2160_));
 sg13g2_nand2_1 _3910_ (.Y(_1148_),
    .A(net322),
    .B(_1146_));
 sg13g2_o21ai_1 _3911_ (.B1(net323),
    .Y(_0191_),
    .A1(_1146_),
    .A2(_1147_));
 sg13g2_nand2_1 _3912_ (.Y(_1149_),
    .A(_2115_),
    .B(_0958_));
 sg13g2_o21ai_1 _3913_ (.B1(_2158_),
    .Y(_1150_),
    .A1(_1984_),
    .A2(_2155_));
 sg13g2_nand2_1 _3914_ (.Y(_1151_),
    .A(_1149_),
    .B(_1150_));
 sg13g2_nor3_1 _3915_ (.A(_1984_),
    .B(_2155_),
    .C(_0958_),
    .Y(_1152_));
 sg13g2_a22oi_1 _3916_ (.Y(_1153_),
    .B1(net639),
    .B2(net731),
    .A2(net636),
    .A1(net512));
 sg13g2_inv_1 _3917_ (.Y(_0192_),
    .A(net513));
 sg13g2_a22oi_1 _3918_ (.Y(_1154_),
    .B1(net639),
    .B2(net415),
    .A2(net636),
    .A1(net452));
 sg13g2_inv_1 _3919_ (.Y(_0193_),
    .A(net453));
 sg13g2_a22oi_1 _3920_ (.Y(_1155_),
    .B1(net639),
    .B2(\measurements.address_counter_reg[2] ),
    .A2(net636),
    .A1(net370));
 sg13g2_inv_1 _3921_ (.Y(_0194_),
    .A(net371));
 sg13g2_a22oi_1 _3922_ (.Y(_1156_),
    .B1(net639),
    .B2(net365),
    .A2(net636),
    .A1(\measurements.n246_q[3] ));
 sg13g2_inv_1 _3923_ (.Y(_0195_),
    .A(net366));
 sg13g2_a22oi_1 _3924_ (.Y(_1157_),
    .B1(net639),
    .B2(\measurements.address_counter_reg[4] ),
    .A2(net636),
    .A1(net235));
 sg13g2_inv_1 _3925_ (.Y(_0196_),
    .A(net236));
 sg13g2_a22oi_1 _3926_ (.Y(_1158_),
    .B1(net639),
    .B2(\measurements.address_counter_reg[5] ),
    .A2(net636),
    .A1(net154));
 sg13g2_inv_1 _3927_ (.Y(_0197_),
    .A(net155));
 sg13g2_a22oi_1 _3928_ (.Y(_1159_),
    .B1(net639),
    .B2(net394),
    .A2(net636),
    .A1(\measurements.n246_q[6] ));
 sg13g2_inv_1 _3929_ (.Y(_0198_),
    .A(net395));
 sg13g2_a22oi_1 _3930_ (.Y(_1160_),
    .B1(net639),
    .B2(net325),
    .A2(net636),
    .A1(\measurements.n246_q[7] ));
 sg13g2_inv_1 _3931_ (.Y(_0199_),
    .A(net326));
 sg13g2_a22oi_1 _3932_ (.Y(_1161_),
    .B1(net640),
    .B2(net207),
    .A2(net637),
    .A1(\measurements.n246_q[8] ));
 sg13g2_inv_1 _3933_ (.Y(_0200_),
    .A(net208));
 sg13g2_a22oi_1 _3934_ (.Y(_1162_),
    .B1(net640),
    .B2(net219),
    .A2(net637),
    .A1(\measurements.n246_q[9] ));
 sg13g2_inv_1 _3935_ (.Y(_0201_),
    .A(net220));
 sg13g2_a22oi_1 _3936_ (.Y(_1163_),
    .B1(net640),
    .B2(net213),
    .A2(net637),
    .A1(\measurements.n246_q[10] ));
 sg13g2_inv_1 _3937_ (.Y(_0202_),
    .A(net214));
 sg13g2_a22oi_1 _3938_ (.Y(_1164_),
    .B1(net640),
    .B2(net101),
    .A2(net637),
    .A1(\measurements.n246_q[11] ));
 sg13g2_inv_1 _3939_ (.Y(_0203_),
    .A(net102));
 sg13g2_a22oi_1 _3940_ (.Y(_1165_),
    .B1(net640),
    .B2(net297),
    .A2(net637),
    .A1(net308));
 sg13g2_inv_1 _3941_ (.Y(_0204_),
    .A(net309));
 sg13g2_a22oi_1 _3942_ (.Y(_1166_),
    .B1(net640),
    .B2(net362),
    .A2(net637),
    .A1(net373));
 sg13g2_inv_1 _3943_ (.Y(_0205_),
    .A(net374));
 sg13g2_a22oi_1 _3944_ (.Y(_1167_),
    .B1(net640),
    .B2(\measurements.address_counter_reg[14] ),
    .A2(net637),
    .A1(net253));
 sg13g2_inv_1 _3945_ (.Y(_0206_),
    .A(net254));
 sg13g2_o21ai_1 _3946_ (.B1(net233),
    .Y(_1168_),
    .A1(_1982_),
    .A2(_0620_));
 sg13g2_o21ai_1 _3947_ (.B1(_1168_),
    .Y(_0207_),
    .A1(net233),
    .A2(_0620_));
 sg13g2_o21ai_1 _3948_ (.B1(net107),
    .Y(_1169_),
    .A1(\measurements.samples_adc.cnt_reg[0] ),
    .A2(_0620_));
 sg13g2_nor2_1 _3949_ (.A(_2159_),
    .B(_0606_),
    .Y(_1170_));
 sg13g2_o21ai_1 _3950_ (.B1(net108),
    .Y(_0208_),
    .A1(_0620_),
    .A2(_1170_));
 sg13g2_nand2_1 _3951_ (.Y(_1171_),
    .A(_2160_),
    .B(_0608_));
 sg13g2_mux2_1 _3952_ (.A0(_1171_),
    .A1(net425),
    .S(_0620_),
    .X(_0209_));
 sg13g2_o21ai_1 _3953_ (.B1(net262),
    .Y(_1172_),
    .A1(_0607_),
    .A2(_0620_));
 sg13g2_o21ai_1 _3954_ (.B1(net263),
    .Y(_0210_),
    .A1(_2160_),
    .A2(_0620_));
 sg13g2_nand2_1 _3955_ (.Y(_1173_),
    .A(\measurements.samples_adc.n84_q[1] ),
    .B(_1982_));
 sg13g2_nand3_1 _3956_ (.B(\measurements.adc_cs ),
    .C(_1173_),
    .A(net79),
    .Y(_1174_));
 sg13g2_nand2_1 _3957_ (.Y(_0211_),
    .A(_0610_),
    .B(net80));
 sg13g2_nor3_1 _3958_ (.A(_1979_),
    .B(_1980_),
    .C(_2157_),
    .Y(_1175_));
 sg13g2_nand2b_1 _3959_ (.Y(_1176_),
    .B(_2165_),
    .A_N(_1175_));
 sg13g2_nor2_1 _3960_ (.A(net118),
    .B(_1176_),
    .Y(_1177_));
 sg13g2_o21ai_1 _3961_ (.B1(net690),
    .Y(_1178_),
    .A1(_0938_),
    .A2(_0955_));
 sg13g2_nand2_1 _3962_ (.Y(_1179_),
    .A(_2102_),
    .B(_1178_));
 sg13g2_a21oi_1 _3963_ (.A1(_2165_),
    .A2(_1175_),
    .Y(_1180_),
    .B1(_0956_));
 sg13g2_a21oi_1 _3964_ (.A1(_2074_),
    .A2(_2162_),
    .Y(_1181_),
    .B1(_2103_));
 sg13g2_a21oi_1 _3965_ (.A1(_2105_),
    .A2(net690),
    .Y(_1182_),
    .B1(_1181_));
 sg13g2_nand2_1 _3966_ (.Y(_1183_),
    .A(_1180_),
    .B(_1182_));
 sg13g2_nor4_1 _3967_ (.A(_2109_),
    .B(_1177_),
    .C(_1179_),
    .D(_1183_),
    .Y(_1184_));
 sg13g2_nand2_1 _3968_ (.Y(_1185_),
    .A(_2076_),
    .B(_0937_));
 sg13g2_mux2_1 _3969_ (.A0(net186),
    .A1(_1185_),
    .S(_1184_),
    .X(_0212_));
 sg13g2_o21ai_1 _3970_ (.B1(_0940_),
    .Y(_1186_),
    .A1(net735),
    .A2(_2163_));
 sg13g2_nor2_1 _3971_ (.A(_2075_),
    .B(_1186_),
    .Y(_1187_));
 sg13g2_nor2_2 _3972_ (.A(net690),
    .B(_1187_),
    .Y(_1188_));
 sg13g2_nor3_2 _3973_ (.A(_2104_),
    .B(net690),
    .C(_2163_),
    .Y(_1189_));
 sg13g2_nand3_1 _3974_ (.B(net757),
    .C(net744),
    .A(\display_x[0] ),
    .Y(_1190_));
 sg13g2_nor2b_1 _3975_ (.A(net755),
    .B_N(_0017_),
    .Y(_1191_));
 sg13g2_a21oi_1 _3976_ (.A1(net755),
    .A2(net737),
    .Y(_1192_),
    .B1(_1191_));
 sg13g2_nor2_1 _3977_ (.A(net755),
    .B(_0015_),
    .Y(_1193_));
 sg13g2_a21oi_1 _3978_ (.A1(net755),
    .A2(_2039_),
    .Y(_1194_),
    .B1(_1193_));
 sg13g2_nor2_1 _3979_ (.A(net705),
    .B(_1194_),
    .Y(_1195_));
 sg13g2_a21oi_2 _3980_ (.B1(_1195_),
    .Y(_1196_),
    .A2(_1192_),
    .A1(net705));
 sg13g2_nor2_2 _3981_ (.A(\display_x[1] ),
    .B(net755),
    .Y(_1197_));
 sg13g2_o21ai_1 _3982_ (.B1(net744),
    .Y(_1198_),
    .A1(net750),
    .A2(_1197_));
 sg13g2_nand2_1 _3983_ (.Y(_1199_),
    .A(net702),
    .B(_1196_));
 sg13g2_nand3_1 _3984_ (.B(_1198_),
    .C(_1199_),
    .A(_1190_),
    .Y(_1200_));
 sg13g2_mux2_1 _3985_ (.A0(\measurements.address_counter_reg[1] ),
    .A1(net731),
    .S(net759),
    .X(_1201_));
 sg13g2_mux4_1 _3986_ (.S0(net759),
    .A0(\measurements.address_counter_reg[3] ),
    .A1(\measurements.address_counter_reg[2] ),
    .A2(\measurements.address_counter_reg[1] ),
    .A3(net731),
    .S1(net753),
    .X(_1202_));
 sg13g2_nand2_1 _3987_ (.Y(_1203_),
    .A(net703),
    .B(_1202_));
 sg13g2_nand2_1 _3988_ (.Y(_1204_),
    .A(\measurements.n246_q[3] ),
    .B(_1203_));
 sg13g2_mux2_1 _3989_ (.A0(\measurements.address_counter_reg[4] ),
    .A1(\measurements.address_counter_reg[3] ),
    .S(net759),
    .X(_1205_));
 sg13g2_mux2_1 _3990_ (.A0(\measurements.address_counter_reg[2] ),
    .A1(\measurements.address_counter_reg[1] ),
    .S(net759),
    .X(_1206_));
 sg13g2_mux2_1 _3991_ (.A0(_1205_),
    .A1(_1206_),
    .S(net753),
    .X(_1207_));
 sg13g2_inv_1 _3992_ (.Y(_1208_),
    .A(_1207_));
 sg13g2_nand2_1 _3993_ (.Y(_1209_),
    .A(net744),
    .B(_0917_));
 sg13g2_nand3_1 _3994_ (.B(net748),
    .C(_0917_),
    .A(net731),
    .Y(_1210_));
 sg13g2_o21ai_1 _3995_ (.B1(_1210_),
    .Y(_1211_),
    .A1(net748),
    .A2(_1208_));
 sg13g2_or2_1 _3996_ (.X(_1212_),
    .B(_1211_),
    .A(_2004_));
 sg13g2_xnor2_1 _3997_ (.Y(_1213_),
    .A(_2004_),
    .B(_1211_));
 sg13g2_or2_1 _3998_ (.X(_1214_),
    .B(_1213_),
    .A(_1204_));
 sg13g2_xor2_1 _3999_ (.B(_1203_),
    .A(\measurements.n246_q[3] ),
    .X(_1215_));
 sg13g2_inv_1 _4000_ (.Y(_1216_),
    .A(_1215_));
 sg13g2_nor2b_2 _4001_ (.A(net757),
    .B_N(net751),
    .Y(_1217_));
 sg13g2_a22oi_1 _4002_ (.Y(_1218_),
    .B1(_1217_),
    .B2(net731),
    .A2(_1206_),
    .A1(net706));
 sg13g2_o21ai_1 _4003_ (.B1(\measurements.n246_q[2] ),
    .Y(_1219_),
    .A1(net746),
    .A2(_1218_));
 sg13g2_nor2_1 _4004_ (.A(_1216_),
    .B(_1219_),
    .Y(_1220_));
 sg13g2_or3_1 _4005_ (.A(\measurements.n246_q[2] ),
    .B(net746),
    .C(_1218_),
    .X(_1221_));
 sg13g2_nand3_1 _4006_ (.B(net703),
    .C(_1201_),
    .A(net706),
    .Y(_1222_));
 sg13g2_and2_1 _4007_ (.A(\measurements.n246_q[1] ),
    .B(_1222_),
    .X(_1223_));
 sg13g2_and3_1 _4008_ (.X(_1224_),
    .A(_1219_),
    .B(_1221_),
    .C(_1223_));
 sg13g2_nand3_1 _4009_ (.B(_1221_),
    .C(_1223_),
    .A(_1219_),
    .Y(_1225_));
 sg13g2_nand3_1 _4010_ (.B(net702),
    .C(_0917_),
    .A(net732),
    .Y(_1226_));
 sg13g2_nor2_1 _4011_ (.A(\measurements.n246_q[0] ),
    .B(_1226_),
    .Y(_1227_));
 sg13g2_xor2_1 _4012_ (.B(_1222_),
    .A(\measurements.n246_q[1] ),
    .X(_1228_));
 sg13g2_nor2b_1 _4013_ (.A(_1227_),
    .B_N(_1228_),
    .Y(_1229_));
 sg13g2_a21o_1 _4014_ (.A2(_1221_),
    .A1(_1219_),
    .B1(_1223_),
    .X(_1230_));
 sg13g2_nand3_1 _4015_ (.B(_1229_),
    .C(_1230_),
    .A(_1225_),
    .Y(_1231_));
 sg13g2_a21o_1 _4016_ (.A2(_1230_),
    .A1(_1229_),
    .B1(_1224_),
    .X(_1232_));
 sg13g2_xnor2_1 _4017_ (.Y(_1233_),
    .A(_1215_),
    .B(_1219_));
 sg13g2_a21oi_2 _4018_ (.B1(_1220_),
    .Y(_1234_),
    .A2(_1233_),
    .A1(_1232_));
 sg13g2_xnor2_1 _4019_ (.Y(_1235_),
    .A(_1204_),
    .B(_1213_));
 sg13g2_o21ai_1 _4020_ (.B1(_1214_),
    .Y(_1236_),
    .A1(_1234_),
    .A2(_1235_));
 sg13g2_nand3_1 _4021_ (.B(net748),
    .C(_1201_),
    .A(net706),
    .Y(_1237_));
 sg13g2_mux4_1 _4022_ (.S0(net760),
    .A0(\measurements.address_counter_reg[5] ),
    .A1(\measurements.address_counter_reg[4] ),
    .A2(\measurements.address_counter_reg[3] ),
    .A3(\measurements.address_counter_reg[2] ),
    .S1(net753),
    .X(_1238_));
 sg13g2_nand2_1 _4023_ (.Y(_1239_),
    .A(net703),
    .B(_1238_));
 sg13g2_nand2_1 _4024_ (.Y(_1240_),
    .A(_1237_),
    .B(_1239_));
 sg13g2_nand3_1 _4025_ (.B(_1237_),
    .C(_1239_),
    .A(\measurements.memoryShift[0] ),
    .Y(_1241_));
 sg13g2_xnor2_1 _4026_ (.Y(_1242_),
    .A(_2020_),
    .B(_1240_));
 sg13g2_xnor2_1 _4027_ (.Y(_1243_),
    .A(_2005_),
    .B(_1242_));
 sg13g2_nor2_1 _4028_ (.A(_1212_),
    .B(_1243_),
    .Y(_1244_));
 sg13g2_xor2_1 _4029_ (.B(_1243_),
    .A(_1212_),
    .X(_1245_));
 sg13g2_xor2_1 _4030_ (.B(_1245_),
    .A(_1236_),
    .X(_1246_));
 sg13g2_nand2b_1 _4031_ (.Y(_1247_),
    .B(_1246_),
    .A_N(_1200_));
 sg13g2_o21ai_1 _4032_ (.B1(_1247_),
    .Y(_1248_),
    .A1(net751),
    .A2(_1190_));
 sg13g2_a21oi_2 _4033_ (.B1(_1244_),
    .Y(_1249_),
    .A2(_1245_),
    .A1(_1236_));
 sg13g2_o21ai_1 _4034_ (.B1(_1241_),
    .Y(_1250_),
    .A1(_2005_),
    .A2(_1242_));
 sg13g2_nor2b_1 _4035_ (.A(net760),
    .B_N(\measurements.address_counter_reg[6] ),
    .Y(_1251_));
 sg13g2_a21oi_2 _4036_ (.B1(_1251_),
    .Y(_1252_),
    .A2(net759),
    .A1(\measurements.address_counter_reg[5] ));
 sg13g2_nor2_1 _4037_ (.A(net706),
    .B(_1205_),
    .Y(_1253_));
 sg13g2_a21oi_2 _4038_ (.B1(_1253_),
    .Y(_1254_),
    .A2(_1252_),
    .A1(net706));
 sg13g2_nand2_1 _4039_ (.Y(_1255_),
    .A(net748),
    .B(_1218_));
 sg13g2_o21ai_1 _4040_ (.B1(_1255_),
    .Y(_1256_),
    .A1(net748),
    .A2(_1254_));
 sg13g2_and2_1 _4041_ (.A(\measurements.memoryShift[1] ),
    .B(_1256_),
    .X(_1257_));
 sg13g2_xnor2_1 _4042_ (.Y(_1258_),
    .A(_2019_),
    .B(_1256_));
 sg13g2_xnor2_1 _4043_ (.Y(_1259_),
    .A(\measurements.n246_q[6] ),
    .B(_1258_));
 sg13g2_nand2b_1 _4044_ (.Y(_1260_),
    .B(_1250_),
    .A_N(_1259_));
 sg13g2_xor2_1 _4045_ (.B(_1259_),
    .A(_1250_),
    .X(_1261_));
 sg13g2_xor2_1 _4046_ (.B(_1261_),
    .A(_1249_),
    .X(_1262_));
 sg13g2_nor2b_1 _4047_ (.A(net756),
    .B_N(_0018_),
    .Y(_1263_));
 sg13g2_a21oi_1 _4048_ (.A1(net755),
    .A2(_0017_),
    .Y(_1264_),
    .B1(_1263_));
 sg13g2_mux2_1 _4049_ (.A0(_0016_),
    .A1(_0015_),
    .S(net755),
    .X(_1265_));
 sg13g2_nor2_1 _4050_ (.A(net705),
    .B(_1265_),
    .Y(_1266_));
 sg13g2_a21oi_2 _4051_ (.B1(_1266_),
    .Y(_1267_),
    .A2(_1264_),
    .A1(net705));
 sg13g2_mux2_1 _4052_ (.A0(\display_x[2] ),
    .A1(\display_x[1] ),
    .S(net755),
    .X(_1268_));
 sg13g2_o21ai_1 _4053_ (.B1(_0913_),
    .Y(_1269_),
    .A1(net750),
    .A2(_1268_));
 sg13g2_a21oi_1 _4054_ (.A1(net738),
    .A2(_1217_),
    .Y(_1270_),
    .B1(_1269_));
 sg13g2_inv_1 _4055_ (.Y(_1271_),
    .A(_1270_));
 sg13g2_nor2_1 _4056_ (.A(net702),
    .B(_1270_),
    .Y(_1272_));
 sg13g2_nand3_1 _4057_ (.B(net744),
    .C(_1217_),
    .A(net738),
    .Y(_1273_));
 sg13g2_a21oi_1 _4058_ (.A1(net702),
    .A2(_1267_),
    .Y(_1274_),
    .B1(_1272_));
 sg13g2_nand2_1 _4059_ (.Y(_1275_),
    .A(_1262_),
    .B(_1274_));
 sg13g2_xnor2_1 _4060_ (.Y(_1276_),
    .A(_1262_),
    .B(_1274_));
 sg13g2_nand2b_1 _4061_ (.Y(_1277_),
    .B(_1248_),
    .A_N(_1276_));
 sg13g2_nand2_1 _4062_ (.Y(_1278_),
    .A(net750),
    .B(_1268_));
 sg13g2_o21ai_1 _4063_ (.B1(_1278_),
    .Y(_1279_),
    .A1(net750),
    .A2(_1265_));
 sg13g2_nand2_1 _4064_ (.Y(_1280_),
    .A(net702),
    .B(_1279_));
 sg13g2_o21ai_1 _4065_ (.B1(_1280_),
    .Y(_1281_),
    .A1(net738),
    .A2(_1209_));
 sg13g2_xor2_1 _4066_ (.B(_1235_),
    .A(_1234_),
    .X(_1282_));
 sg13g2_nand2_1 _4067_ (.Y(_1283_),
    .A(_1281_),
    .B(_1282_));
 sg13g2_o21ai_1 _4068_ (.B1(_1283_),
    .Y(_1284_),
    .A1(_1999_),
    .A2(_1209_));
 sg13g2_xnor2_1 _4069_ (.Y(_1285_),
    .A(_1200_),
    .B(_1246_));
 sg13g2_nand2_1 _4070_ (.Y(_1286_),
    .A(_1284_),
    .B(_1285_));
 sg13g2_nor2_2 _4071_ (.A(_1999_),
    .B(net744),
    .Y(_1287_));
 sg13g2_nor2b_1 _4072_ (.A(_0913_),
    .B_N(_1287_),
    .Y(_1288_));
 sg13g2_nand2_1 _4073_ (.Y(_1289_),
    .A(net705),
    .B(_1194_));
 sg13g2_nand2_1 _4074_ (.Y(_1290_),
    .A(net750),
    .B(_1197_));
 sg13g2_a21oi_2 _4075_ (.B1(_0914_),
    .Y(_1291_),
    .A2(_1290_),
    .A1(_1289_));
 sg13g2_nor3_1 _4076_ (.A(net744),
    .B(_1288_),
    .C(_1291_),
    .Y(_1292_));
 sg13g2_xnor2_1 _4077_ (.Y(_1293_),
    .A(_1232_),
    .B(_1233_));
 sg13g2_nor4_1 _4078_ (.A(net744),
    .B(_1288_),
    .C(_1291_),
    .D(_1293_),
    .Y(_1294_));
 sg13g2_nor2_1 _4079_ (.A(_1288_),
    .B(_1294_),
    .Y(_1295_));
 sg13g2_xnor2_1 _4080_ (.Y(_1296_),
    .A(_1281_),
    .B(_1282_));
 sg13g2_or2_1 _4081_ (.X(_1297_),
    .B(_1296_),
    .A(_1295_));
 sg13g2_nor2_1 _4082_ (.A(net744),
    .B(_1271_),
    .Y(_1298_));
 sg13g2_a21o_1 _4083_ (.A2(_1230_),
    .A1(_1225_),
    .B1(_1229_),
    .X(_1299_));
 sg13g2_and2_1 _4084_ (.A(_1231_),
    .B(_1299_),
    .X(_1300_));
 sg13g2_nand3_1 _4085_ (.B(_1298_),
    .C(_1299_),
    .A(_1231_),
    .Y(_1301_));
 sg13g2_a22oi_1 _4086_ (.Y(_1302_),
    .B1(_1298_),
    .B2(_1300_),
    .A2(_1287_),
    .A1(_1217_));
 sg13g2_xor2_1 _4087_ (.B(_1293_),
    .A(_1292_),
    .X(_1303_));
 sg13g2_or2_1 _4088_ (.X(_1304_),
    .B(_1303_),
    .A(_1302_));
 sg13g2_and2_1 _4089_ (.A(_0923_),
    .B(_1287_),
    .X(_1305_));
 sg13g2_or4_1 _4090_ (.A(net752),
    .B(net745),
    .C(_1197_),
    .D(_1305_),
    .X(_1306_));
 sg13g2_xnor2_1 _4091_ (.Y(_1307_),
    .A(_1227_),
    .B(_1228_));
 sg13g2_nor2b_1 _4092_ (.A(_1306_),
    .B_N(_1307_),
    .Y(_1308_));
 sg13g2_or2_1 _4093_ (.X(_1309_),
    .B(_1308_),
    .A(_1305_));
 sg13g2_a21o_1 _4094_ (.A2(_1299_),
    .A1(_1231_),
    .B1(_1298_),
    .X(_1310_));
 sg13g2_and3_1 _4095_ (.X(_1311_),
    .A(_1301_),
    .B(_1309_),
    .C(_1310_));
 sg13g2_xnor2_1 _4096_ (.Y(_1312_),
    .A(_1306_),
    .B(_1307_));
 sg13g2_nand2_1 _4097_ (.Y(_1313_),
    .A(_0917_),
    .B(_1287_));
 sg13g2_nand2_1 _4098_ (.Y(_1314_),
    .A(_0918_),
    .B(_1313_));
 sg13g2_nand3_1 _4099_ (.B(_0917_),
    .C(_1287_),
    .A(_0002_),
    .Y(_1315_));
 sg13g2_xor2_1 _4100_ (.B(_1226_),
    .A(\measurements.n246_q[0] ),
    .X(_1316_));
 sg13g2_nand2_1 _4101_ (.Y(_1317_),
    .A(_1315_),
    .B(_1316_));
 sg13g2_nand3_1 _4102_ (.B(_1314_),
    .C(_1317_),
    .A(_1312_),
    .Y(_1318_));
 sg13g2_a21oi_1 _4103_ (.A1(_1301_),
    .A2(_1310_),
    .Y(_1319_),
    .B1(_1309_));
 sg13g2_nor2_1 _4104_ (.A(_1311_),
    .B(_1319_),
    .Y(_1320_));
 sg13g2_nor3_1 _4105_ (.A(_1311_),
    .B(_1318_),
    .C(_1319_),
    .Y(_1321_));
 sg13g2_xor2_1 _4106_ (.B(_1303_),
    .A(_1302_),
    .X(_1322_));
 sg13g2_o21ai_1 _4107_ (.B1(_1322_),
    .Y(_1323_),
    .A1(_1311_),
    .A2(_1321_));
 sg13g2_xnor2_1 _4108_ (.Y(_1324_),
    .A(_1295_),
    .B(_1296_));
 sg13g2_a21o_1 _4109_ (.A2(_1323_),
    .A1(_1304_),
    .B1(_1324_),
    .X(_1325_));
 sg13g2_xnor2_1 _4110_ (.Y(_1326_),
    .A(_1284_),
    .B(_1285_));
 sg13g2_a21o_1 _4111_ (.A2(_1325_),
    .A1(_1297_),
    .B1(_1326_),
    .X(_1327_));
 sg13g2_xor2_1 _4112_ (.B(_1276_),
    .A(_1248_),
    .X(_1328_));
 sg13g2_a21o_1 _4113_ (.A2(_1327_),
    .A1(_1286_),
    .B1(_1328_),
    .X(_1329_));
 sg13g2_nand2_1 _4114_ (.Y(_1330_),
    .A(_1273_),
    .B(_1275_));
 sg13g2_o21ai_1 _4115_ (.B1(_1260_),
    .Y(_1331_),
    .A1(_1249_),
    .A2(_1261_));
 sg13g2_a21oi_1 _4116_ (.A1(\measurements.n246_q[6] ),
    .A2(_1258_),
    .Y(_1332_),
    .B1(_1257_));
 sg13g2_nor2_1 _4117_ (.A(\measurements.address_counter_reg[7] ),
    .B(net759),
    .Y(_1333_));
 sg13g2_nor2b_1 _4118_ (.A(\measurements.address_counter_reg[6] ),
    .B_N(net759),
    .Y(_1334_));
 sg13g2_mux4_1 _4119_ (.S0(net760),
    .A0(\measurements.address_counter_reg[7] ),
    .A1(\measurements.address_counter_reg[6] ),
    .A2(\measurements.address_counter_reg[5] ),
    .A3(\measurements.address_counter_reg[4] ),
    .S1(net753),
    .X(_1335_));
 sg13g2_mux2_1 _4120_ (.A0(_1202_),
    .A1(_1335_),
    .S(net703),
    .X(_1336_));
 sg13g2_xnor2_1 _4121_ (.Y(_1337_),
    .A(\measurements.memoryShift[2] ),
    .B(_1336_));
 sg13g2_xnor2_1 _4122_ (.Y(_1338_),
    .A(\measurements.n246_q[7] ),
    .B(_1337_));
 sg13g2_nor2_1 _4123_ (.A(_1332_),
    .B(_1338_),
    .Y(_1339_));
 sg13g2_xor2_1 _4124_ (.B(_1338_),
    .A(_1332_),
    .X(_1340_));
 sg13g2_xnor2_1 _4125_ (.Y(_1341_),
    .A(_1331_),
    .B(_1340_));
 sg13g2_inv_1 _4126_ (.Y(_1342_),
    .A(_1341_));
 sg13g2_nand2_1 _4127_ (.Y(_1343_),
    .A(net745),
    .B(_1291_));
 sg13g2_nand4_1 _4128_ (.B(net757),
    .C(net751),
    .A(net738),
    .Y(_1344_),
    .D(net745));
 sg13g2_mux2_1 _4129_ (.A0(_0019_),
    .A1(_0018_),
    .S(net756),
    .X(_1345_));
 sg13g2_nor2_1 _4130_ (.A(net751),
    .B(_1345_),
    .Y(_1346_));
 sg13g2_a21oi_1 _4131_ (.A1(net750),
    .A2(_1192_),
    .Y(_1347_),
    .B1(_1346_));
 sg13g2_nand2_1 _4132_ (.Y(_1348_),
    .A(net704),
    .B(_1347_));
 sg13g2_nand3_1 _4133_ (.B(_1344_),
    .C(_1348_),
    .A(_1343_),
    .Y(_1349_));
 sg13g2_xor2_1 _4134_ (.B(_1349_),
    .A(_1341_),
    .X(_1350_));
 sg13g2_and2_1 _4135_ (.A(_1330_),
    .B(_1350_),
    .X(_1351_));
 sg13g2_xnor2_1 _4136_ (.Y(_1352_),
    .A(_1330_),
    .B(_1350_));
 sg13g2_a21oi_2 _4137_ (.B1(_1352_),
    .Y(_1353_),
    .A2(_1329_),
    .A1(_1277_));
 sg13g2_nand3_1 _4138_ (.B(_1329_),
    .C(_1352_),
    .A(_1277_),
    .Y(_1354_));
 sg13g2_nand2_1 _4139_ (.Y(_1355_),
    .A(net656),
    .B(_1354_));
 sg13g2_nor2b_1 _4140_ (.A(_2167_),
    .B_N(_2067_),
    .Y(_1356_));
 sg13g2_nand2b_1 _4141_ (.Y(_1357_),
    .B(_2067_),
    .A_N(_2167_));
 sg13g2_a21oi_1 _4142_ (.A1(net658),
    .A2(_1342_),
    .Y(_1358_),
    .B1(net662));
 sg13g2_o21ai_1 _4143_ (.B1(_1358_),
    .Y(_1359_),
    .A1(_1353_),
    .A2(_1355_));
 sg13g2_a21oi_1 _4144_ (.A1(net1008),
    .A2(net665),
    .Y(_1360_),
    .B1(_0942_));
 sg13g2_a22oi_1 _4145_ (.Y(_1361_),
    .B1(_1359_),
    .B2(_1360_),
    .A2(_1189_),
    .A1(net345));
 sg13g2_nand2b_1 _4146_ (.Y(_1362_),
    .B(_1188_),
    .A_N(_1361_));
 sg13g2_o21ai_1 _4147_ (.B1(_0954_),
    .Y(_1363_),
    .A1(net525),
    .A2(_1117_));
 sg13g2_a22oi_1 _4148_ (.Y(_0215_),
    .B1(_1362_),
    .B2(_1363_),
    .A2(net633),
    .A1(net618));
 sg13g2_mux2_1 _4149_ (.A0(\measurements.address_counter_reg[8] ),
    .A1(\measurements.address_counter_reg[7] ),
    .S(net759),
    .X(_1364_));
 sg13g2_mux2_1 _4150_ (.A0(\measurements.address_counter_reg[10] ),
    .A1(\measurements.address_counter_reg[9] ),
    .S(net760),
    .X(_1365_));
 sg13g2_mux2_1 _4151_ (.A0(_1364_),
    .A1(_1365_),
    .S(net706),
    .X(_1366_));
 sg13g2_inv_1 _4152_ (.Y(_1367_),
    .A(_1366_));
 sg13g2_nand2_1 _4153_ (.Y(_1368_),
    .A(net703),
    .B(_1367_));
 sg13g2_o21ai_1 _4154_ (.B1(_1368_),
    .Y(_1369_),
    .A1(net703),
    .A2(_1254_));
 sg13g2_and2_1 _4155_ (.A(\measurements.memoryShift[5] ),
    .B(_1369_),
    .X(_1370_));
 sg13g2_xnor2_1 _4156_ (.Y(_1371_),
    .A(_2022_),
    .B(_1369_));
 sg13g2_a21oi_2 _4157_ (.B1(_1370_),
    .Y(_1372_),
    .A2(_1371_),
    .A1(\measurements.n246_q[10] ));
 sg13g2_nand2b_1 _4158_ (.Y(_1373_),
    .B(net748),
    .A_N(_1335_));
 sg13g2_mux2_1 _4159_ (.A0(\measurements.address_counter_reg[9] ),
    .A1(\measurements.address_counter_reg[8] ),
    .S(net761),
    .X(_1374_));
 sg13g2_nand2_1 _4160_ (.Y(_1375_),
    .A(\measurements.address_counter_reg[10] ),
    .B(net761));
 sg13g2_o21ai_1 _4161_ (.B1(_1375_),
    .Y(_1376_),
    .A1(_2006_),
    .A2(net760));
 sg13g2_mux2_1 _4162_ (.A0(_1374_),
    .A1(_1376_),
    .S(net705),
    .X(_1377_));
 sg13g2_o21ai_1 _4163_ (.B1(_1373_),
    .Y(_1378_),
    .A1(net749),
    .A2(_1377_));
 sg13g2_xor2_1 _4164_ (.B(_1378_),
    .A(\measurements.memoryShift[6] ),
    .X(_1379_));
 sg13g2_xnor2_1 _4165_ (.Y(_1380_),
    .A(\measurements.n246_q[11] ),
    .B(_1379_));
 sg13g2_or2_1 _4166_ (.X(_1381_),
    .B(_1380_),
    .A(_1372_));
 sg13g2_o21ai_1 _4167_ (.B1(net753),
    .Y(_1382_),
    .A1(_1333_),
    .A2(_1334_));
 sg13g2_o21ai_1 _4168_ (.B1(_1382_),
    .Y(_1383_),
    .A1(net754),
    .A2(_1374_));
 sg13g2_nor2_1 _4169_ (.A(net703),
    .B(_1238_),
    .Y(_1384_));
 sg13g2_a21oi_1 _4170_ (.A1(net704),
    .A2(_1383_),
    .Y(_1385_),
    .B1(_1384_));
 sg13g2_nor2_1 _4171_ (.A(_0028_),
    .B(_1385_),
    .Y(_1386_));
 sg13g2_xnor2_1 _4172_ (.Y(_1387_),
    .A(\measurements.memoryShift[4] ),
    .B(_1385_));
 sg13g2_a21oi_1 _4173_ (.A1(\measurements.n246_q[9] ),
    .A2(_1387_),
    .Y(_1388_),
    .B1(_1386_));
 sg13g2_xnor2_1 _4174_ (.Y(_1389_),
    .A(\measurements.n246_q[10] ),
    .B(_1371_));
 sg13g2_nor2_1 _4175_ (.A(_1388_),
    .B(_1389_),
    .Y(_1390_));
 sg13g2_nor2_1 _4176_ (.A(net753),
    .B(_1364_),
    .Y(_1391_));
 sg13g2_a21oi_1 _4177_ (.A1(net753),
    .A2(_1252_),
    .Y(_1392_),
    .B1(_1391_));
 sg13g2_nand2_1 _4178_ (.Y(_1393_),
    .A(net704),
    .B(_1392_));
 sg13g2_o21ai_1 _4179_ (.B1(_1393_),
    .Y(_1394_),
    .A1(net703),
    .A2(_1208_));
 sg13g2_nor2_1 _4180_ (.A(_2021_),
    .B(_1394_),
    .Y(_1395_));
 sg13g2_xnor2_1 _4181_ (.Y(_1396_),
    .A(\measurements.memoryShift[3] ),
    .B(_1394_));
 sg13g2_a21oi_1 _4182_ (.A1(\measurements.n246_q[8] ),
    .A2(_1396_),
    .Y(_1397_),
    .B1(_1395_));
 sg13g2_xnor2_1 _4183_ (.Y(_1398_),
    .A(\measurements.n246_q[9] ),
    .B(_1387_));
 sg13g2_nor2_1 _4184_ (.A(_1397_),
    .B(_1398_),
    .Y(_1399_));
 sg13g2_nor2_1 _4185_ (.A(_0027_),
    .B(_1336_),
    .Y(_1400_));
 sg13g2_a21oi_2 _4186_ (.B1(_1400_),
    .Y(_1401_),
    .A2(_1337_),
    .A1(\measurements.n246_q[7] ));
 sg13g2_xnor2_1 _4187_ (.Y(_1402_),
    .A(\measurements.n246_q[8] ),
    .B(_1396_));
 sg13g2_or2_1 _4188_ (.X(_1403_),
    .B(_1402_),
    .A(_1401_));
 sg13g2_a21oi_2 _4189_ (.B1(_1339_),
    .Y(_1404_),
    .A2(_1340_),
    .A1(_1331_));
 sg13g2_and2_1 _4190_ (.A(_1401_),
    .B(_1402_),
    .X(_1405_));
 sg13g2_xor2_1 _4191_ (.B(_1402_),
    .A(_1401_),
    .X(_1406_));
 sg13g2_o21ai_1 _4192_ (.B1(_1403_),
    .Y(_1407_),
    .A1(_1404_),
    .A2(_1405_));
 sg13g2_xor2_1 _4193_ (.B(_1398_),
    .A(_1397_),
    .X(_1408_));
 sg13g2_a21o_1 _4194_ (.A2(_1408_),
    .A1(_1407_),
    .B1(_1399_),
    .X(_1409_));
 sg13g2_xor2_1 _4195_ (.B(_1389_),
    .A(_1388_),
    .X(_1410_));
 sg13g2_a21oi_1 _4196_ (.A1(_1409_),
    .A2(_1410_),
    .Y(_1411_),
    .B1(_1390_));
 sg13g2_and2_1 _4197_ (.A(_1372_),
    .B(_1380_),
    .X(_1412_));
 sg13g2_xor2_1 _4198_ (.B(_1380_),
    .A(_1372_),
    .X(_1413_));
 sg13g2_o21ai_1 _4199_ (.B1(_1381_),
    .Y(_1414_),
    .A1(_1411_),
    .A2(_1412_));
 sg13g2_a22oi_1 _4200_ (.Y(_1415_),
    .B1(_1379_),
    .B2(\measurements.n246_q[11] ),
    .A2(_1378_),
    .A1(_2042_));
 sg13g2_nor2_1 _4201_ (.A(\measurements.address_counter_reg[12] ),
    .B(net760),
    .Y(_1416_));
 sg13g2_a21oi_1 _4202_ (.A1(_2006_),
    .A2(net761),
    .Y(_1417_),
    .B1(_1416_));
 sg13g2_nor3_1 _4203_ (.A(net754),
    .B(net749),
    .C(_1417_),
    .Y(_1418_));
 sg13g2_nor3_1 _4204_ (.A(net705),
    .B(net749),
    .C(_1365_),
    .Y(_1419_));
 sg13g2_nor2_1 _4205_ (.A(_1418_),
    .B(_1419_),
    .Y(_1420_));
 sg13g2_o21ai_1 _4206_ (.B1(_1420_),
    .Y(_1421_),
    .A1(net704),
    .A2(_1392_));
 sg13g2_xor2_1 _4207_ (.B(_1421_),
    .A(\measurements.memoryShift[7] ),
    .X(_1422_));
 sg13g2_nand2_1 _4208_ (.Y(_1423_),
    .A(net308),
    .B(_1422_));
 sg13g2_xor2_1 _4209_ (.B(_1422_),
    .A(\measurements.n246_q[12] ),
    .X(_1424_));
 sg13g2_nor2b_1 _4210_ (.A(_1415_),
    .B_N(_1424_),
    .Y(_1425_));
 sg13g2_xnor2_1 _4211_ (.Y(_1426_),
    .A(_1415_),
    .B(_1424_));
 sg13g2_xnor2_1 _4212_ (.Y(_1427_),
    .A(_1414_),
    .B(_1426_));
 sg13g2_nand2_1 _4213_ (.Y(_1428_),
    .A(\display_x[9] ),
    .B(net758));
 sg13g2_nand4_1 _4214_ (.B(net758),
    .C(net752),
    .A(\display_x[9] ),
    .Y(_1429_),
    .D(net704));
 sg13g2_nand2_1 _4215_ (.Y(_1430_),
    .A(net756),
    .B(_0019_));
 sg13g2_o21ai_1 _4216_ (.B1(_1430_),
    .Y(_1431_),
    .A1(net756),
    .A2(_2040_));
 sg13g2_nor2_1 _4217_ (.A(net750),
    .B(_1431_),
    .Y(_1432_));
 sg13g2_a21oi_1 _4218_ (.A1(net750),
    .A2(_1264_),
    .Y(_1433_),
    .B1(_1432_));
 sg13g2_o21ai_1 _4219_ (.B1(_1429_),
    .Y(_1434_),
    .A1(net704),
    .A2(_1433_));
 sg13g2_nand2b_1 _4220_ (.Y(_1435_),
    .B(_1434_),
    .A_N(_1427_));
 sg13g2_nand2_1 _4221_ (.Y(_1436_),
    .A(net758),
    .B(_0020_));
 sg13g2_o21ai_1 _4222_ (.B1(_1436_),
    .Y(_1437_),
    .A1(_2002_),
    .A2(net758));
 sg13g2_mux2_1 _4223_ (.A0(_1345_),
    .A1(_1437_),
    .S(net705),
    .X(_1438_));
 sg13g2_nand2b_1 _4224_ (.Y(_1439_),
    .B(net747),
    .A_N(_1438_));
 sg13g2_a21oi_1 _4225_ (.A1(_1414_),
    .A2(_1426_),
    .Y(_1440_),
    .B1(_1425_));
 sg13g2_nand2b_1 _4226_ (.Y(_1441_),
    .B(_1421_),
    .A_N(_0031_));
 sg13g2_nand2_1 _4227_ (.Y(_1442_),
    .A(net754),
    .B(_1376_));
 sg13g2_a221oi_1 _4228_ (.B2(\measurements.address_counter_reg[12] ),
    .C1(net749),
    .B1(_0923_),
    .A1(\measurements.address_counter_reg[13] ),
    .Y(_1443_),
    .A2(_0917_));
 sg13g2_a22oi_1 _4229_ (.Y(_1444_),
    .B1(_1442_),
    .B2(_1443_),
    .A2(_1383_),
    .A1(net749));
 sg13g2_xnor2_1 _4230_ (.Y(_1445_),
    .A(net343),
    .B(_1444_));
 sg13g2_xnor2_1 _4231_ (.Y(_1446_),
    .A(net373),
    .B(_1445_));
 sg13g2_a21oi_1 _4232_ (.A1(_1423_),
    .A2(_1441_),
    .Y(_1447_),
    .B1(_1446_));
 sg13g2_nand3_1 _4233_ (.B(_1441_),
    .C(_1446_),
    .A(_1423_),
    .Y(_1448_));
 sg13g2_nor2b_1 _4234_ (.A(_1447_),
    .B_N(_1448_),
    .Y(_1449_));
 sg13g2_nor2b_1 _4235_ (.A(_1440_),
    .B_N(_1449_),
    .Y(_1450_));
 sg13g2_xnor2_1 _4236_ (.Y(_1451_),
    .A(_1440_),
    .B(_1449_));
 sg13g2_nor2b_1 _4237_ (.A(_1439_),
    .B_N(_1451_),
    .Y(_1452_));
 sg13g2_xnor2_1 _4238_ (.Y(_1453_),
    .A(_1439_),
    .B(_1451_));
 sg13g2_nor2b_1 _4239_ (.A(_1435_),
    .B_N(_1453_),
    .Y(_1454_));
 sg13g2_xnor2_1 _4240_ (.Y(_1455_),
    .A(_1411_),
    .B(_1413_));
 sg13g2_or3_1 _4241_ (.A(net747),
    .B(_0008_),
    .C(_1437_),
    .X(_1456_));
 sg13g2_o21ai_1 _4242_ (.B1(_1456_),
    .Y(_1457_),
    .A1(net702),
    .A2(_1347_));
 sg13g2_nand2_1 _4243_ (.Y(_1458_),
    .A(_1455_),
    .B(_1457_));
 sg13g2_xor2_1 _4244_ (.B(_1434_),
    .A(_1427_),
    .X(_1459_));
 sg13g2_or2_1 _4245_ (.X(_1460_),
    .B(_1459_),
    .A(_1458_));
 sg13g2_xor2_1 _4246_ (.B(_1410_),
    .A(_1409_),
    .X(_1461_));
 sg13g2_mux2_1 _4247_ (.A0(_1428_),
    .A1(_1431_),
    .S(net752),
    .X(_1462_));
 sg13g2_and2_1 _4248_ (.A(net702),
    .B(_1462_),
    .X(_1463_));
 sg13g2_a21oi_2 _4249_ (.B1(_1463_),
    .Y(_1464_),
    .A2(_1267_),
    .A1(net747));
 sg13g2_nand2_1 _4250_ (.Y(_1465_),
    .A(_1461_),
    .B(_1464_));
 sg13g2_xor2_1 _4251_ (.B(_1457_),
    .A(_1455_),
    .X(_1466_));
 sg13g2_nor2b_1 _4252_ (.A(_1465_),
    .B_N(_1466_),
    .Y(_1467_));
 sg13g2_xnor2_1 _4253_ (.Y(_1468_),
    .A(_1407_),
    .B(_1408_));
 sg13g2_mux2_1 _4254_ (.A0(_1196_),
    .A1(_1438_),
    .S(net702),
    .X(_1469_));
 sg13g2_nor2_1 _4255_ (.A(_1468_),
    .B(_1469_),
    .Y(_1470_));
 sg13g2_xor2_1 _4256_ (.B(_1464_),
    .A(_1461_),
    .X(_1471_));
 sg13g2_nand2_1 _4257_ (.Y(_1472_),
    .A(_1470_),
    .B(_1471_));
 sg13g2_xnor2_1 _4258_ (.Y(_1473_),
    .A(_1404_),
    .B(_1406_));
 sg13g2_nand2_1 _4259_ (.Y(_1474_),
    .A(net745),
    .B(_1279_));
 sg13g2_o21ai_1 _4260_ (.B1(_1474_),
    .Y(_1475_),
    .A1(net747),
    .A2(_1433_));
 sg13g2_and2_1 _4261_ (.A(_1473_),
    .B(_1475_),
    .X(_1476_));
 sg13g2_xor2_1 _4262_ (.B(_1469_),
    .A(_1468_),
    .X(_1477_));
 sg13g2_and2_1 _4263_ (.A(_1476_),
    .B(_1477_),
    .X(_1478_));
 sg13g2_o21ai_1 _4264_ (.B1(_1344_),
    .Y(_1479_),
    .A1(_1341_),
    .A2(_1349_));
 sg13g2_xor2_1 _4265_ (.B(_1475_),
    .A(_1473_),
    .X(_1480_));
 sg13g2_nand2_1 _4266_ (.Y(_1481_),
    .A(_1479_),
    .B(_1480_));
 sg13g2_xor2_1 _4267_ (.B(_1480_),
    .A(_1479_),
    .X(_1482_));
 sg13g2_o21ai_1 _4268_ (.B1(_1482_),
    .Y(_1483_),
    .A1(_1351_),
    .A2(_1353_));
 sg13g2_xnor2_1 _4269_ (.Y(_1484_),
    .A(_1476_),
    .B(_1477_));
 sg13g2_a21oi_2 _4270_ (.B1(_1484_),
    .Y(_1485_),
    .A2(_1483_),
    .A1(_1481_));
 sg13g2_xor2_1 _4271_ (.B(_1471_),
    .A(_1470_),
    .X(_1486_));
 sg13g2_o21ai_1 _4272_ (.B1(_1486_),
    .Y(_1487_),
    .A1(_1478_),
    .A2(_1485_));
 sg13g2_xor2_1 _4273_ (.B(_1466_),
    .A(_1465_),
    .X(_1488_));
 sg13g2_a21oi_1 _4274_ (.A1(_1472_),
    .A2(_1487_),
    .Y(_1489_),
    .B1(_1488_));
 sg13g2_xor2_1 _4275_ (.B(_1459_),
    .A(_1458_),
    .X(_1490_));
 sg13g2_o21ai_1 _4276_ (.B1(_1490_),
    .Y(_1491_),
    .A1(_1467_),
    .A2(_1489_));
 sg13g2_xor2_1 _4277_ (.B(_1453_),
    .A(_1435_),
    .X(_1492_));
 sg13g2_a21oi_1 _4278_ (.A1(_1460_),
    .A2(_1491_),
    .Y(_1493_),
    .B1(_1492_));
 sg13g2_nor2_1 _4279_ (.A(_1447_),
    .B(_1450_),
    .Y(_1494_));
 sg13g2_nor2_1 _4280_ (.A(_0030_),
    .B(_1444_),
    .Y(_1495_));
 sg13g2_a21oi_1 _4281_ (.A1(net373),
    .A2(_1445_),
    .Y(_1496_),
    .B1(_1495_));
 sg13g2_xor2_1 _4282_ (.B(net343),
    .A(net253),
    .X(_1497_));
 sg13g2_nand2_1 _4283_ (.Y(_1498_),
    .A(net754),
    .B(_1417_));
 sg13g2_a221oi_1 _4284_ (.B2(\measurements.address_counter_reg[13] ),
    .C1(net748),
    .B1(_0923_),
    .A1(\measurements.address_counter_reg[14] ),
    .Y(_1499_),
    .A2(_0917_));
 sg13g2_a22oi_1 _4285_ (.Y(_1500_),
    .B1(_1498_),
    .B2(_1499_),
    .A2(_1367_),
    .A1(net748));
 sg13g2_xnor2_1 _4286_ (.Y(_1501_),
    .A(_1497_),
    .B(_1500_));
 sg13g2_xnor2_1 _4287_ (.Y(_1502_),
    .A(_1496_),
    .B(_1501_));
 sg13g2_xnor2_1 _4288_ (.Y(_1503_),
    .A(_1494_),
    .B(_1502_));
 sg13g2_nor2_1 _4289_ (.A(_0002_),
    .B(_1462_),
    .Y(_1504_));
 sg13g2_xnor2_1 _4290_ (.Y(_1505_),
    .A(_1452_),
    .B(_1504_));
 sg13g2_xnor2_1 _4291_ (.Y(_1506_),
    .A(_1503_),
    .B(_1505_));
 sg13g2_o21ai_1 _4292_ (.B1(_1506_),
    .Y(_1507_),
    .A1(_1454_),
    .A2(_1493_));
 sg13g2_or3_1 _4293_ (.A(_1454_),
    .B(_1493_),
    .C(_1506_),
    .X(_1508_));
 sg13g2_nand3_1 _4294_ (.B(_1507_),
    .C(_1508_),
    .A(net657),
    .Y(_1509_));
 sg13g2_a21oi_1 _4295_ (.A1(net660),
    .A2(_1503_),
    .Y(_1510_),
    .B1(net664));
 sg13g2_o21ai_1 _4296_ (.B1(_0939_),
    .Y(_1511_),
    .A1(net949),
    .A2(net667));
 sg13g2_a21oi_2 _4297_ (.B1(_1511_),
    .Y(_1512_),
    .A2(_1510_),
    .A1(_1509_));
 sg13g2_nand3_1 _4298_ (.B(_1327_),
    .C(_1328_),
    .A(_1286_),
    .Y(_1513_));
 sg13g2_nand3_1 _4299_ (.B(_1329_),
    .C(_1513_),
    .A(net656),
    .Y(_1514_));
 sg13g2_a21oi_1 _4300_ (.A1(net658),
    .A2(_1262_),
    .Y(_1515_),
    .B1(net661));
 sg13g2_nand2_2 _4301_ (.Y(_1516_),
    .A(net504),
    .B(_0941_));
 sg13g2_a221oi_1 _4302_ (.B2(_1515_),
    .C1(_1516_),
    .B1(_1514_),
    .A1(net432),
    .Y(_1517_),
    .A2(net661));
 sg13g2_a21o_1 _4303_ (.A2(_1189_),
    .A1(net894),
    .B1(_1517_),
    .X(_1518_));
 sg13g2_o21ai_1 _4304_ (.B1(_1188_),
    .Y(_1519_),
    .A1(_1512_),
    .A2(_1518_));
 sg13g2_o21ai_1 _4305_ (.B1(_0954_),
    .Y(_1520_),
    .A1(net528),
    .A2(_1117_));
 sg13g2_a22oi_1 _4306_ (.Y(_0216_),
    .B1(_1519_),
    .B2(_1520_),
    .A2(net633),
    .A1(net526));
 sg13g2_nand3_1 _4307_ (.B(_1491_),
    .C(_1492_),
    .A(_1460_),
    .Y(_1521_));
 sg13g2_nand2b_1 _4308_ (.Y(_1522_),
    .B(_1521_),
    .A_N(_1493_));
 sg13g2_a21oi_1 _4309_ (.A1(net659),
    .A2(_1451_),
    .Y(_1523_),
    .B1(net663));
 sg13g2_o21ai_1 _4310_ (.B1(_1523_),
    .Y(_1524_),
    .A1(net660),
    .A2(_1522_));
 sg13g2_a21oi_1 _4311_ (.A1(net903),
    .A2(net664),
    .Y(_1525_),
    .B1(_0940_));
 sg13g2_nand3_1 _4312_ (.B(_1325_),
    .C(_1326_),
    .A(_1297_),
    .Y(_1526_));
 sg13g2_nand3_1 _4313_ (.B(_1327_),
    .C(_1526_),
    .A(net656),
    .Y(_1527_));
 sg13g2_a21oi_1 _4314_ (.A1(net658),
    .A2(_1246_),
    .Y(_1528_),
    .B1(net661));
 sg13g2_a221oi_1 _4315_ (.B2(_1528_),
    .C1(_1516_),
    .B1(_1527_),
    .A1(net476),
    .Y(_1529_),
    .A2(net662));
 sg13g2_a221oi_1 _4316_ (.B2(_1525_),
    .C1(_1529_),
    .B1(_1524_),
    .A1(net357),
    .Y(_1530_),
    .A2(_1189_));
 sg13g2_nand2b_1 _4317_ (.Y(_1531_),
    .B(_1188_),
    .A_N(_1530_));
 sg13g2_o21ai_1 _4318_ (.B1(_0954_),
    .Y(_1532_),
    .A1(net456),
    .A2(_1117_));
 sg13g2_a22oi_1 _4319_ (.Y(_0217_),
    .B1(_1531_),
    .B2(_1532_),
    .A2(net633),
    .A1(net529));
 sg13g2_or3_1 _4320_ (.A(_1467_),
    .B(_1489_),
    .C(_1490_),
    .X(_1533_));
 sg13g2_nand3_1 _4321_ (.B(_1491_),
    .C(_1533_),
    .A(net657),
    .Y(_1534_));
 sg13g2_nor2_1 _4322_ (.A(net657),
    .B(_1427_),
    .Y(_1535_));
 sg13g2_nor2_1 _4323_ (.A(net665),
    .B(_1535_),
    .Y(_1536_));
 sg13g2_a22oi_1 _4324_ (.Y(_1537_),
    .B1(_1534_),
    .B2(_1536_),
    .A2(net664),
    .A1(net909));
 sg13g2_nand3_1 _4325_ (.B(_1323_),
    .C(_1324_),
    .A(_1304_),
    .Y(_1538_));
 sg13g2_nand3_1 _4326_ (.B(_1325_),
    .C(_1538_),
    .A(net656),
    .Y(_1539_));
 sg13g2_a21oi_1 _4327_ (.A1(net658),
    .A2(_1282_),
    .Y(_1540_),
    .B1(net661));
 sg13g2_a221oi_1 _4328_ (.B2(_1540_),
    .C1(_1516_),
    .B1(_1539_),
    .A1(_0059_),
    .Y(_1541_),
    .A2(net661));
 sg13g2_a221oi_1 _4329_ (.B2(_0939_),
    .C1(_1541_),
    .B1(_1537_),
    .A1(net479),
    .Y(_1542_),
    .A2(_1189_));
 sg13g2_nand2b_1 _4330_ (.Y(_1543_),
    .B(_1188_),
    .A_N(_1542_));
 sg13g2_o21ai_1 _4331_ (.B1(_0954_),
    .Y(_1544_),
    .A1(net316),
    .A2(_1117_));
 sg13g2_a22oi_1 _4332_ (.Y(_0218_),
    .B1(_1543_),
    .B2(_1544_),
    .A2(net633),
    .A1(net457));
 sg13g2_nand3_1 _4333_ (.B(_1487_),
    .C(_1488_),
    .A(_1472_),
    .Y(_1545_));
 sg13g2_nand2b_1 _4334_ (.Y(_1546_),
    .B(_1545_),
    .A_N(_1489_));
 sg13g2_a21oi_1 _4335_ (.A1(net658),
    .A2(_1455_),
    .Y(_1547_),
    .B1(net663));
 sg13g2_o21ai_1 _4336_ (.B1(_1547_),
    .Y(_1548_),
    .A1(net659),
    .A2(_1546_));
 sg13g2_a21oi_1 _4337_ (.A1(net1004),
    .A2(net663),
    .Y(_1549_),
    .B1(_0940_));
 sg13g2_nand2_1 _4338_ (.Y(_1550_),
    .A(_1548_),
    .B(_1549_));
 sg13g2_nand2_1 _4339_ (.Y(_1551_),
    .A(net305),
    .B(_1189_));
 sg13g2_or3_1 _4340_ (.A(_1311_),
    .B(_1321_),
    .C(_1322_),
    .X(_1552_));
 sg13g2_nand3_1 _4341_ (.B(_1323_),
    .C(_1552_),
    .A(net656),
    .Y(_1553_));
 sg13g2_o21ai_1 _4342_ (.B1(_1553_),
    .Y(_1554_),
    .A1(net656),
    .A2(_1293_));
 sg13g2_a21oi_1 _4343_ (.A1(_0058_),
    .A2(net661),
    .Y(_1555_),
    .B1(_1516_));
 sg13g2_o21ai_1 _4344_ (.B1(_1555_),
    .Y(_1556_),
    .A1(net661),
    .A2(_1554_));
 sg13g2_nand3_1 _4345_ (.B(_1551_),
    .C(_1556_),
    .A(_1550_),
    .Y(_1557_));
 sg13g2_a221oi_1 _4346_ (.B2(_1557_),
    .C1(net634),
    .B1(_1188_),
    .A1(net375),
    .Y(_1558_),
    .A2(_0954_));
 sg13g2_a21oi_1 _4347_ (.A1(net317),
    .A2(net634),
    .Y(_0219_),
    .B1(_1558_));
 sg13g2_nor3_1 _4348_ (.A(_1478_),
    .B(_1485_),
    .C(_1486_),
    .Y(_1559_));
 sg13g2_nand2_1 _4349_ (.Y(_1560_),
    .A(net657),
    .B(_1487_));
 sg13g2_a21oi_1 _4350_ (.A1(net659),
    .A2(_1461_),
    .Y(_1561_),
    .B1(net663));
 sg13g2_o21ai_1 _4351_ (.B1(_1561_),
    .Y(_1562_),
    .A1(_1559_),
    .A2(_1560_));
 sg13g2_a21oi_1 _4352_ (.A1(net285),
    .A2(net663),
    .Y(_1563_),
    .B1(_0940_));
 sg13g2_nand2_1 _4353_ (.Y(_1564_),
    .A(_1562_),
    .B(_1563_));
 sg13g2_xor2_1 _4354_ (.B(_1320_),
    .A(_1318_),
    .X(_1565_));
 sg13g2_a21oi_1 _4355_ (.A1(net658),
    .A2(_1300_),
    .Y(_1566_),
    .B1(net661));
 sg13g2_o21ai_1 _4356_ (.B1(_1566_),
    .Y(_1567_),
    .A1(_2097_),
    .A2(_1565_));
 sg13g2_a21oi_1 _4357_ (.A1(_0057_),
    .A2(net665),
    .Y(_1568_),
    .B1(_1516_));
 sg13g2_a221oi_1 _4358_ (.B2(_1568_),
    .C1(_2116_),
    .B1(_1567_),
    .A1(net399),
    .Y(_1569_),
    .A2(_1189_));
 sg13g2_nand2_2 _4359_ (.Y(_1570_),
    .A(_1564_),
    .B(_1569_));
 sg13g2_a221oi_1 _4360_ (.B2(_1570_),
    .C1(net633),
    .B1(_1188_),
    .A1(net467),
    .Y(_1571_),
    .A2(net690));
 sg13g2_a21oi_1 _4361_ (.A1(net376),
    .A2(net633),
    .Y(_0220_),
    .B1(_1571_));
 sg13g2_nand3_1 _4362_ (.B(_1483_),
    .C(_1484_),
    .A(_1481_),
    .Y(_1572_));
 sg13g2_nor2_1 _4363_ (.A(net659),
    .B(_1485_),
    .Y(_1573_));
 sg13g2_o21ai_1 _4364_ (.B1(net667),
    .Y(_1574_),
    .A1(net657),
    .A2(_1468_));
 sg13g2_a21oi_1 _4365_ (.A1(_1572_),
    .A2(_1573_),
    .Y(_1575_),
    .B1(_1574_));
 sg13g2_a21oi_1 _4366_ (.A1(net302),
    .A2(net663),
    .Y(_1576_),
    .B1(_0940_));
 sg13g2_nor2b_2 _4367_ (.A(_1575_),
    .B_N(_1576_),
    .Y(_1577_));
 sg13g2_a21o_1 _4368_ (.A2(_1317_),
    .A1(_1314_),
    .B1(_1312_),
    .X(_1578_));
 sg13g2_nand3_1 _4369_ (.B(_1318_),
    .C(_1578_),
    .A(net656),
    .Y(_1579_));
 sg13g2_a21oi_1 _4370_ (.A1(net658),
    .A2(_1307_),
    .Y(_1580_),
    .B1(net662));
 sg13g2_a221oi_1 _4371_ (.B2(_1580_),
    .C1(_1516_),
    .B1(_1579_),
    .A1(_0056_),
    .Y(_1581_),
    .A2(net662));
 sg13g2_a22oi_1 _4372_ (.Y(_1582_),
    .B1(_1189_),
    .B2(net427),
    .A2(_0943_),
    .A1(_2111_));
 sg13g2_o21ai_1 _4373_ (.B1(_1582_),
    .Y(_1583_),
    .A1(_2071_),
    .A2(_2076_));
 sg13g2_nor4_2 _4374_ (.A(_2109_),
    .B(_1577_),
    .C(_1581_),
    .Y(_1584_),
    .D(_1583_));
 sg13g2_nand2b_1 _4375_ (.Y(_1585_),
    .B(_1188_),
    .A_N(_1584_));
 sg13g2_o21ai_1 _4376_ (.B1(_0954_),
    .Y(_1586_),
    .A1(net244),
    .A2(_1117_));
 sg13g2_a22oi_1 _4377_ (.Y(_0221_),
    .B1(_1585_),
    .B2(_1586_),
    .A2(net633),
    .A1(net468));
 sg13g2_nor3_1 _4378_ (.A(_1351_),
    .B(_1353_),
    .C(_1482_),
    .Y(_1587_));
 sg13g2_nand2_1 _4379_ (.Y(_1588_),
    .A(net657),
    .B(_1483_));
 sg13g2_a21oi_1 _4380_ (.A1(net658),
    .A2(_1473_),
    .Y(_1589_),
    .B1(net662));
 sg13g2_o21ai_1 _4381_ (.B1(_1589_),
    .Y(_1590_),
    .A1(_1587_),
    .A2(_1588_));
 sg13g2_a21oi_1 _4382_ (.A1(net289),
    .A2(net663),
    .Y(_1591_),
    .B1(_0940_));
 sg13g2_nand2_2 _4383_ (.Y(_1592_),
    .A(_1590_),
    .B(_1591_));
 sg13g2_and3_1 _4384_ (.X(_1593_),
    .A(net657),
    .B(_1314_),
    .C(_1315_));
 sg13g2_a21oi_1 _4385_ (.A1(_1316_),
    .A2(_1593_),
    .Y(_1594_),
    .B1(net663));
 sg13g2_o21ai_1 _4386_ (.B1(_1594_),
    .Y(_1595_),
    .A1(_1316_),
    .A2(_1593_));
 sg13g2_a21oi_1 _4387_ (.A1(net1007),
    .A2(net664),
    .Y(_1596_),
    .B1(_1516_));
 sg13g2_a221oi_1 _4388_ (.B2(_1596_),
    .C1(_2109_),
    .B1(_1595_),
    .A1(net322),
    .Y(_1597_),
    .A2(_1189_));
 sg13g2_nand2_1 _4389_ (.Y(_1598_),
    .A(_1592_),
    .B(_1597_));
 sg13g2_a221oi_1 _4390_ (.B2(_1598_),
    .C1(net633),
    .B1(_1188_),
    .A1(net340),
    .Y(_1599_),
    .A2(net691));
 sg13g2_a21oi_1 _4391_ (.A1(net245),
    .A2(net634),
    .Y(_0222_),
    .B1(_1599_));
 sg13g2_nor2b_1 _4392_ (.A(net225),
    .B_N(net186),
    .Y(_1600_));
 sg13g2_a21oi_1 _4393_ (.A1(_0955_),
    .A2(_1600_),
    .Y(_1601_),
    .B1(net690));
 sg13g2_a21oi_1 _4394_ (.A1(net690),
    .A2(_0944_),
    .Y(_1602_),
    .B1(_1601_));
 sg13g2_or4_2 _4395_ (.A(_2117_),
    .B(_1177_),
    .C(_1179_),
    .D(_1602_),
    .X(_1603_));
 sg13g2_a21oi_1 _4396_ (.A1(_2011_),
    .A2(_0941_),
    .Y(_1604_),
    .B1(_2075_));
 sg13g2_nand3_1 _4397_ (.B(_0957_),
    .C(_1604_),
    .A(_2166_),
    .Y(_1605_));
 sg13g2_mux2_1 _4398_ (.A0(_1605_),
    .A1(net548),
    .S(_1603_),
    .X(_0223_));
 sg13g2_a21oi_1 _4399_ (.A1(net333),
    .A2(_0941_),
    .Y(_1606_),
    .B1(_0956_));
 sg13g2_nand3_1 _4400_ (.B(_2074_),
    .C(_2164_),
    .A(net604),
    .Y(_1607_));
 sg13g2_nand3b_1 _4401_ (.B(_1606_),
    .C(net605),
    .Y(_1608_),
    .A_N(_2109_));
 sg13g2_mux2_1 _4402_ (.A0(net606),
    .A1(net734),
    .S(_1603_),
    .X(_0224_));
 sg13g2_nand3_1 _4403_ (.B(net610),
    .C(_1180_),
    .A(_0940_),
    .Y(_1609_));
 sg13g2_mux2_1 _4404_ (.A0(net611),
    .A1(net733),
    .S(_1603_),
    .X(_0225_));
 sg13g2_nand2_1 _4405_ (.Y(_1610_),
    .A(_0937_),
    .B(_1176_));
 sg13g2_nor2_1 _4406_ (.A(_1603_),
    .B(_1610_),
    .Y(_1611_));
 sg13g2_a21oi_1 _4407_ (.A1(net589),
    .A2(_1603_),
    .Y(_0226_),
    .B1(_1611_));
 sg13g2_o21ai_1 _4408_ (.B1(net634),
    .Y(_1612_),
    .A1(net506),
    .A2(net692));
 sg13g2_inv_1 _4409_ (.Y(_0227_),
    .A(net507));
 sg13g2_nand2_1 _4410_ (.Y(_1613_),
    .A(net238),
    .B(net634));
 sg13g2_o21ai_1 _4411_ (.B1(net239),
    .Y(_0228_),
    .A1(net238),
    .A2(_1117_));
 sg13g2_a21oi_1 _4412_ (.A1(net506),
    .A2(net238),
    .Y(_1614_),
    .B1(net160));
 sg13g2_or3_1 _4413_ (.A(net504),
    .B(_0952_),
    .C(_1614_),
    .X(_1615_));
 sg13g2_o21ai_1 _4414_ (.B1(_1615_),
    .Y(_0229_),
    .A1(net161),
    .A2(_0951_));
 sg13g2_a21oi_1 _4415_ (.A1(net210),
    .A2(_0950_),
    .Y(_1616_),
    .B1(net692));
 sg13g2_nor2_1 _4416_ (.A(net210),
    .B(_0952_),
    .Y(_1617_));
 sg13g2_nor3_1 _4417_ (.A(_0953_),
    .B(_1616_),
    .C(net211),
    .Y(_0230_));
 sg13g2_a21oi_1 _4418_ (.A1(_1979_),
    .A2(net576),
    .Y(_1618_),
    .B1(_2157_));
 sg13g2_and2_1 _4419_ (.A(_2066_),
    .B(_1618_),
    .X(_1619_));
 sg13g2_nand2_1 _4420_ (.Y(_1620_),
    .A(_2166_),
    .B(_1619_));
 sg13g2_and2_1 _4421_ (.A(net576),
    .B(_2067_),
    .X(_1621_));
 sg13g2_a21oi_1 _4422_ (.A1(_2076_),
    .A2(_1621_),
    .Y(_1622_),
    .B1(_2180_));
 sg13g2_nand3b_1 _4423_ (.B(_1620_),
    .C(_1622_),
    .Y(_1623_),
    .A_N(_2161_));
 sg13g2_a21o_1 _4424_ (.A2(_2099_),
    .A1(_2077_),
    .B1(_1623_),
    .X(_1624_));
 sg13g2_o21ai_1 _4425_ (.B1(_2158_),
    .Y(_1625_),
    .A1(net348),
    .A2(_1011_));
 sg13g2_a21oi_1 _4426_ (.A1(net413),
    .A2(_0831_),
    .Y(_1626_),
    .B1(_2066_));
 sg13g2_nor2b_1 _4427_ (.A(_1626_),
    .B_N(_2067_),
    .Y(_1627_));
 sg13g2_nor4_1 _4428_ (.A(net673),
    .B(_1619_),
    .C(_1624_),
    .D(_1627_),
    .Y(_1628_));
 sg13g2_a22oi_1 _4429_ (.Y(_0231_),
    .B1(_1625_),
    .B2(_1628_),
    .A2(_1624_),
    .A1(net621));
 sg13g2_nor3_1 _4430_ (.A(net945),
    .B(_2174_),
    .C(_1623_),
    .Y(_1629_));
 sg13g2_a22oi_1 _4431_ (.Y(_0232_),
    .B1(_1625_),
    .B2(_1629_),
    .A2(_1624_),
    .A1(net577));
 sg13g2_a21oi_1 _4432_ (.A1(_2077_),
    .A2(_2099_),
    .Y(_1630_),
    .B1(_2070_));
 sg13g2_nor3_1 _4433_ (.A(_2070_),
    .B(_1618_),
    .C(_1624_),
    .Y(_1631_));
 sg13g2_a22oi_1 _4434_ (.Y(_0233_),
    .B1(_1625_),
    .B2(_1631_),
    .A2(_1624_),
    .A1(net580));
 sg13g2_nand2_1 _4435_ (.Y(_1632_),
    .A(net732),
    .B(net415));
 sg13g2_nand4_1 _4436_ (.B(net415),
    .C(\measurements.address_counter_reg[2] ),
    .A(net731),
    .Y(_1633_),
    .D(net365));
 sg13g2_inv_1 _4437_ (.Y(_1634_),
    .A(_1633_));
 sg13g2_nand3_1 _4438_ (.B(\measurements.address_counter_reg[5] ),
    .C(_1634_),
    .A(net459),
    .Y(_1635_));
 sg13g2_nand2_1 _4439_ (.Y(_1636_),
    .A(\measurements.address_counter_reg[6] ),
    .B(net325));
 sg13g2_nor2_2 _4440_ (.A(_1635_),
    .B(_1636_),
    .Y(_1637_));
 sg13g2_nand3_1 _4441_ (.B(net219),
    .C(_1637_),
    .A(net207),
    .Y(_1638_));
 sg13g2_inv_1 _4442_ (.Y(_1639_),
    .A(_1638_));
 sg13g2_nand3_1 _4443_ (.B(net101),
    .C(_1639_),
    .A(net213),
    .Y(_1640_));
 sg13g2_inv_1 _4444_ (.Y(_1641_),
    .A(_1640_));
 sg13g2_nand3_1 _4445_ (.B(net362),
    .C(_1641_),
    .A(net297),
    .Y(_1642_));
 sg13g2_nor4_1 _4446_ (.A(\measurements.alreadytriggered_reg ),
    .B(\measurements.address_counter_reg[14] ),
    .C(_0958_),
    .D(_1642_),
    .Y(_1643_));
 sg13g2_nor2_1 _4447_ (.A(net134),
    .B(_1643_),
    .Y(_1644_));
 sg13g2_nor3_1 _4448_ (.A(net347),
    .B(_2155_),
    .C(_0958_),
    .Y(_1645_));
 sg13g2_nor2_1 _4449_ (.A(net135),
    .B(_1645_),
    .Y(_0235_));
 sg13g2_nand2_1 _4450_ (.Y(_1646_),
    .A(_2077_),
    .B(_0831_));
 sg13g2_nand3_1 _4451_ (.B(_0438_),
    .C(_0532_),
    .A(_2213_),
    .Y(_1647_));
 sg13g2_nand2_1 _4452_ (.Y(_1648_),
    .A(_1979_),
    .B(_1647_));
 sg13g2_a21o_1 _4453_ (.A2(_1648_),
    .A1(_1621_),
    .B1(_2068_),
    .X(_1649_));
 sg13g2_nand4_1 _4454_ (.B(_1630_),
    .C(_1646_),
    .A(_1622_),
    .Y(_1650_),
    .D(_1649_));
 sg13g2_nand2_1 _4455_ (.Y(_1651_),
    .A(_2049_),
    .B(net666));
 sg13g2_o21ai_1 _4456_ (.B1(_1651_),
    .Y(_1652_),
    .A1(net322),
    .A2(net666));
 sg13g2_nand2_1 _4457_ (.Y(_1653_),
    .A(net119),
    .B(net644));
 sg13g2_o21ai_1 _4458_ (.B1(net120),
    .Y(_0236_),
    .A1(net644),
    .A2(_1652_));
 sg13g2_nand2_1 _4459_ (.Y(_1654_),
    .A(_2048_),
    .B(net666));
 sg13g2_o21ai_1 _4460_ (.B1(_1654_),
    .Y(_1655_),
    .A1(net427),
    .A2(net666));
 sg13g2_nand2_1 _4461_ (.Y(_1656_),
    .A(net173),
    .B(net644));
 sg13g2_o21ai_1 _4462_ (.B1(net174),
    .Y(_0237_),
    .A1(net644),
    .A2(_1655_));
 sg13g2_nand2_1 _4463_ (.Y(_1657_),
    .A(_2047_),
    .B(net667));
 sg13g2_o21ai_1 _4464_ (.B1(_1657_),
    .Y(_1658_),
    .A1(net399),
    .A2(net667));
 sg13g2_nand2_1 _4465_ (.Y(_1659_),
    .A(net192),
    .B(net644));
 sg13g2_o21ai_1 _4466_ (.B1(net193),
    .Y(_0238_),
    .A1(net644),
    .A2(_1658_));
 sg13g2_nand2_1 _4467_ (.Y(_1660_),
    .A(net317),
    .B(net666));
 sg13g2_o21ai_1 _4468_ (.B1(_1660_),
    .Y(_1661_),
    .A1(net305),
    .A2(net666));
 sg13g2_nand2_1 _4469_ (.Y(_1662_),
    .A(net387),
    .B(net644));
 sg13g2_o21ai_1 _4470_ (.B1(net388),
    .Y(_0239_),
    .A1(net644),
    .A2(_1661_));
 sg13g2_mux2_1 _4471_ (.A0(_1985_),
    .A1(_2045_),
    .S(net666),
    .X(_1663_));
 sg13g2_nand2_1 _4472_ (.Y(_1664_),
    .A(net429),
    .B(net643));
 sg13g2_o21ai_1 _4473_ (.B1(net430),
    .Y(_0240_),
    .A1(net643),
    .A2(_1663_));
 sg13g2_nand2_1 _4474_ (.Y(_1665_),
    .A(net357),
    .B(net664));
 sg13g2_o21ai_1 _4475_ (.B1(_1665_),
    .Y(_1666_),
    .A1(_2044_),
    .A2(net664));
 sg13g2_nor2_1 _4476_ (.A(net643),
    .B(_1666_),
    .Y(_1667_));
 sg13g2_a21oi_1 _4477_ (.A1(net329),
    .A2(net643),
    .Y(_0241_),
    .B1(_1667_));
 sg13g2_nor2_1 _4478_ (.A(net525),
    .B(net664),
    .Y(_1668_));
 sg13g2_a21oi_1 _4479_ (.A1(_1988_),
    .A2(net664),
    .Y(_1669_),
    .B1(_1668_));
 sg13g2_nor2_1 _4480_ (.A(net643),
    .B(_1669_),
    .Y(_1670_));
 sg13g2_a21oi_1 _4481_ (.A1(net379),
    .A2(net643),
    .Y(_0242_),
    .B1(_1670_));
 sg13g2_nand2_1 _4482_ (.Y(_1671_),
    .A(_2050_),
    .B(net666));
 sg13g2_o21ai_1 _4483_ (.B1(_1671_),
    .Y(_1672_),
    .A1(net345),
    .A2(net667));
 sg13g2_nand2_1 _4484_ (.Y(_1673_),
    .A(net446),
    .B(net643));
 sg13g2_o21ai_1 _4485_ (.B1(net447),
    .Y(_0243_),
    .A1(net643),
    .A2(_1672_));
 sg13g2_a21o_1 _4486_ (.A2(_2155_),
    .A1(net117),
    .B1(_0958_),
    .X(_1674_));
 sg13g2_o21ai_1 _4487_ (.B1(_1674_),
    .Y(_0244_),
    .A1(net348),
    .A2(_1149_));
 sg13g2_nor2_1 _4488_ (.A(net532),
    .B(_0615_),
    .Y(_1675_));
 sg13g2_a21oi_1 _4489_ (.A1(net532),
    .A2(_0614_),
    .Y(_0245_),
    .B1(_1675_));
 sg13g2_a21oi_1 _4490_ (.A1(_2174_),
    .A2(_1632_),
    .Y(_1676_),
    .B1(net648));
 sg13g2_a21oi_1 _4491_ (.A1(net732),
    .A2(_0614_),
    .Y(_1677_),
    .B1(net415));
 sg13g2_nor2_1 _4492_ (.A(_1676_),
    .B(net416),
    .Y(_0246_));
 sg13g2_nor2_1 _4493_ (.A(_0057_),
    .B(_1632_),
    .Y(_1678_));
 sg13g2_xnor2_1 _4494_ (.Y(_1679_),
    .A(net934),
    .B(_1632_));
 sg13g2_a22oi_1 _4495_ (.Y(_1680_),
    .B1(net648),
    .B2(\measurements.address_counter_reg[2] ),
    .A2(net673),
    .A1(net313));
 sg13g2_o21ai_1 _4496_ (.B1(net314),
    .Y(_0247_),
    .A1(net645),
    .A2(_1679_));
 sg13g2_xor2_1 _4497_ (.B(_1678_),
    .A(net449),
    .X(_1681_));
 sg13g2_a22oi_1 _4498_ (.Y(_1682_),
    .B1(net648),
    .B2(net365),
    .A2(net673),
    .A1(_0447_));
 sg13g2_o21ai_1 _4499_ (.B1(_1682_),
    .Y(_0248_),
    .A1(net645),
    .A2(net450));
 sg13g2_nor2_1 _4500_ (.A(net473),
    .B(_1633_),
    .Y(_1683_));
 sg13g2_xnor2_1 _4501_ (.Y(_1684_),
    .A(net473),
    .B(_1633_));
 sg13g2_a22oi_1 _4502_ (.Y(_1685_),
    .B1(net648),
    .B2(net459),
    .A2(net673),
    .A1(_0453_));
 sg13g2_o21ai_1 _4503_ (.B1(_1685_),
    .Y(_0249_),
    .A1(net645),
    .A2(net474));
 sg13g2_xor2_1 _4504_ (.B(_1683_),
    .A(net476),
    .X(_1686_));
 sg13g2_a22oi_1 _4505_ (.Y(_1687_),
    .B1(net648),
    .B2(net898),
    .A2(net673),
    .A1(_0450_));
 sg13g2_o21ai_1 _4506_ (.B1(net899),
    .Y(_0250_),
    .A1(net645),
    .A2(net477));
 sg13g2_nor2_1 _4507_ (.A(net432),
    .B(_1635_),
    .Y(_1688_));
 sg13g2_xnor2_1 _4508_ (.Y(_1689_),
    .A(net432),
    .B(net460));
 sg13g2_a22oi_1 _4509_ (.Y(_1690_),
    .B1(net648),
    .B2(net394),
    .A2(net673),
    .A1(_0455_));
 sg13g2_o21ai_1 _4510_ (.B1(_1690_),
    .Y(_0251_),
    .A1(net645),
    .A2(net461));
 sg13g2_xor2_1 _4511_ (.B(net433),
    .A(_0062_),
    .X(_1691_));
 sg13g2_a22oi_1 _4512_ (.Y(_1692_),
    .B1(net648),
    .B2(net325),
    .A2(net673),
    .A1(_0458_));
 sg13g2_o21ai_1 _4513_ (.B1(_1692_),
    .Y(_0252_),
    .A1(net645),
    .A2(net434));
 sg13g2_nand2b_1 _4514_ (.Y(_1693_),
    .B(_1637_),
    .A_N(net289));
 sg13g2_xor2_1 _4515_ (.B(_1637_),
    .A(net289),
    .X(_1694_));
 sg13g2_a22oi_1 _4516_ (.Y(_1695_),
    .B1(net648),
    .B2(net207),
    .A2(net673),
    .A1(_0452_));
 sg13g2_o21ai_1 _4517_ (.B1(_1695_),
    .Y(_0253_),
    .A1(net645),
    .A2(net290));
 sg13g2_o21ai_1 _4518_ (.B1(_0615_),
    .Y(_1696_),
    .A1(net302),
    .A2(_1693_));
 sg13g2_a21oi_1 _4519_ (.A1(net302),
    .A2(_1693_),
    .Y(_1697_),
    .B1(_1696_));
 sg13g2_a21o_1 _4520_ (.A2(net649),
    .A1(net219),
    .B1(net303),
    .X(_0254_));
 sg13g2_or2_1 _4521_ (.X(_1698_),
    .B(_1638_),
    .A(net285));
 sg13g2_a21oi_1 _4522_ (.A1(net285),
    .A2(_1638_),
    .Y(_1699_),
    .B1(net645));
 sg13g2_a22oi_1 _4523_ (.Y(_1700_),
    .B1(_1698_),
    .B2(net286),
    .A2(net649),
    .A1(net213));
 sg13g2_inv_1 _4524_ (.Y(_0255_),
    .A(net287));
 sg13g2_a21oi_1 _4525_ (.A1(net390),
    .A2(_1698_),
    .Y(_1701_),
    .B1(net646));
 sg13g2_o21ai_1 _4526_ (.B1(net391),
    .Y(_1702_),
    .A1(net390),
    .A2(_1698_));
 sg13g2_o21ai_1 _4527_ (.B1(net392),
    .Y(_0256_),
    .A1(_2006_),
    .A2(_0614_));
 sg13g2_nand2_1 _4528_ (.Y(_1703_),
    .A(net297),
    .B(net649));
 sg13g2_nor2_1 _4529_ (.A(net909),
    .B(_1640_),
    .Y(_1704_));
 sg13g2_a21o_1 _4530_ (.A2(_1640_),
    .A1(net909),
    .B1(net646),
    .X(_1705_));
 sg13g2_o21ai_1 _4531_ (.B1(net298),
    .Y(_0257_),
    .A1(_1704_),
    .A2(_1705_));
 sg13g2_nand2_1 _4532_ (.Y(_1706_),
    .A(net362),
    .B(net649));
 sg13g2_xor2_1 _4533_ (.B(_1704_),
    .A(net903),
    .X(_1707_));
 sg13g2_o21ai_1 _4534_ (.B1(net363),
    .Y(_0258_),
    .A1(net646),
    .A2(net904));
 sg13g2_xnor2_1 _4535_ (.Y(_1708_),
    .A(net949),
    .B(_1642_));
 sg13g2_a22oi_1 _4536_ (.Y(_0259_),
    .B1(_0615_),
    .B2(_1708_),
    .A2(net649),
    .A1(net129));
 sg13g2_nand2_1 _4537_ (.Y(_1709_),
    .A(net256),
    .B(_0605_));
 sg13g2_nor2_1 _4538_ (.A(net971),
    .B(\siggen.da_cs ),
    .Y(_1710_));
 sg13g2_a21oi_1 _4539_ (.A1(_1709_),
    .A2(_1710_),
    .Y(_1711_),
    .B1(_0843_));
 sg13g2_a21o_2 _4540_ (.A2(_1710_),
    .A1(_1709_),
    .B1(_0843_),
    .X(_1712_));
 sg13g2_nand2_2 _4541_ (.Y(_1713_),
    .A(net714),
    .B(net715));
 sg13g2_a21oi_1 _4542_ (.A1(net721),
    .A2(_2054_),
    .Y(_1714_),
    .B1(_1713_));
 sg13g2_nor2b_2 _4543_ (.A(net729),
    .B_N(net727),
    .Y(_1715_));
 sg13g2_nor2b_2 _4544_ (.A(net727),
    .B_N(net729),
    .Y(_1716_));
 sg13g2_nor2_1 _4545_ (.A(_1715_),
    .B(_1716_),
    .Y(_1717_));
 sg13g2_o21ai_1 _4546_ (.B1(_1714_),
    .Y(_1718_),
    .A1(net721),
    .A2(_1717_));
 sg13g2_nor2_2 _4547_ (.A(net714),
    .B(net718),
    .Y(_1719_));
 sg13g2_nand2_1 _4548_ (.Y(_1720_),
    .A(net723),
    .B(net726));
 sg13g2_nor2b_1 _4549_ (.A(net714),
    .B_N(net716),
    .Y(_1721_));
 sg13g2_and2_1 _4550_ (.A(net728),
    .B(net681),
    .X(_1722_));
 sg13g2_nand2b_2 _4551_ (.Y(_1723_),
    .B(net722),
    .A_N(net728));
 sg13g2_and2_2 _4552_ (.A(net724),
    .B(_1715_),
    .X(_1724_));
 sg13g2_nand2b_2 _4553_ (.Y(_1725_),
    .B(net714),
    .A_N(net715));
 sg13g2_nor2_1 _4554_ (.A(net721),
    .B(_0036_),
    .Y(_1726_));
 sg13g2_nor3_2 _4555_ (.A(_1724_),
    .B(_1725_),
    .C(_1726_),
    .Y(_1727_));
 sg13g2_nor2b_2 _4556_ (.A(net721),
    .B_N(net728),
    .Y(_1728_));
 sg13g2_nor2b_1 _4557_ (.A(net721),
    .B_N(net725),
    .Y(_1729_));
 sg13g2_nor3_1 _4558_ (.A(_1713_),
    .B(_1728_),
    .C(_1729_),
    .Y(_1730_));
 sg13g2_and2_2 _4559_ (.A(net728),
    .B(net725),
    .X(_1731_));
 sg13g2_nand2_2 _4560_ (.Y(_1732_),
    .A(net728),
    .B(net725));
 sg13g2_nand3_1 _4561_ (.B(_1723_),
    .C(_1732_),
    .A(net681),
    .Y(_1733_));
 sg13g2_a221oi_1 _4562_ (.B2(_1722_),
    .C1(net711),
    .B1(_1720_),
    .A1(_0036_),
    .Y(_1734_),
    .A2(_1719_));
 sg13g2_nor2_1 _4563_ (.A(net694),
    .B(_1730_),
    .Y(_1735_));
 sg13g2_a22oi_1 _4564_ (.Y(_1736_),
    .B1(_1735_),
    .B2(_1733_),
    .A2(_1734_),
    .A1(_1718_));
 sg13g2_nor3_1 _4565_ (.A(_2055_),
    .B(_1727_),
    .C(_1736_),
    .Y(_1737_));
 sg13g2_nor2_1 _4566_ (.A(net267),
    .B(_1737_),
    .Y(_1738_));
 sg13g2_nor2_2 _4567_ (.A(net724),
    .B(_1716_),
    .Y(_1739_));
 sg13g2_inv_1 _4568_ (.Y(_1740_),
    .A(_1739_));
 sg13g2_a21o_1 _4569_ (.A2(net720),
    .A1(net728),
    .B1(_1739_),
    .X(_1741_));
 sg13g2_o21ai_1 _4570_ (.B1(_1719_),
    .Y(_1742_),
    .A1(_0038_),
    .A2(_1731_));
 sg13g2_nor2_1 _4571_ (.A(net728),
    .B(net725),
    .Y(_1743_));
 sg13g2_nor3_1 _4572_ (.A(_1725_),
    .B(_1728_),
    .C(_1743_),
    .Y(_1744_));
 sg13g2_a21oi_1 _4573_ (.A1(net681),
    .A2(_1741_),
    .Y(_1745_),
    .B1(_1744_));
 sg13g2_a21oi_1 _4574_ (.A1(_1742_),
    .A2(_1745_),
    .Y(_1746_),
    .B1(net710));
 sg13g2_nor2_1 _4575_ (.A(net725),
    .B(_1728_),
    .Y(_1747_));
 sg13g2_o21ai_1 _4576_ (.B1(_1741_),
    .Y(_1748_),
    .A1(net717),
    .A2(net725));
 sg13g2_nor2b_2 _4577_ (.A(net717),
    .B_N(net721),
    .Y(_1749_));
 sg13g2_a21oi_1 _4578_ (.A1(_1743_),
    .A2(_1749_),
    .Y(_1750_),
    .B1(net712));
 sg13g2_a21o_1 _4579_ (.A2(net715),
    .A1(net729),
    .B1(net693),
    .X(_1751_));
 sg13g2_nor2_1 _4580_ (.A(net720),
    .B(_1715_),
    .Y(_1752_));
 sg13g2_nor2b_1 _4581_ (.A(_0036_),
    .B_N(net720),
    .Y(_1753_));
 sg13g2_nor2_1 _4582_ (.A(net719),
    .B(net723),
    .Y(_1754_));
 sg13g2_or2_1 _4583_ (.X(_1755_),
    .B(net723),
    .A(net718));
 sg13g2_nand2b_1 _4584_ (.Y(_1756_),
    .B(_1715_),
    .A_N(net717));
 sg13g2_nor3_1 _4585_ (.A(net715),
    .B(_1752_),
    .C(_1753_),
    .Y(_1757_));
 sg13g2_o21ai_1 _4586_ (.B1(net710),
    .Y(_1758_),
    .A1(_1751_),
    .A2(_1757_));
 sg13g2_a21oi_1 _4587_ (.A1(_1748_),
    .A2(_1750_),
    .Y(_1759_),
    .B1(_1758_));
 sg13g2_o21ai_1 _4588_ (.B1(net709),
    .Y(_1760_),
    .A1(_1746_),
    .A2(_1759_));
 sg13g2_or2_2 _4589_ (.X(_1761_),
    .B(\oscilloscope_control.n220_q[1] ),
    .A(net980));
 sg13g2_nor2_1 _4590_ (.A(net267),
    .B(net708),
    .Y(_1762_));
 sg13g2_nor2b_1 _4591_ (.A(_1737_),
    .B_N(_1762_),
    .Y(_1763_));
 sg13g2_nor2_1 _4592_ (.A(_1761_),
    .B(_1763_),
    .Y(_1764_));
 sg13g2_xnor2_1 _4593_ (.Y(_1765_),
    .A(_2056_),
    .B(_1760_));
 sg13g2_o21ai_1 _4594_ (.B1(_1764_),
    .Y(_1766_),
    .A1(_1738_),
    .A2(_1765_));
 sg13g2_or2_1 _4595_ (.X(_1767_),
    .B(_0930_),
    .A(_2056_));
 sg13g2_nor2b_2 _4596_ (.A(net980),
    .B_N(\oscilloscope_control.n220_q[1] ),
    .Y(_1768_));
 sg13g2_o21ai_1 _4597_ (.B1(_1768_),
    .Y(_1769_),
    .A1(_2051_),
    .A2(_2056_));
 sg13g2_a21oi_1 _4598_ (.A1(_1767_),
    .A2(_1769_),
    .Y(_1770_),
    .B1(_1762_));
 sg13g2_nand2_2 _4599_ (.Y(_1771_),
    .A(net558),
    .B(net515));
 sg13g2_o21ai_1 _4600_ (.B1(_1766_),
    .Y(_1772_),
    .A1(net920),
    .A2(_1771_));
 sg13g2_o21ai_1 _4601_ (.B1(_0843_),
    .Y(_1773_),
    .A1(_1770_),
    .A2(_1772_));
 sg13g2_o21ai_1 _4602_ (.B1(_1773_),
    .Y(_0260_),
    .A1(net138),
    .A2(_1712_));
 sg13g2_nand2_1 _4603_ (.Y(_1774_),
    .A(net76),
    .B(net654));
 sg13g2_o21ai_1 _4604_ (.B1(_1719_),
    .Y(_1775_),
    .A1(_1724_),
    .A2(_1728_));
 sg13g2_a21oi_1 _4605_ (.A1(net720),
    .A2(net727),
    .Y(_1776_),
    .B1(_1739_));
 sg13g2_o21ai_1 _4606_ (.B1(_1775_),
    .Y(_1777_),
    .A1(_1725_),
    .A2(_1776_));
 sg13g2_o21ai_1 _4607_ (.B1(net723),
    .Y(_1778_),
    .A1(net729),
    .A2(net726));
 sg13g2_o21ai_1 _4608_ (.B1(_1740_),
    .Y(_1779_),
    .A1(_1731_),
    .A2(_1778_));
 sg13g2_nor2_1 _4609_ (.A(net717),
    .B(_2054_),
    .Y(_1780_));
 sg13g2_o21ai_1 _4610_ (.B1(net712),
    .Y(_1781_),
    .A1(net721),
    .A2(_1780_));
 sg13g2_a21oi_1 _4611_ (.A1(_1731_),
    .A2(_1749_),
    .Y(_1782_),
    .B1(_1781_));
 sg13g2_nor2_2 _4612_ (.A(net709),
    .B(_2055_),
    .Y(_1783_));
 sg13g2_o21ai_1 _4613_ (.B1(net718),
    .Y(_1784_),
    .A1(net725),
    .A2(_1728_));
 sg13g2_nor2b_1 _4614_ (.A(net717),
    .B_N(_0038_),
    .Y(_1785_));
 sg13g2_nor2_1 _4615_ (.A(net712),
    .B(_1785_),
    .Y(_1786_));
 sg13g2_nor2_1 _4616_ (.A(_1715_),
    .B(_1740_),
    .Y(_1787_));
 sg13g2_nor3_1 _4617_ (.A(net715),
    .B(_1724_),
    .C(_1787_),
    .Y(_1788_));
 sg13g2_nor2_1 _4618_ (.A(_1751_),
    .B(_1788_),
    .Y(_1789_));
 sg13g2_a21oi_1 _4619_ (.A1(_1784_),
    .A2(_1786_),
    .Y(_1790_),
    .B1(_1789_));
 sg13g2_nor3_1 _4620_ (.A(_1713_),
    .B(_1739_),
    .C(_1753_),
    .Y(_1791_));
 sg13g2_nand2_2 _4621_ (.Y(_1792_),
    .A(net718),
    .B(net723));
 sg13g2_nand2_2 _4622_ (.Y(_1793_),
    .A(net722),
    .B(net681));
 sg13g2_nor2b_2 _4623_ (.A(net722),
    .B_N(net718),
    .Y(_1794_));
 sg13g2_nand3_1 _4624_ (.B(_0039_),
    .C(_1794_),
    .A(_2053_),
    .Y(_1795_));
 sg13g2_or2_1 _4625_ (.X(_1796_),
    .B(_1716_),
    .A(net715));
 sg13g2_a21oi_1 _4626_ (.A1(_1793_),
    .A2(_1796_),
    .Y(_1797_),
    .B1(_1715_));
 sg13g2_o21ai_1 _4627_ (.B1(_1795_),
    .Y(_1798_),
    .A1(_1723_),
    .A2(_1725_));
 sg13g2_nor3_1 _4628_ (.A(_1791_),
    .B(_1797_),
    .C(_1798_),
    .Y(_1799_));
 sg13g2_a221oi_1 _4629_ (.B2(_1779_),
    .C1(_1782_),
    .B1(_1721_),
    .A1(_0036_),
    .Y(_1800_),
    .A2(_1719_));
 sg13g2_mux2_1 _4630_ (.A0(_1799_),
    .A1(_1800_),
    .S(net710),
    .X(_1801_));
 sg13g2_a221oi_1 _4631_ (.B2(_1752_),
    .C1(_1777_),
    .B1(net681),
    .A1(net715),
    .Y(_1802_),
    .A2(_1717_));
 sg13g2_o21ai_1 _4632_ (.B1(net709),
    .Y(_1803_),
    .A1(net694),
    .A2(_1802_));
 sg13g2_a21oi_1 _4633_ (.A1(net694),
    .A2(_1790_),
    .Y(_1804_),
    .B1(_1803_));
 sg13g2_a21oi_1 _4634_ (.A1(_1783_),
    .A2(_1801_),
    .Y(_1805_),
    .B1(_1804_));
 sg13g2_or2_2 _4635_ (.X(_1806_),
    .B(_1761_),
    .A(_2056_));
 sg13g2_nor2b_1 _4636_ (.A(_1806_),
    .B_N(_1805_),
    .Y(_1807_));
 sg13g2_nor2_2 _4637_ (.A(net708),
    .B(_1761_),
    .Y(_1808_));
 sg13g2_nor2b_1 _4638_ (.A(_1805_),
    .B_N(_1808_),
    .Y(_1809_));
 sg13g2_and2_2 _4639_ (.A(net682),
    .B(_1767_),
    .X(_1810_));
 sg13g2_o21ai_1 _4640_ (.B1(_1768_),
    .Y(_1811_),
    .A1(net729),
    .A2(net707));
 sg13g2_a21oi_1 _4641_ (.A1(net728),
    .A2(net707),
    .Y(_1812_),
    .B1(_1811_));
 sg13g2_o21ai_1 _4642_ (.B1(_1810_),
    .Y(_1813_),
    .A1(net979),
    .A2(_1771_));
 sg13g2_nor4_1 _4643_ (.A(_1807_),
    .B(_1809_),
    .C(_1812_),
    .D(_1813_),
    .Y(_1814_));
 sg13g2_o21ai_1 _4644_ (.B1(_1712_),
    .Y(_1815_),
    .A1(net137),
    .A2(net682));
 sg13g2_o21ai_1 _4645_ (.B1(net77),
    .Y(_0261_),
    .A1(_1814_),
    .A2(_1815_));
 sg13g2_nand2_1 _4646_ (.Y(_1816_),
    .A(net87),
    .B(net654));
 sg13g2_o21ai_1 _4647_ (.B1(net715),
    .Y(_1817_),
    .A1(net714),
    .A2(_1716_));
 sg13g2_o21ai_1 _4648_ (.B1(_1817_),
    .Y(_1818_),
    .A1(_1724_),
    .A2(_1752_));
 sg13g2_o21ai_1 _4649_ (.B1(_1714_),
    .Y(_1819_),
    .A1(_1715_),
    .A2(_1740_));
 sg13g2_nand3_1 _4650_ (.B(_1716_),
    .C(net681),
    .A(net720),
    .Y(_1820_));
 sg13g2_and2_1 _4651_ (.A(_1818_),
    .B(_1820_),
    .X(_1821_));
 sg13g2_a21oi_2 _4652_ (.B1(net710),
    .Y(_1822_),
    .A2(_1821_),
    .A1(_1819_));
 sg13g2_nor2_1 _4653_ (.A(_1743_),
    .B(_1792_),
    .Y(_1823_));
 sg13g2_a21oi_1 _4654_ (.A1(_0039_),
    .A2(_1794_),
    .Y(_1824_),
    .B1(_1823_));
 sg13g2_nor2_2 _4655_ (.A(_1749_),
    .B(_1794_),
    .Y(_1825_));
 sg13g2_nor2_1 _4656_ (.A(net712),
    .B(_1780_),
    .Y(_1826_));
 sg13g2_a221oi_1 _4657_ (.B2(_1824_),
    .C1(net694),
    .B1(_1826_),
    .A1(net712),
    .Y(_1827_),
    .A2(_1825_));
 sg13g2_or3_1 _4658_ (.A(_2055_),
    .B(_1822_),
    .C(_1827_),
    .X(_1828_));
 sg13g2_nand2_1 _4659_ (.Y(_1829_),
    .A(_2051_),
    .B(_1828_));
 sg13g2_a21oi_1 _4660_ (.A1(_1723_),
    .A2(_1747_),
    .Y(_1830_),
    .B1(_1729_));
 sg13g2_a22oi_1 _4661_ (.Y(_1831_),
    .B1(_1756_),
    .B2(_1830_),
    .A2(_1754_),
    .A1(_1715_));
 sg13g2_nor3_1 _4662_ (.A(net694),
    .B(net693),
    .C(_1831_),
    .Y(_1832_));
 sg13g2_nor2b_1 _4663_ (.A(_1830_),
    .B_N(net718),
    .Y(_1833_));
 sg13g2_nor2_1 _4664_ (.A(net717),
    .B(_1729_),
    .Y(_1834_));
 sg13g2_o21ai_1 _4665_ (.B1(_1834_),
    .Y(_1835_),
    .A1(_1731_),
    .A2(_1778_));
 sg13g2_nand3_1 _4666_ (.B(net693),
    .C(_1835_),
    .A(net711),
    .Y(_1836_));
 sg13g2_nand2_1 _4667_ (.Y(_1837_),
    .A(net718),
    .B(net726));
 sg13g2_nand2_1 _4668_ (.Y(_1838_),
    .A(net713),
    .B(_1837_));
 sg13g2_nand2b_1 _4669_ (.Y(_1839_),
    .B(_1732_),
    .A_N(net721));
 sg13g2_a21oi_1 _4670_ (.A1(_1720_),
    .A2(_1839_),
    .Y(_1840_),
    .B1(net719));
 sg13g2_nor2_1 _4671_ (.A(net712),
    .B(_1749_),
    .Y(_1841_));
 sg13g2_nand2_1 _4672_ (.Y(_1842_),
    .A(net693),
    .B(_1825_));
 sg13g2_a21oi_1 _4673_ (.A1(net693),
    .A2(_1825_),
    .Y(_1843_),
    .B1(net710));
 sg13g2_o21ai_1 _4674_ (.B1(_1843_),
    .Y(_1844_),
    .A1(_1838_),
    .A2(_1840_));
 sg13g2_o21ai_1 _4675_ (.B1(_1844_),
    .Y(_1845_),
    .A1(_1833_),
    .A2(_1836_));
 sg13g2_o21ai_1 _4676_ (.B1(net709),
    .Y(_1846_),
    .A1(_1832_),
    .A2(_1845_));
 sg13g2_xnor2_1 _4677_ (.Y(_1847_),
    .A(net707),
    .B(_1846_));
 sg13g2_a221oi_1 _4678_ (.B2(_1847_),
    .C1(_1761_),
    .B1(_1829_),
    .A1(_1762_),
    .Y(_1848_),
    .A2(_1828_));
 sg13g2_o21ai_1 _4679_ (.B1(_1768_),
    .Y(_1849_),
    .A1(net726),
    .A2(net707));
 sg13g2_a21oi_1 _4680_ (.A1(net726),
    .A2(net707),
    .Y(_1850_),
    .B1(_1849_));
 sg13g2_o21ai_1 _4681_ (.B1(_1810_),
    .Y(_1851_),
    .A1(net976),
    .A2(_1771_));
 sg13g2_nor3_1 _4682_ (.A(_1848_),
    .B(_1850_),
    .C(_1851_),
    .Y(_1852_));
 sg13g2_o21ai_1 _4683_ (.B1(_1712_),
    .Y(_1853_),
    .A1(net76),
    .A2(net682));
 sg13g2_o21ai_1 _4684_ (.B1(net88),
    .Y(_0262_),
    .A1(net977),
    .A2(_1853_));
 sg13g2_nand2_1 _4685_ (.Y(_1854_),
    .A(net98),
    .B(_1711_));
 sg13g2_nand2_1 _4686_ (.Y(_1855_),
    .A(_1778_),
    .B(_1839_));
 sg13g2_or2_1 _4687_ (.X(_1856_),
    .B(_1855_),
    .A(_1725_));
 sg13g2_nand4_1 _4688_ (.B(_1742_),
    .C(_1824_),
    .A(net711),
    .Y(_1857_),
    .D(_1856_));
 sg13g2_nor2_1 _4689_ (.A(net717),
    .B(_1732_),
    .Y(_1858_));
 sg13g2_nand2_1 _4690_ (.Y(_1859_),
    .A(net712),
    .B(_0038_));
 sg13g2_o21ai_1 _4691_ (.B1(_1793_),
    .Y(_1860_),
    .A1(_1858_),
    .A2(_1859_));
 sg13g2_o21ai_1 _4692_ (.B1(_1857_),
    .Y(_1861_),
    .A1(net710),
    .A2(_1860_));
 sg13g2_nand2_1 _4693_ (.Y(_1862_),
    .A(net709),
    .B(_1861_));
 sg13g2_and3_1 _4694_ (.X(_1863_),
    .A(net681),
    .B(_1778_),
    .C(_1839_));
 sg13g2_nor3_1 _4695_ (.A(_1730_),
    .B(_1840_),
    .C(_1863_),
    .Y(_1864_));
 sg13g2_a221oi_1 _4696_ (.B2(_1841_),
    .C1(net694),
    .B1(_1778_),
    .A1(net713),
    .Y(_1865_),
    .A2(_1755_));
 sg13g2_nor2b_1 _4697_ (.A(_1865_),
    .B_N(_1783_),
    .Y(_1866_));
 sg13g2_o21ai_1 _4698_ (.B1(_1866_),
    .Y(_1867_),
    .A1(net711),
    .A2(_1864_));
 sg13g2_nand2_1 _4699_ (.Y(_1868_),
    .A(_1862_),
    .B(_1867_));
 sg13g2_o21ai_1 _4700_ (.B1(_1810_),
    .Y(_1869_),
    .A1(net597),
    .A2(_1771_));
 sg13g2_xor2_1 _4701_ (.B(net707),
    .A(net723),
    .X(_1870_));
 sg13g2_a21oi_1 _4702_ (.A1(net981),
    .A2(_1870_),
    .Y(_1871_),
    .B1(_1869_));
 sg13g2_o21ai_1 _4703_ (.B1(_1871_),
    .Y(_1872_),
    .A1(_1806_),
    .A2(_1868_));
 sg13g2_a21oi_1 _4704_ (.A1(_1808_),
    .A2(_1868_),
    .Y(_1873_),
    .B1(_1872_));
 sg13g2_o21ai_1 _4705_ (.B1(_1712_),
    .Y(_1874_),
    .A1(net87),
    .A2(net682));
 sg13g2_o21ai_1 _4706_ (.B1(net99),
    .Y(_0263_),
    .A1(net982),
    .A2(_1874_));
 sg13g2_nor2_1 _4707_ (.A(_1825_),
    .B(_1838_),
    .Y(_1875_));
 sg13g2_nand2_1 _4708_ (.Y(_1876_),
    .A(_1855_),
    .B(_1875_));
 sg13g2_nand2_1 _4709_ (.Y(_1877_),
    .A(net725),
    .B(net681));
 sg13g2_nand4_1 _4710_ (.B(_1842_),
    .C(_1876_),
    .A(net710),
    .Y(_1878_),
    .D(_1877_));
 sg13g2_nand2_1 _4711_ (.Y(_1879_),
    .A(net694),
    .B(_1792_));
 sg13g2_a21o_1 _4712_ (.A2(_1785_),
    .A1(_1732_),
    .B1(_0035_),
    .X(_1880_));
 sg13g2_o21ai_1 _4713_ (.B1(_1878_),
    .Y(_1881_),
    .A1(_1879_),
    .A2(_1880_));
 sg13g2_nor2b_1 _4714_ (.A(net712),
    .B_N(_0038_),
    .Y(_1882_));
 sg13g2_a21oi_1 _4715_ (.A1(_1732_),
    .A2(_1882_),
    .Y(_1883_),
    .B1(_1719_));
 sg13g2_a21oi_1 _4716_ (.A1(net723),
    .A2(net726),
    .Y(_1884_),
    .B1(net717));
 sg13g2_nand2_1 _4717_ (.Y(_1885_),
    .A(net694),
    .B(net693));
 sg13g2_o21ai_1 _4718_ (.B1(_1885_),
    .Y(_1886_),
    .A1(_1879_),
    .A2(_1884_));
 sg13g2_o21ai_1 _4719_ (.B1(_1886_),
    .Y(_1887_),
    .A1(_1883_),
    .A2(_1884_));
 sg13g2_nand2_1 _4720_ (.Y(_1888_),
    .A(net710),
    .B(_1786_));
 sg13g2_o21ai_1 _4721_ (.B1(_1887_),
    .Y(_1889_),
    .A1(_1823_),
    .A2(_1888_));
 sg13g2_a22oi_1 _4722_ (.Y(_1890_),
    .B1(_1889_),
    .B2(_1783_),
    .A2(_1881_),
    .A1(net709));
 sg13g2_o21ai_1 _4723_ (.B1(_1810_),
    .Y(_1891_),
    .A1(_0035_),
    .A2(_1771_));
 sg13g2_xor2_1 _4724_ (.B(net707),
    .A(net719),
    .X(_1892_));
 sg13g2_a221oi_1 _4725_ (.B2(_1768_),
    .C1(_1891_),
    .B1(_1892_),
    .A1(_1808_),
    .Y(_1893_),
    .A2(_1890_));
 sg13g2_o21ai_1 _4726_ (.B1(_1893_),
    .Y(_1894_),
    .A1(_1806_),
    .A2(_1890_));
 sg13g2_a21oi_1 _4727_ (.A1(_2058_),
    .A2(_0842_),
    .Y(_1895_),
    .B1(net654));
 sg13g2_a22oi_1 _4728_ (.Y(_1896_),
    .B1(_1894_),
    .B2(_1895_),
    .A2(net654),
    .A1(net143));
 sg13g2_inv_1 _4729_ (.Y(_0264_),
    .A(net144));
 sg13g2_nand2_1 _4730_ (.Y(_1897_),
    .A(net104),
    .B(net654));
 sg13g2_nand4_1 _4731_ (.B(net713),
    .C(net597),
    .A(net623),
    .Y(_1898_),
    .D(_1778_));
 sg13g2_and4_1 _4732_ (.A(net709),
    .B(_1793_),
    .C(_1877_),
    .D(_1879_),
    .X(_1899_));
 sg13g2_a21oi_1 _4733_ (.A1(_0037_),
    .A2(_1720_),
    .Y(_1900_),
    .B1(net693));
 sg13g2_nor2_1 _4734_ (.A(net623),
    .B(_1900_),
    .Y(_1901_));
 sg13g2_nand2_1 _4735_ (.Y(_1902_),
    .A(net926),
    .B(_1754_));
 sg13g2_a22oi_1 _4736_ (.Y(_1903_),
    .B1(_1902_),
    .B2(net623),
    .A2(_1901_),
    .A1(_1883_));
 sg13g2_a22oi_1 _4737_ (.Y(_1904_),
    .B1(_1903_),
    .B2(_1783_),
    .A2(_1899_),
    .A1(_1898_));
 sg13g2_o21ai_1 _4738_ (.B1(_1810_),
    .Y(_1905_),
    .A1(net961),
    .A2(_1771_));
 sg13g2_xor2_1 _4739_ (.B(net707),
    .A(net713),
    .X(_1906_));
 sg13g2_a21oi_1 _4740_ (.A1(_1768_),
    .A2(_1906_),
    .Y(_1907_),
    .B1(_1905_));
 sg13g2_o21ai_1 _4741_ (.B1(net962),
    .Y(_1908_),
    .A1(_1806_),
    .A2(_1904_));
 sg13g2_a21oi_1 _4742_ (.A1(_1808_),
    .A2(_1904_),
    .Y(_1909_),
    .B1(_1908_));
 sg13g2_o21ai_1 _4743_ (.B1(_1712_),
    .Y(_1910_),
    .A1(net143),
    .A2(net682));
 sg13g2_o21ai_1 _4744_ (.B1(net105),
    .Y(_0265_),
    .A1(net963),
    .A2(_1910_));
 sg13g2_nand3_1 _4745_ (.B(_1792_),
    .C(_1837_),
    .A(_0035_),
    .Y(_1911_));
 sg13g2_nor2_1 _4746_ (.A(_2051_),
    .B(_0034_),
    .Y(_1912_));
 sg13g2_a22oi_1 _4747_ (.Y(_1913_),
    .B1(_1911_),
    .B2(_1912_),
    .A2(_1901_),
    .A1(_1783_));
 sg13g2_o21ai_1 _4748_ (.B1(_1810_),
    .Y(_1914_),
    .A1(_0033_),
    .A2(_1771_));
 sg13g2_xor2_1 _4749_ (.B(net708),
    .A(net711),
    .X(_1915_));
 sg13g2_a221oi_1 _4750_ (.B2(_1768_),
    .C1(_1914_),
    .B1(_1915_),
    .A1(_1808_),
    .Y(_1916_),
    .A2(_1913_));
 sg13g2_o21ai_1 _4751_ (.B1(_1916_),
    .Y(_1917_),
    .A1(_1806_),
    .A2(_1913_));
 sg13g2_a21oi_1 _4752_ (.A1(_2059_),
    .A2(_0842_),
    .Y(_1918_),
    .B1(net654));
 sg13g2_a22oi_1 _4753_ (.Y(_1919_),
    .B1(_1917_),
    .B2(_1918_),
    .A2(net654),
    .A1(net125));
 sg13g2_inv_1 _4754_ (.Y(_0266_),
    .A(net126));
 sg13g2_nor2_1 _4755_ (.A(net914),
    .B(_1771_),
    .Y(_1920_));
 sg13g2_nand2_1 _4756_ (.Y(_1921_),
    .A(net58),
    .B(net654));
 sg13g2_nor4_1 _4757_ (.A(_0842_),
    .B(_1770_),
    .C(_1808_),
    .D(_1920_),
    .Y(_1922_));
 sg13g2_o21ai_1 _4758_ (.B1(_1712_),
    .Y(_1923_),
    .A1(net125),
    .A2(net682));
 sg13g2_o21ai_1 _4759_ (.B1(net59),
    .Y(_0267_),
    .A1(net915),
    .A2(_1923_));
 sg13g2_o21ai_1 _4760_ (.B1(net40),
    .Y(_1924_),
    .A1(\siggen.n22_o ),
    .A2(net682));
 sg13g2_inv_1 _4761_ (.Y(_0268_),
    .A(net41));
 sg13g2_o21ai_1 _4762_ (.B1(_0123_),
    .Y(_1925_),
    .A1(net256),
    .A2(net293));
 sg13g2_nor2_1 _4763_ (.A(_2010_),
    .B(_1925_),
    .Y(_1926_));
 sg13g2_o21ai_1 _4764_ (.B1(net265),
    .Y(_1927_),
    .A1(_2010_),
    .A2(_1925_));
 sg13g2_o21ai_1 _4765_ (.B1(_1927_),
    .Y(_0269_),
    .A1(net265),
    .A2(_1925_));
 sg13g2_o21ai_1 _4766_ (.B1(net148),
    .Y(_1928_),
    .A1(\siggen.dac_pmod.cnt_reg[0] ),
    .A2(_1925_));
 sg13g2_nor2_1 _4767_ (.A(_0841_),
    .B(_0844_),
    .Y(_1929_));
 sg13g2_o21ai_1 _4768_ (.B1(net149),
    .Y(_0270_),
    .A1(_1925_),
    .A2(_1929_));
 sg13g2_nor2_1 _4769_ (.A(net310),
    .B(_0845_),
    .Y(_1930_));
 sg13g2_nor2_1 _4770_ (.A(_0841_),
    .B(_1930_),
    .Y(_1931_));
 sg13g2_nor2_1 _4771_ (.A(_1925_),
    .B(_1931_),
    .Y(_1932_));
 sg13g2_o21ai_1 _4772_ (.B1(net310),
    .Y(_1933_),
    .A1(_0845_),
    .A2(_1925_));
 sg13g2_nand2b_1 _4773_ (.Y(_0271_),
    .B(net311),
    .A_N(_1932_));
 sg13g2_nand3_1 _4774_ (.B(_1926_),
    .C(_1930_),
    .A(net470),
    .Y(_1934_));
 sg13g2_o21ai_1 _4775_ (.B1(_1934_),
    .Y(_1935_),
    .A1(net470),
    .A2(_1932_));
 sg13g2_inv_1 _4776_ (.Y(_0272_),
    .A(net471));
 sg13g2_o21ai_1 _4777_ (.B1(_2010_),
    .Y(_1936_),
    .A1(\siggen.dac_pmod.n85_q[1] ),
    .A2(net40));
 sg13g2_nand3_1 _4778_ (.B(\siggen.da_cs ),
    .C(_1936_),
    .A(net256),
    .Y(_1937_));
 sg13g2_o21ai_1 _4779_ (.B1(net257),
    .Y(_0273_),
    .A1(net256),
    .A2(net293));
 sg13g2_a22oi_1 _4780_ (.Y(_1938_),
    .B1(_0646_),
    .B2(net1010),
    .A2(_0644_),
    .A1(net73));
 sg13g2_inv_1 _4781_ (.Y(_0274_),
    .A(net74));
 sg13g2_nand2_1 _4782_ (.Y(_1939_),
    .A(net55),
    .B(_0644_));
 sg13g2_xnor2_1 _4783_ (.Y(_1940_),
    .A(\settings_uart_printer.uart_tx_module.counter_reg[0] ),
    .B(net870));
 sg13g2_o21ai_1 _4784_ (.B1(net56),
    .Y(_0275_),
    .A1(_0645_),
    .A2(net871));
 sg13g2_o21ai_1 _4785_ (.B1(net688),
    .Y(_1941_),
    .A1(net901),
    .A2(_0637_));
 sg13g2_xnor2_1 _4786_ (.Y(_1942_),
    .A(net90),
    .B(_0629_));
 sg13g2_nor2_1 _4787_ (.A(_1941_),
    .B(net91),
    .Y(_0276_));
 sg13g2_nand2_1 _4788_ (.Y(_1943_),
    .A(net52),
    .B(_0644_));
 sg13g2_xor2_1 _4789_ (.B(_0630_),
    .A(net886),
    .X(_1944_));
 sg13g2_o21ai_1 _4790_ (.B1(net53),
    .Y(_0277_),
    .A1(_0645_),
    .A2(net887));
 sg13g2_xnor2_1 _4791_ (.Y(_1945_),
    .A(net181),
    .B(_0631_));
 sg13g2_nor2_1 _4792_ (.A(_1941_),
    .B(net182),
    .Y(_0278_));
 sg13g2_nand2_1 _4793_ (.Y(_1946_),
    .A(net37),
    .B(_0644_));
 sg13g2_xor2_1 _4794_ (.B(_0632_),
    .A(net882),
    .X(_1947_));
 sg13g2_o21ai_1 _4795_ (.B1(net38),
    .Y(_0279_),
    .A1(_0645_),
    .A2(net883));
 sg13g2_xnor2_1 _4796_ (.Y(_1948_),
    .A(net222),
    .B(_0633_));
 sg13g2_nor2_1 _4797_ (.A(_1941_),
    .B(net223),
    .Y(_0280_));
 sg13g2_nand2b_1 _4798_ (.Y(_1949_),
    .B(net151),
    .A_N(_0634_));
 sg13g2_a21oi_1 _4799_ (.A1(_0635_),
    .A2(net152),
    .Y(_0281_),
    .B1(_1941_));
 sg13g2_xor2_1 _4800_ (.B(_0635_),
    .A(net352),
    .X(_1950_));
 sg13g2_nor2_1 _4801_ (.A(_1941_),
    .B(net353),
    .Y(_0282_));
 sg13g2_nand2_1 _4802_ (.Y(_1951_),
    .A(net31),
    .B(_0644_));
 sg13g2_o21ai_1 _4803_ (.B1(net876),
    .Y(_1952_),
    .A1(net352),
    .A2(_0635_));
 sg13g2_nand2b_1 _4804_ (.Y(_1953_),
    .B(net877),
    .A_N(_0636_));
 sg13g2_o21ai_1 _4805_ (.B1(net32),
    .Y(_0283_),
    .A1(_0645_),
    .A2(_1953_));
 sg13g2_nand2b_1 _4806_ (.Y(_1954_),
    .B(net157),
    .A_N(_0636_));
 sg13g2_a21oi_1 _4807_ (.A1(_0637_),
    .A2(net158),
    .Y(_0284_),
    .B1(_1941_));
 sg13g2_a21oi_1 _4808_ (.A1(net901),
    .A2(_0637_),
    .Y(_1955_),
    .B1(_1941_));
 sg13g2_a21o_1 _4809_ (.A2(_0644_),
    .A1(net110),
    .B1(_1955_),
    .X(_0285_));
 sg13g2_nand2_1 _4810_ (.Y(_1956_),
    .A(net730),
    .B(net920));
 sg13g2_nand2_1 _4811_ (.Y(_1957_),
    .A(_1977_),
    .B(net492));
 sg13g2_o21ai_1 _4812_ (.B1(net493),
    .Y(_0286_),
    .A1(_1086_),
    .A2(_1956_));
 sg13g2_or2_1 _4813_ (.X(_1958_),
    .B(net729),
    .A(net884));
 sg13g2_a21oi_1 _4814_ (.A1(net437),
    .A2(_1958_),
    .Y(_1959_),
    .B1(net360));
 sg13g2_a21o_1 _4815_ (.A2(_1958_),
    .A1(net437),
    .B1(net360),
    .X(_1960_));
 sg13g2_nand2_1 _4816_ (.Y(_1961_),
    .A(net730),
    .B(_1960_));
 sg13g2_a21oi_1 _4817_ (.A1(net730),
    .A2(_1958_),
    .Y(_1962_),
    .B1(net437));
 sg13g2_a21oi_1 _4818_ (.A1(net730),
    .A2(_1960_),
    .Y(_0287_),
    .B1(net438));
 sg13g2_nor2_1 _4819_ (.A(net720),
    .B(_1088_),
    .Y(_1963_));
 sg13g2_mux2_1 _4820_ (.A0(_1963_),
    .A1(net720),
    .S(_1961_),
    .X(_0288_));
 sg13g2_nor2_1 _4821_ (.A(_1959_),
    .B(_1963_),
    .Y(_1964_));
 sg13g2_nor2_1 _4822_ (.A(net730),
    .B(net716),
    .Y(_1965_));
 sg13g2_xor2_1 _4823_ (.B(_1964_),
    .A(net597),
    .X(_1966_));
 sg13g2_a21oi_1 _4824_ (.A1(net730),
    .A2(net598),
    .Y(_0289_),
    .B1(_1965_));
 sg13g2_nor2_1 _4825_ (.A(net384),
    .B(net714),
    .Y(_1967_));
 sg13g2_nor3_1 _4826_ (.A(net597),
    .B(_1088_),
    .C(_1959_),
    .Y(_1968_));
 sg13g2_a22oi_1 _4827_ (.Y(_1969_),
    .B1(_1968_),
    .B2(net720),
    .A2(_1088_),
    .A1(net716));
 sg13g2_xnor2_1 _4828_ (.Y(_1970_),
    .A(net926),
    .B(_1969_));
 sg13g2_a21oi_1 _4829_ (.A1(net730),
    .A2(_1970_),
    .Y(_0290_),
    .B1(net385));
 sg13g2_nor3_2 _4830_ (.A(_1977_),
    .B(net693),
    .C(_1969_),
    .Y(_1971_));
 sg13g2_nand2_1 _4831_ (.Y(_1972_),
    .A(net711),
    .B(_1971_));
 sg13g2_xnor2_1 _4832_ (.Y(_0291_),
    .A(_2052_),
    .B(_1971_));
 sg13g2_xnor2_1 _4833_ (.Y(_0292_),
    .A(net267),
    .B(_1972_));
 sg13g2_nor2_1 _4834_ (.A(net319),
    .B(_1972_),
    .Y(_1973_));
 sg13g2_xnor2_1 _4835_ (.Y(_0293_),
    .A(_2056_),
    .B(net320));
 sg13g2_dfrbp_1 _4836_ (.CLK(clk),
    .RESET_B(net833),
    .D(net428),
    .Q_N(_2500_),
    .Q(\measurements.n98_o[1] ));
 sg13g2_dfrbp_1 _4837_ (.CLK(clk),
    .RESET_B(net831),
    .D(net499),
    .Q_N(_2499_),
    .Q(\measurements.n98_o[2] ));
 sg13g2_dfrbp_1 _4838_ (.CLK(clk),
    .RESET_B(net827),
    .D(net401),
    .Q_N(_2498_),
    .Q(\measurements.n98_o[3] ));
 sg13g2_dfrbp_1 _4839_ (.CLK(clk),
    .RESET_B(net817),
    .D(net307),
    .Q_N(_2497_),
    .Q(\measurements.n244_o[0] ));
 sg13g2_dfrbp_1 _4840_ (.CLK(clk),
    .RESET_B(net826),
    .D(net482),
    .Q_N(_2496_),
    .Q(\measurements.n244_o[1] ));
 sg13g2_dfrbp_1 _4841_ (.CLK(clk),
    .RESET_B(net826),
    .D(net359),
    .Q_N(_2495_),
    .Q(\measurements.n244_o[2] ));
 sg13g2_dfrbp_1 _4842_ (.CLK(clk),
    .RESET_B(net826),
    .D(net346),
    .Q_N(_2494_),
    .Q(\measurements.n244_o[3] ));
 sg13g2_dfrbp_1 _4843_ (.CLK(clk),
    .RESET_B(net809),
    .D(net424),
    .Q_N(_2493_),
    .Q(\settings_uart_printer.uart_tx_module.n88_q[0] ));
 sg13g2_dfrbp_1 _4844_ (.CLK(clk),
    .RESET_B(net807),
    .D(net485),
    .Q_N(_2492_),
    .Q(\settings_uart_printer.uart_tx_module.n88_q[1] ));
 sg13g2_dfrbp_1 _4845_ (.CLK(clk),
    .RESET_B(net804),
    .D(net201),
    .Q_N(_0004_),
    .Q(\settings_uart_printer.n103_q[0] ));
 sg13g2_dfrbp_1 _4846_ (.CLK(clk),
    .RESET_B(net804),
    .D(net596),
    .Q_N(_0003_),
    .Q(\settings_uart_printer.n103_q[1] ));
 sg13g2_dfrbp_1 _4847_ (.CLK(clk),
    .RESET_B(net804),
    .D(net848),
    .Q_N(_0006_),
    .Q(\settings_uart_printer.n103_q[2] ));
 sg13g2_dfrbp_1 _4848_ (.CLK(clk),
    .RESET_B(net803),
    .D(net857),
    .Q_N(_2491_),
    .Q(\settings_uart_printer.n103_q[3] ));
 sg13g2_dfrbp_1 _4849_ (.CLK(clk),
    .RESET_B(net804),
    .D(net142),
    .Q_N(\settings_uart_printer.n103_q[4] ),
    .Q(_0073_));
 sg13g2_dfrbp_1 _4850_ (.CLK(clk),
    .RESET_B(net804),
    .D(net180),
    .Q_N(\settings_uart_printer.n103_q[5] ),
    .Q(_0074_));
 sg13g2_dfrbp_1 _4851_ (.CLK(clk),
    .RESET_B(net808),
    .D(net63),
    .Q_N(\settings_uart_printer.uart_tx_module.datacnt_reg[0] ),
    .Q(_0075_));
 sg13g2_dfrbp_1 _4852_ (.CLK(clk),
    .RESET_B(net808),
    .D(net51),
    .Q_N(\settings_uart_printer.uart_tx_module.datacnt_reg[1] ),
    .Q(_0076_));
 sg13g2_dfrbp_1 _4853_ (.CLK(clk),
    .RESET_B(net808),
    .D(net113),
    .Q_N(\settings_uart_printer.uart_tx_module.datacnt_reg[2] ),
    .Q(_0077_));
 sg13g2_dfrbp_1 _4854_ (.CLK(clk),
    .RESET_B(net808),
    .D(net116),
    .Q_N(_2490_),
    .Q(\settings_uart_printer.uart_tx_module.data_reg[0] ));
 sg13g2_dfrbp_1 _4855_ (.CLK(clk),
    .RESET_B(net807),
    .D(net124),
    .Q_N(_2489_),
    .Q(\settings_uart_printer.uart_tx_module.data_reg[1] ));
 sg13g2_dfrbp_1 _4856_ (.CLK(clk),
    .RESET_B(net807),
    .D(net196),
    .Q_N(_2488_),
    .Q(\settings_uart_printer.uart_tx_module.data_reg[2] ));
 sg13g2_dfrbp_1 _4857_ (.CLK(clk),
    .RESET_B(net808),
    .D(net86),
    .Q_N(_2487_),
    .Q(\settings_uart_printer.uart_tx_module.data_reg[3] ));
 sg13g2_dfrbp_1 _4858_ (.CLK(clk),
    .RESET_B(net807),
    .D(net69),
    .Q_N(_2486_),
    .Q(\settings_uart_printer.uart_tx_module.data_reg[4] ));
 sg13g2_dfrbp_1 _4859_ (.CLK(clk),
    .RESET_B(net807),
    .D(net66),
    .Q_N(_2485_),
    .Q(\settings_uart_printer.uart_tx_module.data_reg[5] ));
 sg13g2_dfrbp_1 _4860_ (.CLK(clk),
    .RESET_B(net807),
    .D(net72),
    .Q_N(_2484_),
    .Q(\settings_uart_printer.uart_tx_module.data_reg[6] ));
 sg13g2_dfrbp_1 _4861_ (.CLK(clk),
    .RESET_B(net838),
    .D(net169),
    .Q_N(\oscilloscope_control.switch_debouncer_n2_debounce_switches.counter_next[0] ),
    .Q(\oscilloscope_control.switch_debouncer_n2_debounce_switches.counter_reg[0] ));
 sg13g2_dfrbp_1 _4862_ (.CLK(clk),
    .RESET_B(net836),
    .D(net185),
    .Q_N(_2483_),
    .Q(\oscilloscope_control.switch_debouncer_n2_debounce_switches.counter_reg[1] ));
 sg13g2_dfrbp_1 _4863_ (.CLK(clk),
    .RESET_B(net836),
    .D(net252),
    .Q_N(_2482_),
    .Q(\oscilloscope_control.switch_debouncer_n2_debounce_switches.counter_reg[2] ));
 sg13g2_dfrbp_1 _4864_ (.CLK(clk),
    .RESET_B(net807),
    .D(_0121_),
    .Q_N(_2481_),
    .Q(\settings_uart_printer.n104_q[0] ));
 sg13g2_dfrbp_1 _4865_ (.CLK(clk),
    .RESET_B(net804),
    .D(net502),
    .Q_N(_2501_),
    .Q(\settings_uart_printer.n104_q[1] ));
 sg13g2_dfrbp_1 _4866_ (.CLK(clk),
    .RESET_B(net824),
    .D(net561),
    .Q_N(_0049_),
    .Q(\videogen.draw_y[0] ));
 sg13g2_dfrbp_1 _4867_ (.CLK(clk),
    .RESET_B(net822),
    .D(net631),
    .Q_N(_0047_),
    .Q(\videogen.draw_y[1] ));
 sg13g2_dfrbp_1 _4868_ (.CLK(clk),
    .RESET_B(net822),
    .D(net339),
    .Q_N(_0021_),
    .Q(\videogen.draw_y[2] ));
 sg13g2_dfrbp_1 _4869_ (.CLK(clk),
    .RESET_B(net820),
    .D(net398),
    .Q_N(_2502_),
    .Q(\videogen.draw_y[3] ));
 sg13g2_dfrbp_1 _4870_ (.CLK(clk),
    .RESET_B(net820),
    .D(net615),
    .Q_N(_0048_),
    .Q(\videogen.draw_y[4] ));
 sg13g2_dfrbp_1 _4871_ (.CLK(clk),
    .RESET_B(net819),
    .D(net496),
    .Q_N(_0022_),
    .Q(\videogen.draw_y[5] ));
 sg13g2_dfrbp_1 _4872_ (.CLK(clk),
    .RESET_B(net820),
    .D(net466),
    .Q_N(_0023_),
    .Q(\videogen.draw_y[6] ));
 sg13g2_dfrbp_1 _4873_ (.CLK(clk),
    .RESET_B(net819),
    .D(net575),
    .Q_N(_0024_),
    .Q(\videogen.draw_y[7] ));
 sg13g2_dfrbp_1 _4874_ (.CLK(clk),
    .RESET_B(net819),
    .D(net27),
    .Q_N(_0025_),
    .Q(\videogen.draw_y[8] ));
 sg13g2_dfrbp_1 _4875_ (.CLK(clk),
    .RESET_B(net820),
    .D(net539),
    .Q_N(_0026_),
    .Q(\videogen.draw_y[9] ));
 sg13g2_dfrbp_1 _4876_ (.CLK(clk),
    .RESET_B(net823),
    .D(net572),
    .Q_N(_2480_),
    .Q(\siggen.dac_pmod.n85_q[0] ));
 sg13g2_dfrbp_1 _4877_ (.CLK(clk),
    .RESET_B(net823),
    .D(net294),
    .Q_N(_2479_),
    .Q(\siggen.dac_pmod.n85_q[1] ));
 sg13g2_dfrbp_1 _4878_ (.CLK(clk),
    .RESET_B(net835),
    .D(net336),
    .Q_N(\measurements.samples_storage.n101_o ),
    .Q(_0078_));
 sg13g2_dfrbp_1 _4879_ (.CLK(clk),
    .RESET_B(net827),
    .D(net227),
    .Q_N(_2478_),
    .Q(\measurements.samples_storage.n170_o ));
 sg13g2_dfrbp_1 _4880_ (.CLK(clk),
    .RESET_B(net836),
    .D(net230),
    .Q_N(_2477_),
    .Q(\oscilloscope_control.switch_debouncer_n2_debounce_switches.debounced ));
 sg13g2_dfrbp_1 _4881_ (.CLK(clk),
    .RESET_B(net837),
    .D(net83),
    .Q_N(\oscilloscope_control.switch_debouncer_n1_debounce_switches.counter_next[0] ),
    .Q(\oscilloscope_control.switch_debouncer_n1_debounce_switches.counter_reg[0] ));
 sg13g2_dfrbp_1 _4882_ (.CLK(clk),
    .RESET_B(net837),
    .D(net356),
    .Q_N(_2476_),
    .Q(\oscilloscope_control.switch_debouncer_n1_debounce_switches.counter_reg[1] ));
 sg13g2_dfrbp_1 _4883_ (.CLK(clk),
    .RESET_B(net837),
    .D(net191),
    .Q_N(_2475_),
    .Q(\oscilloscope_control.switch_debouncer_n1_debounce_switches.counter_reg[2] ));
 sg13g2_dfrbp_1 _4884_ (.CLK(clk),
    .RESET_B(net835),
    .D(net490),
    .Q_N(_2474_),
    .Q(\oscilloscope_control.switch_debouncer_n1_debounce_switches.debounced ));
 sg13g2_dfrbp_1 _4885_ (.CLK(clk),
    .RESET_B(net837),
    .D(net189),
    .Q_N(\oscilloscope_control.button_debouncer_n4_debounce_buttons.counter_next[0] ),
    .Q(\oscilloscope_control.button_debouncer_n4_debounce_buttons.counter_reg[0] ));
 sg13g2_dfrbp_1 _4886_ (.CLK(clk),
    .RESET_B(net837),
    .D(net301),
    .Q_N(_2473_),
    .Q(\oscilloscope_control.button_debouncer_n4_debounce_buttons.counter_reg[1] ));
 sg13g2_dfrbp_1 _4887_ (.CLK(clk),
    .RESET_B(net837),
    .D(net248),
    .Q_N(_2472_),
    .Q(\oscilloscope_control.button_debouncer_n4_debounce_buttons.counter_reg[2] ));
 sg13g2_dfrbp_1 _4888_ (.CLK(clk),
    .RESET_B(net835),
    .D(net165),
    .Q_N(_2471_),
    .Q(\oscilloscope_control.button_debouncer_n4_debounce_buttons.debounced ));
 sg13g2_dfrbp_1 _4889_ (.CLK(clk),
    .RESET_B(net816),
    .D(net94),
    .Q_N(\oscilloscope_control.button_debouncer_n3_debounce_buttons.counter_next[0] ),
    .Q(\oscilloscope_control.button_debouncer_n3_debounce_buttons.counter_reg[0] ));
 sg13g2_dfrbp_1 _4890_ (.CLK(clk),
    .RESET_B(net815),
    .D(net279),
    .Q_N(_2470_),
    .Q(\oscilloscope_control.button_debouncer_n3_debounce_buttons.counter_reg[1] ));
 sg13g2_dfrbp_1 _4891_ (.CLK(clk),
    .RESET_B(net815),
    .D(net232),
    .Q_N(_2469_),
    .Q(\oscilloscope_control.button_debouncer_n3_debounce_buttons.counter_reg[2] ));
 sg13g2_dfrbp_1 _4892_ (.CLK(clk),
    .RESET_B(net816),
    .D(net172),
    .Q_N(_2468_),
    .Q(\oscilloscope_control.button_debouncer_n3_debounce_buttons.debounced ));
 sg13g2_dfrbp_1 _4893_ (.CLK(clk),
    .RESET_B(net839),
    .D(net167),
    .Q_N(\oscilloscope_control.button_debouncer_n2_debounce_buttons.counter_next[0] ),
    .Q(\oscilloscope_control.button_debouncer_n2_debounce_buttons.counter_reg[0] ));
 sg13g2_dfrbp_1 _4894_ (.CLK(clk),
    .RESET_B(net839),
    .D(net284),
    .Q_N(_2467_),
    .Q(\oscilloscope_control.button_debouncer_n2_debounce_buttons.counter_reg[1] ));
 sg13g2_dfrbp_1 _4895_ (.CLK(clk),
    .RESET_B(net835),
    .D(net351),
    .Q_N(_2466_),
    .Q(\oscilloscope_control.button_debouncer_n2_debounce_buttons.counter_reg[2] ));
 sg13g2_dfrbp_1 _4896_ (.CLK(clk),
    .RESET_B(net839),
    .D(net206),
    .Q_N(_2465_),
    .Q(\oscilloscope_control.button_debouncer_n2_debounce_buttons.debounced ));
 sg13g2_dfrbp_1 _4897_ (.CLK(clk),
    .RESET_B(net829),
    .D(net203),
    .Q_N(\oscilloscope_control.button_debouncer_n1_debounce_buttons.counter_next[0] ),
    .Q(\oscilloscope_control.button_debouncer_n1_debounce_buttons.counter_reg[0] ));
 sg13g2_dfrbp_1 _4898_ (.CLK(clk),
    .RESET_B(net829),
    .D(net296),
    .Q_N(_2464_),
    .Q(\oscilloscope_control.button_debouncer_n1_debounce_buttons.counter_reg[1] ));
 sg13g2_dfrbp_1 _4899_ (.CLK(clk),
    .RESET_B(net829),
    .D(net369),
    .Q_N(_2463_),
    .Q(\oscilloscope_control.button_debouncer_n1_debounce_buttons.counter_reg[2] ));
 sg13g2_dfrbp_1 _4900_ (.CLK(clk),
    .RESET_B(net829),
    .D(net271),
    .Q_N(_2462_),
    .Q(\oscilloscope_control.button_debouncer_n1_debounce_buttons.debounced ));
 sg13g2_dfrbp_1 _4901_ (.CLK(clk),
    .RESET_B(net824),
    .D(net602),
    .Q_N(\oscilloscope_control.n114_o[0] ),
    .Q(\champlitude[0] ));
 sg13g2_dfrbp_1 _4902_ (.CLK(clk),
    .RESET_B(net824),
    .D(net851),
    .Q_N(_0009_),
    .Q(\champlitude[1] ));
 sg13g2_dfrbp_1 _4903_ (.CLK(clk),
    .RESET_B(net824),
    .D(net844),
    .Q_N(_0042_),
    .Q(\champlitude[2] ));
 sg13g2_dfrbp_1 _4904_ (.CLK(clk),
    .RESET_B(net810),
    .D(net332),
    .Q_N(\oscilloscope_control.n146_o[0] ),
    .Q(\measurements.n200_o[0] ));
 sg13g2_dfrbp_1 _4905_ (.CLK(clk),
    .RESET_B(net810),
    .D(net511),
    .Q_N(_0008_),
    .Q(\measurements.n200_o[1] ));
 sg13g2_dfrbp_1 _4906_ (.CLK(clk),
    .RESET_B(net810),
    .D(net587),
    .Q_N(_0002_),
    .Q(\measurements.n200_o[2] ));
 sg13g2_dfrbp_1 _4907_ (.CLK(clk),
    .RESET_B(net808),
    .D(net559),
    .Q_N(_2461_),
    .Q(\oscilloscope_control.n220_q[0] ));
 sg13g2_dfrbp_1 _4908_ (.CLK(clk),
    .RESET_B(net808),
    .D(net517),
    .Q_N(_2460_),
    .Q(\oscilloscope_control.n220_q[1] ));
 sg13g2_dfrbp_1 _4909_ (.CLK(clk),
    .RESET_B(net810),
    .D(net147),
    .Q_N(\measurements.trigger.sample_on_rising_edge ),
    .Q(_0079_));
 sg13g2_dfrbp_1 _4910_ (.CLK(clk),
    .RESET_B(net831),
    .D(net505),
    .Q_N(_2459_),
    .Q(\measurements.samples_storage.spi_master_inst.n100_q[0] ));
 sg13g2_dfrbp_1 _4911_ (.CLK(clk),
    .RESET_B(net835),
    .D(net554),
    .Q_N(_2458_),
    .Q(\measurements.samples_storage.spi_master_inst.n100_q[1] ));
 sg13g2_dfrbp_1 _4912_ (.CLK(clk),
    .RESET_B(net810),
    .D(net36),
    .Q_N(\measurements.trigger.trigger_threshold[0] ),
    .Q(_0080_));
 sg13g2_dfrbp_1 _4913_ (.CLK(clk),
    .RESET_B(net817),
    .D(net30),
    .Q_N(\measurements.trigger.trigger_threshold[1] ),
    .Q(_0081_));
 sg13g2_dfrbp_1 _4914_ (.CLK(clk),
    .RESET_B(net810),
    .D(net412),
    .Q_N(_0010_),
    .Q(\measurements.trigger.trigger_threshold[2] ));
 sg13g2_dfrbp_1 _4915_ (.CLK(clk),
    .RESET_B(net811),
    .D(net536),
    .Q_N(_0011_),
    .Q(\measurements.trigger.trigger_threshold[3] ));
 sg13g2_dfrbp_1 _4916_ (.CLK(clk),
    .RESET_B(net838),
    .D(net2),
    .Q_N(_2503_),
    .Q(\oscilloscope_control.button_ff_stage_1_reg[0] ));
 sg13g2_dfrbp_1 _4917_ (.CLK(clk),
    .RESET_B(net836),
    .D(net6),
    .Q_N(_2504_),
    .Q(\oscilloscope_control.button_ff_stage_1_reg[1] ));
 sg13g2_dfrbp_1 _4918_ (.CLK(clk),
    .RESET_B(net837),
    .D(net3),
    .Q_N(_2505_),
    .Q(\oscilloscope_control.button_ff_stage_1_reg[2] ));
 sg13g2_dfrbp_1 _4919_ (.CLK(clk),
    .RESET_B(net836),
    .D(net7),
    .Q_N(_2457_),
    .Q(\oscilloscope_control.button_ff_stage_1_reg[3] ));
 sg13g2_dfrbp_1 _4920_ (.CLK(clk),
    .RESET_B(net813),
    .D(net566),
    .Q_N(_2456_),
    .Q(\measurements.memoryShift[0] ));
 sg13g2_dfrbp_1 _4921_ (.CLK(clk),
    .RESET_B(net813),
    .D(net568),
    .Q_N(_2455_),
    .Q(\measurements.memoryShift[1] ));
 sg13g2_dfrbp_1 _4922_ (.CLK(clk),
    .RESET_B(net813),
    .D(net455),
    .Q_N(_0027_),
    .Q(\measurements.memoryShift[2] ));
 sg13g2_dfrbp_1 _4923_ (.CLK(clk),
    .RESET_B(net813),
    .D(net404),
    .Q_N(_2454_),
    .Q(\measurements.memoryShift[3] ));
 sg13g2_dfrbp_1 _4924_ (.CLK(clk),
    .RESET_B(net814),
    .D(net487),
    .Q_N(_0028_),
    .Q(\measurements.memoryShift[4] ));
 sg13g2_dfrbp_1 _4925_ (.CLK(clk),
    .RESET_B(net814),
    .D(net420),
    .Q_N(_2453_),
    .Q(\measurements.memoryShift[5] ));
 sg13g2_dfrbp_1 _4926_ (.CLK(clk),
    .RESET_B(net816),
    .D(net441),
    .Q_N(_0029_),
    .Q(\measurements.memoryShift[6] ));
 sg13g2_dfrbp_1 _4927_ (.CLK(clk),
    .RESET_B(net816),
    .D(net464),
    .Q_N(_0031_),
    .Q(\measurements.memoryShift[7] ));
 sg13g2_dfrbp_1 _4928_ (.CLK(clk),
    .RESET_B(net816),
    .D(net344),
    .Q_N(_0030_),
    .Q(\measurements.memoryShift[8] ));
 sg13g2_dfrbp_1 _4929_ (.CLK(clk),
    .RESET_B(net829),
    .D(net869),
    .Q_N(_0071_),
    .Q(\oscilloscope_control.button_debouncer_n1_debounce_buttons.in_raw ));
 sg13g2_dfrbp_1 _4930_ (.CLK(clk),
    .RESET_B(net835),
    .D(net861),
    .Q_N(_0069_),
    .Q(\oscilloscope_control.button_debouncer_n2_debounce_buttons.in_raw ));
 sg13g2_dfrbp_1 _4931_ (.CLK(clk),
    .RESET_B(net830),
    .D(net867),
    .Q_N(_2506_),
    .Q(\oscilloscope_control.button_debouncer_n3_debounce_buttons.in_raw ));
 sg13g2_dfrbp_1 _4932_ (.CLK(clk),
    .RESET_B(net837),
    .D(net865),
    .Q_N(_0072_),
    .Q(\oscilloscope_control.button_debouncer_n4_debounce_buttons.in_raw ));
 sg13g2_dfrbp_1 _4933_ (.CLK(clk),
    .RESET_B(net803),
    .D(net48),
    .Q_N(_0005_),
    .Q(\measurements.n163_o[0] ));
 sg13g2_dfrbp_1 _4934_ (.CLK(clk),
    .RESET_B(net805),
    .D(net551),
    .Q_N(_2452_),
    .Q(\measurements.n163_o[1] ));
 sg13g2_dfrbp_1 _4935_ (.CLK(clk),
    .RESET_B(net803),
    .D(net45),
    .Q_N(\measurements.n163_o[2] ),
    .Q(_0082_));
 sg13g2_dfrbp_1 _4936_ (.CLK(clk),
    .RESET_B(net836),
    .D(net4),
    .Q_N(_2507_),
    .Q(\oscilloscope_control.n223_q[0] ));
 sg13g2_dfrbp_1 _4937_ (.CLK(clk),
    .RESET_B(net836),
    .D(net8),
    .Q_N(_2451_),
    .Q(\oscilloscope_control.n223_q[1] ));
 sg13g2_dfrbp_1 _4938_ (.CLK(clk),
    .RESET_B(net809),
    .D(net177),
    .Q_N(\oscilloscope_control.n171_o[0] ),
    .Q(\dsgfreqshift[0] ));
 sg13g2_dfrbp_1 _4939_ (.CLK(clk),
    .RESET_B(net808),
    .D(net361),
    .Q_N(_2508_),
    .Q(\dsgfreqshift[1] ));
 sg13g2_dfrbp_1 _4940_ (.CLK(clk),
    .RESET_B(net838),
    .D(net859),
    .Q_N(_0001_),
    .Q(\oscilloscope_control.n206_o ));
 sg13g2_dfrbp_1 _4941_ (.CLK(clk),
    .RESET_B(net836),
    .D(net863),
    .Q_N(_0070_),
    .Q(\oscilloscope_control.n208_o ));
 sg13g2_dfrbp_1 _4942_ (.CLK(clk),
    .RESET_B(net810),
    .D(net557),
    .Q_N(\oscilloscope_control.n111_o[0] ),
    .Q(\choffset[0] ));
 sg13g2_dfrbp_1 _4943_ (.CLK(clk),
    .RESET_B(net810),
    .D(net584),
    .Q_N(_0007_),
    .Q(\choffset[1] ));
 sg13g2_dfrbp_1 _4944_ (.CLK(clk),
    .RESET_B(net809),
    .D(net97),
    .Q_N(\choffset[2] ),
    .Q(_0083_));
 sg13g2_dfrbp_1 _4945_ (.CLK(clk),
    .RESET_B(net811),
    .D(net593),
    .Q_N(_0041_),
    .Q(\choffset[3] ));
 sg13g2_dfrbp_1 _4946_ (.CLK(clk),
    .RESET_B(net811),
    .D(net547),
    .Q_N(_0043_),
    .Q(\choffset[4] ));
 sg13g2_dfrbp_1 _4947_ (.CLK(clk),
    .RESET_B(net832),
    .D(net342),
    .Q_N(_2450_),
    .Q(\measurements.samples_storage.spi_master_inst.n96_o ));
 sg13g2_dfrbp_1 _4948_ (.CLK(clk),
    .RESET_B(net805),
    .D(net628),
    .Q_N(_2449_),
    .Q(\display_x[0] ));
 sg13g2_dfrbp_1 _4949_ (.CLK(clk),
    .RESET_B(net805),
    .D(net406),
    .Q_N(_2448_),
    .Q(\display_x[1] ));
 sg13g2_dfrbp_1 _4950_ (.CLK(clk),
    .RESET_B(net805),
    .D(net445),
    .Q_N(_0014_),
    .Q(\display_x[2] ));
 sg13g2_dfrbp_1 _4951_ (.CLK(clk),
    .RESET_B(net805),
    .D(net409),
    .Q_N(_0015_),
    .Q(\display_x[3] ));
 sg13g2_dfrbp_1 _4952_ (.CLK(clk),
    .RESET_B(net805),
    .D(net520),
    .Q_N(_0016_),
    .Q(\display_x[4] ));
 sg13g2_dfrbp_1 _4953_ (.CLK(clk),
    .RESET_B(net805),
    .D(net524),
    .Q_N(_0017_),
    .Q(\display_x[5] ));
 sg13g2_dfrbp_1 _4954_ (.CLK(clk),
    .RESET_B(net806),
    .D(net277),
    .Q_N(_0018_),
    .Q(\display_x[6] ));
 sg13g2_dfrbp_1 _4955_ (.CLK(clk),
    .RESET_B(net806),
    .D(net261),
    .Q_N(_0019_),
    .Q(\display_x[7] ));
 sg13g2_dfrbp_1 _4956_ (.CLK(clk),
    .RESET_B(net806),
    .D(net383),
    .Q_N(_0020_),
    .Q(\display_x[8] ));
 sg13g2_dfrbp_1 _4957_ (.CLK(clk),
    .RESET_B(net805),
    .D(net543),
    .Q_N(_0055_),
    .Q(\display_x[9] ));
 sg13g2_dfrbp_1 _4958_ (.CLK(clk),
    .RESET_B(net832),
    .D(net324),
    .Q_N(_2447_),
    .Q(\measurements.n98_o[0] ));
 sg13g2_dfrbp_1 _4959_ (.CLK(clk),
    .RESET_B(net812),
    .D(net514),
    .Q_N(_2446_),
    .Q(\measurements.n246_q[0] ));
 sg13g2_dfrbp_1 _4960_ (.CLK(clk),
    .RESET_B(net812),
    .D(_0193_),
    .Q_N(_2445_),
    .Q(\measurements.n246_q[1] ));
 sg13g2_dfrbp_1 _4961_ (.CLK(clk),
    .RESET_B(net812),
    .D(net372),
    .Q_N(_2444_),
    .Q(\measurements.n246_q[2] ));
 sg13g2_dfrbp_1 _4962_ (.CLK(clk),
    .RESET_B(net812),
    .D(net367),
    .Q_N(_2443_),
    .Q(\measurements.n246_q[3] ));
 sg13g2_dfrbp_1 _4963_ (.CLK(clk),
    .RESET_B(net813),
    .D(net237),
    .Q_N(_2442_),
    .Q(\measurements.n246_q[4] ));
 sg13g2_dfrbp_1 _4964_ (.CLK(clk),
    .RESET_B(net813),
    .D(net156),
    .Q_N(_2441_),
    .Q(\measurements.n246_q[5] ));
 sg13g2_dfrbp_1 _4965_ (.CLK(clk),
    .RESET_B(net814),
    .D(net396),
    .Q_N(_2440_),
    .Q(\measurements.n246_q[6] ));
 sg13g2_dfrbp_1 _4966_ (.CLK(clk),
    .RESET_B(net814),
    .D(net327),
    .Q_N(_2439_),
    .Q(\measurements.n246_q[7] ));
 sg13g2_dfrbp_1 _4967_ (.CLK(clk),
    .RESET_B(net814),
    .D(net209),
    .Q_N(_2438_),
    .Q(\measurements.n246_q[8] ));
 sg13g2_dfrbp_1 _4968_ (.CLK(clk),
    .RESET_B(net814),
    .D(net221),
    .Q_N(_2437_),
    .Q(\measurements.n246_q[9] ));
 sg13g2_dfrbp_1 _4969_ (.CLK(clk),
    .RESET_B(net816),
    .D(net215),
    .Q_N(_2436_),
    .Q(\measurements.n246_q[10] ));
 sg13g2_dfrbp_1 _4970_ (.CLK(clk),
    .RESET_B(net815),
    .D(net103),
    .Q_N(_2435_),
    .Q(\measurements.n246_q[11] ));
 sg13g2_dfrbp_1 _4971_ (.CLK(clk),
    .RESET_B(net815),
    .D(_0204_),
    .Q_N(_2434_),
    .Q(\measurements.n246_q[12] ));
 sg13g2_dfrbp_1 _4972_ (.CLK(clk),
    .RESET_B(net815),
    .D(_0205_),
    .Q_N(_2433_),
    .Q(\measurements.n246_q[13] ));
 sg13g2_dfrbp_1 _4973_ (.CLK(clk),
    .RESET_B(net815),
    .D(net255),
    .Q_N(_2432_),
    .Q(\measurements.n246_q[14] ));
 sg13g2_dfrbp_1 _4974_ (.CLK(clk),
    .RESET_B(net832),
    .D(net234),
    .Q_N(_2431_),
    .Q(\measurements.samples_adc.cnt_reg[0] ));
 sg13g2_dfrbp_1 _4975_ (.CLK(clk),
    .RESET_B(net832),
    .D(net109),
    .Q_N(_2430_),
    .Q(\measurements.samples_adc.cnt_reg[1] ));
 sg13g2_dfrbp_1 _4976_ (.CLK(clk),
    .RESET_B(net832),
    .D(net426),
    .Q_N(_2429_),
    .Q(\measurements.samples_adc.cnt_reg[2] ));
 sg13g2_dfrbp_1 _4977_ (.CLK(clk),
    .RESET_B(net832),
    .D(net264),
    .Q_N(_2428_),
    .Q(\measurements.samples_adc.cnt_reg[3] ));
 sg13g2_dfrbp_1 _4978_ (.CLK(clk),
    .RESET_B(net823),
    .D(net81),
    .Q_N(\measurements.adc_sclk ),
    .Q(_0084_));
 sg13g2_dfrbp_1 _4979_ (.CLK(clk),
    .RESET_B(net835),
    .D(net187),
    .Q_N(_2427_),
    .Q(\measurements.samples_storage.n232_q ));
 sg13g2_dfrbp_1 _4980_ (.CLK(clk),
    .RESET_B(net832),
    .D(net564),
    .Q_N(_2426_),
    .Q(\measurements.samples_adc.n84_q[0] ));
 sg13g2_dfrbp_1 _4981_ (.CLK(clk),
    .RESET_B(net832),
    .D(net198),
    .Q_N(_2425_),
    .Q(\measurements.samples_adc.n84_q[1] ));
 sg13g2_dfrbp_1 _4982_ (.CLK(clk),
    .RESET_B(net824),
    .D(net619),
    .Q_N(_0050_),
    .Q(\measurements.fram_mosi ));
 sg13g2_dfrbp_1 _4983_ (.CLK(clk),
    .RESET_B(net827),
    .D(net527),
    .Q_N(_0051_),
    .Q(\measurements.samples_storage.spi_master_inst.n30_o ));
 sg13g2_dfrbp_1 _4984_ (.CLK(clk),
    .RESET_B(net827),
    .D(net530),
    .Q_N(_0052_),
    .Q(\measurements.samples_storage.spi_master_inst.n28_o ));
 sg13g2_dfrbp_1 _4985_ (.CLK(clk),
    .RESET_B(net827),
    .D(net458),
    .Q_N(_2424_),
    .Q(\measurements.samples_storage.spi_master_inst.n26_o ));
 sg13g2_dfrbp_1 _4986_ (.CLK(clk),
    .RESET_B(net827),
    .D(net318),
    .Q_N(_2423_),
    .Q(\measurements.samples_storage.spi_master_inst.n24_o ));
 sg13g2_dfrbp_1 _4987_ (.CLK(clk),
    .RESET_B(net831),
    .D(net377),
    .Q_N(_2422_),
    .Q(\measurements.samples_storage.spi_master_inst.n22_o ));
 sg13g2_dfrbp_1 _4988_ (.CLK(clk),
    .RESET_B(net831),
    .D(net469),
    .Q_N(_2421_),
    .Q(\measurements.samples_storage.spi_master_inst.n20_o ));
 sg13g2_dfrbp_1 _4989_ (.CLK(clk),
    .RESET_B(net834),
    .D(net246),
    .Q_N(_2420_),
    .Q(\measurements.samples_storage.spi_master_inst.n18_o ));
 sg13g2_dfrbp_1 _4990_ (.CLK(clk),
    .RESET_B(net830),
    .D(net549),
    .Q_N(_2419_),
    .Q(\measurements.samples_storage.n230_q[0] ));
 sg13g2_dfrbp_1 _4991_ (.CLK(clk),
    .RESET_B(net829),
    .D(net607),
    .Q_N(_2418_),
    .Q(\measurements.samples_storage.n230_q[1] ));
 sg13g2_dfrbp_1 _4992_ (.CLK(clk),
    .RESET_B(net829),
    .D(net612),
    .Q_N(_2417_),
    .Q(\measurements.samples_storage.n230_q[2] ));
 sg13g2_dfrbp_1 _4993_ (.CLK(clk),
    .RESET_B(net829),
    .D(net590),
    .Q_N(_2416_),
    .Q(\measurements.samples_storage.n230_q[3] ));
 sg13g2_dfrbp_1 _4994_ (.CLK(clk),
    .RESET_B(net833),
    .D(net508),
    .Q_N(_2415_),
    .Q(\measurements.fram_sclk ));
 sg13g2_dfrbp_1 _4995_ (.CLK(clk),
    .RESET_B(net833),
    .D(net240),
    .Q_N(_2414_),
    .Q(\measurements.samples_storage.spi_master_inst.n103_q[1] ));
 sg13g2_dfrbp_1 _4996_ (.CLK(clk),
    .RESET_B(net833),
    .D(net162),
    .Q_N(_2413_),
    .Q(\measurements.samples_storage.spi_master_inst.n103_q[2] ));
 sg13g2_dfrbp_1 _4997_ (.CLK(clk),
    .RESET_B(net835),
    .D(net212),
    .Q_N(_2412_),
    .Q(\measurements.samples_storage.spi_master_inst.n103_q[3] ));
 sg13g2_dfrbp_1 _4998_ (.CLK(clk),
    .RESET_B(net828),
    .D(net622),
    .Q_N(_2411_),
    .Q(\measurements.n250_q[0] ));
 sg13g2_dfrbp_1 _4999_ (.CLK(clk),
    .RESET_B(net828),
    .D(net578),
    .Q_N(_2410_),
    .Q(\measurements.n250_q[1] ));
 sg13g2_dfrbp_1 _5000_ (.CLK(clk),
    .RESET_B(net828),
    .D(net581),
    .Q_N(_2409_),
    .Q(\measurements.n250_q[2] ));
 sg13g2_dfrbp_1 _5001_ (.CLK(clk),
    .RESET_B(net828),
    .D(net118),
    .Q_N(_2408_),
    .Q(\measurements.n250_q[3] ));
 sg13g2_dfrbp_1 _5002_ (.CLK(clk),
    .RESET_B(net817),
    .D(net136),
    .Q_N(_2509_),
    .Q(\measurements.enough_samples_in_fram_reg ));
 sg13g2_dfrbp_1 _5003_ (.CLK(clk),
    .RESET_B(net828),
    .D(net25),
    .Q_N(_0013_),
    .Q(\measurements.n249_q[0] ));
 sg13g2_dfrbp_1 _5004_ (.CLK(clk),
    .RESET_B(net830),
    .D(net243),
    .Q_N(_2510_),
    .Q(\measurements.n249_q[1] ));
 sg13g2_dfrbp_1 _5005_ (.CLK(clk),
    .RESET_B(net830),
    .D(net133),
    .Q_N(_2511_),
    .Q(\measurements.n249_q[2] ));
 sg13g2_dfrbp_1 _5006_ (.CLK(clk),
    .RESET_B(net828),
    .D(net218),
    .Q_N(_2512_),
    .Q(\measurements.n249_q[3] ));
 sg13g2_dfrbp_1 _5007_ (.CLK(clk),
    .RESET_B(net828),
    .D(net282),
    .Q_N(_2513_),
    .Q(\measurements.n249_q[4] ));
 sg13g2_dfrbp_1 _5008_ (.CLK(clk),
    .RESET_B(net828),
    .D(net274),
    .Q_N(_2407_),
    .Q(\measurements.n249_q[5] ));
 sg13g2_dfrbp_1 _5009_ (.CLK(clk),
    .RESET_B(net831),
    .D(net121),
    .Q_N(_2406_),
    .Q(\lastsample[0] ));
 sg13g2_dfrbp_1 _5010_ (.CLK(clk),
    .RESET_B(net831),
    .D(net175),
    .Q_N(_2405_),
    .Q(\lastsample[1] ));
 sg13g2_dfrbp_1 _5011_ (.CLK(clk),
    .RESET_B(net831),
    .D(net194),
    .Q_N(_2404_),
    .Q(\lastsample[2] ));
 sg13g2_dfrbp_1 _5012_ (.CLK(clk),
    .RESET_B(net831),
    .D(net389),
    .Q_N(_2403_),
    .Q(\lastsample[3] ));
 sg13g2_dfrbp_1 _5013_ (.CLK(clk),
    .RESET_B(net826),
    .D(net431),
    .Q_N(_2402_),
    .Q(\lastsample[4] ));
 sg13g2_dfrbp_1 _5014_ (.CLK(clk),
    .RESET_B(net826),
    .D(net330),
    .Q_N(_0046_),
    .Q(\lastsample[5] ));
 sg13g2_dfrbp_1 _5015_ (.CLK(clk),
    .RESET_B(net826),
    .D(net380),
    .Q_N(_0045_),
    .Q(\lastsample[6] ));
 sg13g2_dfrbp_1 _5016_ (.CLK(clk),
    .RESET_B(net825),
    .D(net448),
    .Q_N(_0044_),
    .Q(\lastsample[7] ));
 sg13g2_dfrbp_1 _5017_ (.CLK(clk),
    .RESET_B(net826),
    .D(net414),
    .Q_N(_0054_),
    .Q(\measurements.n253_q ));
 sg13g2_dfrbp_1 _5018_ (.CLK(clk),
    .RESET_B(net826),
    .D(net349),
    .Q_N(_0053_),
    .Q(\measurements.alreadytriggered_reg ));
 sg13g2_dfrbp_1 _5019_ (.CLK(clk),
    .RESET_B(net817),
    .D(net533),
    .Q_N(_0032_),
    .Q(\measurements.address_counter_reg[0] ));
 sg13g2_dfrbp_1 _5020_ (.CLK(clk),
    .RESET_B(net812),
    .D(net417),
    .Q_N(_0056_),
    .Q(\measurements.address_counter_reg[1] ));
 sg13g2_dfrbp_1 _5021_ (.CLK(clk),
    .RESET_B(net812),
    .D(net315),
    .Q_N(_0057_),
    .Q(\measurements.address_counter_reg[2] ));
 sg13g2_dfrbp_1 _5022_ (.CLK(clk),
    .RESET_B(net812),
    .D(net451),
    .Q_N(_0058_),
    .Q(\measurements.address_counter_reg[3] ));
 sg13g2_dfrbp_1 _5023_ (.CLK(clk),
    .RESET_B(net812),
    .D(net475),
    .Q_N(_0059_),
    .Q(\measurements.address_counter_reg[4] ));
 sg13g2_dfrbp_1 _5024_ (.CLK(clk),
    .RESET_B(net813),
    .D(net478),
    .Q_N(_0060_),
    .Q(\measurements.address_counter_reg[5] ));
 sg13g2_dfrbp_1 _5025_ (.CLK(clk),
    .RESET_B(net813),
    .D(net462),
    .Q_N(_0061_),
    .Q(\measurements.address_counter_reg[6] ));
 sg13g2_dfrbp_1 _5026_ (.CLK(clk),
    .RESET_B(net814),
    .D(net435),
    .Q_N(_0062_),
    .Q(\measurements.address_counter_reg[7] ));
 sg13g2_dfrbp_1 _5027_ (.CLK(clk),
    .RESET_B(net818),
    .D(net291),
    .Q_N(_0063_),
    .Q(\measurements.address_counter_reg[8] ));
 sg13g2_dfrbp_1 _5028_ (.CLK(clk),
    .RESET_B(net817),
    .D(net304),
    .Q_N(_0064_),
    .Q(\measurements.address_counter_reg[9] ));
 sg13g2_dfrbp_1 _5029_ (.CLK(clk),
    .RESET_B(net817),
    .D(net288),
    .Q_N(_0065_),
    .Q(\measurements.address_counter_reg[10] ));
 sg13g2_dfrbp_1 _5030_ (.CLK(clk),
    .RESET_B(net816),
    .D(net393),
    .Q_N(_0066_),
    .Q(\measurements.address_counter_reg[11] ));
 sg13g2_dfrbp_1 _5031_ (.CLK(clk),
    .RESET_B(net815),
    .D(net299),
    .Q_N(_0067_),
    .Q(\measurements.address_counter_reg[12] ));
 sg13g2_dfrbp_1 _5032_ (.CLK(clk),
    .RESET_B(net815),
    .D(net364),
    .Q_N(_0068_),
    .Q(\measurements.address_counter_reg[13] ));
 sg13g2_dfrbp_1 _5033_ (.CLK(clk),
    .RESET_B(net817),
    .D(net130),
    .Q_N(\measurements.address_counter_reg[14] ),
    .Q(_0085_));
 sg13g2_dfrbp_1 _5034_ (.CLK(clk),
    .RESET_B(net822),
    .D(net139),
    .Q_N(_2401_),
    .Q(\siggen.dac_pmod.n50_o[0] ));
 sg13g2_dfrbp_1 _5035_ (.CLK(clk),
    .RESET_B(net822),
    .D(net78),
    .Q_N(_2400_),
    .Q(\siggen.dac_pmod.n50_o[1] ));
 sg13g2_dfrbp_1 _5036_ (.CLK(clk),
    .RESET_B(net822),
    .D(net89),
    .Q_N(_2399_),
    .Q(\siggen.dac_pmod.n50_o[2] ));
 sg13g2_dfrbp_1 _5037_ (.CLK(clk),
    .RESET_B(net821),
    .D(net100),
    .Q_N(_2398_),
    .Q(\siggen.dac_pmod.n50_o[3] ));
 sg13g2_dfrbp_1 _5038_ (.CLK(clk),
    .RESET_B(net821),
    .D(net145),
    .Q_N(_2397_),
    .Q(\siggen.dac_pmod.n50_o[4] ));
 sg13g2_dfrbp_1 _5039_ (.CLK(clk),
    .RESET_B(net821),
    .D(net106),
    .Q_N(_2396_),
    .Q(\siggen.dac_pmod.n50_o[5] ));
 sg13g2_dfrbp_1 _5040_ (.CLK(clk),
    .RESET_B(net821),
    .D(net127),
    .Q_N(_2395_),
    .Q(\siggen.dac_pmod.n50_o[6] ));
 sg13g2_dfrbp_1 _5041_ (.CLK(clk),
    .RESET_B(net821),
    .D(net60),
    .Q_N(_2394_),
    .Q(\siggen.dac_pmod.n66_o ));
 sg13g2_dfrbp_1 _5042_ (.CLK(clk),
    .RESET_B(net822),
    .D(net42),
    .Q_N(\siggen.n20_o ),
    .Q(\siggen.n22_o ));
 sg13g2_dfrbp_1 _5043_ (.CLK(clk),
    .RESET_B(net823),
    .D(net266),
    .Q_N(_2393_),
    .Q(\siggen.dac_pmod.cnt_reg[0] ));
 sg13g2_dfrbp_1 _5044_ (.CLK(clk),
    .RESET_B(net823),
    .D(net150),
    .Q_N(_2392_),
    .Q(\siggen.dac_pmod.cnt_reg[1] ));
 sg13g2_dfrbp_1 _5045_ (.CLK(clk),
    .RESET_B(net823),
    .D(net312),
    .Q_N(_2391_),
    .Q(\siggen.dac_pmod.cnt_reg[2] ));
 sg13g2_dfrbp_1 _5046_ (.CLK(clk),
    .RESET_B(net823),
    .D(net472),
    .Q_N(_2390_),
    .Q(\siggen.dac_pmod.cnt_reg[3] ));
 sg13g2_dfrbp_1 _5047_ (.CLK(clk),
    .RESET_B(net823),
    .D(net258),
    .Q_N(\siggen.da_sclk ),
    .Q(\siggen.dac_pmod.n88_q ));
 sg13g2_dfrbp_1 _5048_ (.CLK(clk),
    .RESET_B(net802),
    .D(net75),
    .Q_N(\settings_uart_printer.uart_tx_module.counter_reg[0] ),
    .Q(_0086_));
 sg13g2_dfrbp_1 _5049_ (.CLK(clk),
    .RESET_B(net802),
    .D(net57),
    .Q_N(\settings_uart_printer.uart_tx_module.counter_reg[1] ),
    .Q(_0087_));
 sg13g2_dfrbp_1 _5050_ (.CLK(clk),
    .RESET_B(net802),
    .D(net92),
    .Q_N(_0012_),
    .Q(\settings_uart_printer.uart_tx_module.counter_reg[2] ));
 sg13g2_dfrbp_1 _5051_ (.CLK(clk),
    .RESET_B(net802),
    .D(net54),
    .Q_N(\settings_uart_printer.uart_tx_module.counter_reg[3] ),
    .Q(_0088_));
 sg13g2_dfrbp_1 _5052_ (.CLK(clk),
    .RESET_B(net802),
    .D(net183),
    .Q_N(_2389_),
    .Q(\settings_uart_printer.uart_tx_module.counter_reg[4] ));
 sg13g2_dfrbp_1 _5053_ (.CLK(clk),
    .RESET_B(net802),
    .D(net39),
    .Q_N(\settings_uart_printer.uart_tx_module.counter_reg[5] ),
    .Q(_0089_));
 sg13g2_dfrbp_1 _5054_ (.CLK(clk),
    .RESET_B(net803),
    .D(net224),
    .Q_N(_2388_),
    .Q(\settings_uart_printer.uart_tx_module.counter_reg[6] ));
 sg13g2_dfrbp_1 _5055_ (.CLK(clk),
    .RESET_B(net803),
    .D(net153),
    .Q_N(_2387_),
    .Q(\settings_uart_printer.uart_tx_module.counter_reg[7] ));
 sg13g2_dfrbp_1 _5056_ (.CLK(clk),
    .RESET_B(net802),
    .D(net354),
    .Q_N(_2386_),
    .Q(\settings_uart_printer.uart_tx_module.counter_reg[8] ));
 sg13g2_dfrbp_1 _5057_ (.CLK(clk),
    .RESET_B(net802),
    .D(net33),
    .Q_N(\settings_uart_printer.uart_tx_module.counter_reg[9] ),
    .Q(_0090_));
 sg13g2_dfrbp_1 _5058_ (.CLK(clk),
    .RESET_B(net806),
    .D(net159),
    .Q_N(_2385_),
    .Q(\settings_uart_printer.uart_tx_module.counter_reg[10] ));
 sg13g2_dfrbp_1 _5059_ (.CLK(clk),
    .RESET_B(net807),
    .D(net111),
    .Q_N(\settings_uart_printer.uart_tx_module.counter_reg[11] ),
    .Q(_0091_));
 sg13g2_dfrbp_1 _5060_ (.CLK(clk),
    .RESET_B(net819),
    .D(net494),
    .Q_N(_0036_),
    .Q(\siggen.n66_q[0] ));
 sg13g2_dfrbp_1 _5061_ (.CLK(clk),
    .RESET_B(net819),
    .D(net439),
    .Q_N(_0039_),
    .Q(\siggen.n66_q[1] ));
 sg13g2_dfrbp_1 _5062_ (.CLK(clk),
    .RESET_B(net819),
    .D(net854),
    .Q_N(_0038_),
    .Q(\siggen.n66_q[2] ));
 sg13g2_dfrbp_1 _5063_ (.CLK(clk),
    .RESET_B(net819),
    .D(net599),
    .Q_N(_0037_),
    .Q(\siggen.n49_o[3] ));
 sg13g2_dfrbp_1 _5064_ (.CLK(clk),
    .RESET_B(net819),
    .D(net386),
    .Q_N(_0035_),
    .Q(\siggen.n49_o[4] ));
 sg13g2_dfrbp_1 _5065_ (.CLK(clk),
    .RESET_B(net821),
    .D(net625),
    .Q_N(_0034_),
    .Q(\siggen.n49_o[5] ));
 sg13g2_dfrbp_1 _5066_ (.CLK(clk),
    .RESET_B(net821),
    .D(net268),
    .Q_N(_0033_),
    .Q(\siggen.n49_o[6] ));
 sg13g2_dfrbp_1 _5067_ (.CLK(clk),
    .RESET_B(net821),
    .D(net321),
    .Q_N(_0040_),
    .Q(\siggen.n49_o[7] ));
 sg13g2_tiehi tt_um_gfcwfzkm_scope_bfh_mht1_3_10 (.L_HI(net10));
 sg13g2_tiehi tt_um_gfcwfzkm_scope_bfh_mht1_3_11 (.L_HI(net11));
 sg13g2_tiehi tt_um_gfcwfzkm_scope_bfh_mht1_3_12 (.L_HI(net12));
 sg13g2_tiehi tt_um_gfcwfzkm_scope_bfh_mht1_3_13 (.L_HI(net13));
 sg13g2_tiehi tt_um_gfcwfzkm_scope_bfh_mht1_3_14 (.L_HI(net14));
 sg13g2_tiehi tt_um_gfcwfzkm_scope_bfh_mht1_3_15 (.L_HI(net15));
 sg13g2_tiehi tt_um_gfcwfzkm_scope_bfh_mht1_3_16 (.L_HI(net16));
 sg13g2_dlygate4sd3_1 hold1 (.A(net860),
    .X(net17));
 sg13g2_buf_1 _5076_ (.A(\measurements.adc_cs ),
    .X(uio_out[0]));
 sg13g2_buf_1 _5077_ (.A(\siggen.da_mosi ),
    .X(uio_out[1]));
 sg13g2_buf_1 _5078_ (.A(\measurements.adc_sclk ),
    .X(uio_out[2]));
 sg13g2_buf_1 _5079_ (.A(\measurements.fram_sclk ),
    .X(uio_out[3]));
 sg13g2_buf_1 _5080_ (.A(\siggen.da_cs ),
    .X(uio_out[4]));
 sg13g2_buf_1 _5081_ (.A(\siggen.da_sclk ),
    .X(uio_out[5]));
 sg13g2_buf_2 _5082_ (.A(\measurements.fram_cs ),
    .X(uio_out[6]));
 sg13g2_buf_1 _5083_ (.A(\measurements.fram_mosi ),
    .X(uio_out[7]));
 sg13g2_buf_4 _5084_ (.X(uo_out[0]),
    .A(\videogen.g ));
 sg13g2_buf_1 _5085_ (.A(clk),
    .X(uo_out[1]));
 sg13g2_buf_2 _5086_ (.A(\videogen.hsync ),
    .X(uo_out[2]));
 sg13g2_buf_4 _5087_ (.X(uo_out[3]),
    .A(\settings_uart_printer.tx ));
 sg13g2_buf_4 _5088_ (.X(uo_out[4]),
    .A(\videogen.r ));
 sg13g2_buf_4 _5089_ (.X(uo_out[5]),
    .A(\videogen.b ));
 sg13g2_buf_4 _5090_ (.X(uo_out[6]),
    .A(\videogen.de ));
 sg13g2_buf_4 _5091_ (.X(uo_out[7]),
    .A(\videogen.video_timing_generator.hdmi_vsync ));
 sg13g2_buf_2 fanout633 (.A(net634),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_1118_),
    .X(net634));
 sg13g2_buf_4 fanout635 (.X(net635),
    .A(_0621_));
 sg13g2_buf_4 fanout636 (.X(net636),
    .A(net637));
 sg13g2_buf_4 fanout637 (.X(net637),
    .A(_1151_));
 sg13g2_buf_2 fanout638 (.A(_0339_),
    .X(net638));
 sg13g2_buf_4 fanout639 (.X(net639),
    .A(net640));
 sg13g2_buf_4 fanout640 (.X(net640),
    .A(_1152_));
 sg13g2_buf_2 fanout641 (.A(_0674_),
    .X(net641));
 sg13g2_buf_1 fanout642 (.A(_0674_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_1650_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_1650_),
    .X(net644));
 sg13g2_buf_4 fanout645 (.X(net645),
    .A(net646));
 sg13g2_buf_4 fanout646 (.X(net646),
    .A(_0616_));
 sg13g2_buf_4 fanout647 (.X(net647),
    .A(_1041_));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(net649));
 sg13g2_buf_4 fanout649 (.X(net649),
    .A(_0613_));
 sg13g2_buf_2 fanout650 (.A(_1098_),
    .X(net650));
 sg13g2_buf_4 fanout651 (.X(net651),
    .A(_1040_));
 sg13g2_buf_2 fanout652 (.A(_0662_),
    .X(net652));
 sg13g2_buf_4 fanout653 (.X(net653),
    .A(_2195_));
 sg13g2_buf_2 fanout654 (.A(_1711_),
    .X(net654));
 sg13g2_buf_4 fanout655 (.X(net655),
    .A(_2123_));
 sg13g2_buf_2 fanout656 (.A(_2095_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_2095_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(net660),
    .X(net658));
 sg13g2_buf_1 fanout659 (.A(net660),
    .X(net659));
 sg13g2_buf_4 fanout660 (.X(net660),
    .A(_2094_));
 sg13g2_buf_2 fanout661 (.A(net662),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(net665),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(net665),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net665),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_1357_),
    .X(net665));
 sg13g2_buf_4 fanout666 (.X(net666),
    .A(net667));
 sg13g2_buf_4 fanout667 (.X(net667),
    .A(_1356_));
 sg13g2_buf_4 fanout668 (.X(net668),
    .A(_0934_));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(_0933_));
 sg13g2_buf_4 fanout670 (.X(net670),
    .A(net671));
 sg13g2_buf_1 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_0933_),
    .X(net672));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(_0611_));
 sg13g2_buf_4 fanout674 (.X(net674),
    .A(_2247_));
 sg13g2_buf_2 fanout675 (.A(_2247_),
    .X(net675));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(_2245_));
 sg13g2_buf_1 fanout677 (.A(_2245_),
    .X(net677));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(_2244_));
 sg13g2_buf_1 fanout679 (.A(_2244_),
    .X(net679));
 sg13g2_buf_4 fanout680 (.X(net680),
    .A(_2235_));
 sg13g2_buf_4 fanout681 (.X(net681),
    .A(_1721_));
 sg13g2_buf_2 fanout682 (.A(_0841_),
    .X(net682));
 sg13g2_buf_4 fanout683 (.X(net683),
    .A(_0655_));
 sg13g2_buf_4 fanout684 (.X(net684),
    .A(_2253_));
 sg13g2_buf_2 fanout685 (.A(_2236_),
    .X(net685));
 sg13g2_buf_4 fanout686 (.X(net686),
    .A(_2223_));
 sg13g2_buf_2 fanout687 (.A(_2223_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_2172_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_2172_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_1 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(_2110_),
    .X(net692));
 sg13g2_buf_4 fanout693 (.X(net693),
    .A(_2053_));
 sg13g2_buf_2 fanout694 (.A(_2052_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_2033_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(net701),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(net701),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(net701),
    .X(net699));
 sg13g2_buf_1 fanout700 (.A(net701),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_2028_),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(net704),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(net704),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(_2025_),
    .X(net704));
 sg13g2_buf_4 fanout705 (.X(net705),
    .A(_2024_));
 sg13g2_buf_2 fanout706 (.A(_2024_),
    .X(net706));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(net941));
 sg13g2_buf_2 fanout708 (.A(net941),
    .X(net708));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(net267));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(net711));
 sg13g2_buf_2 fanout711 (.A(net623),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(\siggen.n49_o[4] ),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(net714),
    .X(net713));
 sg13g2_buf_4 fanout714 (.X(net714),
    .A(net1009));
 sg13g2_buf_2 fanout715 (.A(net716),
    .X(net715));
 sg13g2_buf_1 fanout716 (.A(net719),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(net718),
    .X(net717));
 sg13g2_buf_4 fanout718 (.X(net718),
    .A(net719));
 sg13g2_buf_2 fanout719 (.A(net983),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(net853),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(net722),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(net723),
    .X(net722));
 sg13g2_buf_4 fanout723 (.X(net723),
    .A(net724));
 sg13g2_buf_1 fanout724 (.A(net852),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(net727),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(net727),
    .X(net726));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(net436));
 sg13g2_buf_2 fanout728 (.A(net729),
    .X(net728));
 sg13g2_buf_4 fanout729 (.X(net729),
    .A(net491));
 sg13g2_buf_2 fanout730 (.A(net384),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(net732),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(net531),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(net603),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(net735),
    .X(net734));
 sg13g2_buf_1 fanout735 (.A(net608),
    .X(net735));
 sg13g2_buf_4 fanout736 (.X(net736),
    .A(net521));
 sg13g2_buf_2 fanout737 (.A(net957),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(net626),
    .X(net738));
 sg13g2_buf_4 fanout739 (.X(net739),
    .A(net591));
 sg13g2_buf_2 fanout740 (.A(\choffset[3] ),
    .X(net740));
 sg13g2_buf_4 fanout741 (.X(net741),
    .A(net995));
 sg13g2_buf_2 fanout742 (.A(\choffset[2] ),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(net313),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(net746),
    .X(net744));
 sg13g2_buf_1 fanout745 (.A(net746),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(net747),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(net585),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(\measurements.n200_o[2] ),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(\measurements.n200_o[2] ),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(net751),
    .X(net750));
 sg13g2_buf_1 fanout751 (.A(net752),
    .X(net751));
 sg13g2_buf_4 fanout752 (.X(net752),
    .A(net509));
 sg13g2_buf_4 fanout753 (.X(net753),
    .A(net509));
 sg13g2_buf_1 fanout754 (.A(\measurements.n200_o[1] ),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(net757),
    .X(net755));
 sg13g2_buf_1 fanout756 (.A(net757),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(net758),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(net761),
    .X(net758));
 sg13g2_buf_4 fanout759 (.X(net759),
    .A(net760));
 sg13g2_buf_4 fanout760 (.X(net760),
    .A(net761));
 sg13g2_buf_2 fanout761 (.A(net985),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(net769),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(net765),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(net765),
    .X(net764));
 sg13g2_buf_1 fanout765 (.A(net769),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(net768),
    .X(net766));
 sg13g2_buf_1 fanout767 (.A(net768),
    .X(net767));
 sg13g2_buf_1 fanout768 (.A(net842),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(net632),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(net771),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(net776),
    .X(net771));
 sg13g2_buf_4 fanout772 (.X(net772),
    .A(net775));
 sg13g2_buf_2 fanout773 (.A(net775),
    .X(net773));
 sg13g2_buf_1 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(net776),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(\champlitude[1] ),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(net778),
    .X(net777));
 sg13g2_buf_1 fanout778 (.A(net779),
    .X(net778));
 sg13g2_buf_4 fanout779 (.X(net779),
    .A(\champlitude[0] ));
 sg13g2_buf_2 fanout780 (.A(net781),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(net784),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(net783),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(net784),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(\champlitude[0] ),
    .X(net784));
 sg13g2_buf_4 fanout785 (.X(net785),
    .A(\videogen.draw_y[9] ));
 sg13g2_buf_4 fanout786 (.X(net786),
    .A(net573));
 sg13g2_buf_2 fanout787 (.A(net924),
    .X(net787));
 sg13g2_buf_1 fanout788 (.A(net924),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(net855),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(net791),
    .X(net790));
 sg13g2_buf_1 fanout791 (.A(net846),
    .X(net791));
 sg13g2_buf_4 fanout792 (.X(net792),
    .A(net845));
 sg13g2_buf_4 fanout793 (.X(net793),
    .A(net795));
 sg13g2_buf_1 fanout794 (.A(net795),
    .X(net794));
 sg13g2_buf_1 fanout795 (.A(net797),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(net797),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(net998),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(\settings_uart_printer.n103_q[0] ),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(net969),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(net801),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(net969),
    .X(net801));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(net804));
 sg13g2_buf_4 fanout803 (.X(net803),
    .A(net804));
 sg13g2_buf_4 fanout804 (.X(net804),
    .A(net806));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(net806));
 sg13g2_buf_4 fanout806 (.X(net806),
    .A(net841));
 sg13g2_buf_4 fanout807 (.X(net807),
    .A(net809));
 sg13g2_buf_4 fanout808 (.X(net808),
    .A(net809));
 sg13g2_buf_2 fanout809 (.A(net811),
    .X(net809));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(net811));
 sg13g2_buf_2 fanout811 (.A(net841),
    .X(net811));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(net818));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(net814));
 sg13g2_buf_4 fanout814 (.X(net814),
    .A(net818));
 sg13g2_buf_4 fanout815 (.X(net815),
    .A(net816));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(net817));
 sg13g2_buf_4 fanout817 (.X(net817),
    .A(net818));
 sg13g2_buf_2 fanout818 (.A(net841),
    .X(net818));
 sg13g2_buf_4 fanout819 (.X(net819),
    .A(net820));
 sg13g2_buf_4 fanout820 (.X(net820),
    .A(net825));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(net822));
 sg13g2_buf_4 fanout822 (.X(net822),
    .A(net825));
 sg13g2_buf_4 fanout823 (.X(net823),
    .A(net824));
 sg13g2_buf_4 fanout824 (.X(net824),
    .A(net825));
 sg13g2_buf_2 fanout825 (.A(net841),
    .X(net825));
 sg13g2_buf_4 fanout826 (.X(net826),
    .A(net840));
 sg13g2_buf_4 fanout827 (.X(net827),
    .A(net840));
 sg13g2_buf_4 fanout828 (.X(net828),
    .A(net830));
 sg13g2_buf_4 fanout829 (.X(net829),
    .A(net830));
 sg13g2_buf_2 fanout830 (.A(net840),
    .X(net830));
 sg13g2_buf_4 fanout831 (.X(net831),
    .A(net834));
 sg13g2_buf_4 fanout832 (.X(net832),
    .A(net834));
 sg13g2_buf_2 fanout833 (.A(net834),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(net840),
    .X(net834));
 sg13g2_buf_4 fanout835 (.X(net835),
    .A(net839));
 sg13g2_buf_4 fanout836 (.X(net836),
    .A(net838));
 sg13g2_buf_4 fanout837 (.X(net837),
    .A(net838));
 sg13g2_buf_2 fanout838 (.A(net839),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(net840),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_4 fanout841 (.X(net841),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tiehi tt_um_gfcwfzkm_scope_bfh_mht1_3_9 (.L_HI(net9));
 sg13g2_dlygate4sd3_1 hold2 (.A(net862),
    .X(net18));
 sg13g2_dlygate4sd3_1 hold3 (.A(net858),
    .X(net19));
 sg13g2_dlygate4sd3_1 hold4 (.A(net866),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold5 (.A(net864),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold6 (.A(net868),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0013_),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold8 (.A(_2176_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold9 (.A(net879),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0025_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold11 (.A(net908),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0081_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold13 (.A(_1023_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold14 (.A(net992),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0090_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold16 (.A(_1951_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0283_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0080_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold19 (.A(_1019_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0157_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0089_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold22 (.A(_1946_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0279_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold24 (.A(\siggen.n20_o ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold25 (.A(_1924_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0268_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0082_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold28 (.A(_1085_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0172_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0005_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold31 (.A(_1082_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0170_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0076_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0670_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold35 (.A(net897),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0088_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold37 (.A(_1943_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0277_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0087_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold40 (.A(_1939_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0275_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold42 (.A(\siggen.dac_pmod.n66_o ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold43 (.A(_1921_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold44 (.A(net916),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0075_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0669_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0108_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold48 (.A(\settings_uart_printer.uart_tx_module.data_reg[5] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0819_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0116_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold51 (.A(\settings_uart_printer.uart_tx_module.data_reg[4] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0806_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0115_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold54 (.A(\settings_uart_printer.uart_tx_module.data_reg[6] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0820_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0117_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0086_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold58 (.A(_1938_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0274_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold60 (.A(\siggen.dac_pmod.n50_o[1] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold61 (.A(_1774_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0261_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0084_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold64 (.A(_1174_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0211_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold66 (.A(\oscilloscope_control.switch_debouncer_n1_debounce_switches.counter_next[0] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold67 (.A(net891),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold68 (.A(\settings_uart_printer.uart_tx_module.data_reg[3] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0790_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0114_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold71 (.A(\siggen.dac_pmod.n50_o[2] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold72 (.A(_1816_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0262_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0012_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold75 (.A(_1942_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0276_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold77 (.A(\oscilloscope_control.button_debouncer_n3_debounce_buttons.counter_next[0] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold78 (.A(net889),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0083_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold80 (.A(_1975_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0177_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold82 (.A(\siggen.dac_pmod.n50_o[3] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold83 (.A(_1854_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0263_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold85 (.A(\measurements.address_counter_reg[11] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold86 (.A(_1164_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0203_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold88 (.A(\siggen.dac_pmod.n50_o[5] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold89 (.A(_1897_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold90 (.A(net964),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold91 (.A(\measurements.samples_adc.cnt_reg[1] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold92 (.A(_1169_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0208_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0091_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold95 (.A(net902),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0077_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold97 (.A(net938),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold98 (.A(\settings_uart_printer.uart_tx_module.data_reg[0] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold99 (.A(_2038_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0111_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0053_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0234_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold103 (.A(\lastsample[0] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold104 (.A(_1653_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0236_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold106 (.A(\settings_uart_printer.uart_tx_module.data_reg[1] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0747_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0112_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold109 (.A(\siggen.dac_pmod.n50_o[6] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold110 (.A(_1919_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0266_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0085_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold113 (.A(_1974_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold114 (.A(net950),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold115 (.A(\measurements.n249_q[2] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold116 (.A(_2185_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold117 (.A(\measurements.n175_o[2] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold118 (.A(\measurements.enough_samples_in_fram_reg ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold119 (.A(_1644_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0235_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold121 (.A(\siggen.dac_pmod.n50_o[0] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold122 (.A(_2057_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold123 (.A(net972),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0073_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold125 (.A(_1976_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0106_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold127 (.A(\siggen.dac_pmod.n50_o[4] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold128 (.A(_1896_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0264_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0079_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold131 (.A(net918),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold132 (.A(\siggen.dac_pmod.cnt_reg[1] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold133 (.A(_1928_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0270_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold135 (.A(\settings_uart_printer.uart_tx_module.counter_reg[7] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold136 (.A(_1949_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0281_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold138 (.A(\measurements.n246_q[5] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold139 (.A(_1158_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0197_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold141 (.A(\settings_uart_printer.uart_tx_module.counter_reg[10] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold142 (.A(_1954_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0284_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold144 (.A(\measurements.samples_storage.spi_master_inst.n103_q[2] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold145 (.A(_2031_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0229_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold147 (.A(\oscilloscope_control.button_debouncer_n4_debounce_buttons.debounced ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold148 (.A(_2014_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0133_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold150 (.A(\oscilloscope_control.button_debouncer_n2_debounce_buttons.counter_next[0] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold151 (.A(net873),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold152 (.A(\oscilloscope_control.switch_debouncer_n2_debounce_switches.counter_next[0] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0118_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold154 (.A(\oscilloscope_control.button_debouncer_n3_debounce_buttons.debounced ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0880_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0137_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold157 (.A(\lastsample[1] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold158 (.A(_1656_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0237_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold160 (.A(\oscilloscope_control.n171_o[0] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold161 (.A(net885),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0074_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0664_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0107_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold165 (.A(\settings_uart_printer.uart_tx_module.counter_reg[4] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold166 (.A(_1945_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0278_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold168 (.A(\oscilloscope_control.switch_debouncer_n2_debounce_switches.counter_reg[1] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0119_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold170 (.A(\measurements.samples_storage.n232_q ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0212_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold172 (.A(\oscilloscope_control.button_debouncer_n4_debounce_buttons.counter_next[0] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold173 (.A(net875),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold174 (.A(\oscilloscope_control.switch_debouncer_n1_debounce_switches.counter_reg[2] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0128_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold176 (.A(\lastsample[2] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold177 (.A(_1659_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0238_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold179 (.A(\settings_uart_printer.uart_tx_module.data_reg[2] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0113_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold181 (.A(\measurements.samples_adc.n84_q[1] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0214_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0004_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0654_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0102_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold186 (.A(\oscilloscope_control.button_debouncer_n1_debounce_buttons.counter_next[0] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold187 (.A(net881),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold188 (.A(\oscilloscope_control.button_debouncer_n2_debounce_buttons.debounced ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold189 (.A(_2017_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0141_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold191 (.A(\measurements.address_counter_reg[8] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold192 (.A(_1161_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0200_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold194 (.A(\measurements.samples_storage.spi_master_inst.n103_q[3] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold195 (.A(_1617_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0230_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold197 (.A(\measurements.address_counter_reg[10] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold198 (.A(_1163_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0202_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold200 (.A(\measurements.n249_q[3] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold201 (.A(_2187_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold202 (.A(\measurements.n175_o[3] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold203 (.A(\measurements.address_counter_reg[9] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold204 (.A(_1162_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0201_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold206 (.A(\settings_uart_printer.uart_tx_module.counter_reg[6] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold207 (.A(_1948_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0280_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold209 (.A(\measurements.samples_storage.n170_o ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold210 (.A(_2119_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0000_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold212 (.A(\oscilloscope_control.switch_debouncer_n2_debounce_switches.counter_reg[2] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0834_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0125_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold215 (.A(\oscilloscope_control.button_debouncer_n3_debounce_buttons.counter_reg[2] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0136_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold217 (.A(\measurements.samples_adc.cnt_reg[0] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0207_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold219 (.A(\measurements.n246_q[4] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold220 (.A(_1157_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0196_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold222 (.A(\measurements.samples_storage.spi_master_inst.n103_q[1] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold223 (.A(_1613_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0228_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold225 (.A(\measurements.n249_q[1] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold226 (.A(_2182_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold227 (.A(\measurements.n175_o[1] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold228 (.A(\measurements.samples_storage.spi_master_inst.n18_o ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold229 (.A(_2049_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0222_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold231 (.A(\oscilloscope_control.button_debouncer_n4_debounce_buttons.counter_reg[2] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0132_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold233 (.A(\oscilloscope_control.switch_debouncer_n2_debounce_switches.counter_reg[0] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0835_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0840_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0120_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold237 (.A(\measurements.n246_q[14] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold238 (.A(_1167_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0206_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold240 (.A(\siggen.dac_pmod.n88_q ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold241 (.A(_1937_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0273_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold243 (.A(\display_x[7] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold244 (.A(_1138_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0188_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold246 (.A(\measurements.samples_adc.cnt_reg[3] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold247 (.A(_1172_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0210_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold249 (.A(\siggen.dac_pmod.cnt_reg[0] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0269_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold251 (.A(\siggen.n49_o[6] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0292_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold253 (.A(\oscilloscope_control.button_debouncer_n1_debounce_buttons.debounced ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold254 (.A(_2015_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0145_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold256 (.A(\measurements.n249_q[5] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold257 (.A(_2190_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold258 (.A(\measurements.n175_o[5] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold259 (.A(\display_x[6] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold260 (.A(_1134_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0187_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold262 (.A(\oscilloscope_control.button_debouncer_n3_debounce_buttons.counter_reg[1] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0135_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold264 (.A(\measurements.n249_q[4] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold265 (.A(_2189_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold266 (.A(\measurements.n175_o[4] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold267 (.A(\oscilloscope_control.button_debouncer_n2_debounce_buttons.counter_reg[1] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0139_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0065_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold270 (.A(_1699_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold271 (.A(_1700_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0255_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0063_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold274 (.A(_1694_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0253_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold276 (.A(\siggen.dac_pmod.n85_q[0] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold277 (.A(\siggen.da_cs ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0124_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold279 (.A(\oscilloscope_control.button_debouncer_n1_debounce_buttons.counter_reg[1] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0143_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold281 (.A(\measurements.address_counter_reg[12] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold282 (.A(_1703_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0257_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold284 (.A(\oscilloscope_control.button_debouncer_n4_debounce_buttons.counter_reg[1] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0131_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0064_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold287 (.A(_1697_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0254_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold289 (.A(\measurements.n98_o[3] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0625_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0096_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold292 (.A(\measurements.n246_q[12] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold293 (.A(_1165_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold294 (.A(\siggen.dac_pmod.cnt_reg[2] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold295 (.A(_1933_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0271_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold297 (.A(\measurements.n163_o[0] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold298 (.A(_1680_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0247_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold300 (.A(\measurements.samples_storage.spi_master_inst.n24_o ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold301 (.A(_2046_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0219_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0033_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold304 (.A(_1973_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0293_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold306 (.A(\measurements.n98_o[0] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold307 (.A(_1148_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0191_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold309 (.A(\measurements.address_counter_reg[7] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold310 (.A(_1160_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0199_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold312 (.A(\lastsample[5] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold313 (.A(_1991_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0241_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold315 (.A(\oscilloscope_control.n146_o[0] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold316 (.A(net986),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold317 (.A(\measurements.samples_storage.n101_o ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold318 (.A(_2113_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold319 (.A(_2114_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0092_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0021_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold322 (.A(_2196_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold323 (.A(\videogen.video_timing_generator.n21_o[2] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold324 (.A(\measurements.samples_storage.spi_master_inst.n96_o ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold325 (.A(_1119_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0180_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold327 (.A(\measurements.memoryShift[8] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0169_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold329 (.A(\measurements.n244_o[3] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0099_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold331 (.A(\measurements.alreadytriggered_reg ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold332 (.A(_1983_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0244_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold334 (.A(\oscilloscope_control.button_debouncer_n2_debounce_buttons.counter_reg[2] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0140_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold336 (.A(\settings_uart_printer.uart_tx_module.counter_reg[8] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold337 (.A(_1950_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0282_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold339 (.A(\oscilloscope_control.switch_debouncer_n1_debounce_switches.counter_reg[1] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0127_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold341 (.A(\measurements.n244_o[1] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0627_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0098_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold344 (.A(\dsgfreqshift[1] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0174_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold346 (.A(\measurements.address_counter_reg[13] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold347 (.A(_1706_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0258_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold349 (.A(\measurements.address_counter_reg[3] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold350 (.A(_1156_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0195_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold352 (.A(\oscilloscope_control.button_debouncer_n1_debounce_buttons.counter_reg[2] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold353 (.A(_0144_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold354 (.A(\measurements.n246_q[2] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold355 (.A(_1155_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0194_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold357 (.A(\measurements.n246_q[13] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold358 (.A(_1166_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold359 (.A(\measurements.samples_storage.spi_master_inst.n22_o ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold360 (.A(_2047_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0220_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold362 (.A(\lastsample[6] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold363 (.A(_1990_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0242_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold365 (.A(\display_x[8] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold366 (.A(_1140_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0189_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold368 (.A(\siggen.n22_o ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold369 (.A(_1967_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0290_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold371 (.A(\lastsample[3] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold372 (.A(_1662_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0239_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0066_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold375 (.A(_1701_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold376 (.A(_1702_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0256_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold378 (.A(\measurements.address_counter_reg[6] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold379 (.A(_1159_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0198_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold381 (.A(\videogen.draw_y[3] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold382 (.A(\videogen.video_timing_generator.n21_o[3] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold383 (.A(\measurements.n98_o[2] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0624_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0095_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold386 (.A(\measurements.memoryShift[3] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold387 (.A(_1054_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0164_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold389 (.A(\display_x[1] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0182_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold391 (.A(\display_x[3] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold392 (.A(_1127_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0184_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold394 (.A(\measurements.trigger.trigger_threshold[2] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold395 (.A(_1024_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0159_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0054_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold398 (.A(\measurements.n182_o ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold399 (.A(\measurements.address_counter_reg[1] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold400 (.A(_1677_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0246_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold402 (.A(\measurements.memoryShift[5] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold403 (.A(_1064_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0166_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold405 (.A(\settings_uart_printer.uart_tx_module.datacnt_reg[2] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0639_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0641_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold408 (.A(_0100_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold409 (.A(\measurements.samples_adc.cnt_reg[2] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0209_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold411 (.A(\measurements.n98_o[1] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0093_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold413 (.A(\lastsample[4] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold414 (.A(_1664_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0240_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0061_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold417 (.A(_1688_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold418 (.A(_1691_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0252_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold420 (.A(\siggen.n66_q[1] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold421 (.A(net727),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold422 (.A(_1962_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0287_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold424 (.A(\measurements.memoryShift[6] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold425 (.A(net1002),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold426 (.A(_0014_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold427 (.A(_2039_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold428 (.A(_1123_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold429 (.A(_0183_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold430 (.A(\lastsample[7] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold431 (.A(_1673_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold432 (.A(_0243_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold433 (.A(_0058_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold434 (.A(_1681_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold435 (.A(_0248_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold436 (.A(\measurements.n246_q[1] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold437 (.A(_1154_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold438 (.A(\measurements.memoryShift[2] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold439 (.A(_0163_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold440 (.A(\measurements.samples_storage.spi_master_inst.n26_o ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold441 (.A(_2045_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold442 (.A(_0218_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold443 (.A(\measurements.address_counter_reg[4] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold444 (.A(_1635_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold445 (.A(_1689_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0251_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold447 (.A(\measurements.memoryShift[7] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0168_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold449 (.A(_0023_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold450 (.A(\videogen.video_timing_generator.n21_o[6] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold451 (.A(\measurements.samples_storage.spi_master_inst.n20_o ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold452 (.A(_2048_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold453 (.A(_0221_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold454 (.A(\siggen.dac_pmod.cnt_reg[3] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold455 (.A(_1935_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0272_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold457 (.A(_0059_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold458 (.A(_1684_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold459 (.A(_0249_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0060_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold461 (.A(_1686_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold462 (.A(_0250_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold463 (.A(\measurements.n244_o[0] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold464 (.A(_1985_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold465 (.A(_0626_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0097_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold467 (.A(\settings_uart_printer.uart_tx_module.n88_q[1] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold468 (.A(_0647_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold469 (.A(_0101_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold470 (.A(\measurements.memoryShift[4] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold471 (.A(_0165_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold472 (.A(\oscilloscope_control.n206_o ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold473 (.A(_2018_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold474 (.A(_0129_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold475 (.A(\siggen.n66_q[0] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold476 (.A(net729),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold477 (.A(_1957_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold478 (.A(_0286_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold479 (.A(_0022_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold480 (.A(\videogen.video_timing_generator.n21_o[5] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold481 (.A(\measurements.samples_adc.n84_q[0] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold482 (.A(_0621_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold483 (.A(_0094_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold484 (.A(\settings_uart_printer.n103_q[5] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold485 (.A(_0652_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold486 (.A(_0122_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold487 (.A(\measurements.samples_storage.spi_master_inst.n100_q[0] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold488 (.A(_2111_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold489 (.A(_0155_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold490 (.A(\measurements.fram_sclk ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold491 (.A(_1612_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold492 (.A(_0227_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold493 (.A(\measurements.n200_o[1] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold494 (.A(net752),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold495 (.A(_0150_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold496 (.A(\measurements.n246_q[0] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold497 (.A(_1153_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold498 (.A(_0192_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold499 (.A(\oscilloscope_control.n220_q[1] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold500 (.A(_0929_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold501 (.A(_0153_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold502 (.A(\display_x[4] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold503 (.A(_1129_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold504 (.A(_0185_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold505 (.A(\display_x[5] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold506 (.A(net736),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold507 (.A(_1132_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold508 (.A(_0186_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold509 (.A(\measurements.samples_storage.spi_master_inst.n30_o ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold510 (.A(_2043_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold511 (.A(_0216_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold512 (.A(\measurements.samples_storage.spi_master_inst.n28_o ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold513 (.A(_2044_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold514 (.A(_0217_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold515 (.A(\measurements.address_counter_reg[0] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold516 (.A(net732),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold517 (.A(_0245_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold518 (.A(\measurements.trigger.trigger_threshold[3] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold519 (.A(_1987_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold520 (.A(_0160_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold521 (.A(_0026_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold522 (.A(_2207_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold523 (.A(\videogen.video_timing_generator.n21_o[9] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold524 (.A(_0055_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold525 (.A(_1144_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold526 (.A(_1145_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold527 (.A(_0190_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold528 (.A(_0041_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold529 (.A(_1115_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold530 (.A(_1116_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold531 (.A(_0179_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold532 (.A(\measurements.samples_storage.n230_q[0] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold533 (.A(_0223_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold534 (.A(\measurements.n163_o[1] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold535 (.A(_0171_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold536 (.A(\measurements.samples_storage.spi_master_inst.n100_q[1] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0949_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold538 (.A(_0156_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold539 (.A(\oscilloscope_control.n111_o[0] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold540 (.A(_1099_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold541 (.A(_0175_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold542 (.A(\oscilloscope_control.n220_q[0] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold543 (.A(_0152_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold544 (.A(\videogen.draw_y[0] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold545 (.A(\videogen.video_timing_generator.n21_o[0] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold546 (.A(\measurements.adc_sclk ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold547 (.A(_0619_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0213_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold549 (.A(\measurements.memoryShift[0] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold550 (.A(_0161_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold551 (.A(\measurements.memoryShift[1] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold552 (.A(_0162_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold553 (.A(\siggen.dac_pmod.n85_q[1] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold554 (.A(_0841_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold555 (.A(_0843_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold556 (.A(_0123_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold557 (.A(_0024_),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold558 (.A(net786),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold559 (.A(\videogen.video_timing_generator.n21_o[7] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold560 (.A(\measurements.n250_q[1] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold561 (.A(_1980_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold562 (.A(_0232_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold563 (.A(\measurements.n250_q[2] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold564 (.A(_1981_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold565 (.A(_0233_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold566 (.A(\choffset[1] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold567 (.A(_2026_),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold568 (.A(_0176_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold569 (.A(\measurements.n200_o[2] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold570 (.A(net747),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold571 (.A(_0151_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold572 (.A(\measurements.samples_storage.n230_q[3] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold573 (.A(_1992_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold574 (.A(_0226_),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold575 (.A(\choffset[3] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold576 (.A(net739),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold577 (.A(_0178_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold578 (.A(\settings_uart_printer.n104_q[0] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold579 (.A(_0642_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold580 (.A(_0103_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold581 (.A(_0037_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold582 (.A(_1966_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold583 (.A(_0289_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold584 (.A(\oscilloscope_control.n114_o[0] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold585 (.A(_0906_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold586 (.A(_0146_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold587 (.A(\measurements.samples_storage.n230_q[2] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold588 (.A(_2072_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold589 (.A(_1607_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold590 (.A(_1608_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold591 (.A(_0224_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold592 (.A(\measurements.samples_storage.n230_q[1] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold593 (.A(_2073_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold594 (.A(_0942_),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold595 (.A(_1609_),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold596 (.A(_0225_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold597 (.A(\videogen.draw_y[4] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold598 (.A(_2197_),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold599 (.A(\videogen.video_timing_generator.n21_o[4] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold600 (.A(\settings_uart_printer.uart_tx_module.n88_q[0] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold601 (.A(\measurements.fram_mosi ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold602 (.A(_2050_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold603 (.A(_0215_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold604 (.A(\measurements.n250_q[0] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold605 (.A(_1979_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold606 (.A(_0231_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold607 (.A(\siggen.n49_o[5] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold608 (.A(net711),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold609 (.A(_0291_),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold610 (.A(\display_x[0] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold611 (.A(net738),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold612 (.A(_0181_),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold613 (.A(\videogen.draw_y[1] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold614 (.A(_2078_),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold615 (.A(\videogen.video_timing_generator.n21_o[1] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold616 (.A(\champlitude[2] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold617 (.A(net769),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold618 (.A(_0909_),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold619 (.A(_0148_),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold620 (.A(\settings_uart_printer.n103_q[2] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold621 (.A(net792),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold622 (.A(_0659_),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold623 (.A(_0104_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold624 (.A(\oscilloscope_control.switch_debouncer_n1_debounce_switches.debounced ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold625 (.A(_0902_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold626 (.A(_0147_),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold627 (.A(\siggen.n66_q[2] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold628 (.A(net724),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold629 (.A(_0288_),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold630 (.A(\settings_uart_printer.n103_q[3] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold631 (.A(net789),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold632 (.A(_0105_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold633 (.A(\oscilloscope_control.n223_q[0] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold634 (.A(net19),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold635 (.A(\oscilloscope_control.button_ff_stage_1_reg[1] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold636 (.A(net17),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold637 (.A(\oscilloscope_control.n223_q[1] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold638 (.A(net18),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold639 (.A(\oscilloscope_control.button_ff_stage_1_reg[3] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold640 (.A(net21),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold641 (.A(\oscilloscope_control.button_ff_stage_1_reg[2] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold642 (.A(net20),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold643 (.A(\oscilloscope_control.button_ff_stage_1_reg[0] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold644 (.A(net22),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold645 (.A(\settings_uart_printer.uart_tx_module.counter_reg[1] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold646 (.A(_1940_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold647 (.A(\oscilloscope_control.button_debouncer_n2_debounce_buttons.counter_reg[0] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold648 (.A(_0138_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold649 (.A(\oscilloscope_control.button_debouncer_n4_debounce_buttons.counter_reg[0] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold650 (.A(_0130_),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold651 (.A(\settings_uart_printer.uart_tx_module.counter_reg[9] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold652 (.A(_1952_),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold653 (.A(\measurements.n249_q[0] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold654 (.A(\measurements.n175_o[0] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold655 (.A(\oscilloscope_control.button_debouncer_n1_debounce_buttons.counter_reg[0] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold656 (.A(_0142_),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold657 (.A(\settings_uart_printer.uart_tx_module.counter_reg[5] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold658 (.A(_1947_),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold659 (.A(\dsgfreqshift[0] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold660 (.A(_0173_),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold661 (.A(\settings_uart_printer.uart_tx_module.counter_reg[3] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold662 (.A(_1944_),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold663 (.A(\oscilloscope_control.button_debouncer_n3_debounce_buttons.counter_reg[0] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold664 (.A(_0134_),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold665 (.A(\oscilloscope_control.switch_debouncer_n1_debounce_switches.counter_reg[0] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold666 (.A(_0126_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold667 (.A(_0020_),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold668 (.A(\oscilloscope_control.button_debouncer_n4_debounce_buttons.in_raw ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold669 (.A(\measurements.n244_o[2] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold670 (.A(\settings_uart_printer.uart_tx_module.datacnt_reg[1] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold671 (.A(_0671_),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold672 (.A(_0109_),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold673 (.A(\measurements.address_counter_reg[5] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold674 (.A(_1687_),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold675 (.A(\display_x[2] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold676 (.A(\settings_uart_printer.uart_tx_module.counter_reg[11] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold677 (.A(_0285_),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold678 (.A(_0068_),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold679 (.A(_1707_),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold680 (.A(\oscilloscope_control.button_debouncer_n3_debounce_buttons.in_raw ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold681 (.A(\videogen.draw_y[7] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold682 (.A(_2203_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold683 (.A(\videogen.video_timing_generator.n21_o[8] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold684 (.A(_0067_),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold685 (.A(_0015_),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold686 (.A(_0069_),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold687 (.A(_0885_),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold688 (.A(_0887_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold689 (.A(_0040_),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold690 (.A(_1922_),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold691 (.A(_0267_),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold692 (.A(\measurements.trigger.sample_on_rising_edge ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold693 (.A(_0154_),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold694 (.A(_0072_),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold695 (.A(_0036_),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold696 (.A(\oscilloscope_control.button_debouncer_n1_debounce_buttons.in_raw ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold697 (.A(_0899_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold698 (.A(\oscilloscope_control.button_debouncer_n2_debounce_buttons.in_raw ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold699 (.A(\settings_uart_printer.n104_q[1] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold700 (.A(\videogen.draw_y[5] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold701 (.A(_0035_),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold702 (.A(\oscilloscope_control.switch_debouncer_n2_debounce_switches.debounced ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold703 (.A(\choffset[4] ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold704 (.A(\measurements.n163_o[2] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold705 (.A(\oscilloscope_control.n208_o ),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold706 (.A(_0839_),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold707 (.A(\display_x[9] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold708 (.A(\choffset[0] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold709 (.A(_0057_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold710 (.A(_0030_),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold711 (.A(_1079_),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold712 (.A(\settings_uart_printer.uart_tx_module.datacnt_reg[0] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold713 (.A(_0110_),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold714 (.A(_0071_),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold715 (.A(\videogen.draw_y[2] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold716 (.A(\siggen.n49_o[7] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold717 (.A(\settings_uart_printer.uart_tx_module.counter_reg[2] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold718 (.A(\videogen.draw_y[6] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold719 (.A(\measurements.n253_q ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold720 (.A(_2077_),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold721 (.A(_0001_),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold722 (.A(_0017_),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold723 (.A(_1133_),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold724 (.A(\measurements.address_counter_reg[14] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold725 (.A(_0259_),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold726 (.A(_0018_),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold727 (.A(_0019_),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold728 (.A(\measurements.n250_q[3] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold729 (.A(\measurements.n249_q[1] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold730 (.A(\videogen.draw_y[8] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold731 (.A(_2083_),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold732 (.A(_0016_),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold733 (.A(\measurements.n246_q[11] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold734 (.A(_1008_),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold735 (.A(_0070_),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold736 (.A(_0034_),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold737 (.A(_1907_),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold738 (.A(_1909_),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold739 (.A(_0265_),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold740 (.A(_0029_),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold741 (.A(_0008_),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold742 (.A(_0926_),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold743 (.A(_0927_),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold744 (.A(\settings_uart_printer.n103_q[0] ),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold745 (.A(_0829_),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold746 (.A(\siggen.da_sclk ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold747 (.A(_0260_),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold748 (.A(_0010_),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold749 (.A(_1031_),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold750 (.A(\measurements.trigger.trigger_threshold[0] ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold751 (.A(_0038_),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold752 (.A(_1852_),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold753 (.A(\measurements.n249_q[0] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold754 (.A(_0039_),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold755 (.A(\oscilloscope_control.n220_q[0] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold756 (.A(_1768_),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold757 (.A(_1873_),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold758 (.A(\siggen.n49_o[3] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold759 (.A(\settings_uart_printer.n103_q[4] ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold760 (.A(\measurements.n200_o[0] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold761 (.A(_0149_),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold762 (.A(_0004_),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold763 (.A(_0812_),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold764 (.A(_0011_),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold765 (.A(_0002_),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold766 (.A(\measurements.trigger.trigger_threshold[1] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold767 (.A(_0158_),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold768 (.A(\measurements.n163_o[1] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold769 (.A(_0744_),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold770 (.A(\choffset[2] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold771 (.A(\dsgfreqshift[0] ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold772 (.A(_0720_),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold773 (.A(\settings_uart_printer.n103_q[1] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold774 (.A(\measurements.trigger.trigger_threshold[1] ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold775 (.A(_0027_),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold776 (.A(_0028_),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold777 (.A(_0167_),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold778 (.A(\settings_uart_printer.n103_q[5] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold779 (.A(_0066_),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold780 (.A(_0009_),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold781 (.A(_0910_),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold782 (.A(_0032_),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold783 (.A(_0062_),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold784 (.A(\siggen.n49_o[4] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold785 (.A(\settings_uart_printer.uart_tx_module.counter_reg[0] ),
    .X(net1010));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_4 FILLER_0_7 ();
 sg13g2_fill_2 FILLER_0_135 ();
 sg13g2_fill_2 FILLER_0_158 ();
 sg13g2_decap_8 FILLER_0_164 ();
 sg13g2_fill_2 FILLER_0_171 ();
 sg13g2_decap_8 FILLER_0_178 ();
 sg13g2_decap_8 FILLER_0_185 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_decap_8 FILLER_0_213 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_227 ();
 sg13g2_decap_8 FILLER_0_234 ();
 sg13g2_decap_8 FILLER_0_241 ();
 sg13g2_decap_8 FILLER_0_248 ();
 sg13g2_decap_8 FILLER_0_255 ();
 sg13g2_fill_2 FILLER_0_262 ();
 sg13g2_fill_1 FILLER_0_264 ();
 sg13g2_decap_8 FILLER_0_276 ();
 sg13g2_fill_1 FILLER_0_283 ();
 sg13g2_decap_8 FILLER_0_296 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_fill_1 FILLER_0_310 ();
 sg13g2_decap_8 FILLER_0_314 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_fill_2 FILLER_0_336 ();
 sg13g2_fill_1 FILLER_0_338 ();
 sg13g2_decap_8 FILLER_0_347 ();
 sg13g2_decap_4 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_4 FILLER_0_404 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_4 FILLER_1_7 ();
 sg13g2_fill_2 FILLER_1_11 ();
 sg13g2_fill_2 FILLER_1_84 ();
 sg13g2_decap_4 FILLER_1_221 ();
 sg13g2_fill_1 FILLER_1_225 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_4 FILLER_1_238 ();
 sg13g2_fill_1 FILLER_1_242 ();
 sg13g2_decap_4 FILLER_1_253 ();
 sg13g2_fill_1 FILLER_1_257 ();
 sg13g2_fill_2 FILLER_1_265 ();
 sg13g2_fill_1 FILLER_1_267 ();
 sg13g2_fill_2 FILLER_1_284 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_4 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_4 ();
 sg13g2_fill_2 FILLER_2_42 ();
 sg13g2_fill_1 FILLER_2_44 ();
 sg13g2_fill_2 FILLER_2_89 ();
 sg13g2_fill_1 FILLER_2_114 ();
 sg13g2_fill_1 FILLER_2_124 ();
 sg13g2_fill_2 FILLER_2_180 ();
 sg13g2_fill_1 FILLER_2_182 ();
 sg13g2_fill_1 FILLER_2_262 ();
 sg13g2_fill_2 FILLER_2_279 ();
 sg13g2_fill_1 FILLER_2_382 ();
 sg13g2_fill_2 FILLER_3_91 ();
 sg13g2_fill_1 FILLER_3_93 ();
 sg13g2_fill_1 FILLER_3_143 ();
 sg13g2_fill_1 FILLER_3_179 ();
 sg13g2_fill_2 FILLER_3_241 ();
 sg13g2_fill_1 FILLER_3_255 ();
 sg13g2_fill_1 FILLER_3_280 ();
 sg13g2_fill_2 FILLER_3_325 ();
 sg13g2_decap_4 FILLER_3_381 ();
 sg13g2_decap_4 FILLER_3_394 ();
 sg13g2_fill_2 FILLER_3_398 ();
 sg13g2_fill_1 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_36 ();
 sg13g2_fill_2 FILLER_4_178 ();
 sg13g2_fill_1 FILLER_4_180 ();
 sg13g2_fill_2 FILLER_4_215 ();
 sg13g2_decap_8 FILLER_4_258 ();
 sg13g2_fill_1 FILLER_4_265 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_4 FILLER_4_280 ();
 sg13g2_fill_2 FILLER_4_284 ();
 sg13g2_decap_8 FILLER_4_292 ();
 sg13g2_fill_2 FILLER_4_299 ();
 sg13g2_fill_1 FILLER_4_301 ();
 sg13g2_fill_2 FILLER_4_324 ();
 sg13g2_fill_1 FILLER_4_338 ();
 sg13g2_fill_1 FILLER_4_363 ();
 sg13g2_fill_1 FILLER_4_384 ();
 sg13g2_fill_2 FILLER_4_395 ();
 sg13g2_fill_1 FILLER_4_397 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_fill_2 FILLER_5_68 ();
 sg13g2_fill_1 FILLER_5_70 ();
 sg13g2_fill_2 FILLER_5_103 ();
 sg13g2_fill_1 FILLER_5_105 ();
 sg13g2_fill_2 FILLER_5_127 ();
 sg13g2_fill_1 FILLER_5_129 ();
 sg13g2_fill_2 FILLER_5_161 ();
 sg13g2_decap_4 FILLER_5_182 ();
 sg13g2_fill_1 FILLER_5_186 ();
 sg13g2_decap_4 FILLER_5_192 ();
 sg13g2_fill_2 FILLER_5_196 ();
 sg13g2_decap_4 FILLER_5_207 ();
 sg13g2_fill_2 FILLER_5_214 ();
 sg13g2_fill_1 FILLER_5_219 ();
 sg13g2_fill_2 FILLER_5_225 ();
 sg13g2_decap_4 FILLER_5_231 ();
 sg13g2_decap_4 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_fill_2 FILLER_5_295 ();
 sg13g2_fill_2 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_327 ();
 sg13g2_decap_8 FILLER_5_334 ();
 sg13g2_decap_8 FILLER_5_341 ();
 sg13g2_decap_8 FILLER_5_348 ();
 sg13g2_fill_2 FILLER_5_355 ();
 sg13g2_decap_4 FILLER_5_362 ();
 sg13g2_fill_1 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_fill_1 FILLER_5_382 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_28 ();
 sg13g2_fill_1 FILLER_6_30 ();
 sg13g2_fill_1 FILLER_6_40 ();
 sg13g2_fill_1 FILLER_6_75 ();
 sg13g2_decap_8 FILLER_6_121 ();
 sg13g2_decap_8 FILLER_6_128 ();
 sg13g2_fill_2 FILLER_6_135 ();
 sg13g2_fill_2 FILLER_6_145 ();
 sg13g2_fill_2 FILLER_6_156 ();
 sg13g2_decap_8 FILLER_6_178 ();
 sg13g2_decap_8 FILLER_6_185 ();
 sg13g2_decap_8 FILLER_6_192 ();
 sg13g2_decap_8 FILLER_6_199 ();
 sg13g2_decap_8 FILLER_6_206 ();
 sg13g2_decap_8 FILLER_6_213 ();
 sg13g2_decap_8 FILLER_6_220 ();
 sg13g2_decap_4 FILLER_6_227 ();
 sg13g2_fill_1 FILLER_6_231 ();
 sg13g2_fill_1 FILLER_6_240 ();
 sg13g2_decap_8 FILLER_6_253 ();
 sg13g2_decap_4 FILLER_6_260 ();
 sg13g2_fill_2 FILLER_6_269 ();
 sg13g2_decap_4 FILLER_6_276 ();
 sg13g2_fill_1 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_fill_1 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_328 ();
 sg13g2_decap_8 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_342 ();
 sg13g2_fill_2 FILLER_6_362 ();
 sg13g2_decap_4 FILLER_6_375 ();
 sg13g2_fill_2 FILLER_6_379 ();
 sg13g2_fill_2 FILLER_6_397 ();
 sg13g2_fill_1 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_66 ();
 sg13g2_fill_2 FILLER_7_107 ();
 sg13g2_fill_1 FILLER_7_118 ();
 sg13g2_fill_2 FILLER_7_145 ();
 sg13g2_decap_8 FILLER_7_164 ();
 sg13g2_fill_2 FILLER_7_171 ();
 sg13g2_fill_1 FILLER_7_173 ();
 sg13g2_fill_1 FILLER_7_179 ();
 sg13g2_fill_2 FILLER_7_197 ();
 sg13g2_decap_8 FILLER_7_215 ();
 sg13g2_decap_4 FILLER_7_239 ();
 sg13g2_fill_2 FILLER_7_243 ();
 sg13g2_decap_4 FILLER_7_278 ();
 sg13g2_fill_2 FILLER_7_302 ();
 sg13g2_decap_4 FILLER_7_320 ();
 sg13g2_fill_2 FILLER_7_353 ();
 sg13g2_fill_2 FILLER_7_369 ();
 sg13g2_fill_1 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_377 ();
 sg13g2_fill_2 FILLER_7_384 ();
 sg13g2_fill_1 FILLER_7_386 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_51 ();
 sg13g2_fill_1 FILLER_8_62 ();
 sg13g2_fill_2 FILLER_8_80 ();
 sg13g2_fill_1 FILLER_8_82 ();
 sg13g2_fill_2 FILLER_8_118 ();
 sg13g2_fill_1 FILLER_8_120 ();
 sg13g2_fill_1 FILLER_8_134 ();
 sg13g2_fill_2 FILLER_8_143 ();
 sg13g2_fill_1 FILLER_8_145 ();
 sg13g2_fill_1 FILLER_8_176 ();
 sg13g2_fill_1 FILLER_8_183 ();
 sg13g2_decap_4 FILLER_8_217 ();
 sg13g2_fill_2 FILLER_8_221 ();
 sg13g2_fill_2 FILLER_8_232 ();
 sg13g2_fill_1 FILLER_8_234 ();
 sg13g2_decap_4 FILLER_8_255 ();
 sg13g2_fill_1 FILLER_8_259 ();
 sg13g2_fill_1 FILLER_8_321 ();
 sg13g2_fill_1 FILLER_8_365 ();
 sg13g2_fill_1 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_fill_2 FILLER_9_74 ();
 sg13g2_fill_1 FILLER_9_76 ();
 sg13g2_fill_2 FILLER_9_101 ();
 sg13g2_fill_1 FILLER_9_103 ();
 sg13g2_fill_2 FILLER_9_131 ();
 sg13g2_fill_1 FILLER_9_133 ();
 sg13g2_fill_1 FILLER_9_186 ();
 sg13g2_fill_2 FILLER_9_205 ();
 sg13g2_decap_8 FILLER_9_242 ();
 sg13g2_fill_1 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_255 ();
 sg13g2_decap_4 FILLER_9_262 ();
 sg13g2_fill_1 FILLER_9_276 ();
 sg13g2_fill_1 FILLER_9_282 ();
 sg13g2_fill_1 FILLER_9_351 ();
 sg13g2_fill_1 FILLER_9_365 ();
 sg13g2_decap_4 FILLER_9_374 ();
 sg13g2_fill_2 FILLER_9_378 ();
 sg13g2_fill_2 FILLER_9_390 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_fill_2 FILLER_10_62 ();
 sg13g2_fill_1 FILLER_10_86 ();
 sg13g2_fill_1 FILLER_10_115 ();
 sg13g2_decap_4 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_142 ();
 sg13g2_fill_1 FILLER_10_161 ();
 sg13g2_decap_4 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_199 ();
 sg13g2_decap_8 FILLER_10_206 ();
 sg13g2_decap_8 FILLER_10_213 ();
 sg13g2_fill_1 FILLER_10_220 ();
 sg13g2_fill_2 FILLER_10_226 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_fill_2 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_4 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_374 ();
 sg13g2_fill_2 FILLER_10_381 ();
 sg13g2_fill_1 FILLER_11_26 ();
 sg13g2_fill_2 FILLER_11_83 ();
 sg13g2_fill_1 FILLER_11_85 ();
 sg13g2_fill_2 FILLER_11_105 ();
 sg13g2_fill_1 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_170 ();
 sg13g2_fill_1 FILLER_11_177 ();
 sg13g2_decap_4 FILLER_11_183 ();
 sg13g2_decap_4 FILLER_11_199 ();
 sg13g2_fill_1 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_209 ();
 sg13g2_fill_2 FILLER_11_216 ();
 sg13g2_fill_2 FILLER_11_240 ();
 sg13g2_fill_1 FILLER_11_242 ();
 sg13g2_fill_2 FILLER_11_255 ();
 sg13g2_fill_1 FILLER_11_257 ();
 sg13g2_decap_4 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_330 ();
 sg13g2_decap_8 FILLER_11_337 ();
 sg13g2_decap_8 FILLER_11_344 ();
 sg13g2_decap_8 FILLER_11_351 ();
 sg13g2_decap_8 FILLER_11_358 ();
 sg13g2_decap_8 FILLER_11_365 ();
 sg13g2_decap_4 FILLER_11_372 ();
 sg13g2_fill_1 FILLER_11_376 ();
 sg13g2_fill_2 FILLER_11_381 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_14 ();
 sg13g2_fill_1 FILLER_12_72 ();
 sg13g2_fill_2 FILLER_12_78 ();
 sg13g2_fill_1 FILLER_12_80 ();
 sg13g2_fill_2 FILLER_12_90 ();
 sg13g2_fill_1 FILLER_12_92 ();
 sg13g2_decap_8 FILLER_12_97 ();
 sg13g2_fill_1 FILLER_12_104 ();
 sg13g2_decap_8 FILLER_12_152 ();
 sg13g2_decap_4 FILLER_12_159 ();
 sg13g2_decap_4 FILLER_12_171 ();
 sg13g2_fill_2 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_198 ();
 sg13g2_decap_4 FILLER_12_205 ();
 sg13g2_fill_1 FILLER_12_209 ();
 sg13g2_decap_4 FILLER_12_215 ();
 sg13g2_fill_1 FILLER_12_219 ();
 sg13g2_fill_2 FILLER_12_233 ();
 sg13g2_fill_2 FILLER_12_256 ();
 sg13g2_fill_1 FILLER_12_258 ();
 sg13g2_fill_1 FILLER_12_313 ();
 sg13g2_fill_2 FILLER_12_347 ();
 sg13g2_fill_1 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_360 ();
 sg13g2_fill_1 FILLER_12_367 ();
 sg13g2_fill_2 FILLER_12_388 ();
 sg13g2_fill_1 FILLER_12_390 ();
 sg13g2_fill_2 FILLER_13_44 ();
 sg13g2_fill_1 FILLER_13_77 ();
 sg13g2_fill_2 FILLER_13_82 ();
 sg13g2_fill_2 FILLER_13_120 ();
 sg13g2_fill_1 FILLER_13_122 ();
 sg13g2_fill_2 FILLER_13_137 ();
 sg13g2_fill_2 FILLER_13_147 ();
 sg13g2_fill_2 FILLER_13_160 ();
 sg13g2_fill_2 FILLER_13_196 ();
 sg13g2_fill_1 FILLER_13_198 ();
 sg13g2_decap_4 FILLER_13_204 ();
 sg13g2_decap_8 FILLER_13_220 ();
 sg13g2_decap_8 FILLER_13_227 ();
 sg13g2_fill_2 FILLER_13_234 ();
 sg13g2_fill_1 FILLER_13_236 ();
 sg13g2_decap_8 FILLER_13_250 ();
 sg13g2_fill_1 FILLER_13_257 ();
 sg13g2_fill_2 FILLER_13_271 ();
 sg13g2_fill_1 FILLER_13_320 ();
 sg13g2_fill_2 FILLER_13_342 ();
 sg13g2_fill_1 FILLER_13_352 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_1 FILLER_14_79 ();
 sg13g2_decap_8 FILLER_14_85 ();
 sg13g2_fill_2 FILLER_14_92 ();
 sg13g2_fill_2 FILLER_14_155 ();
 sg13g2_fill_2 FILLER_14_163 ();
 sg13g2_fill_2 FILLER_14_180 ();
 sg13g2_fill_1 FILLER_14_182 ();
 sg13g2_fill_2 FILLER_14_196 ();
 sg13g2_fill_1 FILLER_14_198 ();
 sg13g2_fill_2 FILLER_14_209 ();
 sg13g2_decap_8 FILLER_14_227 ();
 sg13g2_decap_8 FILLER_14_234 ();
 sg13g2_decap_8 FILLER_14_241 ();
 sg13g2_decap_8 FILLER_14_253 ();
 sg13g2_decap_4 FILLER_14_260 ();
 sg13g2_fill_1 FILLER_14_264 ();
 sg13g2_fill_1 FILLER_14_282 ();
 sg13g2_fill_1 FILLER_14_378 ();
 sg13g2_fill_2 FILLER_14_396 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_fill_2 FILLER_15_18 ();
 sg13g2_fill_2 FILLER_15_62 ();
 sg13g2_fill_1 FILLER_15_64 ();
 sg13g2_fill_2 FILLER_15_70 ();
 sg13g2_fill_1 FILLER_15_96 ();
 sg13g2_fill_2 FILLER_15_164 ();
 sg13g2_decap_8 FILLER_15_197 ();
 sg13g2_decap_8 FILLER_15_204 ();
 sg13g2_decap_8 FILLER_15_211 ();
 sg13g2_fill_1 FILLER_15_218 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_4 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_decap_4 FILLER_15_259 ();
 sg13g2_fill_1 FILLER_15_263 ();
 sg13g2_fill_2 FILLER_15_283 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_4 FILLER_15_332 ();
 sg13g2_fill_2 FILLER_15_336 ();
 sg13g2_decap_4 FILLER_15_344 ();
 sg13g2_fill_1 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_4 FILLER_15_379 ();
 sg13g2_fill_1 FILLER_16_39 ();
 sg13g2_fill_2 FILLER_16_63 ();
 sg13g2_fill_1 FILLER_16_65 ();
 sg13g2_fill_2 FILLER_16_76 ();
 sg13g2_decap_8 FILLER_16_83 ();
 sg13g2_fill_2 FILLER_16_90 ();
 sg13g2_fill_2 FILLER_16_112 ();
 sg13g2_fill_1 FILLER_16_114 ();
 sg13g2_decap_8 FILLER_16_124 ();
 sg13g2_fill_2 FILLER_16_157 ();
 sg13g2_fill_2 FILLER_16_181 ();
 sg13g2_fill_1 FILLER_16_192 ();
 sg13g2_decap_4 FILLER_16_202 ();
 sg13g2_fill_1 FILLER_16_206 ();
 sg13g2_decap_4 FILLER_16_216 ();
 sg13g2_fill_1 FILLER_16_230 ();
 sg13g2_fill_1 FILLER_16_240 ();
 sg13g2_fill_1 FILLER_16_293 ();
 sg13g2_fill_1 FILLER_16_309 ();
 sg13g2_fill_1 FILLER_16_319 ();
 sg13g2_decap_8 FILLER_16_340 ();
 sg13g2_fill_2 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_360 ();
 sg13g2_decap_4 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_fill_2 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_17_26 ();
 sg13g2_decap_4 FILLER_17_53 ();
 sg13g2_decap_8 FILLER_17_82 ();
 sg13g2_decap_8 FILLER_17_89 ();
 sg13g2_decap_8 FILLER_17_96 ();
 sg13g2_decap_4 FILLER_17_103 ();
 sg13g2_fill_1 FILLER_17_107 ();
 sg13g2_decap_8 FILLER_17_117 ();
 sg13g2_decap_8 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_131 ();
 sg13g2_fill_1 FILLER_17_133 ();
 sg13g2_fill_2 FILLER_17_147 ();
 sg13g2_fill_2 FILLER_17_157 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_fill_2 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_241 ();
 sg13g2_decap_4 FILLER_17_248 ();
 sg13g2_fill_1 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_257 ();
 sg13g2_fill_2 FILLER_17_263 ();
 sg13g2_fill_2 FILLER_17_273 ();
 sg13g2_fill_2 FILLER_17_316 ();
 sg13g2_decap_4 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_fill_1 FILLER_17_395 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_47 ();
 sg13g2_fill_2 FILLER_18_76 ();
 sg13g2_fill_1 FILLER_18_78 ();
 sg13g2_fill_1 FILLER_18_97 ();
 sg13g2_decap_8 FILLER_18_113 ();
 sg13g2_decap_4 FILLER_18_120 ();
 sg13g2_fill_2 FILLER_18_124 ();
 sg13g2_fill_1 FILLER_18_171 ();
 sg13g2_fill_1 FILLER_18_190 ();
 sg13g2_decap_8 FILLER_18_206 ();
 sg13g2_decap_8 FILLER_18_213 ();
 sg13g2_fill_2 FILLER_18_220 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_fill_1 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_251 ();
 sg13g2_decap_4 FILLER_18_265 ();
 sg13g2_fill_2 FILLER_18_390 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_4 ();
 sg13g2_fill_2 FILLER_19_27 ();
 sg13g2_fill_2 FILLER_19_50 ();
 sg13g2_fill_1 FILLER_19_52 ();
 sg13g2_fill_1 FILLER_19_122 ();
 sg13g2_fill_2 FILLER_19_149 ();
 sg13g2_fill_1 FILLER_19_160 ();
 sg13g2_decap_4 FILLER_19_197 ();
 sg13g2_fill_1 FILLER_19_201 ();
 sg13g2_decap_4 FILLER_19_206 ();
 sg13g2_decap_8 FILLER_19_227 ();
 sg13g2_decap_4 FILLER_19_253 ();
 sg13g2_fill_1 FILLER_19_257 ();
 sg13g2_fill_2 FILLER_19_263 ();
 sg13g2_fill_1 FILLER_19_265 ();
 sg13g2_decap_8 FILLER_19_271 ();
 sg13g2_decap_8 FILLER_19_278 ();
 sg13g2_decap_8 FILLER_19_285 ();
 sg13g2_decap_8 FILLER_19_292 ();
 sg13g2_fill_1 FILLER_19_299 ();
 sg13g2_decap_4 FILLER_19_309 ();
 sg13g2_fill_2 FILLER_19_318 ();
 sg13g2_decap_8 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_348 ();
 sg13g2_fill_2 FILLER_19_380 ();
 sg13g2_fill_1 FILLER_19_394 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_34 ();
 sg13g2_fill_2 FILLER_20_46 ();
 sg13g2_fill_2 FILLER_20_79 ();
 sg13g2_decap_8 FILLER_20_96 ();
 sg13g2_fill_2 FILLER_20_103 ();
 sg13g2_fill_2 FILLER_20_110 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_decap_4 FILLER_20_118 ();
 sg13g2_fill_2 FILLER_20_122 ();
 sg13g2_fill_1 FILLER_20_174 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_decap_8 FILLER_20_226 ();
 sg13g2_decap_8 FILLER_20_233 ();
 sg13g2_fill_2 FILLER_20_240 ();
 sg13g2_fill_1 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_248 ();
 sg13g2_fill_2 FILLER_20_255 ();
 sg13g2_fill_1 FILLER_20_257 ();
 sg13g2_fill_1 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_274 ();
 sg13g2_decap_8 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_297 ();
 sg13g2_decap_8 FILLER_20_304 ();
 sg13g2_decap_8 FILLER_20_311 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_8 FILLER_20_325 ();
 sg13g2_decap_8 FILLER_20_332 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_fill_2 FILLER_20_397 ();
 sg13g2_fill_1 FILLER_20_399 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_38 ();
 sg13g2_fill_2 FILLER_21_42 ();
 sg13g2_decap_4 FILLER_21_52 ();
 sg13g2_fill_1 FILLER_21_56 ();
 sg13g2_fill_2 FILLER_21_62 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_4 FILLER_21_112 ();
 sg13g2_fill_2 FILLER_21_116 ();
 sg13g2_decap_8 FILLER_21_125 ();
 sg13g2_fill_2 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_134 ();
 sg13g2_fill_2 FILLER_21_174 ();
 sg13g2_fill_2 FILLER_21_191 ();
 sg13g2_fill_1 FILLER_21_193 ();
 sg13g2_decap_8 FILLER_21_204 ();
 sg13g2_fill_2 FILLER_21_218 ();
 sg13g2_decap_4 FILLER_21_240 ();
 sg13g2_fill_2 FILLER_21_261 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_fill_2 FILLER_21_276 ();
 sg13g2_decap_8 FILLER_21_325 ();
 sg13g2_fill_1 FILLER_21_332 ();
 sg13g2_fill_2 FILLER_21_338 ();
 sg13g2_decap_4 FILLER_21_344 ();
 sg13g2_fill_1 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_fill_2 FILLER_21_379 ();
 sg13g2_fill_1 FILLER_21_381 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_31 ();
 sg13g2_fill_1 FILLER_22_33 ();
 sg13g2_fill_1 FILLER_22_39 ();
 sg13g2_fill_1 FILLER_22_54 ();
 sg13g2_fill_1 FILLER_22_59 ();
 sg13g2_decap_4 FILLER_22_65 ();
 sg13g2_decap_8 FILLER_22_81 ();
 sg13g2_fill_1 FILLER_22_93 ();
 sg13g2_fill_1 FILLER_22_99 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_fill_2 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_121 ();
 sg13g2_decap_8 FILLER_22_128 ();
 sg13g2_decap_4 FILLER_22_135 ();
 sg13g2_fill_1 FILLER_22_139 ();
 sg13g2_fill_2 FILLER_22_160 ();
 sg13g2_fill_1 FILLER_22_162 ();
 sg13g2_decap_8 FILLER_22_181 ();
 sg13g2_fill_2 FILLER_22_188 ();
 sg13g2_decap_4 FILLER_22_203 ();
 sg13g2_fill_1 FILLER_22_207 ();
 sg13g2_decap_4 FILLER_22_217 ();
 sg13g2_fill_1 FILLER_22_238 ();
 sg13g2_decap_4 FILLER_22_244 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_fill_2 FILLER_22_266 ();
 sg13g2_decap_4 FILLER_22_273 ();
 sg13g2_fill_2 FILLER_22_277 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_fill_1 FILLER_22_348 ();
 sg13g2_fill_1 FILLER_22_364 ();
 sg13g2_decap_4 FILLER_22_385 ();
 sg13g2_fill_2 FILLER_22_389 ();
 sg13g2_fill_2 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_15 ();
 sg13g2_fill_1 FILLER_23_75 ();
 sg13g2_fill_1 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_97 ();
 sg13g2_fill_1 FILLER_23_99 ();
 sg13g2_fill_1 FILLER_23_111 ();
 sg13g2_fill_2 FILLER_23_122 ();
 sg13g2_fill_1 FILLER_23_124 ();
 sg13g2_decap_8 FILLER_23_138 ();
 sg13g2_fill_2 FILLER_23_145 ();
 sg13g2_fill_1 FILLER_23_147 ();
 sg13g2_fill_2 FILLER_23_159 ();
 sg13g2_fill_1 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_172 ();
 sg13g2_decap_4 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_191 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_decap_4 FILLER_23_208 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_fill_1 FILLER_23_220 ();
 sg13g2_fill_1 FILLER_23_233 ();
 sg13g2_fill_2 FILLER_23_243 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_fill_1 FILLER_23_253 ();
 sg13g2_decap_8 FILLER_23_269 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_278 ();
 sg13g2_fill_1 FILLER_23_290 ();
 sg13g2_fill_2 FILLER_23_313 ();
 sg13g2_fill_1 FILLER_23_315 ();
 sg13g2_fill_2 FILLER_23_336 ();
 sg13g2_fill_1 FILLER_23_338 ();
 sg13g2_fill_2 FILLER_23_356 ();
 sg13g2_fill_1 FILLER_23_358 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_fill_1 FILLER_24_35 ();
 sg13g2_fill_2 FILLER_24_60 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_decap_4 FILLER_24_114 ();
 sg13g2_decap_8 FILLER_24_145 ();
 sg13g2_decap_4 FILLER_24_152 ();
 sg13g2_fill_2 FILLER_24_156 ();
 sg13g2_decap_8 FILLER_24_166 ();
 sg13g2_decap_4 FILLER_24_173 ();
 sg13g2_fill_2 FILLER_24_177 ();
 sg13g2_decap_4 FILLER_24_188 ();
 sg13g2_fill_2 FILLER_24_249 ();
 sg13g2_fill_1 FILLER_24_280 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_fill_2 FILLER_24_322 ();
 sg13g2_decap_4 FILLER_24_328 ();
 sg13g2_decap_4 FILLER_24_377 ();
 sg13g2_fill_2 FILLER_24_381 ();
 sg13g2_fill_2 FILLER_25_79 ();
 sg13g2_fill_1 FILLER_25_81 ();
 sg13g2_fill_2 FILLER_25_87 ();
 sg13g2_decap_8 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_162 ();
 sg13g2_fill_2 FILLER_25_171 ();
 sg13g2_fill_2 FILLER_25_208 ();
 sg13g2_fill_2 FILLER_25_248 ();
 sg13g2_decap_8 FILLER_25_254 ();
 sg13g2_fill_2 FILLER_25_261 ();
 sg13g2_decap_8 FILLER_25_268 ();
 sg13g2_fill_2 FILLER_25_275 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_fill_2 FILLER_25_309 ();
 sg13g2_decap_8 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_decap_8 FILLER_25_360 ();
 sg13g2_decap_8 FILLER_25_367 ();
 sg13g2_fill_1 FILLER_25_374 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_58 ();
 sg13g2_decap_4 FILLER_26_82 ();
 sg13g2_decap_8 FILLER_26_90 ();
 sg13g2_decap_4 FILLER_26_97 ();
 sg13g2_fill_2 FILLER_26_101 ();
 sg13g2_decap_4 FILLER_26_108 ();
 sg13g2_fill_2 FILLER_26_117 ();
 sg13g2_fill_1 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_124 ();
 sg13g2_decap_4 FILLER_26_135 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_176 ();
 sg13g2_fill_1 FILLER_26_183 ();
 sg13g2_fill_2 FILLER_26_203 ();
 sg13g2_fill_2 FILLER_26_257 ();
 sg13g2_fill_1 FILLER_26_259 ();
 sg13g2_fill_1 FILLER_26_265 ();
 sg13g2_decap_8 FILLER_26_271 ();
 sg13g2_decap_4 FILLER_26_278 ();
 sg13g2_fill_1 FILLER_26_282 ();
 sg13g2_decap_4 FILLER_26_300 ();
 sg13g2_fill_1 FILLER_26_309 ();
 sg13g2_decap_8 FILLER_26_318 ();
 sg13g2_decap_8 FILLER_26_325 ();
 sg13g2_fill_1 FILLER_26_346 ();
 sg13g2_decap_4 FILLER_26_356 ();
 sg13g2_fill_2 FILLER_26_360 ();
 sg13g2_fill_2 FILLER_26_390 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_1 FILLER_27_35 ();
 sg13g2_fill_2 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_95 ();
 sg13g2_decap_8 FILLER_27_102 ();
 sg13g2_decap_8 FILLER_27_109 ();
 sg13g2_decap_8 FILLER_27_116 ();
 sg13g2_decap_4 FILLER_27_123 ();
 sg13g2_fill_2 FILLER_27_136 ();
 sg13g2_fill_2 FILLER_27_154 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_209 ();
 sg13g2_fill_2 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_248 ();
 sg13g2_fill_1 FILLER_27_258 ();
 sg13g2_decap_4 FILLER_27_350 ();
 sg13g2_fill_2 FILLER_27_354 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_4 FILLER_27_391 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_31 ();
 sg13g2_fill_2 FILLER_28_69 ();
 sg13g2_fill_1 FILLER_28_71 ();
 sg13g2_fill_1 FILLER_28_102 ();
 sg13g2_decap_4 FILLER_28_108 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_decap_4 FILLER_28_128 ();
 sg13g2_decap_4 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_160 ();
 sg13g2_fill_2 FILLER_28_175 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_decap_8 FILLER_28_187 ();
 sg13g2_fill_2 FILLER_28_194 ();
 sg13g2_fill_1 FILLER_28_196 ();
 sg13g2_decap_4 FILLER_28_206 ();
 sg13g2_fill_1 FILLER_28_210 ();
 sg13g2_fill_2 FILLER_28_216 ();
 sg13g2_decap_8 FILLER_28_222 ();
 sg13g2_decap_8 FILLER_28_233 ();
 sg13g2_decap_8 FILLER_28_244 ();
 sg13g2_decap_8 FILLER_28_251 ();
 sg13g2_fill_2 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_decap_4 FILLER_28_266 ();
 sg13g2_fill_1 FILLER_28_287 ();
 sg13g2_fill_1 FILLER_28_311 ();
 sg13g2_decap_4 FILLER_28_351 ();
 sg13g2_decap_8 FILLER_28_363 ();
 sg13g2_decap_8 FILLER_28_370 ();
 sg13g2_decap_8 FILLER_28_377 ();
 sg13g2_fill_2 FILLER_28_384 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_29_16 ();
 sg13g2_fill_2 FILLER_29_46 ();
 sg13g2_decap_4 FILLER_29_83 ();
 sg13g2_fill_2 FILLER_29_122 ();
 sg13g2_fill_1 FILLER_29_124 ();
 sg13g2_fill_2 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_153 ();
 sg13g2_decap_8 FILLER_29_167 ();
 sg13g2_fill_1 FILLER_29_218 ();
 sg13g2_fill_1 FILLER_29_232 ();
 sg13g2_fill_2 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_fill_1 FILLER_29_333 ();
 sg13g2_decap_8 FILLER_29_375 ();
 sg13g2_decap_4 FILLER_29_382 ();
 sg13g2_fill_1 FILLER_29_386 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_114 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_fill_2 FILLER_30_252 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_fill_2 FILLER_30_270 ();
 sg13g2_fill_1 FILLER_30_272 ();
 sg13g2_fill_1 FILLER_30_333 ();
 sg13g2_fill_1 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_366 ();
 sg13g2_decap_4 FILLER_30_373 ();
 sg13g2_fill_1 FILLER_30_377 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_decap_8 FILLER_31_64 ();
 sg13g2_decap_4 FILLER_31_71 ();
 sg13g2_fill_2 FILLER_31_80 ();
 sg13g2_fill_1 FILLER_31_82 ();
 sg13g2_fill_1 FILLER_31_88 ();
 sg13g2_fill_2 FILLER_31_99 ();
 sg13g2_fill_1 FILLER_31_106 ();
 sg13g2_fill_1 FILLER_31_111 ();
 sg13g2_decap_4 FILLER_31_158 ();
 sg13g2_fill_1 FILLER_31_162 ();
 sg13g2_fill_1 FILLER_31_203 ();
 sg13g2_fill_1 FILLER_31_264 ();
 sg13g2_fill_2 FILLER_31_284 ();
 sg13g2_fill_1 FILLER_31_322 ();
 sg13g2_fill_2 FILLER_31_329 ();
 sg13g2_fill_1 FILLER_31_356 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_2 FILLER_32_31 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_68 ();
 sg13g2_fill_1 FILLER_32_89 ();
 sg13g2_fill_2 FILLER_32_99 ();
 sg13g2_fill_1 FILLER_32_101 ();
 sg13g2_decap_8 FILLER_32_107 ();
 sg13g2_decap_4 FILLER_32_114 ();
 sg13g2_fill_1 FILLER_32_118 ();
 sg13g2_decap_8 FILLER_32_123 ();
 sg13g2_fill_2 FILLER_32_130 ();
 sg13g2_fill_1 FILLER_32_132 ();
 sg13g2_fill_1 FILLER_32_146 ();
 sg13g2_decap_4 FILLER_32_154 ();
 sg13g2_fill_1 FILLER_32_158 ();
 sg13g2_decap_8 FILLER_32_163 ();
 sg13g2_fill_2 FILLER_32_175 ();
 sg13g2_fill_1 FILLER_32_189 ();
 sg13g2_fill_1 FILLER_32_202 ();
 sg13g2_fill_2 FILLER_32_215 ();
 sg13g2_decap_8 FILLER_32_230 ();
 sg13g2_fill_1 FILLER_32_237 ();
 sg13g2_decap_8 FILLER_32_243 ();
 sg13g2_fill_2 FILLER_32_250 ();
 sg13g2_decap_8 FILLER_32_257 ();
 sg13g2_fill_2 FILLER_32_296 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_4 FILLER_32_357 ();
 sg13g2_fill_2 FILLER_32_372 ();
 sg13g2_fill_1 FILLER_32_379 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_fill_1 FILLER_33_51 ();
 sg13g2_fill_1 FILLER_33_109 ();
 sg13g2_decap_4 FILLER_33_127 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_fill_2 FILLER_33_152 ();
 sg13g2_fill_2 FILLER_33_159 ();
 sg13g2_fill_2 FILLER_33_187 ();
 sg13g2_fill_1 FILLER_33_189 ();
 sg13g2_fill_2 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_399 ();
 sg13g2_fill_1 FILLER_34_50 ();
 sg13g2_fill_1 FILLER_34_82 ();
 sg13g2_fill_2 FILLER_34_127 ();
 sg13g2_fill_2 FILLER_34_149 ();
 sg13g2_fill_1 FILLER_34_151 ();
 sg13g2_fill_2 FILLER_34_158 ();
 sg13g2_fill_1 FILLER_34_160 ();
 sg13g2_fill_2 FILLER_34_171 ();
 sg13g2_fill_1 FILLER_34_173 ();
 sg13g2_fill_2 FILLER_34_189 ();
 sg13g2_fill_2 FILLER_34_255 ();
 sg13g2_fill_2 FILLER_34_310 ();
 sg13g2_decap_8 FILLER_34_351 ();
 sg13g2_decap_4 FILLER_34_358 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_fill_2 FILLER_34_371 ();
 sg13g2_fill_1 FILLER_34_373 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_fill_2 FILLER_35_77 ();
 sg13g2_fill_1 FILLER_35_79 ();
 sg13g2_decap_8 FILLER_35_123 ();
 sg13g2_decap_4 FILLER_35_130 ();
 sg13g2_fill_1 FILLER_35_134 ();
 sg13g2_fill_2 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_156 ();
 sg13g2_fill_2 FILLER_35_165 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_fill_2 FILLER_35_173 ();
 sg13g2_fill_1 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_194 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_decap_4 FILLER_35_206 ();
 sg13g2_fill_2 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_decap_4 FILLER_35_236 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_fill_1 FILLER_35_280 ();
 sg13g2_fill_1 FILLER_35_303 ();
 sg13g2_fill_2 FILLER_35_369 ();
 sg13g2_fill_2 FILLER_35_379 ();
 sg13g2_fill_1 FILLER_35_381 ();
 sg13g2_decap_4 FILLER_36_38 ();
 sg13g2_fill_2 FILLER_36_72 ();
 sg13g2_fill_1 FILLER_36_78 ();
 sg13g2_decap_8 FILLER_36_114 ();
 sg13g2_decap_4 FILLER_36_121 ();
 sg13g2_decap_8 FILLER_36_132 ();
 sg13g2_decap_8 FILLER_36_139 ();
 sg13g2_decap_8 FILLER_36_146 ();
 sg13g2_decap_8 FILLER_36_153 ();
 sg13g2_fill_2 FILLER_36_160 ();
 sg13g2_fill_1 FILLER_36_162 ();
 sg13g2_decap_4 FILLER_36_168 ();
 sg13g2_fill_2 FILLER_36_172 ();
 sg13g2_decap_8 FILLER_36_178 ();
 sg13g2_decap_8 FILLER_36_185 ();
 sg13g2_decap_8 FILLER_36_192 ();
 sg13g2_fill_2 FILLER_36_199 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_decap_8 FILLER_36_206 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_decap_8 FILLER_36_220 ();
 sg13g2_decap_8 FILLER_36_227 ();
 sg13g2_decap_8 FILLER_36_234 ();
 sg13g2_decap_4 FILLER_36_241 ();
 sg13g2_fill_1 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_251 ();
 sg13g2_fill_2 FILLER_36_258 ();
 sg13g2_fill_1 FILLER_36_260 ();
 sg13g2_fill_2 FILLER_36_267 ();
 sg13g2_decap_4 FILLER_36_273 ();
 sg13g2_fill_1 FILLER_36_277 ();
 sg13g2_fill_2 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_304 ();
 sg13g2_fill_1 FILLER_36_336 ();
 sg13g2_fill_2 FILLER_36_346 ();
 sg13g2_fill_2 FILLER_36_357 ();
 sg13g2_fill_1 FILLER_36_359 ();
 sg13g2_fill_2 FILLER_36_380 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_fill_1 FILLER_37_26 ();
 sg13g2_fill_1 FILLER_37_75 ();
 sg13g2_fill_2 FILLER_37_98 ();
 sg13g2_decap_4 FILLER_37_104 ();
 sg13g2_decap_4 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_145 ();
 sg13g2_decap_4 FILLER_37_158 ();
 sg13g2_fill_2 FILLER_37_180 ();
 sg13g2_fill_1 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_201 ();
 sg13g2_decap_8 FILLER_37_208 ();
 sg13g2_fill_2 FILLER_37_215 ();
 sg13g2_fill_1 FILLER_37_217 ();
 sg13g2_decap_4 FILLER_37_222 ();
 sg13g2_fill_2 FILLER_37_226 ();
 sg13g2_decap_8 FILLER_37_233 ();
 sg13g2_decap_8 FILLER_37_240 ();
 sg13g2_decap_8 FILLER_37_247 ();
 sg13g2_fill_1 FILLER_37_254 ();
 sg13g2_decap_8 FILLER_37_260 ();
 sg13g2_decap_8 FILLER_37_267 ();
 sg13g2_decap_8 FILLER_37_274 ();
 sg13g2_decap_8 FILLER_37_281 ();
 sg13g2_fill_1 FILLER_37_288 ();
 sg13g2_fill_1 FILLER_37_310 ();
 sg13g2_decap_8 FILLER_37_346 ();
 sg13g2_decap_4 FILLER_37_353 ();
 sg13g2_fill_1 FILLER_37_357 ();
 sg13g2_fill_2 FILLER_37_362 ();
 sg13g2_fill_1 FILLER_37_364 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_19 ();
 sg13g2_decap_4 FILLER_38_69 ();
 sg13g2_fill_2 FILLER_38_90 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_fill_2 FILLER_38_159 ();
 sg13g2_fill_2 FILLER_38_200 ();
 sg13g2_fill_1 FILLER_38_202 ();
 sg13g2_fill_2 FILLER_38_216 ();
 sg13g2_fill_2 FILLER_38_223 ();
 sg13g2_decap_4 FILLER_38_242 ();
 sg13g2_fill_1 FILLER_38_252 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_decap_8 FILLER_38_281 ();
 sg13g2_fill_1 FILLER_38_288 ();
 sg13g2_fill_2 FILLER_38_340 ();
 sg13g2_decap_4 FILLER_38_370 ();
 sg13g2_fill_2 FILLER_38_374 ();
 sg13g2_decap_4 FILLER_38_394 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_38 ();
 sg13g2_decap_4 FILLER_39_49 ();
 sg13g2_fill_2 FILLER_39_97 ();
 sg13g2_fill_1 FILLER_39_99 ();
 sg13g2_decap_8 FILLER_39_108 ();
 sg13g2_decap_8 FILLER_39_115 ();
 sg13g2_decap_4 FILLER_39_122 ();
 sg13g2_fill_1 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_141 ();
 sg13g2_fill_2 FILLER_39_153 ();
 sg13g2_fill_1 FILLER_39_155 ();
 sg13g2_fill_2 FILLER_39_161 ();
 sg13g2_fill_1 FILLER_39_167 ();
 sg13g2_fill_2 FILLER_39_176 ();
 sg13g2_fill_1 FILLER_39_178 ();
 sg13g2_fill_2 FILLER_39_184 ();
 sg13g2_fill_1 FILLER_39_186 ();
 sg13g2_fill_2 FILLER_39_197 ();
 sg13g2_fill_1 FILLER_39_220 ();
 sg13g2_fill_2 FILLER_39_302 ();
 sg13g2_decap_4 FILLER_39_328 ();
 sg13g2_fill_2 FILLER_39_345 ();
 sg13g2_fill_1 FILLER_39_347 ();
 sg13g2_fill_2 FILLER_39_356 ();
 sg13g2_decap_4 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_9 ();
 sg13g2_fill_2 FILLER_40_13 ();
 sg13g2_decap_8 FILLER_40_19 ();
 sg13g2_fill_2 FILLER_40_26 ();
 sg13g2_decap_8 FILLER_40_37 ();
 sg13g2_decap_4 FILLER_40_44 ();
 sg13g2_fill_1 FILLER_40_48 ();
 sg13g2_fill_1 FILLER_40_75 ();
 sg13g2_fill_2 FILLER_40_81 ();
 sg13g2_fill_1 FILLER_40_83 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_4 FILLER_40_140 ();
 sg13g2_fill_2 FILLER_40_144 ();
 sg13g2_decap_8 FILLER_40_158 ();
 sg13g2_decap_8 FILLER_40_165 ();
 sg13g2_decap_8 FILLER_40_172 ();
 sg13g2_decap_4 FILLER_40_179 ();
 sg13g2_fill_2 FILLER_40_183 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_fill_1 FILLER_40_199 ();
 sg13g2_fill_1 FILLER_40_226 ();
 sg13g2_fill_2 FILLER_40_245 ();
 sg13g2_fill_2 FILLER_40_301 ();
 sg13g2_fill_2 FILLER_40_320 ();
 sg13g2_fill_2 FILLER_40_337 ();
 sg13g2_fill_1 FILLER_40_339 ();
 sg13g2_fill_2 FILLER_40_349 ();
 sg13g2_fill_2 FILLER_40_367 ();
 sg13g2_fill_1 FILLER_40_382 ();
 sg13g2_fill_1 FILLER_40_396 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_fill_2 FILLER_41_39 ();
 sg13g2_fill_1 FILLER_41_59 ();
 sg13g2_decap_4 FILLER_41_71 ();
 sg13g2_fill_1 FILLER_41_75 ();
 sg13g2_decap_4 FILLER_41_113 ();
 sg13g2_fill_1 FILLER_41_117 ();
 sg13g2_decap_8 FILLER_41_127 ();
 sg13g2_decap_8 FILLER_41_134 ();
 sg13g2_fill_2 FILLER_41_141 ();
 sg13g2_fill_1 FILLER_41_143 ();
 sg13g2_fill_2 FILLER_41_149 ();
 sg13g2_fill_2 FILLER_41_156 ();
 sg13g2_fill_2 FILLER_41_163 ();
 sg13g2_fill_1 FILLER_41_165 ();
 sg13g2_decap_8 FILLER_41_171 ();
 sg13g2_decap_4 FILLER_41_178 ();
 sg13g2_fill_2 FILLER_41_193 ();
 sg13g2_fill_1 FILLER_41_195 ();
 sg13g2_decap_8 FILLER_41_214 ();
 sg13g2_decap_4 FILLER_41_221 ();
 sg13g2_fill_1 FILLER_41_225 ();
 sg13g2_decap_4 FILLER_41_230 ();
 sg13g2_fill_2 FILLER_41_234 ();
 sg13g2_fill_2 FILLER_41_280 ();
 sg13g2_fill_1 FILLER_41_282 ();
 sg13g2_fill_2 FILLER_41_294 ();
 sg13g2_fill_2 FILLER_41_312 ();
 sg13g2_fill_1 FILLER_41_314 ();
 sg13g2_fill_2 FILLER_41_332 ();
 sg13g2_decap_4 FILLER_41_352 ();
 sg13g2_decap_8 FILLER_41_365 ();
 sg13g2_fill_1 FILLER_41_372 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_2 ();
 sg13g2_fill_1 FILLER_42_34 ();
 sg13g2_fill_2 FILLER_42_112 ();
 sg13g2_decap_4 FILLER_42_134 ();
 sg13g2_fill_1 FILLER_42_138 ();
 sg13g2_decap_8 FILLER_42_178 ();
 sg13g2_decap_8 FILLER_42_185 ();
 sg13g2_decap_4 FILLER_42_218 ();
 sg13g2_fill_2 FILLER_42_222 ();
 sg13g2_fill_1 FILLER_42_277 ();
 sg13g2_fill_2 FILLER_42_298 ();
 sg13g2_fill_1 FILLER_42_300 ();
 sg13g2_fill_1 FILLER_42_394 ();
 sg13g2_fill_2 FILLER_43_14 ();
 sg13g2_fill_2 FILLER_43_21 ();
 sg13g2_fill_2 FILLER_43_58 ();
 sg13g2_fill_1 FILLER_43_86 ();
 sg13g2_fill_2 FILLER_43_101 ();
 sg13g2_fill_1 FILLER_43_103 ();
 sg13g2_decap_8 FILLER_43_107 ();
 sg13g2_decap_8 FILLER_43_142 ();
 sg13g2_fill_2 FILLER_43_149 ();
 sg13g2_fill_1 FILLER_43_151 ();
 sg13g2_fill_2 FILLER_43_169 ();
 sg13g2_decap_8 FILLER_43_185 ();
 sg13g2_decap_4 FILLER_43_230 ();
 sg13g2_fill_2 FILLER_43_291 ();
 sg13g2_fill_2 FILLER_43_319 ();
 sg13g2_fill_1 FILLER_43_321 ();
 sg13g2_fill_1 FILLER_43_335 ();
 sg13g2_fill_1 FILLER_44_32 ();
 sg13g2_fill_2 FILLER_44_56 ();
 sg13g2_fill_1 FILLER_44_58 ();
 sg13g2_fill_1 FILLER_44_85 ();
 sg13g2_fill_1 FILLER_44_95 ();
 sg13g2_decap_4 FILLER_44_109 ();
 sg13g2_fill_2 FILLER_44_118 ();
 sg13g2_fill_2 FILLER_44_128 ();
 sg13g2_fill_1 FILLER_44_130 ();
 sg13g2_decap_8 FILLER_44_148 ();
 sg13g2_fill_2 FILLER_44_155 ();
 sg13g2_decap_8 FILLER_44_165 ();
 sg13g2_fill_1 FILLER_44_196 ();
 sg13g2_fill_1 FILLER_44_215 ();
 sg13g2_fill_2 FILLER_44_225 ();
 sg13g2_fill_2 FILLER_44_278 ();
 sg13g2_fill_2 FILLER_44_291 ();
 sg13g2_fill_1 FILLER_44_293 ();
 sg13g2_decap_4 FILLER_44_324 ();
 sg13g2_fill_1 FILLER_44_334 ();
 sg13g2_fill_2 FILLER_44_353 ();
 sg13g2_fill_1 FILLER_44_355 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_2 ();
 sg13g2_fill_2 FILLER_45_17 ();
 sg13g2_fill_2 FILLER_45_46 ();
 sg13g2_fill_1 FILLER_45_99 ();
 sg13g2_fill_1 FILLER_45_113 ();
 sg13g2_decap_4 FILLER_45_127 ();
 sg13g2_fill_2 FILLER_45_139 ();
 sg13g2_decap_8 FILLER_45_146 ();
 sg13g2_decap_8 FILLER_45_153 ();
 sg13g2_fill_2 FILLER_45_160 ();
 sg13g2_fill_1 FILLER_45_162 ();
 sg13g2_fill_2 FILLER_45_178 ();
 sg13g2_fill_1 FILLER_45_180 ();
 sg13g2_fill_1 FILLER_45_188 ();
 sg13g2_fill_1 FILLER_45_194 ();
 sg13g2_fill_1 FILLER_45_202 ();
 sg13g2_fill_1 FILLER_45_213 ();
 sg13g2_fill_1 FILLER_45_235 ();
 sg13g2_decap_4 FILLER_45_274 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_fill_2 FILLER_45_301 ();
 sg13g2_fill_1 FILLER_45_303 ();
 sg13g2_fill_2 FILLER_45_313 ();
 sg13g2_fill_1 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_342 ();
 sg13g2_decap_8 FILLER_45_349 ();
 sg13g2_fill_1 FILLER_45_382 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_14 ();
 sg13g2_fill_2 FILLER_46_65 ();
 sg13g2_fill_1 FILLER_46_67 ();
 sg13g2_fill_2 FILLER_46_77 ();
 sg13g2_fill_1 FILLER_46_112 ();
 sg13g2_fill_1 FILLER_46_127 ();
 sg13g2_fill_2 FILLER_46_167 ();
 sg13g2_decap_4 FILLER_46_176 ();
 sg13g2_decap_8 FILLER_46_195 ();
 sg13g2_decap_4 FILLER_46_212 ();
 sg13g2_fill_2 FILLER_46_216 ();
 sg13g2_fill_2 FILLER_46_227 ();
 sg13g2_fill_2 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_262 ();
 sg13g2_fill_2 FILLER_46_285 ();
 sg13g2_fill_1 FILLER_46_287 ();
 sg13g2_fill_2 FILLER_46_309 ();
 sg13g2_fill_1 FILLER_46_349 ();
 sg13g2_fill_2 FILLER_47_4 ();
 sg13g2_fill_2 FILLER_47_25 ();
 sg13g2_fill_1 FILLER_47_27 ();
 sg13g2_fill_1 FILLER_47_71 ();
 sg13g2_decap_8 FILLER_47_109 ();
 sg13g2_decap_8 FILLER_47_116 ();
 sg13g2_decap_8 FILLER_47_123 ();
 sg13g2_decap_8 FILLER_47_130 ();
 sg13g2_fill_2 FILLER_47_137 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_4 FILLER_47_166 ();
 sg13g2_fill_2 FILLER_47_170 ();
 sg13g2_fill_1 FILLER_47_177 ();
 sg13g2_fill_1 FILLER_47_192 ();
 sg13g2_decap_4 FILLER_47_206 ();
 sg13g2_fill_2 FILLER_47_210 ();
 sg13g2_fill_2 FILLER_47_231 ();
 sg13g2_fill_1 FILLER_47_233 ();
 sg13g2_decap_8 FILLER_47_283 ();
 sg13g2_fill_1 FILLER_47_290 ();
 sg13g2_fill_2 FILLER_47_329 ();
 sg13g2_fill_2 FILLER_47_339 ();
 sg13g2_fill_1 FILLER_47_355 ();
 sg13g2_fill_2 FILLER_47_373 ();
 sg13g2_fill_2 FILLER_47_383 ();
 sg13g2_fill_1 FILLER_47_385 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_2 ();
 sg13g2_fill_2 FILLER_48_81 ();
 sg13g2_fill_1 FILLER_48_83 ();
 sg13g2_fill_1 FILLER_48_98 ();
 sg13g2_fill_2 FILLER_48_108 ();
 sg13g2_fill_1 FILLER_48_110 ();
 sg13g2_decap_4 FILLER_48_119 ();
 sg13g2_fill_1 FILLER_48_123 ();
 sg13g2_decap_4 FILLER_48_132 ();
 sg13g2_fill_2 FILLER_48_136 ();
 sg13g2_fill_2 FILLER_48_143 ();
 sg13g2_fill_1 FILLER_48_145 ();
 sg13g2_fill_1 FILLER_48_155 ();
 sg13g2_fill_2 FILLER_48_164 ();
 sg13g2_fill_1 FILLER_48_166 ();
 sg13g2_fill_2 FILLER_48_200 ();
 sg13g2_fill_1 FILLER_48_202 ();
 sg13g2_fill_2 FILLER_48_215 ();
 sg13g2_fill_1 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_262 ();
 sg13g2_fill_1 FILLER_48_269 ();
 sg13g2_fill_1 FILLER_48_279 ();
 sg13g2_fill_2 FILLER_48_298 ();
 sg13g2_fill_1 FILLER_48_300 ();
 sg13g2_fill_2 FILLER_48_321 ();
 sg13g2_fill_1 FILLER_48_323 ();
 sg13g2_fill_2 FILLER_48_384 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_16 ();
 sg13g2_fill_2 FILLER_49_92 ();
 sg13g2_fill_1 FILLER_49_104 ();
 sg13g2_decap_8 FILLER_49_124 ();
 sg13g2_decap_8 FILLER_49_131 ();
 sg13g2_fill_2 FILLER_49_146 ();
 sg13g2_fill_1 FILLER_49_148 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_fill_1 FILLER_49_166 ();
 sg13g2_decap_8 FILLER_49_172 ();
 sg13g2_decap_4 FILLER_49_179 ();
 sg13g2_fill_1 FILLER_49_183 ();
 sg13g2_fill_1 FILLER_49_231 ();
 sg13g2_fill_2 FILLER_49_242 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_fill_2 FILLER_49_259 ();
 sg13g2_fill_1 FILLER_49_261 ();
 sg13g2_decap_4 FILLER_49_271 ();
 sg13g2_fill_2 FILLER_49_275 ();
 sg13g2_fill_2 FILLER_49_285 ();
 sg13g2_fill_1 FILLER_49_287 ();
 sg13g2_fill_2 FILLER_49_303 ();
 sg13g2_fill_1 FILLER_49_305 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_9 ();
 sg13g2_decap_8 FILLER_50_15 ();
 sg13g2_decap_8 FILLER_50_22 ();
 sg13g2_fill_1 FILLER_50_29 ();
 sg13g2_decap_4 FILLER_50_86 ();
 sg13g2_fill_1 FILLER_50_111 ();
 sg13g2_decap_8 FILLER_50_135 ();
 sg13g2_decap_4 FILLER_50_142 ();
 sg13g2_decap_8 FILLER_50_151 ();
 sg13g2_decap_4 FILLER_50_168 ();
 sg13g2_decap_8 FILLER_50_178 ();
 sg13g2_decap_8 FILLER_50_185 ();
 sg13g2_decap_8 FILLER_50_192 ();
 sg13g2_fill_2 FILLER_50_199 ();
 sg13g2_decap_8 FILLER_50_211 ();
 sg13g2_decap_8 FILLER_50_218 ();
 sg13g2_decap_8 FILLER_50_239 ();
 sg13g2_decap_8 FILLER_50_246 ();
 sg13g2_fill_1 FILLER_50_284 ();
 sg13g2_fill_2 FILLER_50_297 ();
 sg13g2_fill_1 FILLER_50_299 ();
 sg13g2_fill_2 FILLER_50_306 ();
 sg13g2_fill_1 FILLER_50_362 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_4 ();
 sg13g2_fill_2 FILLER_51_29 ();
 sg13g2_fill_1 FILLER_51_62 ();
 sg13g2_decap_8 FILLER_51_68 ();
 sg13g2_decap_8 FILLER_51_75 ();
 sg13g2_decap_8 FILLER_51_82 ();
 sg13g2_fill_2 FILLER_51_104 ();
 sg13g2_decap_8 FILLER_51_111 ();
 sg13g2_fill_2 FILLER_51_118 ();
 sg13g2_fill_2 FILLER_51_130 ();
 sg13g2_fill_1 FILLER_51_132 ();
 sg13g2_decap_4 FILLER_51_147 ();
 sg13g2_fill_1 FILLER_51_156 ();
 sg13g2_fill_2 FILLER_51_161 ();
 sg13g2_fill_1 FILLER_51_163 ();
 sg13g2_fill_2 FILLER_51_168 ();
 sg13g2_fill_1 FILLER_51_170 ();
 sg13g2_fill_2 FILLER_51_180 ();
 sg13g2_fill_1 FILLER_51_182 ();
 sg13g2_decap_8 FILLER_51_198 ();
 sg13g2_fill_2 FILLER_51_205 ();
 sg13g2_fill_1 FILLER_51_207 ();
 sg13g2_decap_8 FILLER_51_213 ();
 sg13g2_fill_2 FILLER_51_220 ();
 sg13g2_fill_1 FILLER_51_222 ();
 sg13g2_decap_4 FILLER_51_226 ();
 sg13g2_fill_1 FILLER_51_230 ();
 sg13g2_decap_8 FILLER_51_235 ();
 sg13g2_fill_2 FILLER_51_242 ();
 sg13g2_decap_8 FILLER_51_262 ();
 sg13g2_fill_1 FILLER_51_269 ();
 sg13g2_fill_2 FILLER_51_303 ();
 sg13g2_fill_2 FILLER_51_367 ();
 sg13g2_decap_4 FILLER_52_0 ();
 sg13g2_decap_4 FILLER_52_24 ();
 sg13g2_fill_1 FILLER_52_44 ();
 sg13g2_decap_4 FILLER_52_68 ();
 sg13g2_fill_2 FILLER_52_72 ();
 sg13g2_fill_1 FILLER_52_93 ();
 sg13g2_fill_1 FILLER_52_102 ();
 sg13g2_fill_1 FILLER_52_110 ();
 sg13g2_decap_8 FILLER_52_118 ();
 sg13g2_fill_1 FILLER_52_125 ();
 sg13g2_fill_2 FILLER_52_152 ();
 sg13g2_fill_1 FILLER_52_194 ();
 sg13g2_decap_4 FILLER_52_212 ();
 sg13g2_fill_2 FILLER_52_273 ();
 sg13g2_fill_1 FILLER_52_275 ();
 sg13g2_fill_2 FILLER_52_282 ();
 sg13g2_fill_1 FILLER_52_284 ();
 sg13g2_fill_2 FILLER_52_291 ();
 sg13g2_fill_1 FILLER_52_293 ();
 sg13g2_fill_1 FILLER_52_310 ();
 sg13g2_fill_1 FILLER_52_342 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_4 FILLER_53_7 ();
 sg13g2_fill_2 FILLER_53_25 ();
 sg13g2_decap_4 FILLER_53_32 ();
 sg13g2_fill_2 FILLER_53_78 ();
 sg13g2_fill_2 FILLER_53_93 ();
 sg13g2_fill_1 FILLER_53_95 ();
 sg13g2_fill_2 FILLER_53_106 ();
 sg13g2_decap_8 FILLER_53_115 ();
 sg13g2_decap_4 FILLER_53_122 ();
 sg13g2_fill_2 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_136 ();
 sg13g2_decap_8 FILLER_53_143 ();
 sg13g2_decap_8 FILLER_53_150 ();
 sg13g2_fill_2 FILLER_53_157 ();
 sg13g2_decap_8 FILLER_53_166 ();
 sg13g2_fill_2 FILLER_53_189 ();
 sg13g2_fill_1 FILLER_53_191 ();
 sg13g2_decap_4 FILLER_53_205 ();
 sg13g2_fill_1 FILLER_53_292 ();
 sg13g2_decap_8 FILLER_53_302 ();
 sg13g2_fill_1 FILLER_53_309 ();
 sg13g2_decap_8 FILLER_53_314 ();
 sg13g2_decap_8 FILLER_53_321 ();
 sg13g2_decap_8 FILLER_53_328 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_25 ();
 sg13g2_fill_2 FILLER_54_32 ();
 sg13g2_fill_1 FILLER_54_34 ();
 sg13g2_fill_2 FILLER_54_53 ();
 sg13g2_decap_4 FILLER_54_60 ();
 sg13g2_fill_2 FILLER_54_64 ();
 sg13g2_decap_8 FILLER_54_75 ();
 sg13g2_fill_2 FILLER_54_96 ();
 sg13g2_fill_1 FILLER_54_98 ();
 sg13g2_fill_2 FILLER_54_111 ();
 sg13g2_fill_1 FILLER_54_113 ();
 sg13g2_fill_1 FILLER_54_119 ();
 sg13g2_fill_1 FILLER_54_130 ();
 sg13g2_fill_1 FILLER_54_136 ();
 sg13g2_decap_4 FILLER_54_141 ();
 sg13g2_fill_2 FILLER_54_145 ();
 sg13g2_decap_4 FILLER_54_174 ();
 sg13g2_decap_8 FILLER_54_182 ();
 sg13g2_fill_2 FILLER_54_189 ();
 sg13g2_fill_1 FILLER_54_218 ();
 sg13g2_fill_1 FILLER_54_266 ();
 sg13g2_decap_8 FILLER_54_290 ();
 sg13g2_decap_8 FILLER_54_297 ();
 sg13g2_decap_8 FILLER_54_313 ();
 sg13g2_decap_8 FILLER_54_320 ();
 sg13g2_decap_8 FILLER_54_327 ();
 sg13g2_decap_8 FILLER_54_334 ();
 sg13g2_fill_1 FILLER_54_373 ();
 sg13g2_decap_4 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_4 ();
 sg13g2_fill_1 FILLER_55_23 ();
 sg13g2_fill_1 FILLER_55_51 ();
 sg13g2_fill_2 FILLER_55_57 ();
 sg13g2_fill_2 FILLER_55_110 ();
 sg13g2_fill_1 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_147 ();
 sg13g2_fill_1 FILLER_55_154 ();
 sg13g2_decap_8 FILLER_55_167 ();
 sg13g2_fill_2 FILLER_55_174 ();
 sg13g2_fill_1 FILLER_55_176 ();
 sg13g2_decap_8 FILLER_55_181 ();
 sg13g2_decap_8 FILLER_55_188 ();
 sg13g2_decap_8 FILLER_55_195 ();
 sg13g2_decap_4 FILLER_55_202 ();
 sg13g2_fill_1 FILLER_55_206 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_fill_2 FILLER_55_224 ();
 sg13g2_fill_2 FILLER_55_244 ();
 sg13g2_fill_1 FILLER_55_246 ();
 sg13g2_fill_2 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_284 ();
 sg13g2_decap_4 FILLER_55_291 ();
 sg13g2_fill_2 FILLER_55_311 ();
 sg13g2_fill_1 FILLER_55_324 ();
 sg13g2_decap_8 FILLER_55_334 ();
 sg13g2_decap_8 FILLER_55_341 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_4 ();
 sg13g2_fill_2 FILLER_56_20 ();
 sg13g2_fill_2 FILLER_56_31 ();
 sg13g2_fill_1 FILLER_56_33 ();
 sg13g2_fill_1 FILLER_56_41 ();
 sg13g2_fill_2 FILLER_56_66 ();
 sg13g2_fill_1 FILLER_56_77 ();
 sg13g2_fill_2 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_115 ();
 sg13g2_decap_4 FILLER_56_122 ();
 sg13g2_fill_1 FILLER_56_126 ();
 sg13g2_fill_2 FILLER_56_132 ();
 sg13g2_fill_1 FILLER_56_134 ();
 sg13g2_decap_8 FILLER_56_144 ();
 sg13g2_decap_8 FILLER_56_151 ();
 sg13g2_decap_8 FILLER_56_162 ();
 sg13g2_fill_1 FILLER_56_169 ();
 sg13g2_decap_4 FILLER_56_187 ();
 sg13g2_fill_1 FILLER_56_196 ();
 sg13g2_fill_2 FILLER_56_206 ();
 sg13g2_decap_8 FILLER_56_213 ();
 sg13g2_fill_1 FILLER_56_220 ();
 sg13g2_decap_8 FILLER_56_275 ();
 sg13g2_decap_4 FILLER_56_282 ();
 sg13g2_fill_1 FILLER_56_324 ();
 sg13g2_fill_2 FILLER_56_356 ();
 sg13g2_fill_1 FILLER_56_358 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_16 ();
 sg13g2_decap_4 FILLER_57_22 ();
 sg13g2_fill_2 FILLER_57_43 ();
 sg13g2_fill_2 FILLER_57_50 ();
 sg13g2_fill_1 FILLER_57_52 ();
 sg13g2_decap_8 FILLER_57_58 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_fill_1 FILLER_57_98 ();
 sg13g2_decap_4 FILLER_57_104 ();
 sg13g2_fill_2 FILLER_57_112 ();
 sg13g2_decap_4 FILLER_57_117 ();
 sg13g2_fill_2 FILLER_57_152 ();
 sg13g2_fill_1 FILLER_57_154 ();
 sg13g2_fill_2 FILLER_57_183 ();
 sg13g2_fill_1 FILLER_57_185 ();
 sg13g2_fill_1 FILLER_57_193 ();
 sg13g2_fill_2 FILLER_57_220 ();
 sg13g2_fill_2 FILLER_57_262 ();
 sg13g2_decap_8 FILLER_57_272 ();
 sg13g2_decap_4 FILLER_57_283 ();
 sg13g2_fill_1 FILLER_57_287 ();
 sg13g2_decap_4 FILLER_57_305 ();
 sg13g2_fill_2 FILLER_57_328 ();
 sg13g2_fill_2 FILLER_57_383 ();
 sg13g2_fill_1 FILLER_57_399 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_12 ();
 sg13g2_decap_8 FILLER_58_19 ();
 sg13g2_decap_8 FILLER_58_26 ();
 sg13g2_fill_1 FILLER_58_33 ();
 sg13g2_fill_2 FILLER_58_38 ();
 sg13g2_decap_8 FILLER_58_44 ();
 sg13g2_decap_8 FILLER_58_51 ();
 sg13g2_decap_8 FILLER_58_58 ();
 sg13g2_decap_8 FILLER_58_65 ();
 sg13g2_fill_1 FILLER_58_72 ();
 sg13g2_fill_2 FILLER_58_99 ();
 sg13g2_fill_1 FILLER_58_101 ();
 sg13g2_decap_8 FILLER_58_121 ();
 sg13g2_fill_2 FILLER_58_132 ();
 sg13g2_decap_8 FILLER_58_144 ();
 sg13g2_decap_8 FILLER_58_151 ();
 sg13g2_decap_8 FILLER_58_158 ();
 sg13g2_fill_2 FILLER_58_165 ();
 sg13g2_fill_2 FILLER_58_173 ();
 sg13g2_fill_1 FILLER_58_175 ();
 sg13g2_fill_2 FILLER_58_181 ();
 sg13g2_decap_4 FILLER_58_189 ();
 sg13g2_fill_2 FILLER_58_209 ();
 sg13g2_decap_8 FILLER_58_221 ();
 sg13g2_decap_8 FILLER_58_228 ();
 sg13g2_fill_1 FILLER_58_235 ();
 sg13g2_fill_1 FILLER_58_241 ();
 sg13g2_decap_4 FILLER_58_247 ();
 sg13g2_fill_2 FILLER_58_251 ();
 sg13g2_decap_8 FILLER_58_258 ();
 sg13g2_decap_8 FILLER_58_265 ();
 sg13g2_fill_1 FILLER_58_272 ();
 sg13g2_fill_2 FILLER_58_279 ();
 sg13g2_fill_1 FILLER_58_281 ();
 sg13g2_fill_2 FILLER_58_287 ();
 sg13g2_fill_2 FILLER_58_294 ();
 sg13g2_fill_1 FILLER_58_296 ();
 sg13g2_fill_2 FILLER_58_318 ();
 sg13g2_fill_1 FILLER_58_320 ();
 sg13g2_decap_4 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_4 ();
 sg13g2_decap_4 FILLER_59_24 ();
 sg13g2_fill_1 FILLER_59_28 ();
 sg13g2_fill_2 FILLER_59_34 ();
 sg13g2_fill_2 FILLER_59_55 ();
 sg13g2_fill_1 FILLER_59_57 ();
 sg13g2_decap_8 FILLER_59_72 ();
 sg13g2_decap_4 FILLER_59_79 ();
 sg13g2_fill_1 FILLER_59_83 ();
 sg13g2_fill_2 FILLER_59_93 ();
 sg13g2_fill_1 FILLER_59_95 ();
 sg13g2_fill_1 FILLER_59_101 ();
 sg13g2_decap_8 FILLER_59_123 ();
 sg13g2_decap_8 FILLER_59_130 ();
 sg13g2_decap_4 FILLER_59_146 ();
 sg13g2_fill_2 FILLER_59_150 ();
 sg13g2_fill_1 FILLER_59_165 ();
 sg13g2_fill_1 FILLER_59_171 ();
 sg13g2_decap_8 FILLER_59_182 ();
 sg13g2_fill_2 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_196 ();
 sg13g2_decap_4 FILLER_59_203 ();
 sg13g2_decap_4 FILLER_59_217 ();
 sg13g2_fill_1 FILLER_59_221 ();
 sg13g2_decap_4 FILLER_59_261 ();
 sg13g2_fill_2 FILLER_59_277 ();
 sg13g2_fill_1 FILLER_59_279 ();
 sg13g2_fill_2 FILLER_59_334 ();
 sg13g2_fill_2 FILLER_59_350 ();
 sg13g2_fill_1 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_21 ();
 sg13g2_fill_2 FILLER_60_28 ();
 sg13g2_fill_1 FILLER_60_30 ();
 sg13g2_decap_8 FILLER_60_48 ();
 sg13g2_decap_8 FILLER_60_55 ();
 sg13g2_fill_2 FILLER_60_73 ();
 sg13g2_fill_1 FILLER_60_75 ();
 sg13g2_fill_1 FILLER_60_106 ();
 sg13g2_fill_2 FILLER_60_125 ();
 sg13g2_fill_2 FILLER_60_142 ();
 sg13g2_fill_2 FILLER_60_154 ();
 sg13g2_fill_1 FILLER_60_161 ();
 sg13g2_fill_2 FILLER_60_166 ();
 sg13g2_fill_1 FILLER_60_173 ();
 sg13g2_decap_4 FILLER_60_180 ();
 sg13g2_fill_1 FILLER_60_184 ();
 sg13g2_fill_1 FILLER_60_202 ();
 sg13g2_fill_2 FILLER_60_223 ();
 sg13g2_fill_2 FILLER_60_293 ();
 sg13g2_fill_1 FILLER_60_295 ();
 sg13g2_fill_1 FILLER_60_322 ();
 sg13g2_fill_2 FILLER_60_336 ();
 sg13g2_fill_1 FILLER_60_346 ();
 sg13g2_fill_2 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_4 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_4 ();
 sg13g2_fill_2 FILLER_61_20 ();
 sg13g2_fill_2 FILLER_61_27 ();
 sg13g2_decap_4 FILLER_61_35 ();
 sg13g2_fill_1 FILLER_61_39 ();
 sg13g2_fill_2 FILLER_61_50 ();
 sg13g2_fill_1 FILLER_61_52 ();
 sg13g2_decap_4 FILLER_61_66 ();
 sg13g2_fill_2 FILLER_61_113 ();
 sg13g2_fill_1 FILLER_61_115 ();
 sg13g2_decap_4 FILLER_61_126 ();
 sg13g2_fill_1 FILLER_61_130 ();
 sg13g2_fill_2 FILLER_61_146 ();
 sg13g2_fill_2 FILLER_61_168 ();
 sg13g2_fill_2 FILLER_61_194 ();
 sg13g2_fill_1 FILLER_61_196 ();
 sg13g2_fill_2 FILLER_61_217 ();
 sg13g2_fill_1 FILLER_61_219 ();
 sg13g2_fill_1 FILLER_61_234 ();
 sg13g2_fill_1 FILLER_61_249 ();
 sg13g2_fill_1 FILLER_61_264 ();
 sg13g2_decap_4 FILLER_61_279 ();
 sg13g2_fill_2 FILLER_61_297 ();
 sg13g2_fill_1 FILLER_61_299 ();
 sg13g2_fill_1 FILLER_61_326 ();
 sg13g2_fill_2 FILLER_61_362 ();
 sg13g2_fill_1 FILLER_61_382 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_fill_1 FILLER_62_35 ();
 sg13g2_fill_1 FILLER_62_46 ();
 sg13g2_decap_4 FILLER_62_71 ();
 sg13g2_fill_2 FILLER_62_88 ();
 sg13g2_fill_1 FILLER_62_90 ();
 sg13g2_decap_8 FILLER_62_124 ();
 sg13g2_fill_2 FILLER_62_131 ();
 sg13g2_fill_1 FILLER_62_138 ();
 sg13g2_decap_8 FILLER_62_143 ();
 sg13g2_decap_8 FILLER_62_150 ();
 sg13g2_decap_8 FILLER_62_157 ();
 sg13g2_decap_8 FILLER_62_169 ();
 sg13g2_fill_1 FILLER_62_176 ();
 sg13g2_decap_8 FILLER_62_182 ();
 sg13g2_decap_4 FILLER_62_189 ();
 sg13g2_fill_2 FILLER_62_198 ();
 sg13g2_fill_1 FILLER_62_215 ();
 sg13g2_fill_2 FILLER_62_293 ();
 sg13g2_fill_1 FILLER_62_300 ();
 sg13g2_fill_2 FILLER_62_311 ();
 sg13g2_fill_1 FILLER_62_322 ();
 sg13g2_fill_1 FILLER_62_358 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_20 ();
 sg13g2_fill_2 FILLER_63_40 ();
 sg13g2_decap_4 FILLER_63_56 ();
 sg13g2_fill_1 FILLER_63_60 ();
 sg13g2_decap_8 FILLER_63_71 ();
 sg13g2_fill_2 FILLER_63_78 ();
 sg13g2_fill_1 FILLER_63_80 ();
 sg13g2_decap_4 FILLER_63_137 ();
 sg13g2_decap_4 FILLER_63_146 ();
 sg13g2_fill_1 FILLER_63_150 ();
 sg13g2_fill_1 FILLER_63_158 ();
 sg13g2_fill_2 FILLER_63_168 ();
 sg13g2_decap_4 FILLER_63_206 ();
 sg13g2_decap_8 FILLER_63_220 ();
 sg13g2_decap_4 FILLER_63_274 ();
 sg13g2_fill_1 FILLER_63_295 ();
 sg13g2_fill_1 FILLER_63_336 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_27 ();
 sg13g2_fill_1 FILLER_64_29 ();
 sg13g2_fill_1 FILLER_64_38 ();
 sg13g2_decap_8 FILLER_64_44 ();
 sg13g2_decap_8 FILLER_64_51 ();
 sg13g2_decap_8 FILLER_64_58 ();
 sg13g2_decap_8 FILLER_64_65 ();
 sg13g2_decap_8 FILLER_64_72 ();
 sg13g2_decap_8 FILLER_64_79 ();
 sg13g2_decap_8 FILLER_64_86 ();
 sg13g2_fill_2 FILLER_64_93 ();
 sg13g2_decap_4 FILLER_64_104 ();
 sg13g2_fill_1 FILLER_64_108 ();
 sg13g2_fill_1 FILLER_64_127 ();
 sg13g2_fill_1 FILLER_64_136 ();
 sg13g2_fill_2 FILLER_64_147 ();
 sg13g2_fill_2 FILLER_64_166 ();
 sg13g2_fill_2 FILLER_64_181 ();
 sg13g2_fill_1 FILLER_64_183 ();
 sg13g2_decap_4 FILLER_64_195 ();
 sg13g2_decap_8 FILLER_64_209 ();
 sg13g2_decap_4 FILLER_64_216 ();
 sg13g2_fill_1 FILLER_64_220 ();
 sg13g2_fill_2 FILLER_64_253 ();
 sg13g2_fill_2 FILLER_64_281 ();
 sg13g2_fill_1 FILLER_64_283 ();
 sg13g2_fill_2 FILLER_64_289 ();
 sg13g2_fill_2 FILLER_64_301 ();
 sg13g2_fill_1 FILLER_64_326 ();
 sg13g2_fill_2 FILLER_64_398 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_31 ();
 sg13g2_fill_2 FILLER_65_35 ();
 sg13g2_decap_4 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_90 ();
 sg13g2_decap_8 FILLER_65_97 ();
 sg13g2_decap_8 FILLER_65_104 ();
 sg13g2_decap_4 FILLER_65_111 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_fill_1 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_139 ();
 sg13g2_decap_4 FILLER_65_146 ();
 sg13g2_decap_8 FILLER_65_179 ();
 sg13g2_decap_8 FILLER_65_186 ();
 sg13g2_decap_8 FILLER_65_193 ();
 sg13g2_decap_8 FILLER_65_200 ();
 sg13g2_decap_8 FILLER_65_207 ();
 sg13g2_fill_2 FILLER_65_214 ();
 sg13g2_fill_2 FILLER_65_279 ();
 sg13g2_fill_2 FILLER_65_309 ();
 sg13g2_fill_1 FILLER_65_372 ();
 sg13g2_fill_1 FILLER_65_382 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_26 ();
 sg13g2_fill_2 FILLER_66_48 ();
 sg13g2_decap_8 FILLER_66_103 ();
 sg13g2_decap_8 FILLER_66_110 ();
 sg13g2_fill_1 FILLER_66_129 ();
 sg13g2_fill_2 FILLER_66_139 ();
 sg13g2_fill_1 FILLER_66_141 ();
 sg13g2_decap_4 FILLER_66_147 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_4 FILLER_66_175 ();
 sg13g2_fill_2 FILLER_66_179 ();
 sg13g2_decap_4 FILLER_66_186 ();
 sg13g2_fill_2 FILLER_66_194 ();
 sg13g2_fill_1 FILLER_66_205 ();
 sg13g2_fill_2 FILLER_66_233 ();
 sg13g2_fill_1 FILLER_66_256 ();
 sg13g2_fill_2 FILLER_66_297 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_4 FILLER_67_21 ();
 sg13g2_fill_1 FILLER_67_25 ();
 sg13g2_decap_4 FILLER_67_40 ();
 sg13g2_decap_8 FILLER_67_103 ();
 sg13g2_decap_4 FILLER_67_110 ();
 sg13g2_fill_2 FILLER_67_140 ();
 sg13g2_decap_4 FILLER_67_156 ();
 sg13g2_fill_1 FILLER_67_160 ();
 sg13g2_fill_1 FILLER_67_172 ();
 sg13g2_fill_2 FILLER_67_176 ();
 sg13g2_fill_2 FILLER_67_241 ();
 sg13g2_fill_2 FILLER_67_284 ();
 sg13g2_fill_1 FILLER_67_286 ();
 sg13g2_fill_2 FILLER_67_309 ();
 sg13g2_fill_1 FILLER_67_384 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_4 ();
 sg13g2_fill_1 FILLER_68_20 ();
 sg13g2_fill_2 FILLER_68_33 ();
 sg13g2_fill_2 FILLER_68_67 ();
 sg13g2_decap_4 FILLER_68_116 ();
 sg13g2_fill_2 FILLER_68_120 ();
 sg13g2_fill_1 FILLER_68_148 ();
 sg13g2_fill_1 FILLER_68_197 ();
 sg13g2_fill_1 FILLER_68_210 ();
 sg13g2_fill_2 FILLER_68_277 ();
 sg13g2_fill_1 FILLER_68_279 ();
 sg13g2_fill_1 FILLER_68_320 ();
 sg13g2_fill_1 FILLER_68_382 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_2 ();
 sg13g2_fill_2 FILLER_69_30 ();
 sg13g2_fill_1 FILLER_69_87 ();
 sg13g2_decap_8 FILLER_69_124 ();
 sg13g2_decap_4 FILLER_69_131 ();
 sg13g2_fill_2 FILLER_69_135 ();
 sg13g2_fill_1 FILLER_69_151 ();
 sg13g2_decap_8 FILLER_69_169 ();
 sg13g2_fill_2 FILLER_69_176 ();
 sg13g2_fill_1 FILLER_69_178 ();
 sg13g2_fill_2 FILLER_69_188 ();
 sg13g2_decap_8 FILLER_69_198 ();
 sg13g2_fill_2 FILLER_69_262 ();
 sg13g2_fill_1 FILLER_69_341 ();
 sg13g2_fill_2 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_2 ();
 sg13g2_fill_2 FILLER_70_23 ();
 sg13g2_fill_1 FILLER_70_25 ();
 sg13g2_fill_2 FILLER_70_30 ();
 sg13g2_fill_1 FILLER_70_32 ();
 sg13g2_decap_4 FILLER_70_51 ();
 sg13g2_fill_2 FILLER_70_55 ();
 sg13g2_decap_4 FILLER_70_130 ();
 sg13g2_fill_1 FILLER_70_134 ();
 sg13g2_fill_2 FILLER_70_141 ();
 sg13g2_decap_8 FILLER_70_180 ();
 sg13g2_decap_8 FILLER_70_187 ();
 sg13g2_decap_8 FILLER_70_194 ();
 sg13g2_decap_8 FILLER_70_201 ();
 sg13g2_decap_8 FILLER_70_208 ();
 sg13g2_fill_1 FILLER_70_246 ();
 sg13g2_fill_1 FILLER_70_252 ();
 sg13g2_fill_2 FILLER_70_311 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_4 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_fill_2 FILLER_71_35 ();
 sg13g2_fill_1 FILLER_71_37 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_fill_2 FILLER_71_49 ();
 sg13g2_fill_1 FILLER_71_98 ();
 sg13g2_fill_1 FILLER_71_108 ();
 sg13g2_fill_1 FILLER_71_144 ();
 sg13g2_fill_2 FILLER_71_169 ();
 sg13g2_fill_1 FILLER_71_171 ();
 sg13g2_decap_8 FILLER_71_198 ();
 sg13g2_decap_8 FILLER_71_205 ();
 sg13g2_decap_8 FILLER_71_212 ();
 sg13g2_decap_8 FILLER_71_219 ();
 sg13g2_decap_4 FILLER_71_226 ();
 sg13g2_fill_2 FILLER_71_230 ();
 sg13g2_fill_2 FILLER_71_360 ();
 sg13g2_decap_4 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_72_4 ();
 sg13g2_fill_2 FILLER_72_13 ();
 sg13g2_fill_1 FILLER_72_15 ();
 sg13g2_decap_4 FILLER_72_21 ();
 sg13g2_fill_1 FILLER_72_25 ();
 sg13g2_fill_1 FILLER_72_33 ();
 sg13g2_fill_2 FILLER_72_37 ();
 sg13g2_fill_1 FILLER_72_99 ();
 sg13g2_fill_1 FILLER_72_187 ();
 sg13g2_decap_8 FILLER_72_214 ();
 sg13g2_fill_2 FILLER_72_221 ();
 sg13g2_fill_2 FILLER_72_231 ();
 sg13g2_fill_2 FILLER_72_296 ();
 sg13g2_fill_1 FILLER_72_307 ();
 sg13g2_fill_2 FILLER_72_326 ();
 sg13g2_fill_2 FILLER_73_14 ();
 sg13g2_fill_1 FILLER_73_24 ();
 sg13g2_fill_2 FILLER_73_61 ();
 sg13g2_fill_2 FILLER_73_74 ();
 sg13g2_fill_1 FILLER_73_146 ();
 sg13g2_decap_4 FILLER_73_173 ();
 sg13g2_fill_2 FILLER_73_221 ();
 sg13g2_fill_2 FILLER_73_236 ();
 sg13g2_fill_1 FILLER_73_248 ();
 sg13g2_fill_1 FILLER_74_34 ();
 sg13g2_fill_2 FILLER_74_78 ();
 sg13g2_fill_1 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_164 ();
 sg13g2_fill_2 FILLER_74_171 ();
 sg13g2_fill_1 FILLER_74_173 ();
 sg13g2_fill_2 FILLER_74_179 ();
 sg13g2_fill_2 FILLER_74_276 ();
 sg13g2_fill_1 FILLER_74_345 ();
 sg13g2_fill_1 FILLER_74_360 ();
 sg13g2_fill_1 FILLER_74_394 ();
 sg13g2_fill_2 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_23 ();
 sg13g2_fill_1 FILLER_75_38 ();
 sg13g2_fill_1 FILLER_75_47 ();
 sg13g2_fill_1 FILLER_75_74 ();
 sg13g2_fill_1 FILLER_75_94 ();
 sg13g2_fill_1 FILLER_75_134 ();
 sg13g2_decap_8 FILLER_75_158 ();
 sg13g2_decap_8 FILLER_75_165 ();
 sg13g2_fill_1 FILLER_75_172 ();
 sg13g2_fill_1 FILLER_75_240 ();
 sg13g2_fill_1 FILLER_75_303 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_32 ();
 sg13g2_fill_1 FILLER_76_46 ();
 sg13g2_fill_2 FILLER_76_125 ();
 sg13g2_fill_1 FILLER_76_127 ();
 sg13g2_fill_1 FILLER_76_216 ();
 sg13g2_fill_2 FILLER_76_236 ();
 sg13g2_fill_2 FILLER_76_314 ();
 sg13g2_fill_1 FILLER_76_344 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_4 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_4 ();
 sg13g2_fill_1 FILLER_77_115 ();
 sg13g2_fill_2 FILLER_77_166 ();
 sg13g2_fill_1 FILLER_77_190 ();
 sg13g2_fill_1 FILLER_77_200 ();
 sg13g2_fill_2 FILLER_77_271 ();
 sg13g2_fill_1 FILLER_77_356 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_28 ();
 sg13g2_fill_2 FILLER_78_64 ();
 sg13g2_fill_2 FILLER_78_107 ();
 sg13g2_fill_1 FILLER_78_109 ();
 sg13g2_fill_2 FILLER_78_123 ();
 sg13g2_fill_1 FILLER_78_148 ();
 sg13g2_fill_1 FILLER_78_167 ();
 sg13g2_fill_2 FILLER_78_194 ();
 sg13g2_fill_2 FILLER_78_289 ();
 sg13g2_fill_1 FILLER_78_300 ();
 sg13g2_fill_2 FILLER_78_345 ();
 sg13g2_fill_1 FILLER_78_347 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_2 ();
 sg13g2_fill_1 FILLER_79_79 ();
 sg13g2_fill_2 FILLER_79_132 ();
 sg13g2_fill_1 FILLER_79_169 ();
 sg13g2_fill_2 FILLER_79_196 ();
 sg13g2_fill_1 FILLER_79_198 ();
 sg13g2_fill_2 FILLER_79_283 ();
 sg13g2_fill_1 FILLER_79_285 ();
 sg13g2_fill_1 FILLER_79_317 ();
 sg13g2_fill_2 FILLER_79_353 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_7 ();
 sg13g2_fill_2 FILLER_80_73 ();
 sg13g2_fill_2 FILLER_80_84 ();
 sg13g2_fill_2 FILLER_80_90 ();
 sg13g2_fill_1 FILLER_80_121 ();
 sg13g2_fill_2 FILLER_80_148 ();
 sg13g2_fill_1 FILLER_80_150 ();
 sg13g2_fill_2 FILLER_80_214 ();
 sg13g2_fill_2 FILLER_80_243 ();
 sg13g2_fill_2 FILLER_80_249 ();
 sg13g2_fill_1 FILLER_80_279 ();
 sg13g2_fill_2 FILLER_80_292 ();
 sg13g2_fill_1 FILLER_80_294 ();
 sg13g2_fill_1 FILLER_80_313 ();
 sg13g2_fill_1 FILLER_80_336 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
endmodule

module tt_um_flummer_ltc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire \ltc.bit_clk ;
 wire \ltc.bit_counter[0] ;
 wire \ltc.bit_counter[10] ;
 wire \ltc.bit_counter[11] ;
 wire \ltc.bit_counter[1] ;
 wire \ltc.bit_counter[2] ;
 wire \ltc.bit_counter[3] ;
 wire \ltc.bit_counter[4] ;
 wire \ltc.bit_counter[5] ;
 wire \ltc.bit_counter[6] ;
 wire \ltc.bit_counter[7] ;
 wire \ltc.bit_counter[8] ;
 wire \ltc.bit_counter[9] ;
 wire \ltc.frm_counter[0] ;
 wire \ltc.frm_counter[10] ;
 wire \ltc.frm_counter[11] ;
 wire \ltc.frm_counter[12] ;
 wire \ltc.frm_counter[13] ;
 wire \ltc.frm_counter[14] ;
 wire \ltc.frm_counter[15] ;
 wire \ltc.frm_counter[16] ;
 wire \ltc.frm_counter[17] ;
 wire \ltc.frm_counter[18] ;
 wire \ltc.frm_counter[19] ;
 wire \ltc.frm_counter[1] ;
 wire \ltc.frm_counter[20] ;
 wire \ltc.frm_counter[21] ;
 wire \ltc.frm_counter[22] ;
 wire \ltc.frm_counter[23] ;
 wire \ltc.frm_counter[2] ;
 wire \ltc.frm_counter[3] ;
 wire \ltc.frm_counter[4] ;
 wire \ltc.frm_counter[5] ;
 wire \ltc.frm_counter[6] ;
 wire \ltc.frm_counter[7] ;
 wire \ltc.frm_counter[8] ;
 wire \ltc.frm_counter[9] ;
 wire \ltc.frm_d[0] ;
 wire \ltc.frm_d[1] ;
 wire \ltc.frm_u[0] ;
 wire \ltc.frm_u[1] ;
 wire \ltc.frm_u[2] ;
 wire \ltc.frm_u[3] ;
 wire \ltc.hrs_d[0] ;
 wire \ltc.hrs_d[1] ;
 wire \ltc.hrs_u[0] ;
 wire \ltc.hrs_u[1] ;
 wire \ltc.hrs_u[2] ;
 wire \ltc.hrs_u[3] ;
 wire \ltc.min_d[0] ;
 wire \ltc.min_d[1] ;
 wire \ltc.min_d[2] ;
 wire \ltc.min_u[0] ;
 wire \ltc.min_u[1] ;
 wire \ltc.min_u[2] ;
 wire \ltc.min_u[3] ;
 wire \ltc.output_buffer[0] ;
 wire \ltc.output_buffer[10] ;
 wire \ltc.output_buffer[11] ;
 wire \ltc.output_buffer[12] ;
 wire \ltc.output_buffer[13] ;
 wire \ltc.output_buffer[14] ;
 wire \ltc.output_buffer[15] ;
 wire \ltc.output_buffer[16] ;
 wire \ltc.output_buffer[17] ;
 wire \ltc.output_buffer[18] ;
 wire \ltc.output_buffer[19] ;
 wire \ltc.output_buffer[1] ;
 wire \ltc.output_buffer[20] ;
 wire \ltc.output_buffer[21] ;
 wire \ltc.output_buffer[22] ;
 wire \ltc.output_buffer[23] ;
 wire \ltc.output_buffer[24] ;
 wire \ltc.output_buffer[25] ;
 wire \ltc.output_buffer[26] ;
 wire \ltc.output_buffer[27] ;
 wire \ltc.output_buffer[28] ;
 wire \ltc.output_buffer[29] ;
 wire \ltc.output_buffer[2] ;
 wire \ltc.output_buffer[30] ;
 wire \ltc.output_buffer[31] ;
 wire \ltc.output_buffer[32] ;
 wire \ltc.output_buffer[33] ;
 wire \ltc.output_buffer[34] ;
 wire \ltc.output_buffer[35] ;
 wire \ltc.output_buffer[36] ;
 wire \ltc.output_buffer[37] ;
 wire \ltc.output_buffer[38] ;
 wire \ltc.output_buffer[39] ;
 wire \ltc.output_buffer[3] ;
 wire \ltc.output_buffer[40] ;
 wire \ltc.output_buffer[41] ;
 wire \ltc.output_buffer[42] ;
 wire \ltc.output_buffer[43] ;
 wire \ltc.output_buffer[44] ;
 wire \ltc.output_buffer[45] ;
 wire \ltc.output_buffer[46] ;
 wire \ltc.output_buffer[47] ;
 wire \ltc.output_buffer[48] ;
 wire \ltc.output_buffer[49] ;
 wire \ltc.output_buffer[4] ;
 wire \ltc.output_buffer[50] ;
 wire \ltc.output_buffer[51] ;
 wire \ltc.output_buffer[52] ;
 wire \ltc.output_buffer[53] ;
 wire \ltc.output_buffer[54] ;
 wire \ltc.output_buffer[55] ;
 wire \ltc.output_buffer[56] ;
 wire \ltc.output_buffer[57] ;
 wire \ltc.output_buffer[58] ;
 wire \ltc.output_buffer[59] ;
 wire \ltc.output_buffer[5] ;
 wire \ltc.output_buffer[60] ;
 wire \ltc.output_buffer[61] ;
 wire \ltc.output_buffer[62] ;
 wire \ltc.output_buffer[63] ;
 wire \ltc.output_buffer[64] ;
 wire \ltc.output_buffer[65] ;
 wire \ltc.output_buffer[66] ;
 wire \ltc.output_buffer[67] ;
 wire \ltc.output_buffer[68] ;
 wire \ltc.output_buffer[69] ;
 wire \ltc.output_buffer[6] ;
 wire \ltc.output_buffer[70] ;
 wire \ltc.output_buffer[71] ;
 wire \ltc.output_buffer[72] ;
 wire \ltc.output_buffer[73] ;
 wire \ltc.output_buffer[74] ;
 wire \ltc.output_buffer[75] ;
 wire \ltc.output_buffer[76] ;
 wire \ltc.output_buffer[77] ;
 wire \ltc.output_buffer[78] ;
 wire \ltc.output_buffer[79] ;
 wire \ltc.output_buffer[7] ;
 wire \ltc.output_buffer[8] ;
 wire \ltc.output_buffer[9] ;
 wire \ltc.sec_d[0] ;
 wire \ltc.sec_d[1] ;
 wire \ltc.sec_d[2] ;
 wire \ltc.sec_u[0] ;
 wire \ltc.sec_u[1] ;
 wire \ltc.sec_u[2] ;
 wire \ltc.sec_u[3] ;
 wire \ltc.timecode ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_0_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;

 sg13g2_inv_1 _0875_ (.Y(_0155_),
    .A(\ltc.bit_clk ));
 sg13g2_inv_1 _0876_ (.Y(_0156_),
    .A(net384));
 sg13g2_inv_1 _0877_ (.Y(_0157_),
    .A(net415));
 sg13g2_inv_1 _0878_ (.Y(_0158_),
    .A(net212));
 sg13g2_inv_1 _0879_ (.Y(_0159_),
    .A(\ltc.frm_d[0] ));
 sg13g2_inv_1 _0880_ (.Y(_0160_),
    .A(net373));
 sg13g2_inv_1 _0881_ (.Y(_0161_),
    .A(net409));
 sg13g2_inv_1 _0882_ (.Y(_0162_),
    .A(net448));
 sg13g2_inv_1 _0883_ (.Y(_0163_),
    .A(\ltc.frm_counter[12] ));
 sg13g2_inv_1 _0884_ (.Y(_0164_),
    .A(\ltc.frm_counter[14] ));
 sg13g2_inv_1 _0885_ (.Y(_0165_),
    .A(\ltc.bit_counter[10] ));
 sg13g2_inv_2 _0886_ (.Y(_0166_),
    .A(net227));
 sg13g2_inv_1 _0887_ (.Y(_0167_),
    .A(net170));
 sg13g2_inv_1 _0888_ (.Y(_0168_),
    .A(\ltc.output_buffer[79] ));
 sg13g2_inv_1 _0889_ (.Y(_0169_),
    .A(net238));
 sg13g2_inv_1 _0890_ (.Y(_0170_),
    .A(net282));
 sg13g2_inv_1 _0891_ (.Y(_0171_),
    .A(net280));
 sg13g2_inv_1 _0892_ (.Y(_0172_),
    .A(net275));
 sg13g2_inv_1 _0893_ (.Y(_0173_),
    .A(net287));
 sg13g2_inv_1 _0894_ (.Y(_0174_),
    .A(net262));
 sg13g2_inv_1 _0895_ (.Y(_0175_),
    .A(net277));
 sg13g2_inv_1 _0896_ (.Y(_0176_),
    .A(net289));
 sg13g2_inv_1 _0897_ (.Y(_0177_),
    .A(net260));
 sg13g2_inv_1 _0898_ (.Y(_0178_),
    .A(net266));
 sg13g2_inv_1 _0899_ (.Y(_0179_),
    .A(net286));
 sg13g2_inv_1 _0900_ (.Y(_0180_),
    .A(net302));
 sg13g2_inv_1 _0901_ (.Y(_0181_),
    .A(net251));
 sg13g2_nand2_1 _0902_ (.Y(_0182_),
    .A(net7),
    .B(net8));
 sg13g2_nand4_1 _0903_ (.B(net5),
    .C(net2),
    .A(net6),
    .Y(_0183_),
    .D(net1));
 sg13g2_nor2_2 _0904_ (.A(_0182_),
    .B(_0183_),
    .Y(uo_out[0]));
 sg13g2_nor2_1 _0905_ (.A(\ltc.bit_counter[1] ),
    .B(net391),
    .Y(_0184_));
 sg13g2_nor4_2 _0906_ (.A(\ltc.bit_counter[1] ),
    .B(\ltc.bit_counter[0] ),
    .C(\ltc.bit_counter[6] ),
    .Y(_0185_),
    .D(\ltc.bit_counter[7] ));
 sg13g2_nor4_1 _0907_ (.A(\ltc.bit_counter[8] ),
    .B(\ltc.bit_counter[9] ),
    .C(\ltc.bit_counter[10] ),
    .D(\ltc.bit_counter[11] ),
    .Y(_0186_));
 sg13g2_nor4_1 _0908_ (.A(\ltc.bit_counter[5] ),
    .B(\ltc.bit_counter[4] ),
    .C(\ltc.bit_counter[3] ),
    .D(\ltc.bit_counter[2] ),
    .Y(_0187_));
 sg13g2_nand3_1 _0909_ (.B(_0186_),
    .C(_0187_),
    .A(_0185_),
    .Y(_0188_));
 sg13g2_nor2_2 _0910_ (.A(\ltc.bit_clk ),
    .B(_0188_),
    .Y(_0189_));
 sg13g2_nor2_2 _0911_ (.A(net216),
    .B(net204),
    .Y(_0190_));
 sg13g2_nor3_1 _0912_ (.A(\ltc.frm_counter[16] ),
    .B(\ltc.frm_counter[17] ),
    .C(\ltc.frm_counter[18] ),
    .Y(_0191_));
 sg13g2_nor4_1 _0913_ (.A(\ltc.frm_counter[10] ),
    .B(\ltc.frm_counter[11] ),
    .C(\ltc.frm_counter[12] ),
    .D(\ltc.frm_counter[13] ),
    .Y(_0192_));
 sg13g2_nor4_1 _0914_ (.A(\ltc.frm_counter[3] ),
    .B(\ltc.frm_counter[2] ),
    .C(\ltc.frm_counter[6] ),
    .D(\ltc.frm_counter[7] ),
    .Y(_0193_));
 sg13g2_nand3_1 _0915_ (.B(_0192_),
    .C(_0193_),
    .A(_0191_),
    .Y(_0194_));
 sg13g2_nor2_1 _0916_ (.A(\ltc.frm_counter[19] ),
    .B(\ltc.frm_counter[20] ),
    .Y(_0195_));
 sg13g2_nor3_1 _0917_ (.A(\ltc.frm_counter[21] ),
    .B(\ltc.frm_counter[22] ),
    .C(\ltc.frm_counter[23] ),
    .Y(_0196_));
 sg13g2_nand2_1 _0918_ (.Y(_0197_),
    .A(_0195_),
    .B(_0196_));
 sg13g2_nor2_1 _0919_ (.A(\ltc.frm_counter[14] ),
    .B(\ltc.frm_counter[15] ),
    .Y(_0198_));
 sg13g2_nor2_1 _0920_ (.A(\ltc.frm_counter[9] ),
    .B(\ltc.frm_counter[8] ),
    .Y(_0199_));
 sg13g2_nor2_1 _0921_ (.A(\ltc.frm_counter[5] ),
    .B(\ltc.frm_counter[4] ),
    .Y(_0200_));
 sg13g2_nand3_1 _0922_ (.B(_0199_),
    .C(_0200_),
    .A(_0198_),
    .Y(_0201_));
 sg13g2_nor3_2 _0923_ (.A(_0194_),
    .B(_0197_),
    .C(_0201_),
    .Y(_0202_));
 sg13g2_nor2b_1 _0924_ (.A(\ltc.frm_counter[1] ),
    .B_N(net422),
    .Y(_0203_));
 sg13g2_and2_1 _0925_ (.A(_0202_),
    .B(_0203_),
    .X(_0204_));
 sg13g2_nand2_2 _0926_ (.Y(_0205_),
    .A(_0202_),
    .B(_0203_));
 sg13g2_o21ai_1 _0927_ (.B1(net198),
    .Y(_0206_),
    .A1(net388),
    .A2(net193));
 sg13g2_inv_1 _0928_ (.Y(_0011_),
    .A(_0206_));
 sg13g2_nor2_1 _0929_ (.A(net203),
    .B(net192),
    .Y(_0207_));
 sg13g2_a22oi_1 _0930_ (.Y(_0208_),
    .B1(net180),
    .B2(net238),
    .A2(net206),
    .A1(\ltc.output_buffer[0] ));
 sg13g2_nor2_1 _0931_ (.A(net217),
    .B(net239),
    .Y(_0012_));
 sg13g2_a221oi_1 _0932_ (.B2(_0170_),
    .C1(net217),
    .B1(net180),
    .A1(_0169_),
    .Y(_0013_),
    .A2(net206));
 sg13g2_a221oi_1 _0933_ (.B2(_0171_),
    .C1(net217),
    .B1(net180),
    .A1(_0170_),
    .Y(_0014_),
    .A2(net206));
 sg13g2_a221oi_1 _0934_ (.B2(_0172_),
    .C1(net217),
    .B1(net181),
    .A1(_0171_),
    .Y(_0015_),
    .A2(net206));
 sg13g2_a221oi_1 _0935_ (.B2(_0173_),
    .C1(net217),
    .B1(net180),
    .A1(_0172_),
    .Y(_0016_),
    .A2(net206));
 sg13g2_a221oi_1 _0936_ (.B2(_0174_),
    .C1(net219),
    .B1(net182),
    .A1(_0173_),
    .Y(_0017_),
    .A2(net207));
 sg13g2_a221oi_1 _0937_ (.B2(_0175_),
    .C1(net219),
    .B1(net182),
    .A1(_0174_),
    .Y(_0018_),
    .A2(net207));
 sg13g2_a221oi_1 _0938_ (.B2(_0176_),
    .C1(net219),
    .B1(net183),
    .A1(_0175_),
    .Y(_0019_),
    .A2(net208));
 sg13g2_a221oi_1 _0939_ (.B2(_0177_),
    .C1(net220),
    .B1(net183),
    .A1(_0176_),
    .Y(_0020_),
    .A2(net208));
 sg13g2_a221oi_1 _0940_ (.B2(_0178_),
    .C1(net219),
    .B1(net183),
    .A1(_0177_),
    .Y(_0021_),
    .A2(net207));
 sg13g2_a221oi_1 _0941_ (.B2(_0179_),
    .C1(net219),
    .B1(net183),
    .A1(_0178_),
    .Y(_0022_),
    .A2(net207));
 sg13g2_a221oi_1 _0942_ (.B2(_0180_),
    .C1(net219),
    .B1(net183),
    .A1(_0179_),
    .Y(_0023_),
    .A2(net207));
 sg13g2_a221oi_1 _0943_ (.B2(_0181_),
    .C1(net219),
    .B1(net182),
    .A1(_0180_),
    .Y(_0024_),
    .A2(net207));
 sg13g2_a22oi_1 _0944_ (.Y(_0209_),
    .B1(net182),
    .B2(net240),
    .A2(net207),
    .A1(\ltc.output_buffer[13] ));
 sg13g2_nor2_1 _0945_ (.A(net219),
    .B(net241),
    .Y(_0025_));
 sg13g2_a22oi_1 _0946_ (.Y(_0210_),
    .B1(net180),
    .B2(net236),
    .A2(net207),
    .A1(\ltc.output_buffer[14] ));
 sg13g2_nor2_1 _0947_ (.A(net217),
    .B(net237),
    .Y(_0026_));
 sg13g2_a22oi_1 _0948_ (.Y(_0211_),
    .B1(net180),
    .B2(net257),
    .A2(net206),
    .A1(net236));
 sg13g2_nor2_1 _0949_ (.A(net217),
    .B(_0211_),
    .Y(_0027_));
 sg13g2_a22oi_1 _0950_ (.Y(_0212_),
    .B1(net180),
    .B2(net285),
    .A2(net206),
    .A1(net257));
 sg13g2_nor2_1 _0951_ (.A(net217),
    .B(_0212_),
    .Y(_0028_));
 sg13g2_a22oi_1 _0952_ (.Y(_0213_),
    .B1(net180),
    .B2(net288),
    .A2(net209),
    .A1(net285));
 sg13g2_nor2_1 _0953_ (.A(net218),
    .B(_0213_),
    .Y(_0029_));
 sg13g2_a22oi_1 _0954_ (.Y(_0214_),
    .B1(net179),
    .B2(net290),
    .A2(net209),
    .A1(net288));
 sg13g2_nor2_1 _0955_ (.A(net215),
    .B(_0214_),
    .Y(_0030_));
 sg13g2_nand2_1 _0956_ (.Y(_0215_),
    .A(net290),
    .B(net201));
 sg13g2_nor2b_1 _0957_ (.A(net422),
    .B_N(\ltc.frm_counter[1] ),
    .Y(_0216_));
 sg13g2_and2_1 _0958_ (.A(_0202_),
    .B(_0216_),
    .X(_0217_));
 sg13g2_nor2b_2 _0959_ (.A(net4),
    .B_N(net3),
    .Y(_0218_));
 sg13g2_nand2b_1 _0960_ (.Y(_0219_),
    .B(net3),
    .A_N(net4));
 sg13g2_nand2_1 _0961_ (.Y(_0220_),
    .A(_0217_),
    .B(_0218_));
 sg13g2_xnor2_1 _0962_ (.Y(_0221_),
    .A(\ltc.output_buffer[35] ),
    .B(\ltc.output_buffer[34] ));
 sg13g2_xnor2_1 _0963_ (.Y(_0222_),
    .A(\ltc.output_buffer[37] ),
    .B(\ltc.output_buffer[36] ));
 sg13g2_xnor2_1 _0964_ (.Y(_0223_),
    .A(_0221_),
    .B(_0222_));
 sg13g2_xor2_1 _0965_ (.B(\ltc.output_buffer[32] ),
    .A(\ltc.output_buffer[33] ),
    .X(_0224_));
 sg13g2_xnor2_1 _0966_ (.Y(_0225_),
    .A(\ltc.output_buffer[39] ),
    .B(\ltc.output_buffer[38] ));
 sg13g2_xnor2_1 _0967_ (.Y(_0226_),
    .A(_0224_),
    .B(_0225_));
 sg13g2_xnor2_1 _0968_ (.Y(_0227_),
    .A(_0223_),
    .B(_0226_));
 sg13g2_xor2_1 _0969_ (.B(\ltc.output_buffer[46] ),
    .A(\ltc.output_buffer[47] ),
    .X(_0228_));
 sg13g2_xor2_1 _0970_ (.B(\ltc.output_buffer[44] ),
    .A(\ltc.output_buffer[45] ),
    .X(_0229_));
 sg13g2_xnor2_1 _0971_ (.Y(_0230_),
    .A(_0228_),
    .B(_0229_));
 sg13g2_xnor2_1 _0972_ (.Y(_0231_),
    .A(\ltc.output_buffer[31] ),
    .B(\ltc.output_buffer[30] ));
 sg13g2_xor2_1 _0973_ (.B(\ltc.output_buffer[28] ),
    .A(\ltc.output_buffer[29] ),
    .X(_0232_));
 sg13g2_xnor2_1 _0974_ (.Y(_0233_),
    .A(_0231_),
    .B(_0232_));
 sg13g2_xnor2_1 _0975_ (.Y(_0234_),
    .A(_0230_),
    .B(_0233_));
 sg13g2_xnor2_1 _0976_ (.Y(_0235_),
    .A(_0227_),
    .B(_0234_));
 sg13g2_xor2_1 _0977_ (.B(\ltc.output_buffer[18] ),
    .A(\ltc.output_buffer[19] ),
    .X(_0236_));
 sg13g2_xor2_1 _0978_ (.B(\ltc.output_buffer[16] ),
    .A(\ltc.output_buffer[17] ),
    .X(_0237_));
 sg13g2_xnor2_1 _0979_ (.Y(_0238_),
    .A(_0236_),
    .B(_0237_));
 sg13g2_xnor2_1 _0980_ (.Y(_0239_),
    .A(\ltc.output_buffer[23] ),
    .B(\ltc.output_buffer[22] ));
 sg13g2_xor2_1 _0981_ (.B(\ltc.output_buffer[20] ),
    .A(\ltc.output_buffer[21] ),
    .X(_0240_));
 sg13g2_xnor2_1 _0982_ (.Y(_0241_),
    .A(_0239_),
    .B(_0240_));
 sg13g2_xnor2_1 _0983_ (.Y(_0242_),
    .A(_0238_),
    .B(_0241_));
 sg13g2_xor2_1 _0984_ (.B(\ltc.output_buffer[26] ),
    .A(\ltc.output_buffer[27] ),
    .X(_0243_));
 sg13g2_xnor2_1 _0985_ (.Y(_0244_),
    .A(\ltc.output_buffer[41] ),
    .B(\ltc.output_buffer[40] ));
 sg13g2_xnor2_1 _0986_ (.Y(_0245_),
    .A(_0243_),
    .B(_0244_));
 sg13g2_xor2_1 _0987_ (.B(\ltc.output_buffer[24] ),
    .A(\ltc.output_buffer[25] ),
    .X(_0246_));
 sg13g2_xnor2_1 _0988_ (.Y(_0247_),
    .A(\ltc.output_buffer[43] ),
    .B(\ltc.output_buffer[42] ));
 sg13g2_xnor2_1 _0989_ (.Y(_0248_),
    .A(_0246_),
    .B(_0247_));
 sg13g2_xnor2_1 _0990_ (.Y(_0249_),
    .A(_0245_),
    .B(_0248_));
 sg13g2_xnor2_1 _0991_ (.Y(_0250_),
    .A(_0242_),
    .B(_0249_));
 sg13g2_xnor2_1 _0992_ (.Y(_0251_),
    .A(_0235_),
    .B(_0250_));
 sg13g2_xor2_1 _0993_ (.B(\ltc.output_buffer[62] ),
    .A(\ltc.output_buffer[63] ),
    .X(_0252_));
 sg13g2_xor2_1 _0994_ (.B(\ltc.output_buffer[60] ),
    .A(\ltc.output_buffer[61] ),
    .X(_0253_));
 sg13g2_xnor2_1 _0995_ (.Y(_0254_),
    .A(_0252_),
    .B(_0253_));
 sg13g2_xnor2_1 _0996_ (.Y(_0255_),
    .A(\ltc.output_buffer[76] ),
    .B(\ltc.output_buffer[78] ));
 sg13g2_xor2_1 _0997_ (.B(\ltc.output_buffer[77] ),
    .A(\ltc.output_buffer[79] ),
    .X(_0256_));
 sg13g2_xnor2_1 _0998_ (.Y(_0257_),
    .A(_0255_),
    .B(_0256_));
 sg13g2_xnor2_1 _0999_ (.Y(_0258_),
    .A(_0254_),
    .B(_0257_));
 sg13g2_xor2_1 _1000_ (.B(\ltc.output_buffer[66] ),
    .A(\ltc.output_buffer[67] ),
    .X(_0259_));
 sg13g2_xor2_1 _1001_ (.B(\ltc.output_buffer[64] ),
    .A(\ltc.output_buffer[65] ),
    .X(_0260_));
 sg13g2_xnor2_1 _1002_ (.Y(_0261_),
    .A(_0259_),
    .B(_0260_));
 sg13g2_xnor2_1 _1003_ (.Y(_0262_),
    .A(\ltc.output_buffer[71] ),
    .B(\ltc.output_buffer[70] ));
 sg13g2_xor2_1 _1004_ (.B(\ltc.output_buffer[68] ),
    .A(\ltc.output_buffer[69] ),
    .X(_0263_));
 sg13g2_xnor2_1 _1005_ (.Y(_0264_),
    .A(_0262_),
    .B(_0263_));
 sg13g2_xnor2_1 _1006_ (.Y(_0265_),
    .A(_0261_),
    .B(_0264_));
 sg13g2_xnor2_1 _1007_ (.Y(_0266_),
    .A(_0258_),
    .B(_0265_));
 sg13g2_xnor2_1 _1008_ (.Y(_0267_),
    .A(\ltc.output_buffer[51] ),
    .B(\ltc.output_buffer[50] ));
 sg13g2_xor2_1 _1009_ (.B(\ltc.output_buffer[48] ),
    .A(\ltc.output_buffer[49] ),
    .X(_0268_));
 sg13g2_xnor2_1 _1010_ (.Y(_0269_),
    .A(_0267_),
    .B(_0268_));
 sg13g2_xnor2_1 _1011_ (.Y(_0270_),
    .A(\ltc.output_buffer[55] ),
    .B(\ltc.output_buffer[54] ));
 sg13g2_xor2_1 _1012_ (.B(\ltc.output_buffer[53] ),
    .A(\ltc.output_buffer[52] ),
    .X(_0271_));
 sg13g2_xnor2_1 _1013_ (.Y(_0272_),
    .A(_0270_),
    .B(_0271_));
 sg13g2_xnor2_1 _1014_ (.Y(_0273_),
    .A(_0269_),
    .B(_0272_));
 sg13g2_xor2_1 _1015_ (.B(\ltc.output_buffer[72] ),
    .A(\ltc.output_buffer[73] ),
    .X(_0274_));
 sg13g2_xor2_1 _1016_ (.B(\ltc.output_buffer[58] ),
    .A(\ltc.output_buffer[59] ),
    .X(_0275_));
 sg13g2_xnor2_1 _1017_ (.Y(_0276_),
    .A(_0274_),
    .B(_0275_));
 sg13g2_xnor2_1 _1018_ (.Y(_0277_),
    .A(\ltc.output_buffer[75] ),
    .B(\ltc.output_buffer[74] ));
 sg13g2_xor2_1 _1019_ (.B(\ltc.output_buffer[56] ),
    .A(\ltc.output_buffer[57] ),
    .X(_0278_));
 sg13g2_xnor2_1 _1020_ (.Y(_0279_),
    .A(_0277_),
    .B(_0278_));
 sg13g2_xnor2_1 _1021_ (.Y(_0280_),
    .A(_0276_),
    .B(_0279_));
 sg13g2_xnor2_1 _1022_ (.Y(_0281_),
    .A(_0273_),
    .B(_0280_));
 sg13g2_xnor2_1 _1023_ (.Y(_0282_),
    .A(_0266_),
    .B(_0281_));
 sg13g2_xnor2_1 _1024_ (.Y(_0283_),
    .A(_0251_),
    .B(_0282_));
 sg13g2_nand2_1 _1025_ (.Y(_0284_),
    .A(\ltc.output_buffer[20] ),
    .B(net189));
 sg13g2_a21oi_1 _1026_ (.A1(_0220_),
    .A2(_0284_),
    .Y(_0285_),
    .B1(net203));
 sg13g2_o21ai_1 _1027_ (.B1(_0285_),
    .Y(_0286_),
    .A1(_0220_),
    .A2(_0283_));
 sg13g2_a21oi_1 _1028_ (.A1(_0215_),
    .A2(_0286_),
    .Y(_0031_),
    .B1(net215));
 sg13g2_a22oi_1 _1029_ (.Y(_0287_),
    .B1(net179),
    .B2(net354),
    .A2(net203),
    .A1(\ltc.output_buffer[20] ));
 sg13g2_nor2_1 _1030_ (.A(net215),
    .B(net355),
    .Y(_0032_));
 sg13g2_nand3_1 _1031_ (.B(net354),
    .C(net201),
    .A(net224),
    .Y(_0288_));
 sg13g2_nor2_1 _1032_ (.A(net373),
    .B(net187),
    .Y(_0289_));
 sg13g2_o21ai_1 _1033_ (.B1(net196),
    .Y(_0290_),
    .A1(\ltc.output_buffer[22] ),
    .A2(net194));
 sg13g2_o21ai_1 _1034_ (.B1(_0288_),
    .Y(_0033_),
    .A1(_0289_),
    .A2(_0290_));
 sg13g2_nor2_1 _1035_ (.A(\ltc.hrs_d[0] ),
    .B(net186),
    .Y(_0291_));
 sg13g2_o21ai_1 _1036_ (.B1(_0190_),
    .Y(_0292_),
    .A1(\ltc.output_buffer[23] ),
    .A2(net194));
 sg13g2_nand3_1 _1037_ (.B(net382),
    .C(net200),
    .A(net224),
    .Y(_0293_));
 sg13g2_o21ai_1 _1038_ (.B1(_0293_),
    .Y(_0034_),
    .A1(_0291_),
    .A2(_0292_));
 sg13g2_a22oi_1 _1039_ (.Y(_0294_),
    .B1(net179),
    .B2(net253),
    .A2(net201),
    .A1(\ltc.output_buffer[23] ));
 sg13g2_nor2_1 _1040_ (.A(net215),
    .B(net254),
    .Y(_0035_));
 sg13g2_a22oi_1 _1041_ (.Y(_0295_),
    .B1(net185),
    .B2(net305),
    .A2(net205),
    .A1(net253));
 sg13g2_nor2_1 _1042_ (.A(net216),
    .B(_0295_),
    .Y(_0036_));
 sg13g2_a22oi_1 _1043_ (.Y(_0296_),
    .B1(net179),
    .B2(net292),
    .A2(net201),
    .A1(\ltc.output_buffer[25] ));
 sg13g2_nor2_1 _1044_ (.A(net215),
    .B(net293),
    .Y(_0037_));
 sg13g2_a22oi_1 _1045_ (.Y(_0297_),
    .B1(net177),
    .B2(net333),
    .A2(net201),
    .A1(net292));
 sg13g2_nor2_1 _1046_ (.A(net214),
    .B(_0297_),
    .Y(_0038_));
 sg13g2_nand3_1 _1047_ (.B(net333),
    .C(net200),
    .A(net224),
    .Y(_0298_));
 sg13g2_nor2_1 _1048_ (.A(net352),
    .B(net186),
    .Y(_0299_));
 sg13g2_o21ai_1 _1049_ (.B1(net195),
    .Y(_0300_),
    .A1(\ltc.output_buffer[28] ),
    .A2(net191));
 sg13g2_o21ai_1 _1050_ (.B1(_0298_),
    .Y(_0039_),
    .A1(_0299_),
    .A2(_0300_));
 sg13g2_nor2_1 _1051_ (.A(net365),
    .B(net191),
    .Y(_0301_));
 sg13g2_o21ai_1 _1052_ (.B1(net195),
    .Y(_0302_),
    .A1(\ltc.hrs_u[2] ),
    .A2(net186));
 sg13g2_nand3_1 _1053_ (.B(net385),
    .C(net202),
    .A(net223),
    .Y(_0303_));
 sg13g2_o21ai_1 _1054_ (.B1(_0303_),
    .Y(_0040_),
    .A1(_0301_),
    .A2(_0302_));
 sg13g2_nor2_1 _1055_ (.A(net342),
    .B(net191),
    .Y(_0304_));
 sg13g2_o21ai_1 _1056_ (.B1(net195),
    .Y(_0305_),
    .A1(\ltc.hrs_u[1] ),
    .A2(net186));
 sg13g2_nand3_1 _1057_ (.B(net365),
    .C(net202),
    .A(net224),
    .Y(_0306_));
 sg13g2_o21ai_1 _1058_ (.B1(_0306_),
    .Y(_0041_),
    .A1(_0304_),
    .A2(_0305_));
 sg13g2_nor2_1 _1059_ (.A(\ltc.hrs_u[0] ),
    .B(net186),
    .Y(_0307_));
 sg13g2_o21ai_1 _1060_ (.B1(net195),
    .Y(_0308_),
    .A1(\ltc.output_buffer[31] ),
    .A2(net191));
 sg13g2_nand3_1 _1061_ (.B(net342),
    .C(net202),
    .A(net223),
    .Y(_0309_));
 sg13g2_o21ai_1 _1062_ (.B1(_0309_),
    .Y(_0042_),
    .A1(_0307_),
    .A2(_0308_));
 sg13g2_a22oi_1 _1063_ (.Y(_0310_),
    .B1(net177),
    .B2(net278),
    .A2(net199),
    .A1(\ltc.output_buffer[31] ));
 sg13g2_nor2_1 _1064_ (.A(net214),
    .B(net279),
    .Y(_0043_));
 sg13g2_a22oi_1 _1065_ (.Y(_0311_),
    .B1(net177),
    .B2(net317),
    .A2(net199),
    .A1(net278));
 sg13g2_nor2_1 _1066_ (.A(net214),
    .B(_0311_),
    .Y(_0044_));
 sg13g2_a22oi_1 _1067_ (.Y(_0312_),
    .B1(net177),
    .B2(net298),
    .A2(net199),
    .A1(\ltc.output_buffer[33] ));
 sg13g2_nor2_1 _1068_ (.A(net214),
    .B(net299),
    .Y(_0045_));
 sg13g2_a22oi_1 _1069_ (.Y(_0313_),
    .B1(net177),
    .B2(net303),
    .A2(net199),
    .A1(net298));
 sg13g2_nor2_1 _1070_ (.A(net214),
    .B(_0313_),
    .Y(_0046_));
 sg13g2_a22oi_1 _1071_ (.Y(_0314_),
    .B1(net177),
    .B2(net325),
    .A2(net199),
    .A1(net303));
 sg13g2_nor2_1 _1072_ (.A(net214),
    .B(_0314_),
    .Y(_0047_));
 sg13g2_nand3_1 _1073_ (.B(net325),
    .C(net200),
    .A(net223),
    .Y(_0315_));
 sg13g2_nor2_1 _1074_ (.A(\ltc.output_buffer[37] ),
    .B(net191),
    .Y(_0316_));
 sg13g2_o21ai_1 _1075_ (.B1(net195),
    .Y(_0317_),
    .A1(\ltc.min_d[2] ),
    .A2(net186));
 sg13g2_o21ai_1 _1076_ (.B1(_0315_),
    .Y(_0048_),
    .A1(_0316_),
    .A2(_0317_));
 sg13g2_nor2_1 _1077_ (.A(net338),
    .B(net191),
    .Y(_0318_));
 sg13g2_o21ai_1 _1078_ (.B1(net195),
    .Y(_0319_),
    .A1(\ltc.min_d[1] ),
    .A2(net186));
 sg13g2_nand3_1 _1079_ (.B(net346),
    .C(net199),
    .A(net223),
    .Y(_0320_));
 sg13g2_o21ai_1 _1080_ (.B1(_0320_),
    .Y(_0049_),
    .A1(_0318_),
    .A2(_0319_));
 sg13g2_nor2_1 _1081_ (.A(\ltc.min_d[0] ),
    .B(net186),
    .Y(_0321_));
 sg13g2_o21ai_1 _1082_ (.B1(net195),
    .Y(_0322_),
    .A1(\ltc.output_buffer[39] ),
    .A2(net191));
 sg13g2_nand3_1 _1083_ (.B(net338),
    .C(net200),
    .A(net223),
    .Y(_0323_));
 sg13g2_o21ai_1 _1084_ (.B1(_0323_),
    .Y(_0050_),
    .A1(_0321_),
    .A2(_0322_));
 sg13g2_a22oi_1 _1085_ (.Y(_0324_),
    .B1(net178),
    .B2(net255),
    .A2(net199),
    .A1(\ltc.output_buffer[39] ));
 sg13g2_nor2_1 _1086_ (.A(net215),
    .B(net256),
    .Y(_0051_));
 sg13g2_a22oi_1 _1087_ (.Y(_0325_),
    .B1(net177),
    .B2(net309),
    .A2(net199),
    .A1(net255));
 sg13g2_nor2_1 _1088_ (.A(net214),
    .B(_0325_),
    .Y(_0052_));
 sg13g2_a22oi_1 _1089_ (.Y(_0326_),
    .B1(net178),
    .B2(net267),
    .A2(net205),
    .A1(\ltc.output_buffer[41] ));
 sg13g2_nor2_1 _1090_ (.A(net215),
    .B(net268),
    .Y(_0053_));
 sg13g2_a22oi_1 _1091_ (.Y(_0327_),
    .B1(net177),
    .B2(net332),
    .A2(net201),
    .A1(net267));
 sg13g2_nor2_1 _1092_ (.A(net214),
    .B(_0327_),
    .Y(_0054_));
 sg13g2_nand3_1 _1093_ (.B(net332),
    .C(net202),
    .A(net224),
    .Y(_0328_));
 sg13g2_nor2_1 _1094_ (.A(net402),
    .B(net187),
    .Y(_0329_));
 sg13g2_o21ai_1 _1095_ (.B1(net196),
    .Y(_0330_),
    .A1(net313),
    .A2(net192));
 sg13g2_o21ai_1 _1096_ (.B1(_0328_),
    .Y(_0055_),
    .A1(_0329_),
    .A2(_0330_));
 sg13g2_nor2_1 _1097_ (.A(\ltc.output_buffer[45] ),
    .B(net192),
    .Y(_0331_));
 sg13g2_o21ai_1 _1098_ (.B1(net196),
    .Y(_0332_),
    .A1(\ltc.min_u[2] ),
    .A2(net187));
 sg13g2_nand3_1 _1099_ (.B(net313),
    .C(net202),
    .A(net223),
    .Y(_0333_));
 sg13g2_o21ai_1 _1100_ (.B1(_0333_),
    .Y(_0056_),
    .A1(_0331_),
    .A2(_0332_));
 sg13g2_nor2_1 _1101_ (.A(\ltc.output_buffer[46] ),
    .B(net192),
    .Y(_0334_));
 sg13g2_o21ai_1 _1102_ (.B1(net196),
    .Y(_0335_),
    .A1(net318),
    .A2(net187));
 sg13g2_nand3_1 _1103_ (.B(net334),
    .C(net202),
    .A(net226),
    .Y(_0336_));
 sg13g2_o21ai_1 _1104_ (.B1(_0336_),
    .Y(_0057_),
    .A1(_0334_),
    .A2(_0335_));
 sg13g2_nor2_1 _1105_ (.A(\ltc.min_u[0] ),
    .B(net187),
    .Y(_0337_));
 sg13g2_o21ai_1 _1106_ (.B1(net195),
    .Y(_0338_),
    .A1(\ltc.output_buffer[47] ),
    .A2(net191));
 sg13g2_nand3_1 _1107_ (.B(net363),
    .C(net202),
    .A(net226),
    .Y(_0339_));
 sg13g2_o21ai_1 _1108_ (.B1(_0339_),
    .Y(_0058_),
    .A1(_0337_),
    .A2(_0338_));
 sg13g2_a22oi_1 _1109_ (.Y(_0340_),
    .B1(net178),
    .B2(net264),
    .A2(net204),
    .A1(\ltc.output_buffer[47] ));
 sg13g2_nor2_1 _1110_ (.A(net216),
    .B(net265),
    .Y(_0059_));
 sg13g2_a22oi_1 _1111_ (.Y(_0341_),
    .B1(net178),
    .B2(net301),
    .A2(net202),
    .A1(net264));
 sg13g2_nor2_1 _1112_ (.A(_0166_),
    .B(_0341_),
    .Y(_0060_));
 sg13g2_a22oi_1 _1113_ (.Y(_0342_),
    .B1(net179),
    .B2(net247),
    .A2(net203),
    .A1(\ltc.output_buffer[49] ));
 sg13g2_nor2_1 _1114_ (.A(net216),
    .B(net248),
    .Y(_0061_));
 sg13g2_a22oi_1 _1115_ (.Y(_0343_),
    .B1(net179),
    .B2(net306),
    .A2(net203),
    .A1(net247));
 sg13g2_nor2_1 _1116_ (.A(net216),
    .B(_0343_),
    .Y(_0062_));
 sg13g2_nand2_1 _1117_ (.Y(_0344_),
    .A(net306),
    .B(net203));
 sg13g2_nor2_2 _1118_ (.A(net4),
    .B(net3),
    .Y(_0345_));
 sg13g2_and2_2 _1119_ (.A(net4),
    .B(net3),
    .X(_0346_));
 sg13g2_o21ai_1 _1120_ (.B1(_0217_),
    .Y(_0347_),
    .A1(_0345_),
    .A2(_0346_));
 sg13g2_nand2_1 _1121_ (.Y(_0348_),
    .A(net370),
    .B(net189));
 sg13g2_a21oi_1 _1122_ (.A1(_0347_),
    .A2(_0348_),
    .Y(_0349_),
    .B1(net203));
 sg13g2_o21ai_1 _1123_ (.B1(_0349_),
    .Y(_0350_),
    .A1(_0283_),
    .A2(_0347_));
 sg13g2_a21oi_1 _1124_ (.A1(_0344_),
    .A2(_0350_),
    .Y(_0063_),
    .B1(net216));
 sg13g2_nor2_1 _1125_ (.A(net340),
    .B(net192),
    .Y(_0351_));
 sg13g2_o21ai_1 _1126_ (.B1(net196),
    .Y(_0352_),
    .A1(net372),
    .A2(net188));
 sg13g2_nand3_1 _1127_ (.B(net370),
    .C(net204),
    .A(net225),
    .Y(_0353_));
 sg13g2_o21ai_1 _1128_ (.B1(_0353_),
    .Y(_0064_),
    .A1(_0351_),
    .A2(_0352_));
 sg13g2_nor2_1 _1129_ (.A(net310),
    .B(net188),
    .Y(_0354_));
 sg13g2_o21ai_1 _1130_ (.B1(net196),
    .Y(_0355_),
    .A1(\ltc.output_buffer[54] ),
    .A2(net192));
 sg13g2_nand3_1 _1131_ (.B(net340),
    .C(net204),
    .A(net225),
    .Y(_0356_));
 sg13g2_o21ai_1 _1132_ (.B1(_0356_),
    .Y(_0065_),
    .A1(_0354_),
    .A2(_0355_));
 sg13g2_nor2_1 _1133_ (.A(\ltc.sec_d[0] ),
    .B(net188),
    .Y(_0357_));
 sg13g2_o21ai_1 _1134_ (.B1(net196),
    .Y(_0358_),
    .A1(\ltc.output_buffer[55] ),
    .A2(net192));
 sg13g2_nand3_1 _1135_ (.B(net367),
    .C(net204),
    .A(net225),
    .Y(_0359_));
 sg13g2_o21ai_1 _1136_ (.B1(_0359_),
    .Y(_0066_),
    .A1(_0357_),
    .A2(_0358_));
 sg13g2_a22oi_1 _1137_ (.Y(_0360_),
    .B1(net179),
    .B2(net273),
    .A2(net203),
    .A1(\ltc.output_buffer[55] ));
 sg13g2_nor2_1 _1138_ (.A(net216),
    .B(net274),
    .Y(_0067_));
 sg13g2_a22oi_1 _1139_ (.Y(_0361_),
    .B1(net181),
    .B2(net304),
    .A2(net211),
    .A1(net273));
 sg13g2_nor2_1 _1140_ (.A(net218),
    .B(_0361_),
    .Y(_0068_));
 sg13g2_a22oi_1 _1141_ (.Y(_0362_),
    .B1(net181),
    .B2(net316),
    .A2(net209),
    .A1(net304));
 sg13g2_nor2_1 _1142_ (.A(net218),
    .B(_0362_),
    .Y(_0069_));
 sg13g2_a22oi_1 _1143_ (.Y(_0363_),
    .B1(net181),
    .B2(net344),
    .A2(net206),
    .A1(net316));
 sg13g2_nor2_1 _1144_ (.A(net218),
    .B(_0363_),
    .Y(_0070_));
 sg13g2_nand3_1 _1145_ (.B(net344),
    .C(net211),
    .A(net227),
    .Y(_0364_));
 sg13g2_nor2_1 _1146_ (.A(net371),
    .B(net189),
    .Y(_0365_));
 sg13g2_o21ai_1 _1147_ (.B1(net198),
    .Y(_0366_),
    .A1(net327),
    .A2(net193));
 sg13g2_o21ai_1 _1148_ (.B1(_0364_),
    .Y(_0071_),
    .A1(_0365_),
    .A2(_0366_));
 sg13g2_nor2_1 _1149_ (.A(\ltc.sec_u[2] ),
    .B(net189),
    .Y(_0367_));
 sg13g2_o21ai_1 _1150_ (.B1(net197),
    .Y(_0368_),
    .A1(\ltc.output_buffer[61] ),
    .A2(net193));
 sg13g2_nand3_1 _1151_ (.B(net327),
    .C(net211),
    .A(net227),
    .Y(_0369_));
 sg13g2_o21ai_1 _1152_ (.B1(_0369_),
    .Y(_0072_),
    .A1(_0367_),
    .A2(_0368_));
 sg13g2_nor2_1 _1153_ (.A(net360),
    .B(net190),
    .Y(_0370_));
 sg13g2_o21ai_1 _1154_ (.B1(net198),
    .Y(_0371_),
    .A1(net321),
    .A2(net194));
 sg13g2_nand3_1 _1155_ (.B(net387),
    .C(net211),
    .A(net227),
    .Y(_0372_));
 sg13g2_o21ai_1 _1156_ (.B1(_0372_),
    .Y(_0073_),
    .A1(_0370_),
    .A2(_0371_));
 sg13g2_nor2_1 _1157_ (.A(\ltc.sec_u[0] ),
    .B(net190),
    .Y(_0373_));
 sg13g2_o21ai_1 _1158_ (.B1(net197),
    .Y(_0374_),
    .A1(\ltc.output_buffer[63] ),
    .A2(net193));
 sg13g2_nand3_1 _1159_ (.B(net321),
    .C(net211),
    .A(net227),
    .Y(_0375_));
 sg13g2_o21ai_1 _1160_ (.B1(_0375_),
    .Y(_0074_),
    .A1(_0373_),
    .A2(_0374_));
 sg13g2_a22oi_1 _1161_ (.Y(_0376_),
    .B1(net184),
    .B2(net296),
    .A2(net208),
    .A1(\ltc.output_buffer[63] ));
 sg13g2_nor2_1 _1162_ (.A(net220),
    .B(net297),
    .Y(_0075_));
 sg13g2_a22oi_1 _1163_ (.Y(_0377_),
    .B1(net182),
    .B2(net300),
    .A2(net208),
    .A1(net296));
 sg13g2_nor2_1 _1164_ (.A(net220),
    .B(_0377_),
    .Y(_0076_));
 sg13g2_a22oi_1 _1165_ (.Y(_0378_),
    .B1(net182),
    .B2(net249),
    .A2(net208),
    .A1(\ltc.output_buffer[65] ));
 sg13g2_nor2_1 _1166_ (.A(net221),
    .B(net250),
    .Y(_0077_));
 sg13g2_a22oi_1 _1167_ (.Y(_0379_),
    .B1(net182),
    .B2(net315),
    .A2(net208),
    .A1(net249));
 sg13g2_nor2_1 _1168_ (.A(net220),
    .B(_0379_),
    .Y(_0078_));
 sg13g2_a22oi_1 _1169_ (.Y(_0380_),
    .B1(net182),
    .B2(net258),
    .A2(net209),
    .A1(\ltc.output_buffer[67] ));
 sg13g2_nor2_1 _1170_ (.A(net220),
    .B(net259),
    .Y(_0079_));
 sg13g2_a22oi_1 _1171_ (.Y(_0381_),
    .B1(net184),
    .B2(net336),
    .A2(net208),
    .A1(net258));
 sg13g2_nor2_1 _1172_ (.A(net221),
    .B(_0381_),
    .Y(_0080_));
 sg13g2_nand3_1 _1173_ (.B(net336),
    .C(net210),
    .A(net227),
    .Y(_0382_));
 sg13g2_nor2_1 _1174_ (.A(\ltc.frm_d[1] ),
    .B(net190),
    .Y(_0383_));
 sg13g2_o21ai_1 _1175_ (.B1(net197),
    .Y(_0384_),
    .A1(net269),
    .A2(net193));
 sg13g2_o21ai_1 _1176_ (.B1(_0382_),
    .Y(_0081_),
    .A1(_0383_),
    .A2(_0384_));
 sg13g2_nor2_1 _1177_ (.A(\ltc.output_buffer[71] ),
    .B(net193),
    .Y(_0385_));
 sg13g2_o21ai_1 _1178_ (.B1(net197),
    .Y(_0386_),
    .A1(\ltc.frm_d[0] ),
    .A2(net190));
 sg13g2_nand3_1 _1179_ (.B(net269),
    .C(net210),
    .A(net229),
    .Y(_0387_));
 sg13g2_o21ai_1 _1180_ (.B1(_0387_),
    .Y(_0082_),
    .A1(_0385_),
    .A2(_0386_));
 sg13g2_a22oi_1 _1181_ (.Y(_0388_),
    .B1(net184),
    .B2(net294),
    .A2(net210),
    .A1(\ltc.output_buffer[71] ));
 sg13g2_nor2_1 _1182_ (.A(net220),
    .B(net295),
    .Y(_0083_));
 sg13g2_a22oi_1 _1183_ (.Y(_0389_),
    .B1(net184),
    .B2(net283),
    .A2(net210),
    .A1(\ltc.output_buffer[72] ));
 sg13g2_nor2_1 _1184_ (.A(net220),
    .B(net284),
    .Y(_0084_));
 sg13g2_a22oi_1 _1185_ (.Y(_0390_),
    .B1(net184),
    .B2(net271),
    .A2(net210),
    .A1(\ltc.output_buffer[73] ));
 sg13g2_nor2_1 _1186_ (.A(net222),
    .B(net272),
    .Y(_0085_));
 sg13g2_a22oi_1 _1187_ (.Y(_0391_),
    .B1(net184),
    .B2(net345),
    .A2(net210),
    .A1(net271));
 sg13g2_nor2_1 _1188_ (.A(net222),
    .B(_0391_),
    .Y(_0086_));
 sg13g2_nand3_1 _1189_ (.B(net345),
    .C(net210),
    .A(net227),
    .Y(_0392_));
 sg13g2_nor2_1 _1190_ (.A(net356),
    .B(net193),
    .Y(_0393_));
 sg13g2_o21ai_1 _1191_ (.B1(net197),
    .Y(_0394_),
    .A1(net384),
    .A2(net189));
 sg13g2_o21ai_1 _1192_ (.B1(_0392_),
    .Y(_0087_),
    .A1(_0393_),
    .A2(_0394_));
 sg13g2_nor2_1 _1193_ (.A(\ltc.frm_u[2] ),
    .B(net189),
    .Y(_0395_));
 sg13g2_o21ai_1 _1194_ (.B1(net197),
    .Y(_0396_),
    .A1(\ltc.output_buffer[77] ),
    .A2(net193));
 sg13g2_nand3_1 _1195_ (.B(net356),
    .C(net210),
    .A(net227),
    .Y(_0397_));
 sg13g2_o21ai_1 _1196_ (.B1(_0397_),
    .Y(_0088_),
    .A1(_0395_),
    .A2(_0396_));
 sg13g2_nor2_1 _1197_ (.A(\ltc.frm_u[1] ),
    .B(net189),
    .Y(_0398_));
 sg13g2_o21ai_1 _1198_ (.B1(net197),
    .Y(_0399_),
    .A1(\ltc.output_buffer[78] ),
    .A2(net194));
 sg13g2_nand3_1 _1199_ (.B(net358),
    .C(net211),
    .A(net229),
    .Y(_0400_));
 sg13g2_o21ai_1 _1200_ (.B1(_0400_),
    .Y(_0089_),
    .A1(_0398_),
    .A2(_0399_));
 sg13g2_nor2_1 _1201_ (.A(\ltc.output_buffer[79] ),
    .B(net194),
    .Y(_0401_));
 sg13g2_o21ai_1 _1202_ (.B1(net197),
    .Y(_0402_),
    .A1(net212),
    .A2(net189));
 sg13g2_nand3_1 _1203_ (.B(net380),
    .C(net211),
    .A(net229),
    .Y(_0403_));
 sg13g2_o21ai_1 _1204_ (.B1(_0403_),
    .Y(_0090_),
    .A1(_0401_),
    .A2(_0402_));
 sg13g2_nand3b_1 _1205_ (.B(net377),
    .C(\ltc.min_d[2] ),
    .Y(_0404_),
    .A_N(\ltc.min_d[0] ));
 sg13g2_nor2_1 _1206_ (.A(_0161_),
    .B(_0404_),
    .Y(_0405_));
 sg13g2_nor4_1 _1207_ (.A(\ltc.hrs_u[1] ),
    .B(_0160_),
    .C(\ltc.hrs_d[0] ),
    .D(\ltc.hrs_u[0] ),
    .Y(_0406_));
 sg13g2_nand3b_1 _1208_ (.B(net459),
    .C(_0406_),
    .Y(_0407_),
    .A_N(net352));
 sg13g2_nand2_1 _1209_ (.Y(_0408_),
    .A(net418),
    .B(\ltc.hrs_u[1] ));
 sg13g2_nor3_2 _1210_ (.A(\ltc.hrs_u[2] ),
    .B(net409),
    .C(_0408_),
    .Y(_0409_));
 sg13g2_nor2_1 _1211_ (.A(_0404_),
    .B(_0409_),
    .Y(_0410_));
 sg13g2_a21oi_1 _1212_ (.A1(_0407_),
    .A2(_0410_),
    .Y(_0411_),
    .B1(net409));
 sg13g2_o21ai_1 _1213_ (.B1(net223),
    .Y(_0091_),
    .A1(_0405_),
    .A2(_0411_));
 sg13g2_and4_2 _1214_ (.A(net416),
    .B(net329),
    .C(\ltc.frm_counter[0] ),
    .D(\ltc.frm_counter[1] ),
    .X(_0412_));
 sg13g2_nand4_1 _1215_ (.B(\ltc.frm_counter[2] ),
    .C(\ltc.frm_counter[0] ),
    .A(net416),
    .Y(_0413_),
    .D(\ltc.frm_counter[1] ));
 sg13g2_nand2_1 _1216_ (.Y(_0414_),
    .A(\ltc.frm_counter[6] ),
    .B(\ltc.frm_counter[7] ));
 sg13g2_and4_1 _1217_ (.A(\ltc.frm_counter[5] ),
    .B(\ltc.frm_counter[4] ),
    .C(\ltc.frm_counter[6] ),
    .D(\ltc.frm_counter[7] ),
    .X(_0415_));
 sg13g2_nand4_1 _1218_ (.B(\ltc.frm_counter[4] ),
    .C(\ltc.frm_counter[6] ),
    .A(\ltc.frm_counter[5] ),
    .Y(_0416_),
    .D(\ltc.frm_counter[7] ));
 sg13g2_nor2_2 _1219_ (.A(_0413_),
    .B(_0416_),
    .Y(_0417_));
 sg13g2_nand4_1 _1220_ (.B(\ltc.frm_counter[8] ),
    .C(\ltc.frm_counter[10] ),
    .A(\ltc.frm_counter[9] ),
    .Y(_0418_),
    .D(\ltc.frm_counter[11] ));
 sg13g2_nor3_1 _1221_ (.A(_0413_),
    .B(_0416_),
    .C(_0418_),
    .Y(_0419_));
 sg13g2_nor4_2 _1222_ (.A(_0163_),
    .B(_0413_),
    .C(_0416_),
    .Y(_0420_),
    .D(_0418_));
 sg13g2_nand3_1 _1223_ (.B(net454),
    .C(_0420_),
    .A(net213),
    .Y(_0421_));
 sg13g2_and4_2 _1224_ (.A(net213),
    .B(\ltc.frm_counter[14] ),
    .C(\ltc.frm_counter[15] ),
    .D(_0420_),
    .X(_0422_));
 sg13g2_and2_1 _1225_ (.A(\ltc.frm_counter[16] ),
    .B(_0422_),
    .X(_0423_));
 sg13g2_nand3_1 _1226_ (.B(\ltc.frm_counter[17] ),
    .C(_0422_),
    .A(\ltc.frm_counter[16] ),
    .Y(_0424_));
 sg13g2_nand3_1 _1227_ (.B(\ltc.frm_counter[18] ),
    .C(_0423_),
    .A(\ltc.frm_counter[17] ),
    .Y(_0425_));
 sg13g2_xor2_1 _1228_ (.B(_0424_),
    .A(net431),
    .X(_0426_));
 sg13g2_or2_1 _1229_ (.X(_0427_),
    .B(_0426_),
    .A(_0197_));
 sg13g2_xor2_1 _1230_ (.B(_0422_),
    .A(\ltc.frm_counter[16] ),
    .X(_0428_));
 sg13g2_xnor2_1 _1231_ (.Y(_0429_),
    .A(net444),
    .B(_0422_));
 sg13g2_and4_1 _1232_ (.A(\ltc.frm_counter[9] ),
    .B(\ltc.frm_counter[8] ),
    .C(_0412_),
    .D(_0415_),
    .X(_0430_));
 sg13g2_a21oi_1 _1233_ (.A1(\ltc.frm_counter[10] ),
    .A2(_0430_),
    .Y(_0431_),
    .B1(net436));
 sg13g2_or2_1 _1234_ (.X(_0432_),
    .B(net437),
    .A(_0419_));
 sg13g2_xnor2_1 _1235_ (.Y(_0433_),
    .A(net438),
    .B(_0430_));
 sg13g2_and4_1 _1236_ (.A(\ltc.frm_counter[17] ),
    .B(_0428_),
    .C(_0432_),
    .D(_0433_),
    .X(_0434_));
 sg13g2_xor2_1 _1237_ (.B(_0421_),
    .A(net452),
    .X(_0435_));
 sg13g2_and3_1 _1238_ (.X(_0436_),
    .A(net407),
    .B(net460),
    .C(_0412_));
 sg13g2_nand4_1 _1239_ (.B(\ltc.frm_counter[4] ),
    .C(\ltc.frm_counter[6] ),
    .A(\ltc.frm_counter[5] ),
    .Y(_0437_),
    .D(_0412_));
 sg13g2_a21o_1 _1240_ (.A2(_0437_),
    .A1(_0162_),
    .B1(_0417_),
    .X(_0438_));
 sg13g2_xnor2_1 _1241_ (.Y(_0439_),
    .A(net453),
    .B(_0419_));
 sg13g2_a21oi_1 _1242_ (.A1(_0412_),
    .A2(_0415_),
    .Y(_0440_),
    .B1(net445));
 sg13g2_or3_1 _1243_ (.A(_0199_),
    .B(_0430_),
    .C(_0440_),
    .X(_0441_));
 sg13g2_or2_1 _1244_ (.X(_0442_),
    .B(_0420_),
    .A(net213));
 sg13g2_nand4_1 _1245_ (.B(_0439_),
    .C(_0441_),
    .A(_0438_),
    .Y(_0443_),
    .D(_0442_));
 sg13g2_a21o_1 _1246_ (.A2(_0420_),
    .A1(net213),
    .B1(net454),
    .X(_0444_));
 sg13g2_xnor2_1 _1247_ (.Y(_0445_),
    .A(net451),
    .B(_0436_));
 sg13g2_xor2_1 _1248_ (.B(_0417_),
    .A(net455),
    .X(_0446_));
 sg13g2_nand2_1 _1249_ (.Y(_0447_),
    .A(\ltc.frm_counter[4] ),
    .B(_0412_));
 sg13g2_nor4_1 _1250_ (.A(\ltc.frm_counter[5] ),
    .B(net4),
    .C(net3),
    .D(_0447_),
    .Y(_0448_));
 sg13g2_nand3_1 _1251_ (.B(_0446_),
    .C(_0448_),
    .A(_0445_),
    .Y(_0449_));
 sg13g2_nor4_1 _1252_ (.A(_0435_),
    .B(_0443_),
    .C(_0444_),
    .D(_0449_),
    .Y(_0450_));
 sg13g2_nor2_1 _1253_ (.A(net213),
    .B(_0439_),
    .Y(_0451_));
 sg13g2_nor2b_2 _1254_ (.A(\ltc.frm_counter[8] ),
    .B_N(\ltc.frm_counter[9] ),
    .Y(_0452_));
 sg13g2_nand4_1 _1255_ (.B(_0417_),
    .C(_0444_),
    .A(_0218_),
    .Y(_0453_),
    .D(_0452_));
 sg13g2_nor4_1 _1256_ (.A(net213),
    .B(\ltc.frm_counter[15] ),
    .C(_0439_),
    .D(_0453_),
    .Y(_0454_));
 sg13g2_o21ai_1 _1257_ (.B1(_0434_),
    .Y(_0455_),
    .A1(_0450_),
    .A2(_0454_));
 sg13g2_xor2_1 _1258_ (.B(_0423_),
    .A(net457),
    .X(_0456_));
 sg13g2_nand3b_1 _1259_ (.B(\ltc.frm_counter[11] ),
    .C(_0198_),
    .Y(_0457_),
    .A_N(\ltc.frm_counter[10] ));
 sg13g2_nand3_1 _1260_ (.B(_0414_),
    .C(_0452_),
    .A(_0346_),
    .Y(_0458_));
 sg13g2_nor3_1 _1261_ (.A(_0437_),
    .B(_0457_),
    .C(_0458_),
    .Y(_0459_));
 sg13g2_nand4_1 _1262_ (.B(_0451_),
    .C(_0456_),
    .A(_0429_),
    .Y(_0460_),
    .D(_0459_));
 sg13g2_a21o_1 _1263_ (.A2(_0460_),
    .A1(_0455_),
    .B1(_0427_),
    .X(_0461_));
 sg13g2_nand2_1 _1264_ (.Y(_0462_),
    .A(_0438_),
    .B(_0442_));
 sg13g2_nand3_1 _1265_ (.B(_0446_),
    .C(_0448_),
    .A(_0445_),
    .Y(_0463_));
 sg13g2_nand3b_1 _1266_ (.B(_0441_),
    .C(_0439_),
    .Y(_0464_),
    .A_N(_0444_));
 sg13g2_nor4_1 _1267_ (.A(_0435_),
    .B(_0462_),
    .C(_0463_),
    .D(_0464_),
    .Y(_0465_));
 sg13g2_nand3_1 _1268_ (.B(_0417_),
    .C(_0452_),
    .A(_0218_),
    .Y(_0466_));
 sg13g2_nor4_1 _1269_ (.A(net213),
    .B(_0164_),
    .C(_0439_),
    .D(_0466_),
    .Y(_0467_));
 sg13g2_nor2b_1 _1270_ (.A(\ltc.frm_counter[15] ),
    .B_N(_0467_),
    .Y(_0468_));
 sg13g2_o21ai_1 _1271_ (.B1(_0434_),
    .Y(_0469_),
    .A1(_0465_),
    .A2(_0468_));
 sg13g2_nand2_1 _1272_ (.Y(_0470_),
    .A(\ltc.frm_counter[11] ),
    .B(_0452_));
 sg13g2_nand3_1 _1273_ (.B(_0346_),
    .C(_0414_),
    .A(_0198_),
    .Y(_0471_));
 sg13g2_nor4_1 _1274_ (.A(\ltc.frm_counter[10] ),
    .B(_0437_),
    .C(_0470_),
    .D(_0471_),
    .Y(_0472_));
 sg13g2_nand4_1 _1275_ (.B(_0451_),
    .C(_0456_),
    .A(_0429_),
    .Y(_0473_),
    .D(_0472_));
 sg13g2_a21oi_2 _1276_ (.B1(_0427_),
    .Y(_0474_),
    .A2(_0473_),
    .A1(_0469_));
 sg13g2_a21o_2 _1277_ (.A2(_0473_),
    .A1(_0469_),
    .B1(_0427_),
    .X(_0475_));
 sg13g2_nand2_1 _1278_ (.Y(_0476_),
    .A(net229),
    .B(_0461_));
 sg13g2_and3_1 _1279_ (.X(_0092_),
    .A(net229),
    .B(net168),
    .C(_0475_));
 sg13g2_nor2_1 _1280_ (.A(_0203_),
    .B(net423),
    .Y(_0477_));
 sg13g2_nor2_1 _1281_ (.A(net174),
    .B(net424),
    .Y(_0093_));
 sg13g2_and3_1 _1282_ (.X(_0478_),
    .A(net329),
    .B(\ltc.frm_counter[0] ),
    .C(\ltc.frm_counter[1] ));
 sg13g2_a21oi_1 _1283_ (.A1(\ltc.frm_counter[0] ),
    .A2(\ltc.frm_counter[1] ),
    .Y(_0479_),
    .B1(net329));
 sg13g2_nor3_1 _1284_ (.A(net174),
    .B(_0478_),
    .C(net330),
    .Y(_0094_));
 sg13g2_o21ai_1 _1285_ (.B1(_0413_),
    .Y(_0480_),
    .A1(net416),
    .A2(_0478_));
 sg13g2_nor2_1 _1286_ (.A(net176),
    .B(net417),
    .Y(_0095_));
 sg13g2_xnor2_1 _1287_ (.Y(_0481_),
    .A(net425),
    .B(_0412_));
 sg13g2_nor2_1 _1288_ (.A(net174),
    .B(net426),
    .Y(_0096_));
 sg13g2_a21oi_1 _1289_ (.A1(\ltc.frm_counter[4] ),
    .A2(_0412_),
    .Y(_0482_),
    .B1(net407));
 sg13g2_nor3_1 _1290_ (.A(_0436_),
    .B(net174),
    .C(net408),
    .Y(_0097_));
 sg13g2_nor2_1 _1291_ (.A(_0445_),
    .B(net174),
    .Y(_0098_));
 sg13g2_nor2_1 _1292_ (.A(_0438_),
    .B(net174),
    .Y(_0099_));
 sg13g2_nor2b_1 _1293_ (.A(net174),
    .B_N(_0446_),
    .Y(_0100_));
 sg13g2_nor2_1 _1294_ (.A(_0441_),
    .B(net176),
    .Y(_0101_));
 sg13g2_nor2_1 _1295_ (.A(net439),
    .B(net175),
    .Y(_0102_));
 sg13g2_nor2_1 _1296_ (.A(_0432_),
    .B(net175),
    .Y(_0103_));
 sg13g2_nor2_1 _1297_ (.A(_0439_),
    .B(net174),
    .Y(_0104_));
 sg13g2_nand3_1 _1298_ (.B(_0442_),
    .C(_0475_),
    .A(net228),
    .Y(_0483_));
 sg13g2_a21oi_1 _1299_ (.A1(net213),
    .A2(_0420_),
    .Y(_0105_),
    .B1(_0483_));
 sg13g2_and4_1 _1300_ (.A(net228),
    .B(_0421_),
    .C(_0444_),
    .D(_0475_),
    .X(_0106_));
 sg13g2_nor2_1 _1301_ (.A(_0435_),
    .B(net175),
    .Y(_0107_));
 sg13g2_nor2_1 _1302_ (.A(_0429_),
    .B(net175),
    .Y(_0108_));
 sg13g2_and3_1 _1303_ (.X(_0109_),
    .A(net228),
    .B(_0456_),
    .C(_0475_));
 sg13g2_nor2_1 _1304_ (.A(net432),
    .B(net175),
    .Y(_0110_));
 sg13g2_and4_1 _1305_ (.A(\ltc.frm_counter[17] ),
    .B(net461),
    .C(net323),
    .D(_0423_),
    .X(_0484_));
 sg13g2_nor2b_1 _1306_ (.A(net323),
    .B_N(_0425_),
    .Y(_0485_));
 sg13g2_nor3_1 _1307_ (.A(net175),
    .B(_0484_),
    .C(net324),
    .Y(_0111_));
 sg13g2_xnor2_1 _1308_ (.Y(_0486_),
    .A(net404),
    .B(_0484_));
 sg13g2_nor2_1 _1309_ (.A(net175),
    .B(net405),
    .Y(_0112_));
 sg13g2_and3_1 _1310_ (.X(_0487_),
    .A(\ltc.frm_counter[20] ),
    .B(net244),
    .C(_0484_));
 sg13g2_a21oi_1 _1311_ (.A1(\ltc.frm_counter[20] ),
    .A2(_0484_),
    .Y(_0488_),
    .B1(net244));
 sg13g2_nor3_1 _1312_ (.A(net176),
    .B(_0487_),
    .C(net245),
    .Y(_0113_));
 sg13g2_nor2_1 _1313_ (.A(net348),
    .B(_0487_),
    .Y(_0489_));
 sg13g2_and2_1 _1314_ (.A(net348),
    .B(_0487_),
    .X(_0490_));
 sg13g2_nor3_1 _1315_ (.A(net175),
    .B(net349),
    .C(_0490_),
    .Y(_0114_));
 sg13g2_nor2_1 _1316_ (.A(net369),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_and2_1 _1317_ (.A(net369),
    .B(_0490_),
    .X(_0492_));
 sg13g2_nor3_1 _1318_ (.A(net176),
    .B(_0491_),
    .C(_0492_),
    .Y(_0115_));
 sg13g2_nand2_1 _1319_ (.Y(_0493_),
    .A(net223),
    .B(_0407_));
 sg13g2_nor2b_1 _1320_ (.A(_0409_),
    .B_N(\ltc.hrs_d[0] ),
    .Y(_0494_));
 sg13g2_a21oi_1 _1321_ (.A1(net172),
    .A2(_0409_),
    .Y(_0495_),
    .B1(_0494_));
 sg13g2_nor2_1 _1322_ (.A(_0493_),
    .B(net173),
    .Y(_0116_));
 sg13g2_nand2_1 _1323_ (.Y(_0496_),
    .A(net420),
    .B(net419));
 sg13g2_xnor2_1 _1324_ (.Y(_0497_),
    .A(_0160_),
    .B(_0496_));
 sg13g2_nor2_1 _1325_ (.A(_0493_),
    .B(_0497_),
    .Y(_0117_));
 sg13g2_or2_1 _1326_ (.X(_0498_),
    .B(_0493_),
    .A(_0409_));
 sg13g2_and2_1 _1327_ (.A(net394),
    .B(_0405_),
    .X(_0499_));
 sg13g2_nor2_1 _1328_ (.A(net394),
    .B(_0405_),
    .Y(_0500_));
 sg13g2_nor3_1 _1329_ (.A(_0498_),
    .B(_0499_),
    .C(net395),
    .Y(_0118_));
 sg13g2_nand2_1 _1330_ (.Y(_0501_),
    .A(net414),
    .B(_0499_));
 sg13g2_xnor2_1 _1331_ (.Y(_0502_),
    .A(net414),
    .B(_0499_));
 sg13g2_nor2_1 _1332_ (.A(_0498_),
    .B(_0502_),
    .Y(_0119_));
 sg13g2_xor2_1 _1333_ (.B(_0501_),
    .A(net352),
    .X(_0503_));
 sg13g2_nor2_1 _1334_ (.A(_0498_),
    .B(_0503_),
    .Y(_0120_));
 sg13g2_nand2_1 _1335_ (.Y(_0504_),
    .A(\ltc.min_u[3] ),
    .B(net318));
 sg13g2_nor3_2 _1336_ (.A(\ltc.min_u[2] ),
    .B(\ltc.min_u[0] ),
    .C(_0504_),
    .Y(_0505_));
 sg13g2_nor2_1 _1337_ (.A(\ltc.min_d[0] ),
    .B(_0505_),
    .Y(_0506_));
 sg13g2_nand2_1 _1338_ (.Y(_0507_),
    .A(net224),
    .B(_0404_));
 sg13g2_nor2b_1 _1339_ (.A(net232),
    .B_N(_0505_),
    .Y(_0508_));
 sg13g2_nor3_1 _1340_ (.A(_0506_),
    .B(_0507_),
    .C(_0508_),
    .Y(_0121_));
 sg13g2_and3_1 _1341_ (.X(_0509_),
    .A(net377),
    .B(\ltc.min_d[0] ),
    .C(_0505_));
 sg13g2_a21oi_1 _1342_ (.A1(\ltc.min_d[0] ),
    .A2(_0505_),
    .Y(_0510_),
    .B1(net377));
 sg13g2_nor3_1 _1343_ (.A(_0507_),
    .B(_0509_),
    .C(net378),
    .Y(_0122_));
 sg13g2_xnor2_1 _1344_ (.Y(_0511_),
    .A(net397),
    .B(_0509_));
 sg13g2_nor2_1 _1345_ (.A(_0507_),
    .B(net398),
    .Y(_0123_));
 sg13g2_nand2_1 _1346_ (.Y(_0512_),
    .A(\ltc.sec_d[2] ),
    .B(net310));
 sg13g2_nor2_2 _1347_ (.A(\ltc.sec_d[0] ),
    .B(_0512_),
    .Y(_0513_));
 sg13g2_nand2b_2 _1348_ (.Y(_0514_),
    .B(net226),
    .A_N(_0505_));
 sg13g2_nand2b_1 _1349_ (.Y(_0515_),
    .B(_0513_),
    .A_N(net307));
 sg13g2_o21ai_1 _1350_ (.B1(_0515_),
    .Y(_0516_),
    .A1(\ltc.min_u[0] ),
    .A2(_0513_));
 sg13g2_nor2_1 _1351_ (.A(_0514_),
    .B(net308),
    .Y(_0124_));
 sg13g2_and3_1 _1352_ (.X(_0517_),
    .A(net318),
    .B(\ltc.min_u[0] ),
    .C(_0513_));
 sg13g2_a21oi_1 _1353_ (.A1(\ltc.min_u[0] ),
    .A2(_0513_),
    .Y(_0518_),
    .B1(net318));
 sg13g2_nor3_1 _1354_ (.A(_0514_),
    .B(_0517_),
    .C(net319),
    .Y(_0125_));
 sg13g2_nand2_1 _1355_ (.Y(_0519_),
    .A(\ltc.min_u[2] ),
    .B(_0517_));
 sg13g2_xnor2_1 _1356_ (.Y(_0520_),
    .A(net410),
    .B(_0517_));
 sg13g2_nor2_1 _1357_ (.A(_0514_),
    .B(net411),
    .Y(_0126_));
 sg13g2_xor2_1 _1358_ (.B(_0519_),
    .A(net402),
    .X(_0521_));
 sg13g2_nor2_1 _1359_ (.A(_0514_),
    .B(net403),
    .Y(_0127_));
 sg13g2_nand2_1 _1360_ (.Y(_0522_),
    .A(\ltc.sec_u[3] ),
    .B(\ltc.sec_u[1] ));
 sg13g2_nor3_2 _1361_ (.A(\ltc.sec_u[2] ),
    .B(\ltc.sec_u[0] ),
    .C(_0522_),
    .Y(_0523_));
 sg13g2_nor2_1 _1362_ (.A(\ltc.sec_d[0] ),
    .B(_0523_),
    .Y(_0524_));
 sg13g2_o21ai_1 _1363_ (.B1(net225),
    .Y(_0525_),
    .A1(net389),
    .A2(_0512_));
 sg13g2_nor2b_1 _1364_ (.A(net230),
    .B_N(_0523_),
    .Y(_0526_));
 sg13g2_nor3_1 _1365_ (.A(_0524_),
    .B(_0525_),
    .C(_0526_),
    .Y(_0128_));
 sg13g2_and3_1 _1366_ (.X(_0527_),
    .A(net310),
    .B(net389),
    .C(_0523_));
 sg13g2_a21oi_1 _1367_ (.A1(\ltc.sec_d[0] ),
    .A2(_0523_),
    .Y(_0528_),
    .B1(net310));
 sg13g2_nor3_1 _1368_ (.A(_0525_),
    .B(_0527_),
    .C(net311),
    .Y(_0129_));
 sg13g2_xnor2_1 _1369_ (.Y(_0529_),
    .A(net372),
    .B(_0527_));
 sg13g2_nor2_1 _1370_ (.A(net390),
    .B(_0529_),
    .Y(_0130_));
 sg13g2_nor2_1 _1371_ (.A(\ltc.frm_u[1] ),
    .B(\ltc.frm_u[0] ),
    .Y(_0530_));
 sg13g2_nor2_1 _1372_ (.A(\ltc.frm_u[1] ),
    .B(_0219_),
    .Y(_0531_));
 sg13g2_a22oi_1 _1373_ (.Y(_0532_),
    .B1(_0531_),
    .B2(net212),
    .A2(_0530_),
    .A1(_0345_));
 sg13g2_nand2_1 _1374_ (.Y(_0533_),
    .A(\ltc.frm_u[2] ),
    .B(_0159_));
 sg13g2_nand4_1 _1375_ (.B(\ltc.frm_d[0] ),
    .C(_0346_),
    .A(_0157_),
    .Y(_0534_),
    .D(_0530_));
 sg13g2_o21ai_1 _1376_ (.B1(_0534_),
    .Y(_0535_),
    .A1(_0532_),
    .A2(_0533_));
 sg13g2_and3_1 _1377_ (.X(_0536_),
    .A(_0156_),
    .B(\ltc.frm_d[1] ),
    .C(_0535_));
 sg13g2_nand3_1 _1378_ (.B(\ltc.frm_d[1] ),
    .C(_0535_),
    .A(_0156_),
    .Y(_0537_));
 sg13g2_nor2_1 _1379_ (.A(net234),
    .B(_0537_),
    .Y(_0538_));
 sg13g2_nand2b_2 _1380_ (.Y(_0539_),
    .B(net228),
    .A_N(_0523_));
 sg13g2_nor2_1 _1381_ (.A(\ltc.sec_u[0] ),
    .B(_0536_),
    .Y(_0540_));
 sg13g2_nor3_1 _1382_ (.A(_0538_),
    .B(_0539_),
    .C(_0540_),
    .Y(_0131_));
 sg13g2_a21oi_1 _1383_ (.A1(\ltc.sec_u[0] ),
    .A2(_0536_),
    .Y(_0541_),
    .B1(net360));
 sg13g2_and3_1 _1384_ (.X(_0542_),
    .A(net360),
    .B(net406),
    .C(_0536_));
 sg13g2_nor3_1 _1385_ (.A(_0539_),
    .B(net361),
    .C(_0542_),
    .Y(_0132_));
 sg13g2_nand2_1 _1386_ (.Y(_0543_),
    .A(net396),
    .B(_0542_));
 sg13g2_xnor2_1 _1387_ (.Y(_0544_),
    .A(net396),
    .B(_0542_));
 sg13g2_nor2_1 _1388_ (.A(_0539_),
    .B(_0544_),
    .Y(_0133_));
 sg13g2_xor2_1 _1389_ (.B(_0543_),
    .A(net371),
    .X(_0545_));
 sg13g2_nor2_1 _1390_ (.A(_0539_),
    .B(_0545_),
    .Y(_0134_));
 sg13g2_nand2_1 _1391_ (.Y(_0546_),
    .A(net228),
    .B(_0537_));
 sg13g2_nand4_1 _1392_ (.B(_0157_),
    .C(\ltc.frm_u[1] ),
    .A(net384),
    .Y(_0547_),
    .D(_0158_));
 sg13g2_mux2_1 _1393_ (.A0(net350),
    .A1(\ltc.frm_d[0] ),
    .S(_0547_),
    .X(_0548_));
 sg13g2_nor2b_1 _1394_ (.A(_0546_),
    .B_N(net351),
    .Y(_0135_));
 sg13g2_nor2_1 _1395_ (.A(_0159_),
    .B(_0547_),
    .Y(_0549_));
 sg13g2_xnor2_1 _1396_ (.Y(_0550_),
    .A(net400),
    .B(_0549_));
 sg13g2_nor2_1 _1397_ (.A(_0546_),
    .B(net401),
    .Y(_0136_));
 sg13g2_nand3_1 _1398_ (.B(_0537_),
    .C(_0547_),
    .A(_0475_),
    .Y(_0551_));
 sg13g2_o21ai_1 _1399_ (.B1(net228),
    .Y(_0552_),
    .A1(net212),
    .A2(_0474_));
 sg13g2_a21oi_1 _1400_ (.A1(net212),
    .A2(_0551_),
    .Y(_0137_),
    .B1(_0552_));
 sg13g2_nand4_1 _1401_ (.B(_0461_),
    .C(_0537_),
    .A(net428),
    .Y(_0553_),
    .D(_0547_));
 sg13g2_nand2_1 _1402_ (.Y(_0554_),
    .A(net428),
    .B(net212));
 sg13g2_nand3b_1 _1403_ (.B(_0554_),
    .C(_0474_),
    .Y(_0555_),
    .A_N(_0530_));
 sg13g2_a21oi_1 _1404_ (.A1(_0553_),
    .A2(_0555_),
    .Y(_0138_),
    .B1(net222));
 sg13g2_nand3_1 _1405_ (.B(net458),
    .C(net212),
    .A(net415),
    .Y(_0556_));
 sg13g2_nand2b_1 _1406_ (.Y(_0557_),
    .B(_0556_),
    .A_N(_0461_));
 sg13g2_nand2_1 _1407_ (.Y(_0558_),
    .A(_0474_),
    .B(_0556_));
 sg13g2_nand4_1 _1408_ (.B(net428),
    .C(net212),
    .A(_0157_),
    .Y(_0559_),
    .D(_0474_));
 sg13g2_a221oi_1 _1409_ (.B2(_0157_),
    .C1(net222),
    .B1(_0559_),
    .A1(_0551_),
    .Y(_0139_),
    .A2(_0558_));
 sg13g2_a21oi_1 _1410_ (.A1(_0475_),
    .A2(_0547_),
    .Y(_0560_),
    .B1(_0156_));
 sg13g2_or2_1 _1411_ (.X(_0561_),
    .B(_0556_),
    .A(_0475_));
 sg13g2_a221oi_1 _1412_ (.B2(_0156_),
    .C1(net222),
    .B1(_0561_),
    .A1(_0557_),
    .Y(_0140_),
    .A2(_0560_));
 sg13g2_a21oi_1 _1413_ (.A1(_0155_),
    .A2(_0168_),
    .Y(_0562_),
    .B1(_0188_));
 sg13g2_o21ai_1 _1414_ (.B1(net226),
    .Y(_0563_),
    .A1(\ltc.timecode ),
    .A2(_0562_));
 sg13g2_a21oi_1 _1415_ (.A1(_0167_),
    .A2(_0562_),
    .Y(_0141_),
    .B1(_0563_));
 sg13g2_and2_1 _1416_ (.A(\ltc.bit_counter[1] ),
    .B(net391),
    .X(_0564_));
 sg13g2_nand2_1 _1417_ (.Y(_0565_),
    .A(\ltc.bit_counter[2] ),
    .B(_0564_));
 sg13g2_and4_2 _1418_ (.A(\ltc.bit_counter[3] ),
    .B(\ltc.bit_counter[2] ),
    .C(\ltc.bit_counter[1] ),
    .D(\ltc.bit_counter[0] ),
    .X(_0566_));
 sg13g2_nand3_1 _1419_ (.B(\ltc.bit_counter[4] ),
    .C(_0566_),
    .A(\ltc.bit_counter[5] ),
    .Y(_0567_));
 sg13g2_and2_1 _1420_ (.A(\ltc.bit_counter[6] ),
    .B(\ltc.bit_counter[7] ),
    .X(_0568_));
 sg13g2_nand4_1 _1421_ (.B(\ltc.bit_counter[4] ),
    .C(net433),
    .A(\ltc.bit_counter[5] ),
    .Y(_0569_),
    .D(_0566_));
 sg13g2_nand4_1 _1422_ (.B(\ltc.bit_counter[4] ),
    .C(_0566_),
    .A(\ltc.bit_counter[5] ),
    .Y(_0570_),
    .D(_0568_));
 sg13g2_nor2_1 _1423_ (.A(net399),
    .B(_0570_),
    .Y(_0571_));
 sg13g2_xnor2_1 _1424_ (.Y(_0572_),
    .A(net399),
    .B(_0570_));
 sg13g2_nand2_1 _1425_ (.Y(_0573_),
    .A(net440),
    .B(\ltc.bit_counter[9] ));
 sg13g2_nor3_1 _1426_ (.A(_0165_),
    .B(_0570_),
    .C(_0573_),
    .Y(_0574_));
 sg13g2_o21ai_1 _1427_ (.B1(_0165_),
    .Y(_0575_),
    .A1(_0570_),
    .A2(net441));
 sg13g2_nand2b_1 _1428_ (.Y(_0576_),
    .B(net442),
    .A_N(_0574_));
 sg13g2_nand2b_1 _1429_ (.Y(_0577_),
    .B(_0576_),
    .A_N(_0572_));
 sg13g2_xnor2_1 _1430_ (.Y(_0578_),
    .A(net443),
    .B(_0571_));
 sg13g2_xnor2_1 _1431_ (.Y(_0579_),
    .A(net449),
    .B(_0569_));
 sg13g2_xor2_1 _1432_ (.B(_0567_),
    .A(net433),
    .X(_0580_));
 sg13g2_xor2_1 _1433_ (.B(_0566_),
    .A(net456),
    .X(_0581_));
 sg13g2_nor3_1 _1434_ (.A(\ltc.bit_counter[3] ),
    .B(_0219_),
    .C(_0565_),
    .Y(_0582_));
 sg13g2_and4_1 _1435_ (.A(\ltc.bit_counter[5] ),
    .B(_0580_),
    .C(_0581_),
    .D(_0582_),
    .X(_0583_));
 sg13g2_a21oi_1 _1436_ (.A1(_0579_),
    .A2(_0583_),
    .Y(_0584_),
    .B1(_0578_));
 sg13g2_nand4_1 _1437_ (.B(_0346_),
    .C(_0564_),
    .A(_0187_),
    .Y(_0585_),
    .D(_0568_));
 sg13g2_a21oi_1 _1438_ (.A1(\ltc.bit_counter[2] ),
    .A2(_0564_),
    .Y(_0586_),
    .B1(net375));
 sg13g2_xnor2_1 _1439_ (.Y(_0587_),
    .A(net427),
    .B(_0564_));
 sg13g2_and2_1 _1440_ (.A(_0578_),
    .B(_0585_),
    .X(_0588_));
 sg13g2_xnor2_1 _1441_ (.Y(_0589_),
    .A(net412),
    .B(_0574_));
 sg13g2_nand4_1 _1442_ (.B(\ltc.bit_counter[11] ),
    .C(_0185_),
    .A(\ltc.bit_counter[10] ),
    .Y(_0590_),
    .D(_0345_));
 sg13g2_nor4_1 _1443_ (.A(_0577_),
    .B(_0584_),
    .C(_0588_),
    .D(_0589_),
    .Y(_0591_));
 sg13g2_nor3_1 _1444_ (.A(\ltc.bit_counter[3] ),
    .B(_0587_),
    .C(_0590_),
    .Y(_0592_));
 sg13g2_and4_1 _1445_ (.A(\ltc.bit_counter[5] ),
    .B(_0572_),
    .C(_0581_),
    .D(_0592_),
    .X(_0593_));
 sg13g2_a21oi_2 _1446_ (.B1(_0591_),
    .Y(_0594_),
    .A2(_0593_),
    .A1(_0578_));
 sg13g2_nand2_2 _1447_ (.Y(_0595_),
    .A(net228),
    .B(_0594_));
 sg13g2_and3_1 _1448_ (.X(_0142_),
    .A(net225),
    .B(net169),
    .C(_0594_));
 sg13g2_nor3_1 _1449_ (.A(net392),
    .B(_0564_),
    .C(_0595_),
    .Y(_0143_));
 sg13g2_nor2_1 _1450_ (.A(_0587_),
    .B(_0595_),
    .Y(_0144_));
 sg13g2_nor3_1 _1451_ (.A(_0566_),
    .B(net376),
    .C(_0595_),
    .Y(_0145_));
 sg13g2_and3_1 _1452_ (.X(_0146_),
    .A(net225),
    .B(_0581_),
    .C(_0594_));
 sg13g2_a21o_1 _1453_ (.A2(_0566_),
    .A1(\ltc.bit_counter[4] ),
    .B1(net446),
    .X(_0596_));
 sg13g2_and4_1 _1454_ (.A(net225),
    .B(_0567_),
    .C(_0594_),
    .D(net447),
    .X(_0147_));
 sg13g2_nor2_1 _1455_ (.A(_0580_),
    .B(_0595_),
    .Y(_0148_));
 sg13g2_and3_1 _1456_ (.X(_0149_),
    .A(net225),
    .B(net450),
    .C(_0594_));
 sg13g2_nor2_1 _1457_ (.A(_0572_),
    .B(_0595_),
    .Y(_0150_));
 sg13g2_nor2_1 _1458_ (.A(_0578_),
    .B(_0595_),
    .Y(_0151_));
 sg13g2_nor2_1 _1459_ (.A(_0576_),
    .B(_0595_),
    .Y(_0152_));
 sg13g2_nor2_1 _1460_ (.A(net413),
    .B(_0595_),
    .Y(_0153_));
 sg13g2_o21ai_1 _1461_ (.B1(net228),
    .Y(_0597_),
    .A1(net242),
    .A2(_0594_));
 sg13g2_a21oi_1 _1462_ (.A1(_0155_),
    .A2(_0594_),
    .Y(_0154_),
    .B1(_0597_));
 sg13g2_dfrbp_1 _1463_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net105),
    .D(_0011_),
    .Q_N(_0730_),
    .Q(\ltc.output_buffer[0] ));
 sg13g2_dfrbp_1 _1464_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net89),
    .D(_0012_),
    .Q_N(_0729_),
    .Q(\ltc.output_buffer[1] ));
 sg13g2_dfrbp_1 _1465_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net88),
    .D(_0013_),
    .Q_N(_0728_),
    .Q(\ltc.output_buffer[2] ));
 sg13g2_dfrbp_1 _1466_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net87),
    .D(net281),
    .Q_N(_0727_),
    .Q(\ltc.output_buffer[3] ));
 sg13g2_dfrbp_1 _1467_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net86),
    .D(net276),
    .Q_N(_0726_),
    .Q(\ltc.output_buffer[4] ));
 sg13g2_dfrbp_1 _1468_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net85),
    .D(_0016_),
    .Q_N(_0725_),
    .Q(\ltc.output_buffer[5] ));
 sg13g2_dfrbp_1 _1469_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net84),
    .D(net263),
    .Q_N(_0724_),
    .Q(\ltc.output_buffer[6] ));
 sg13g2_dfrbp_1 _1470_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net83),
    .D(_0018_),
    .Q_N(_0723_),
    .Q(\ltc.output_buffer[7] ));
 sg13g2_dfrbp_1 _1471_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net82),
    .D(_0019_),
    .Q_N(_0722_),
    .Q(\ltc.output_buffer[8] ));
 sg13g2_dfrbp_1 _1472_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net81),
    .D(net261),
    .Q_N(_0721_),
    .Q(\ltc.output_buffer[9] ));
 sg13g2_dfrbp_1 _1473_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net80),
    .D(_0021_),
    .Q_N(_0720_),
    .Q(\ltc.output_buffer[10] ));
 sg13g2_dfrbp_1 _1474_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net79),
    .D(_0022_),
    .Q_N(_0719_),
    .Q(\ltc.output_buffer[11] ));
 sg13g2_dfrbp_1 _1475_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net78),
    .D(_0023_),
    .Q_N(_0718_),
    .Q(\ltc.output_buffer[12] ));
 sg13g2_dfrbp_1 _1476_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net77),
    .D(net252),
    .Q_N(_0717_),
    .Q(\ltc.output_buffer[13] ));
 sg13g2_dfrbp_1 _1477_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net76),
    .D(_0025_),
    .Q_N(_0716_),
    .Q(\ltc.output_buffer[14] ));
 sg13g2_dfrbp_1 _1478_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net75),
    .D(_0026_),
    .Q_N(_0715_),
    .Q(\ltc.output_buffer[15] ));
 sg13g2_dfrbp_1 _1479_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net74),
    .D(_0027_),
    .Q_N(_0714_),
    .Q(\ltc.output_buffer[16] ));
 sg13g2_dfrbp_1 _1480_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net73),
    .D(_0028_),
    .Q_N(_0713_),
    .Q(\ltc.output_buffer[17] ));
 sg13g2_dfrbp_1 _1481_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net72),
    .D(_0029_),
    .Q_N(_0712_),
    .Q(\ltc.output_buffer[18] ));
 sg13g2_dfrbp_1 _1482_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net71),
    .D(_0030_),
    .Q_N(_0711_),
    .Q(\ltc.output_buffer[19] ));
 sg13g2_dfrbp_1 _1483_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net70),
    .D(net291),
    .Q_N(_0710_),
    .Q(\ltc.output_buffer[20] ));
 sg13g2_dfrbp_1 _1484_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net69),
    .D(_0032_),
    .Q_N(_0709_),
    .Q(\ltc.output_buffer[21] ));
 sg13g2_dfrbp_1 _1485_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net68),
    .D(net374),
    .Q_N(_0708_),
    .Q(\ltc.output_buffer[22] ));
 sg13g2_dfrbp_1 _1486_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net67),
    .D(net383),
    .Q_N(_0707_),
    .Q(\ltc.output_buffer[23] ));
 sg13g2_dfrbp_1 _1487_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net66),
    .D(_0035_),
    .Q_N(_0706_),
    .Q(\ltc.output_buffer[24] ));
 sg13g2_dfrbp_1 _1488_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net65),
    .D(_0036_),
    .Q_N(_0705_),
    .Q(\ltc.output_buffer[25] ));
 sg13g2_dfrbp_1 _1489_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net64),
    .D(_0037_),
    .Q_N(_0704_),
    .Q(\ltc.output_buffer[26] ));
 sg13g2_dfrbp_1 _1490_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net63),
    .D(_0038_),
    .Q_N(_0703_),
    .Q(\ltc.output_buffer[27] ));
 sg13g2_dfrbp_1 _1491_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net62),
    .D(net353),
    .Q_N(_0702_),
    .Q(\ltc.output_buffer[28] ));
 sg13g2_dfrbp_1 _1492_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net61),
    .D(net386),
    .Q_N(_0701_),
    .Q(\ltc.output_buffer[29] ));
 sg13g2_dfrbp_1 _1493_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net60),
    .D(net366),
    .Q_N(_0700_),
    .Q(\ltc.output_buffer[30] ));
 sg13g2_dfrbp_1 _1494_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net59),
    .D(net343),
    .Q_N(_0699_),
    .Q(\ltc.output_buffer[31] ));
 sg13g2_dfrbp_1 _1495_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net58),
    .D(_0043_),
    .Q_N(_0698_),
    .Q(\ltc.output_buffer[32] ));
 sg13g2_dfrbp_1 _1496_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net57),
    .D(_0044_),
    .Q_N(_0697_),
    .Q(\ltc.output_buffer[33] ));
 sg13g2_dfrbp_1 _1497_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net56),
    .D(_0045_),
    .Q_N(_0696_),
    .Q(\ltc.output_buffer[34] ));
 sg13g2_dfrbp_1 _1498_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net55),
    .D(_0046_),
    .Q_N(_0695_),
    .Q(\ltc.output_buffer[35] ));
 sg13g2_dfrbp_1 _1499_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net54),
    .D(_0047_),
    .Q_N(_0694_),
    .Q(\ltc.output_buffer[36] ));
 sg13g2_dfrbp_1 _1500_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net53),
    .D(net326),
    .Q_N(_0693_),
    .Q(\ltc.output_buffer[37] ));
 sg13g2_dfrbp_1 _1501_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net52),
    .D(net347),
    .Q_N(_0692_),
    .Q(\ltc.output_buffer[38] ));
 sg13g2_dfrbp_1 _1502_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net51),
    .D(net339),
    .Q_N(_0691_),
    .Q(\ltc.output_buffer[39] ));
 sg13g2_dfrbp_1 _1503_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net50),
    .D(_0051_),
    .Q_N(_0690_),
    .Q(\ltc.output_buffer[40] ));
 sg13g2_dfrbp_1 _1504_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net49),
    .D(_0052_),
    .Q_N(_0689_),
    .Q(\ltc.output_buffer[41] ));
 sg13g2_dfrbp_1 _1505_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net48),
    .D(_0053_),
    .Q_N(_0688_),
    .Q(\ltc.output_buffer[42] ));
 sg13g2_dfrbp_1 _1506_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net47),
    .D(_0054_),
    .Q_N(_0687_),
    .Q(\ltc.output_buffer[43] ));
 sg13g2_dfrbp_1 _1507_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net46),
    .D(_0055_),
    .Q_N(_0686_),
    .Q(\ltc.output_buffer[44] ));
 sg13g2_dfrbp_1 _1508_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net45),
    .D(net314),
    .Q_N(_0685_),
    .Q(\ltc.output_buffer[45] ));
 sg13g2_dfrbp_1 _1509_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net44),
    .D(net335),
    .Q_N(_0684_),
    .Q(\ltc.output_buffer[46] ));
 sg13g2_dfrbp_1 _1510_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net43),
    .D(net364),
    .Q_N(_0683_),
    .Q(\ltc.output_buffer[47] ));
 sg13g2_dfrbp_1 _1511_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net42),
    .D(_0059_),
    .Q_N(_0682_),
    .Q(\ltc.output_buffer[48] ));
 sg13g2_dfrbp_1 _1512_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net41),
    .D(_0060_),
    .Q_N(_0681_),
    .Q(\ltc.output_buffer[49] ));
 sg13g2_dfrbp_1 _1513_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net40),
    .D(_0061_),
    .Q_N(_0680_),
    .Q(\ltc.output_buffer[50] ));
 sg13g2_dfrbp_1 _1514_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net39),
    .D(_0062_),
    .Q_N(_0679_),
    .Q(\ltc.output_buffer[51] ));
 sg13g2_dfrbp_1 _1515_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net38),
    .D(_0063_),
    .Q_N(_0678_),
    .Q(\ltc.output_buffer[52] ));
 sg13g2_dfrbp_1 _1516_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net37),
    .D(_0064_),
    .Q_N(_0677_),
    .Q(\ltc.output_buffer[53] ));
 sg13g2_dfrbp_1 _1517_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net36),
    .D(net341),
    .Q_N(_0676_),
    .Q(\ltc.output_buffer[54] ));
 sg13g2_dfrbp_1 _1518_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net35),
    .D(net368),
    .Q_N(_0675_),
    .Q(\ltc.output_buffer[55] ));
 sg13g2_dfrbp_1 _1519_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net34),
    .D(_0067_),
    .Q_N(_0674_),
    .Q(\ltc.output_buffer[56] ));
 sg13g2_dfrbp_1 _1520_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net33),
    .D(_0068_),
    .Q_N(_0673_),
    .Q(\ltc.output_buffer[57] ));
 sg13g2_dfrbp_1 _1521_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net32),
    .D(_0069_),
    .Q_N(_0672_),
    .Q(\ltc.output_buffer[58] ));
 sg13g2_dfrbp_1 _1522_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net31),
    .D(_0070_),
    .Q_N(_0671_),
    .Q(\ltc.output_buffer[59] ));
 sg13g2_dfrbp_1 _1523_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net30),
    .D(_0071_),
    .Q_N(_0670_),
    .Q(\ltc.output_buffer[60] ));
 sg13g2_dfrbp_1 _1524_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net29),
    .D(net328),
    .Q_N(_0669_),
    .Q(\ltc.output_buffer[61] ));
 sg13g2_dfrbp_1 _1525_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net28),
    .D(_0073_),
    .Q_N(_0668_),
    .Q(\ltc.output_buffer[62] ));
 sg13g2_dfrbp_1 _1526_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net27),
    .D(net322),
    .Q_N(_0667_),
    .Q(\ltc.output_buffer[63] ));
 sg13g2_dfrbp_1 _1527_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net26),
    .D(_0075_),
    .Q_N(_0666_),
    .Q(\ltc.output_buffer[64] ));
 sg13g2_dfrbp_1 _1528_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net25),
    .D(_0076_),
    .Q_N(_0665_),
    .Q(\ltc.output_buffer[65] ));
 sg13g2_dfrbp_1 _1529_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net24),
    .D(_0077_),
    .Q_N(_0664_),
    .Q(\ltc.output_buffer[66] ));
 sg13g2_dfrbp_1 _1530_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net23),
    .D(_0078_),
    .Q_N(_0663_),
    .Q(\ltc.output_buffer[67] ));
 sg13g2_dfrbp_1 _1531_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net166),
    .D(_0079_),
    .Q_N(_0662_),
    .Q(\ltc.output_buffer[68] ));
 sg13g2_dfrbp_1 _1532_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net165),
    .D(_0080_),
    .Q_N(_0661_),
    .Q(\ltc.output_buffer[69] ));
 sg13g2_dfrbp_1 _1533_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net164),
    .D(net337),
    .Q_N(_0660_),
    .Q(\ltc.output_buffer[70] ));
 sg13g2_dfrbp_1 _1534_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net163),
    .D(net270),
    .Q_N(_0659_),
    .Q(\ltc.output_buffer[71] ));
 sg13g2_dfrbp_1 _1535_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net162),
    .D(_0083_),
    .Q_N(_0658_),
    .Q(\ltc.output_buffer[72] ));
 sg13g2_dfrbp_1 _1536_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net161),
    .D(_0084_),
    .Q_N(_0657_),
    .Q(\ltc.output_buffer[73] ));
 sg13g2_dfrbp_1 _1537_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net160),
    .D(_0085_),
    .Q_N(_0656_),
    .Q(\ltc.output_buffer[74] ));
 sg13g2_dfrbp_1 _1538_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net159),
    .D(_0086_),
    .Q_N(_0655_),
    .Q(\ltc.output_buffer[75] ));
 sg13g2_dfrbp_1 _1539_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net158),
    .D(_0087_),
    .Q_N(_0654_),
    .Q(\ltc.output_buffer[76] ));
 sg13g2_dfrbp_1 _1540_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net157),
    .D(net357),
    .Q_N(_0653_),
    .Q(\ltc.output_buffer[77] ));
 sg13g2_dfrbp_1 _1541_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net156),
    .D(net359),
    .Q_N(_0652_),
    .Q(\ltc.output_buffer[78] ));
 sg13g2_dfrbp_1 _1542_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net155),
    .D(net381),
    .Q_N(_0651_),
    .Q(\ltc.output_buffer[79] ));
 sg13g2_dfrbp_1 _1543_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net154),
    .D(_0091_),
    .Q_N(_0650_),
    .Q(\ltc.hrs_u[0] ));
 sg13g2_dfrbp_1 _1544_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net152),
    .D(_0092_),
    .Q_N(_0010_),
    .Q(\ltc.frm_counter[0] ));
 sg13g2_dfrbp_1 _1545_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net151),
    .D(_0093_),
    .Q_N(_0649_),
    .Q(\ltc.frm_counter[1] ));
 sg13g2_dfrbp_1 _1546_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net150),
    .D(net331),
    .Q_N(_0648_),
    .Q(\ltc.frm_counter[2] ));
 sg13g2_dfrbp_1 _1547_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net149),
    .D(_0095_),
    .Q_N(_0647_),
    .Q(\ltc.frm_counter[3] ));
 sg13g2_dfrbp_1 _1548_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net148),
    .D(_0096_),
    .Q_N(_0646_),
    .Q(\ltc.frm_counter[4] ));
 sg13g2_dfrbp_1 _1549_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net147),
    .D(_0097_),
    .Q_N(_0645_),
    .Q(\ltc.frm_counter[5] ));
 sg13g2_dfrbp_1 _1550_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net146),
    .D(_0098_),
    .Q_N(_0644_),
    .Q(\ltc.frm_counter[6] ));
 sg13g2_dfrbp_1 _1551_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net145),
    .D(_0099_),
    .Q_N(_0643_),
    .Q(\ltc.frm_counter[7] ));
 sg13g2_dfrbp_1 _1552_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net144),
    .D(_0100_),
    .Q_N(_0642_),
    .Q(\ltc.frm_counter[8] ));
 sg13g2_dfrbp_1 _1553_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net143),
    .D(_0101_),
    .Q_N(_0641_),
    .Q(\ltc.frm_counter[9] ));
 sg13g2_dfrbp_1 _1554_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net142),
    .D(_0102_),
    .Q_N(_0640_),
    .Q(\ltc.frm_counter[10] ));
 sg13g2_dfrbp_1 _1555_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net141),
    .D(_0103_),
    .Q_N(_0639_),
    .Q(\ltc.frm_counter[11] ));
 sg13g2_dfrbp_1 _1556_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net140),
    .D(_0104_),
    .Q_N(_0638_),
    .Q(\ltc.frm_counter[12] ));
 sg13g2_dfrbp_1 _1557_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net139),
    .D(net435),
    .Q_N(_0637_),
    .Q(\ltc.frm_counter[13] ));
 sg13g2_dfrbp_1 _1558_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net138),
    .D(_0106_),
    .Q_N(_0636_),
    .Q(\ltc.frm_counter[14] ));
 sg13g2_dfrbp_1 _1559_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net137),
    .D(_0107_),
    .Q_N(_0635_),
    .Q(\ltc.frm_counter[15] ));
 sg13g2_dfrbp_1 _1560_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net136),
    .D(_0108_),
    .Q_N(_0634_),
    .Q(\ltc.frm_counter[16] ));
 sg13g2_dfrbp_1 _1561_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net135),
    .D(_0109_),
    .Q_N(_0633_),
    .Q(\ltc.frm_counter[17] ));
 sg13g2_dfrbp_1 _1562_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net134),
    .D(_0110_),
    .Q_N(_0632_),
    .Q(\ltc.frm_counter[18] ));
 sg13g2_dfrbp_1 _1563_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net133),
    .D(_0111_),
    .Q_N(_0631_),
    .Q(\ltc.frm_counter[19] ));
 sg13g2_dfrbp_1 _1564_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net132),
    .D(_0112_),
    .Q_N(_0630_),
    .Q(\ltc.frm_counter[20] ));
 sg13g2_dfrbp_1 _1565_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net131),
    .D(net246),
    .Q_N(_0629_),
    .Q(\ltc.frm_counter[21] ));
 sg13g2_dfrbp_1 _1566_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net130),
    .D(_0114_),
    .Q_N(_0628_),
    .Q(\ltc.frm_counter[22] ));
 sg13g2_dfrbp_1 _1567_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net129),
    .D(_0115_),
    .Q_N(_0627_),
    .Q(\ltc.frm_counter[23] ));
 sg13g2_dfrbp_1 _1568_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net128),
    .D(_0116_),
    .Q_N(_0009_),
    .Q(\ltc.hrs_d[0] ));
 sg13g2_dfrbp_1 _1569_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net126),
    .D(net421),
    .Q_N(_0626_),
    .Q(\ltc.hrs_d[1] ));
 sg13g2_dfrbp_1 _1570_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net124),
    .D(_0118_),
    .Q_N(_0625_),
    .Q(\ltc.hrs_u[1] ));
 sg13g2_dfrbp_1 _1571_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net122),
    .D(_0119_),
    .Q_N(_0624_),
    .Q(\ltc.hrs_u[2] ));
 sg13g2_dfrbp_1 _1572_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net120),
    .D(_0120_),
    .Q_N(_0623_),
    .Q(\ltc.hrs_u[3] ));
 sg13g2_dfrbp_1 _1573_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net118),
    .D(net233),
    .Q_N(_0008_),
    .Q(\ltc.min_d[0] ));
 sg13g2_dfrbp_1 _1574_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net116),
    .D(net379),
    .Q_N(_0622_),
    .Q(\ltc.min_d[1] ));
 sg13g2_dfrbp_1 _1575_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net114),
    .D(_0123_),
    .Q_N(_0621_),
    .Q(\ltc.min_d[2] ));
 sg13g2_dfrbp_1 _1576_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net112),
    .D(_0124_),
    .Q_N(_0007_),
    .Q(\ltc.min_u[0] ));
 sg13g2_dfrbp_1 _1577_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net110),
    .D(net320),
    .Q_N(_0620_),
    .Q(\ltc.min_u[1] ));
 sg13g2_dfrbp_1 _1578_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net108),
    .D(_0126_),
    .Q_N(_0619_),
    .Q(\ltc.min_u[2] ));
 sg13g2_dfrbp_1 _1579_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net106),
    .D(_0127_),
    .Q_N(_0618_),
    .Q(\ltc.min_u[3] ));
 sg13g2_dfrbp_1 _1580_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net104),
    .D(net231),
    .Q_N(_0006_),
    .Q(\ltc.sec_d[0] ));
 sg13g2_dfrbp_1 _1581_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net102),
    .D(net312),
    .Q_N(_0617_),
    .Q(\ltc.sec_d[1] ));
 sg13g2_dfrbp_1 _1582_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net100),
    .D(_0130_),
    .Q_N(_0616_),
    .Q(\ltc.sec_d[2] ));
 sg13g2_dfrbp_1 _1583_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net98),
    .D(net235),
    .Q_N(_0005_),
    .Q(\ltc.sec_u[0] ));
 sg13g2_dfrbp_1 _1584_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net96),
    .D(net362),
    .Q_N(_0615_),
    .Q(\ltc.sec_u[1] ));
 sg13g2_dfrbp_1 _1585_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net94),
    .D(_0133_),
    .Q_N(_0614_),
    .Q(\ltc.sec_u[2] ));
 sg13g2_dfrbp_1 _1586_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net92),
    .D(_0134_),
    .Q_N(_0613_),
    .Q(\ltc.sec_u[3] ));
 sg13g2_dfrbp_1 _1587_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net90),
    .D(_0135_),
    .Q_N(_0004_),
    .Q(\ltc.frm_d[0] ));
 sg13g2_dfrbp_1 _1588_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net127),
    .D(_0136_),
    .Q_N(_0612_),
    .Q(\ltc.frm_d[1] ));
 sg13g2_dfrbp_1 _1589_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net123),
    .D(_0137_),
    .Q_N(_0611_),
    .Q(\ltc.frm_u[0] ));
 sg13g2_dfrbp_1 _1590_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net119),
    .D(net429),
    .Q_N(_0610_),
    .Q(\ltc.frm_u[1] ));
 sg13g2_dfrbp_1 _1591_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net115),
    .D(_0139_),
    .Q_N(_0609_),
    .Q(\ltc.frm_u[2] ));
 sg13g2_dfrbp_1 _1592_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net111),
    .D(_0140_),
    .Q_N(_0608_),
    .Q(\ltc.frm_u[3] ));
 sg13g2_dfrbp_1 _1593_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net107),
    .D(net171),
    .Q_N(_0002_),
    .Q(\ltc.timecode ));
 sg13g2_dfrbp_1 _1594_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net103),
    .D(_0142_),
    .Q_N(_0003_),
    .Q(\ltc.bit_counter[0] ));
 sg13g2_dfrbp_1 _1595_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net101),
    .D(net393),
    .Q_N(_0607_),
    .Q(\ltc.bit_counter[1] ));
 sg13g2_dfrbp_1 _1596_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net99),
    .D(_0144_),
    .Q_N(_0606_),
    .Q(\ltc.bit_counter[2] ));
 sg13g2_dfrbp_1 _1597_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net97),
    .D(_0145_),
    .Q_N(_0605_),
    .Q(\ltc.bit_counter[3] ));
 sg13g2_dfrbp_1 _1598_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net95),
    .D(_0146_),
    .Q_N(_0604_),
    .Q(\ltc.bit_counter[4] ));
 sg13g2_dfrbp_1 _1599_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net93),
    .D(_0147_),
    .Q_N(_0603_),
    .Q(\ltc.bit_counter[5] ));
 sg13g2_dfrbp_1 _1600_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net91),
    .D(_0148_),
    .Q_N(_0602_),
    .Q(\ltc.bit_counter[6] ));
 sg13g2_dfrbp_1 _1601_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net153),
    .D(_0149_),
    .Q_N(_0601_),
    .Q(\ltc.bit_counter[7] ));
 sg13g2_dfrbp_1 _1602_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net125),
    .D(_0150_),
    .Q_N(_0001_),
    .Q(\ltc.bit_counter[8] ));
 sg13g2_dfrbp_1 _1603_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net121),
    .D(_0151_),
    .Q_N(_0600_),
    .Q(\ltc.bit_counter[9] ));
 sg13g2_dfrbp_1 _1604_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net117),
    .D(_0152_),
    .Q_N(_0599_),
    .Q(\ltc.bit_counter[10] ));
 sg13g2_dfrbp_1 _1605_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net113),
    .D(_0153_),
    .Q_N(_0598_),
    .Q(\ltc.bit_counter[11] ));
 sg13g2_dfrbp_1 _1606_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net109),
    .D(net243),
    .Q_N(_0000_),
    .Q(\ltc.bit_clk ));
 sg13g2_tiehi _1529__24 (.L_HI(net24));
 sg13g2_tiehi _1528__25 (.L_HI(net25));
 sg13g2_tiehi _1527__26 (.L_HI(net26));
 sg13g2_tiehi _1526__27 (.L_HI(net27));
 sg13g2_tiehi _1525__28 (.L_HI(net28));
 sg13g2_tiehi _1524__29 (.L_HI(net29));
 sg13g2_tiehi _1523__30 (.L_HI(net30));
 sg13g2_tiehi _1522__31 (.L_HI(net31));
 sg13g2_tiehi _1521__32 (.L_HI(net32));
 sg13g2_tiehi _1520__33 (.L_HI(net33));
 sg13g2_tiehi _1519__34 (.L_HI(net34));
 sg13g2_tiehi _1518__35 (.L_HI(net35));
 sg13g2_tiehi _1517__36 (.L_HI(net36));
 sg13g2_tiehi _1516__37 (.L_HI(net37));
 sg13g2_tiehi _1515__38 (.L_HI(net38));
 sg13g2_tiehi _1514__39 (.L_HI(net39));
 sg13g2_tiehi _1513__40 (.L_HI(net40));
 sg13g2_tiehi _1512__41 (.L_HI(net41));
 sg13g2_tiehi _1511__42 (.L_HI(net42));
 sg13g2_tiehi _1510__43 (.L_HI(net43));
 sg13g2_tiehi _1509__44 (.L_HI(net44));
 sg13g2_tiehi _1508__45 (.L_HI(net45));
 sg13g2_tiehi _1507__46 (.L_HI(net46));
 sg13g2_tiehi _1506__47 (.L_HI(net47));
 sg13g2_tiehi _1505__48 (.L_HI(net48));
 sg13g2_tiehi _1504__49 (.L_HI(net49));
 sg13g2_tiehi _1503__50 (.L_HI(net50));
 sg13g2_tiehi _1502__51 (.L_HI(net51));
 sg13g2_tiehi _1501__52 (.L_HI(net52));
 sg13g2_tiehi _1500__53 (.L_HI(net53));
 sg13g2_tiehi _1499__54 (.L_HI(net54));
 sg13g2_tiehi _1498__55 (.L_HI(net55));
 sg13g2_tiehi _1497__56 (.L_HI(net56));
 sg13g2_tiehi _1496__57 (.L_HI(net57));
 sg13g2_tiehi _1495__58 (.L_HI(net58));
 sg13g2_tiehi _1494__59 (.L_HI(net59));
 sg13g2_tiehi _1493__60 (.L_HI(net60));
 sg13g2_tiehi _1492__61 (.L_HI(net61));
 sg13g2_tiehi _1491__62 (.L_HI(net62));
 sg13g2_tiehi _1490__63 (.L_HI(net63));
 sg13g2_tiehi _1489__64 (.L_HI(net64));
 sg13g2_tiehi _1488__65 (.L_HI(net65));
 sg13g2_tiehi _1487__66 (.L_HI(net66));
 sg13g2_tiehi _1486__67 (.L_HI(net67));
 sg13g2_tiehi _1485__68 (.L_HI(net68));
 sg13g2_tiehi _1484__69 (.L_HI(net69));
 sg13g2_tiehi _1483__70 (.L_HI(net70));
 sg13g2_tiehi _1482__71 (.L_HI(net71));
 sg13g2_tiehi _1481__72 (.L_HI(net72));
 sg13g2_tiehi _1480__73 (.L_HI(net73));
 sg13g2_tiehi _1479__74 (.L_HI(net74));
 sg13g2_tiehi _1478__75 (.L_HI(net75));
 sg13g2_tiehi _1477__76 (.L_HI(net76));
 sg13g2_tiehi _1476__77 (.L_HI(net77));
 sg13g2_tiehi _1475__78 (.L_HI(net78));
 sg13g2_tiehi _1474__79 (.L_HI(net79));
 sg13g2_tiehi _1473__80 (.L_HI(net80));
 sg13g2_tiehi _1472__81 (.L_HI(net81));
 sg13g2_tiehi _1471__82 (.L_HI(net82));
 sg13g2_tiehi _1470__83 (.L_HI(net83));
 sg13g2_tiehi _1469__84 (.L_HI(net84));
 sg13g2_tiehi _1468__85 (.L_HI(net85));
 sg13g2_tiehi _1467__86 (.L_HI(net86));
 sg13g2_tiehi _1466__87 (.L_HI(net87));
 sg13g2_tiehi _1465__88 (.L_HI(net88));
 sg13g2_tiehi _1464__89 (.L_HI(net89));
 sg13g2_tiehi _1587__90 (.L_HI(net90));
 sg13g2_tiehi _1600__91 (.L_HI(net91));
 sg13g2_tiehi _1586__92 (.L_HI(net92));
 sg13g2_tiehi _1599__93 (.L_HI(net93));
 sg13g2_tiehi _1585__94 (.L_HI(net94));
 sg13g2_tiehi _1598__95 (.L_HI(net95));
 sg13g2_tiehi _1584__96 (.L_HI(net96));
 sg13g2_tiehi _1597__97 (.L_HI(net97));
 sg13g2_tiehi _1583__98 (.L_HI(net98));
 sg13g2_tiehi _1596__99 (.L_HI(net99));
 sg13g2_tiehi _1582__100 (.L_HI(net100));
 sg13g2_tiehi _1595__101 (.L_HI(net101));
 sg13g2_tiehi _1581__102 (.L_HI(net102));
 sg13g2_tiehi _1594__103 (.L_HI(net103));
 sg13g2_tiehi _1580__104 (.L_HI(net104));
 sg13g2_tiehi _1463__105 (.L_HI(net105));
 sg13g2_tiehi _1579__106 (.L_HI(net106));
 sg13g2_tiehi _1593__107 (.L_HI(net107));
 sg13g2_tiehi _1578__108 (.L_HI(net108));
 sg13g2_tiehi _1606__109 (.L_HI(net109));
 sg13g2_tiehi _1577__110 (.L_HI(net110));
 sg13g2_tiehi _1592__111 (.L_HI(net111));
 sg13g2_tiehi _1576__112 (.L_HI(net112));
 sg13g2_tiehi _1605__113 (.L_HI(net113));
 sg13g2_tiehi _1575__114 (.L_HI(net114));
 sg13g2_tiehi _1591__115 (.L_HI(net115));
 sg13g2_tiehi _1574__116 (.L_HI(net116));
 sg13g2_tiehi _1604__117 (.L_HI(net117));
 sg13g2_tiehi _1573__118 (.L_HI(net118));
 sg13g2_tiehi _1590__119 (.L_HI(net119));
 sg13g2_tiehi _1572__120 (.L_HI(net120));
 sg13g2_tiehi _1603__121 (.L_HI(net121));
 sg13g2_tiehi _1571__122 (.L_HI(net122));
 sg13g2_tiehi _1589__123 (.L_HI(net123));
 sg13g2_tiehi _1570__124 (.L_HI(net124));
 sg13g2_tiehi _1602__125 (.L_HI(net125));
 sg13g2_tiehi _1569__126 (.L_HI(net126));
 sg13g2_tiehi _1588__127 (.L_HI(net127));
 sg13g2_tiehi _1568__128 (.L_HI(net128));
 sg13g2_tiehi _1567__129 (.L_HI(net129));
 sg13g2_tiehi _1566__130 (.L_HI(net130));
 sg13g2_tiehi _1565__131 (.L_HI(net131));
 sg13g2_tiehi _1564__132 (.L_HI(net132));
 sg13g2_tiehi _1563__133 (.L_HI(net133));
 sg13g2_tiehi _1562__134 (.L_HI(net134));
 sg13g2_tiehi _1561__135 (.L_HI(net135));
 sg13g2_tiehi _1560__136 (.L_HI(net136));
 sg13g2_tiehi _1559__137 (.L_HI(net137));
 sg13g2_tiehi _1558__138 (.L_HI(net138));
 sg13g2_tiehi _1557__139 (.L_HI(net139));
 sg13g2_tiehi _1556__140 (.L_HI(net140));
 sg13g2_tiehi _1555__141 (.L_HI(net141));
 sg13g2_tiehi _1554__142 (.L_HI(net142));
 sg13g2_tiehi _1553__143 (.L_HI(net143));
 sg13g2_tiehi _1552__144 (.L_HI(net144));
 sg13g2_tiehi _1551__145 (.L_HI(net145));
 sg13g2_tiehi _1550__146 (.L_HI(net146));
 sg13g2_tiehi _1549__147 (.L_HI(net147));
 sg13g2_tiehi _1548__148 (.L_HI(net148));
 sg13g2_tiehi _1547__149 (.L_HI(net149));
 sg13g2_tiehi _1546__150 (.L_HI(net150));
 sg13g2_tiehi _1545__151 (.L_HI(net151));
 sg13g2_tiehi _1544__152 (.L_HI(net152));
 sg13g2_tiehi _1601__153 (.L_HI(net153));
 sg13g2_tiehi _1543__154 (.L_HI(net154));
 sg13g2_tiehi _1542__155 (.L_HI(net155));
 sg13g2_tiehi _1541__156 (.L_HI(net156));
 sg13g2_tiehi _1540__157 (.L_HI(net157));
 sg13g2_tiehi _1539__158 (.L_HI(net158));
 sg13g2_tiehi _1538__159 (.L_HI(net159));
 sg13g2_tiehi _1537__160 (.L_HI(net160));
 sg13g2_tiehi _1536__161 (.L_HI(net161));
 sg13g2_tiehi _1535__162 (.L_HI(net162));
 sg13g2_tiehi _1534__163 (.L_HI(net163));
 sg13g2_tiehi _1533__164 (.L_HI(net164));
 sg13g2_tiehi _1532__165 (.L_HI(net165));
 sg13g2_tiehi _1531__166 (.L_HI(net166));
 sg13g2_tiehi tt_um_flummer_ltc_167 (.L_HI(net167));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_flummer_ltc_10 (.L_LO(net10));
 sg13g2_tielo tt_um_flummer_ltc_11 (.L_LO(net11));
 sg13g2_tielo tt_um_flummer_ltc_12 (.L_LO(net12));
 sg13g2_tielo tt_um_flummer_ltc_13 (.L_LO(net13));
 sg13g2_tielo tt_um_flummer_ltc_14 (.L_LO(net14));
 sg13g2_tielo tt_um_flummer_ltc_15 (.L_LO(net15));
 sg13g2_tielo tt_um_flummer_ltc_16 (.L_LO(net16));
 sg13g2_tielo tt_um_flummer_ltc_17 (.L_LO(net17));
 sg13g2_tielo tt_um_flummer_ltc_18 (.L_LO(net18));
 sg13g2_tielo tt_um_flummer_ltc_19 (.L_LO(net19));
 sg13g2_tielo tt_um_flummer_ltc_20 (.L_LO(net20));
 sg13g2_tielo tt_um_flummer_ltc_21 (.L_LO(net21));
 sg13g2_tielo tt_um_flummer_ltc_22 (.L_LO(net22));
 sg13g2_tiehi _1530__23 (.L_HI(net23));
 sg13g2_buf_1 _1766_ (.A(\ltc.timecode ),
    .X(uio_out[7]));
 sg13g2_buf_1 _1767_ (.A(uio_in[0]),
    .X(uo_out[1]));
 sg13g2_buf_1 _1768_ (.A(uio_in[1]),
    .X(uo_out[2]));
 sg13g2_buf_1 _1769_ (.A(uio_in[2]),
    .X(uo_out[3]));
 sg13g2_buf_1 _1770_ (.A(uio_in[3]),
    .X(uo_out[4]));
 sg13g2_buf_1 _1771_ (.A(uio_in[4]),
    .X(uo_out[5]));
 sg13g2_buf_1 _1772_ (.A(uio_in[5]),
    .X(uo_out[6]));
 sg13g2_buf_1 _1773_ (.A(uio_in[6]),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout174 (.A(net176),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_0476_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(net178),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(net179),
    .X(net178));
 sg13g2_buf_4 fanout179 (.X(net179),
    .A(net185));
 sg13g2_buf_2 fanout180 (.A(net181),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(net185),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(net184),
    .X(net182));
 sg13g2_buf_1 fanout183 (.A(net184),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(net185),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_0207_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(net187),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(net188),
    .X(net187));
 sg13g2_buf_1 fanout188 (.A(_0205_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_0205_),
    .X(net189));
 sg13g2_buf_1 fanout190 (.A(_0205_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(net192),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(net194),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(net194),
    .X(net193));
 sg13g2_buf_4 fanout194 (.X(net194),
    .A(_0204_));
 sg13g2_buf_2 fanout195 (.A(net196),
    .X(net195));
 sg13g2_buf_4 fanout196 (.X(net196),
    .A(_0190_));
 sg13g2_buf_2 fanout197 (.A(net198),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_0190_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(net201),
    .X(net199));
 sg13g2_buf_1 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(net205),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(net204),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(net204),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(net205),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_0189_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(net209),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(net208),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(net209),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_0189_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(net211),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_0189_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(net430),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(net434),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(net215),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(net216),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_0166_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(net221),
    .X(net217));
 sg13g2_buf_1 fanout218 (.A(net221),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(net220),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(net221),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(net222),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_0166_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(net224),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(rst_n),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(net226),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(rst_n),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(net229),
    .X(net227));
 sg13g2_buf_4 fanout228 (.X(net228),
    .A(net229));
 sg13g2_buf_2 fanout229 (.A(rst_n),
    .X(net229));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_flummer_ltc_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0010_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0003_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0002_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0141_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0009_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0495_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0006_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0128_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0008_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0121_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0005_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0131_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold13 (.A(\ltc.output_buffer[15] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0210_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold15 (.A(\ltc.output_buffer[1] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0208_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold17 (.A(\ltc.output_buffer[14] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0209_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0000_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0154_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold21 (.A(\ltc.frm_counter[21] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0488_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0113_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold24 (.A(\ltc.output_buffer[50] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0342_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold26 (.A(\ltc.output_buffer[66] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0378_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold28 (.A(\ltc.output_buffer[13] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0024_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold30 (.A(\ltc.output_buffer[24] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0294_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold32 (.A(\ltc.output_buffer[40] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0324_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold34 (.A(\ltc.output_buffer[16] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold35 (.A(\ltc.output_buffer[68] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0380_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold37 (.A(\ltc.output_buffer[9] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0020_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold39 (.A(\ltc.output_buffer[6] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0017_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold41 (.A(\ltc.output_buffer[48] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0340_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold43 (.A(\ltc.output_buffer[10] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold44 (.A(\ltc.output_buffer[42] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0326_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold46 (.A(\ltc.output_buffer[70] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0082_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold48 (.A(\ltc.output_buffer[74] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0390_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold50 (.A(\ltc.output_buffer[56] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0360_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold52 (.A(\ltc.output_buffer[4] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0015_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold54 (.A(\ltc.output_buffer[7] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold55 (.A(\ltc.output_buffer[32] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0310_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold57 (.A(\ltc.output_buffer[3] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0014_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold59 (.A(\ltc.output_buffer[2] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold60 (.A(\ltc.output_buffer[73] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0389_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold62 (.A(\ltc.output_buffer[17] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold63 (.A(\ltc.output_buffer[11] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold64 (.A(\ltc.output_buffer[5] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold65 (.A(\ltc.output_buffer[18] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold66 (.A(\ltc.output_buffer[8] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold67 (.A(\ltc.output_buffer[19] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0031_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold69 (.A(\ltc.output_buffer[26] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0296_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold71 (.A(\ltc.output_buffer[72] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0388_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold73 (.A(\ltc.output_buffer[64] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0376_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold75 (.A(\ltc.output_buffer[34] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0312_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold77 (.A(\ltc.output_buffer[65] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold78 (.A(\ltc.output_buffer[49] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold79 (.A(\ltc.output_buffer[12] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold80 (.A(\ltc.output_buffer[35] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold81 (.A(\ltc.output_buffer[57] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold82 (.A(\ltc.output_buffer[25] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold83 (.A(\ltc.output_buffer[51] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0007_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0516_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold86 (.A(\ltc.output_buffer[41] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold87 (.A(\ltc.sec_d[1] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0528_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0129_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold90 (.A(\ltc.output_buffer[44] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0056_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold92 (.A(\ltc.output_buffer[67] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold93 (.A(\ltc.output_buffer[58] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold94 (.A(\ltc.output_buffer[33] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold95 (.A(\ltc.min_u[1] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0518_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0125_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold98 (.A(\ltc.output_buffer[62] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0074_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold100 (.A(\ltc.frm_counter[19] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0485_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold102 (.A(\ltc.output_buffer[36] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0048_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold104 (.A(\ltc.output_buffer[60] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0072_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold106 (.A(\ltc.frm_counter[2] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0479_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0094_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold109 (.A(\ltc.output_buffer[43] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold110 (.A(\ltc.output_buffer[27] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold111 (.A(\ltc.output_buffer[45] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0057_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold113 (.A(\ltc.output_buffer[69] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0081_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold115 (.A(\ltc.output_buffer[38] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0050_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold117 (.A(\ltc.output_buffer[53] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0065_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold119 (.A(\ltc.output_buffer[30] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0042_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold121 (.A(\ltc.output_buffer[59] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold122 (.A(\ltc.output_buffer[75] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold123 (.A(\ltc.output_buffer[37] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0049_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold125 (.A(\ltc.frm_counter[22] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0489_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0004_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0548_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold129 (.A(\ltc.hrs_u[3] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0039_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold131 (.A(\ltc.output_buffer[21] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0287_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold133 (.A(\ltc.output_buffer[76] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0088_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold135 (.A(\ltc.output_buffer[77] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0089_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold137 (.A(\ltc.sec_u[1] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0541_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0132_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold140 (.A(\ltc.output_buffer[46] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0058_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold142 (.A(\ltc.output_buffer[29] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0041_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold144 (.A(\ltc.output_buffer[54] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0066_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold146 (.A(\ltc.frm_counter[23] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold147 (.A(\ltc.output_buffer[52] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold148 (.A(\ltc.sec_u[3] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold149 (.A(\ltc.sec_d[2] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold150 (.A(\ltc.hrs_d[1] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0033_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold152 (.A(\ltc.bit_counter[3] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0586_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold154 (.A(\ltc.min_d[1] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0510_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0122_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold157 (.A(\ltc.output_buffer[78] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0090_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold159 (.A(\ltc.output_buffer[22] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0034_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold161 (.A(\ltc.frm_u[3] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold162 (.A(\ltc.output_buffer[28] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0040_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold164 (.A(\ltc.output_buffer[61] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold165 (.A(\ltc.output_buffer[0] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold166 (.A(\ltc.sec_d[0] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0525_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold168 (.A(\ltc.bit_counter[0] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0184_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0143_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold171 (.A(\ltc.hrs_u[1] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0500_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold173 (.A(\ltc.sec_u[2] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold174 (.A(\ltc.min_d[2] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0511_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0001_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold177 (.A(\ltc.frm_d[1] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0550_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold179 (.A(\ltc.min_u[3] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0521_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold181 (.A(\ltc.frm_counter[20] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0486_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold183 (.A(\ltc.sec_u[0] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold184 (.A(\ltc.frm_counter[5] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0482_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold186 (.A(\ltc.hrs_u[0] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold187 (.A(\ltc.min_u[2] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0520_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold189 (.A(\ltc.bit_counter[11] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0589_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold191 (.A(\ltc.hrs_u[2] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold192 (.A(\ltc.frm_u[2] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold193 (.A(\ltc.frm_counter[3] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0480_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold195 (.A(\ltc.hrs_u[3] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0409_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold197 (.A(\ltc.hrs_d[0] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0117_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold199 (.A(\ltc.frm_counter[0] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0216_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0477_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold202 (.A(\ltc.frm_counter[4] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0481_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold204 (.A(\ltc.bit_counter[2] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold205 (.A(\ltc.frm_u[1] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0138_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold207 (.A(\ltc.frm_u[0] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold208 (.A(\ltc.frm_counter[18] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0426_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold210 (.A(\ltc.bit_counter[6] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold211 (.A(\ltc.frm_counter[13] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0105_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold213 (.A(\ltc.frm_counter[11] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0431_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold215 (.A(\ltc.frm_counter[10] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0433_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold217 (.A(\ltc.bit_counter[8] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0573_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0575_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold220 (.A(\ltc.bit_counter[9] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold221 (.A(\ltc.frm_counter[16] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold222 (.A(\ltc.frm_counter[9] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold223 (.A(\ltc.bit_counter[5] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0596_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold225 (.A(\ltc.frm_counter[7] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold226 (.A(\ltc.bit_counter[7] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0579_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold228 (.A(\ltc.frm_counter[6] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold229 (.A(\ltc.frm_counter[15] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold230 (.A(\ltc.frm_counter[12] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold231 (.A(\ltc.frm_counter[14] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold232 (.A(\ltc.frm_counter[8] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold233 (.A(\ltc.bit_counter[4] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold234 (.A(\ltc.frm_counter[17] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold235 (.A(\ltc.frm_u[1] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold236 (.A(\ltc.hrs_u[2] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold237 (.A(\ltc.frm_counter[4] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold238 (.A(\ltc.frm_counter[18] ),
    .X(net461));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_4 FILLER_4_252 ();
 sg13g2_fill_1 FILLER_4_256 ();
 sg13g2_decap_8 FILLER_4_260 ();
 sg13g2_decap_8 FILLER_4_267 ();
 sg13g2_decap_8 FILLER_4_274 ();
 sg13g2_decap_8 FILLER_4_281 ();
 sg13g2_decap_8 FILLER_4_288 ();
 sg13g2_decap_8 FILLER_4_295 ();
 sg13g2_fill_2 FILLER_4_306 ();
 sg13g2_fill_1 FILLER_4_308 ();
 sg13g2_fill_1 FILLER_4_313 ();
 sg13g2_decap_8 FILLER_4_317 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_decap_4 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_339 ();
 sg13g2_decap_8 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_367 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_fill_1 FILLER_5_217 ();
 sg13g2_fill_2 FILLER_5_227 ();
 sg13g2_fill_1 FILLER_5_229 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_decap_8 FILLER_5_277 ();
 sg13g2_fill_2 FILLER_5_284 ();
 sg13g2_decap_4 FILLER_5_290 ();
 sg13g2_fill_1 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_353 ();
 sg13g2_decap_4 FILLER_5_360 ();
 sg13g2_fill_1 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_369 ();
 sg13g2_decap_4 FILLER_5_376 ();
 sg13g2_decap_8 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_390 ();
 sg13g2_decap_8 FILLER_5_397 ();
 sg13g2_decap_4 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_4 FILLER_6_126 ();
 sg13g2_fill_1 FILLER_6_130 ();
 sg13g2_decap_8 FILLER_6_135 ();
 sg13g2_decap_8 FILLER_6_142 ();
 sg13g2_decap_8 FILLER_6_149 ();
 sg13g2_decap_8 FILLER_6_156 ();
 sg13g2_decap_8 FILLER_6_163 ();
 sg13g2_decap_8 FILLER_6_170 ();
 sg13g2_decap_8 FILLER_6_177 ();
 sg13g2_decap_8 FILLER_6_184 ();
 sg13g2_decap_8 FILLER_6_191 ();
 sg13g2_decap_4 FILLER_6_198 ();
 sg13g2_fill_2 FILLER_6_202 ();
 sg13g2_fill_2 FILLER_6_230 ();
 sg13g2_fill_1 FILLER_6_258 ();
 sg13g2_fill_2 FILLER_6_268 ();
 sg13g2_fill_1 FILLER_6_301 ();
 sg13g2_fill_1 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_4 FILLER_6_404 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_4 FILLER_7_49 ();
 sg13g2_fill_1 FILLER_7_53 ();
 sg13g2_decap_8 FILLER_7_58 ();
 sg13g2_fill_1 FILLER_7_65 ();
 sg13g2_fill_2 FILLER_7_74 ();
 sg13g2_fill_1 FILLER_7_76 ();
 sg13g2_decap_8 FILLER_7_81 ();
 sg13g2_decap_4 FILLER_7_88 ();
 sg13g2_fill_1 FILLER_7_92 ();
 sg13g2_fill_2 FILLER_7_96 ();
 sg13g2_fill_1 FILLER_7_98 ();
 sg13g2_fill_2 FILLER_7_125 ();
 sg13g2_fill_1 FILLER_7_131 ();
 sg13g2_decap_8 FILLER_7_158 ();
 sg13g2_decap_8 FILLER_7_165 ();
 sg13g2_decap_8 FILLER_7_172 ();
 sg13g2_decap_8 FILLER_7_179 ();
 sg13g2_decap_8 FILLER_7_186 ();
 sg13g2_decap_8 FILLER_7_193 ();
 sg13g2_decap_8 FILLER_7_200 ();
 sg13g2_decap_8 FILLER_7_207 ();
 sg13g2_fill_1 FILLER_7_214 ();
 sg13g2_fill_2 FILLER_7_219 ();
 sg13g2_fill_1 FILLER_7_221 ();
 sg13g2_fill_1 FILLER_7_226 ();
 sg13g2_fill_2 FILLER_7_291 ();
 sg13g2_fill_2 FILLER_7_351 ();
 sg13g2_fill_1 FILLER_7_353 ();
 sg13g2_decap_4 FILLER_7_362 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_4 FILLER_8_28 ();
 sg13g2_fill_2 FILLER_8_32 ();
 sg13g2_fill_2 FILLER_8_86 ();
 sg13g2_fill_1 FILLER_8_93 ();
 sg13g2_fill_2 FILLER_8_98 ();
 sg13g2_decap_4 FILLER_8_146 ();
 sg13g2_decap_8 FILLER_8_176 ();
 sg13g2_decap_8 FILLER_8_183 ();
 sg13g2_decap_8 FILLER_8_190 ();
 sg13g2_decap_8 FILLER_8_197 ();
 sg13g2_decap_8 FILLER_8_204 ();
 sg13g2_fill_1 FILLER_8_251 ();
 sg13g2_fill_1 FILLER_8_319 ();
 sg13g2_fill_2 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_366 ();
 sg13g2_decap_4 FILLER_8_373 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_fill_1 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_fill_2 FILLER_9_28 ();
 sg13g2_fill_2 FILLER_9_141 ();
 sg13g2_fill_1 FILLER_9_143 ();
 sg13g2_fill_1 FILLER_9_173 ();
 sg13g2_fill_1 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_4 FILLER_10_21 ();
 sg13g2_fill_2 FILLER_10_74 ();
 sg13g2_fill_1 FILLER_10_76 ();
 sg13g2_fill_2 FILLER_10_107 ();
 sg13g2_fill_1 FILLER_10_132 ();
 sg13g2_fill_2 FILLER_10_142 ();
 sg13g2_fill_1 FILLER_10_144 ();
 sg13g2_fill_2 FILLER_10_162 ();
 sg13g2_fill_2 FILLER_10_190 ();
 sg13g2_fill_2 FILLER_10_214 ();
 sg13g2_fill_1 FILLER_10_224 ();
 sg13g2_fill_1 FILLER_10_260 ();
 sg13g2_fill_2 FILLER_10_287 ();
 sg13g2_fill_2 FILLER_10_298 ();
 sg13g2_fill_2 FILLER_10_332 ();
 sg13g2_fill_1 FILLER_10_351 ();
 sg13g2_fill_1 FILLER_10_378 ();
 sg13g2_decap_4 FILLER_10_388 ();
 sg13g2_fill_1 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_4 FILLER_11_21 ();
 sg13g2_fill_2 FILLER_11_25 ();
 sg13g2_fill_2 FILLER_11_76 ();
 sg13g2_fill_1 FILLER_11_78 ();
 sg13g2_fill_2 FILLER_11_101 ();
 sg13g2_fill_1 FILLER_11_103 ();
 sg13g2_fill_1 FILLER_11_147 ();
 sg13g2_fill_1 FILLER_11_157 ();
 sg13g2_fill_2 FILLER_11_166 ();
 sg13g2_fill_1 FILLER_11_168 ();
 sg13g2_fill_2 FILLER_11_177 ();
 sg13g2_fill_1 FILLER_11_179 ();
 sg13g2_fill_2 FILLER_11_229 ();
 sg13g2_fill_1 FILLER_11_254 ();
 sg13g2_fill_2 FILLER_11_261 ();
 sg13g2_fill_1 FILLER_11_263 ();
 sg13g2_fill_1 FILLER_11_278 ();
 sg13g2_fill_1 FILLER_11_377 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_95 ();
 sg13g2_fill_1 FILLER_12_131 ();
 sg13g2_fill_2 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_197 ();
 sg13g2_fill_1 FILLER_12_204 ();
 sg13g2_fill_2 FILLER_12_252 ();
 sg13g2_fill_1 FILLER_12_310 ();
 sg13g2_fill_2 FILLER_12_328 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_11 ();
 sg13g2_fill_1 FILLER_13_52 ();
 sg13g2_fill_2 FILLER_13_71 ();
 sg13g2_fill_1 FILLER_13_73 ();
 sg13g2_fill_2 FILLER_13_114 ();
 sg13g2_fill_1 FILLER_13_129 ();
 sg13g2_fill_2 FILLER_13_138 ();
 sg13g2_fill_2 FILLER_13_189 ();
 sg13g2_fill_1 FILLER_13_191 ();
 sg13g2_fill_2 FILLER_13_201 ();
 sg13g2_fill_1 FILLER_13_203 ();
 sg13g2_fill_2 FILLER_13_230 ();
 sg13g2_fill_1 FILLER_13_232 ();
 sg13g2_decap_8 FILLER_13_241 ();
 sg13g2_decap_8 FILLER_13_248 ();
 sg13g2_fill_1 FILLER_13_261 ();
 sg13g2_fill_1 FILLER_13_322 ();
 sg13g2_fill_2 FILLER_13_349 ();
 sg13g2_fill_2 FILLER_13_361 ();
 sg13g2_fill_1 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_54 ();
 sg13g2_fill_1 FILLER_14_65 ();
 sg13g2_fill_1 FILLER_14_71 ();
 sg13g2_fill_1 FILLER_14_107 ();
 sg13g2_fill_2 FILLER_14_158 ();
 sg13g2_fill_2 FILLER_14_176 ();
 sg13g2_fill_1 FILLER_14_178 ();
 sg13g2_decap_8 FILLER_14_218 ();
 sg13g2_decap_4 FILLER_14_225 ();
 sg13g2_fill_1 FILLER_14_229 ();
 sg13g2_fill_2 FILLER_14_256 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_fill_1 FILLER_14_291 ();
 sg13g2_fill_2 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_57 ();
 sg13g2_fill_2 FILLER_15_108 ();
 sg13g2_fill_2 FILLER_15_142 ();
 sg13g2_fill_2 FILLER_15_157 ();
 sg13g2_fill_1 FILLER_15_159 ();
 sg13g2_fill_1 FILLER_15_165 ();
 sg13g2_fill_2 FILLER_15_175 ();
 sg13g2_fill_1 FILLER_15_190 ();
 sg13g2_decap_4 FILLER_15_237 ();
 sg13g2_fill_2 FILLER_15_245 ();
 sg13g2_fill_1 FILLER_15_247 ();
 sg13g2_decap_4 FILLER_15_287 ();
 sg13g2_fill_1 FILLER_15_291 ();
 sg13g2_fill_2 FILLER_15_339 ();
 sg13g2_fill_2 FILLER_15_359 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_1 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_54 ();
 sg13g2_fill_2 FILLER_16_109 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_fill_1 FILLER_16_151 ();
 sg13g2_fill_2 FILLER_16_179 ();
 sg13g2_fill_1 FILLER_16_181 ();
 sg13g2_fill_1 FILLER_16_186 ();
 sg13g2_fill_1 FILLER_16_204 ();
 sg13g2_fill_1 FILLER_16_214 ();
 sg13g2_fill_2 FILLER_16_241 ();
 sg13g2_fill_2 FILLER_16_290 ();
 sg13g2_fill_2 FILLER_16_301 ();
 sg13g2_fill_2 FILLER_16_308 ();
 sg13g2_fill_1 FILLER_16_310 ();
 sg13g2_fill_1 FILLER_16_321 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_2 FILLER_17_26 ();
 sg13g2_decap_8 FILLER_17_117 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_134 ();
 sg13g2_fill_2 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_142 ();
 sg13g2_fill_2 FILLER_17_147 ();
 sg13g2_fill_1 FILLER_17_176 ();
 sg13g2_fill_1 FILLER_17_225 ();
 sg13g2_fill_2 FILLER_17_234 ();
 sg13g2_decap_4 FILLER_17_267 ();
 sg13g2_fill_2 FILLER_17_271 ();
 sg13g2_fill_2 FILLER_17_278 ();
 sg13g2_fill_1 FILLER_17_280 ();
 sg13g2_fill_1 FILLER_17_290 ();
 sg13g2_fill_1 FILLER_17_302 ();
 sg13g2_fill_2 FILLER_17_312 ();
 sg13g2_fill_1 FILLER_17_314 ();
 sg13g2_fill_1 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_1 FILLER_18_75 ();
 sg13g2_fill_2 FILLER_18_98 ();
 sg13g2_decap_4 FILLER_18_117 ();
 sg13g2_fill_2 FILLER_18_121 ();
 sg13g2_fill_2 FILLER_18_155 ();
 sg13g2_fill_1 FILLER_18_200 ();
 sg13g2_fill_1 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_4 FILLER_18_232 ();
 sg13g2_decap_4 FILLER_18_241 ();
 sg13g2_fill_1 FILLER_18_269 ();
 sg13g2_fill_2 FILLER_18_296 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_fill_2 FILLER_18_343 ();
 sg13g2_fill_1 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_2 FILLER_19_26 ();
 sg13g2_fill_2 FILLER_19_51 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_4 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_130 ();
 sg13g2_fill_2 FILLER_19_163 ();
 sg13g2_decap_8 FILLER_19_173 ();
 sg13g2_fill_2 FILLER_19_180 ();
 sg13g2_decap_4 FILLER_19_198 ();
 sg13g2_decap_4 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_225 ();
 sg13g2_fill_2 FILLER_19_271 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_4 ();
 sg13g2_decap_4 FILLER_20_101 ();
 sg13g2_fill_2 FILLER_20_123 ();
 sg13g2_fill_1 FILLER_20_125 ();
 sg13g2_decap_8 FILLER_20_135 ();
 sg13g2_decap_4 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_176 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_decap_4 FILLER_20_193 ();
 sg13g2_fill_2 FILLER_20_197 ();
 sg13g2_fill_2 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_280 ();
 sg13g2_fill_2 FILLER_20_324 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_4 ();
 sg13g2_fill_2 FILLER_21_48 ();
 sg13g2_fill_2 FILLER_21_74 ();
 sg13g2_fill_1 FILLER_21_141 ();
 sg13g2_fill_2 FILLER_21_187 ();
 sg13g2_decap_4 FILLER_21_197 ();
 sg13g2_fill_2 FILLER_21_201 ();
 sg13g2_fill_1 FILLER_21_233 ();
 sg13g2_decap_4 FILLER_21_265 ();
 sg13g2_fill_2 FILLER_21_295 ();
 sg13g2_fill_1 FILLER_21_297 ();
 sg13g2_fill_2 FILLER_21_302 ();
 sg13g2_fill_1 FILLER_21_304 ();
 sg13g2_fill_1 FILLER_21_326 ();
 sg13g2_decap_4 FILLER_21_341 ();
 sg13g2_fill_1 FILLER_21_345 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_fill_2 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_58 ();
 sg13g2_fill_2 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_123 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_decap_4 FILLER_22_198 ();
 sg13g2_fill_2 FILLER_22_202 ();
 sg13g2_decap_4 FILLER_22_209 ();
 sg13g2_fill_2 FILLER_22_226 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_decap_4 FILLER_22_256 ();
 sg13g2_fill_1 FILLER_22_260 ();
 sg13g2_fill_2 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_360 ();
 sg13g2_decap_8 FILLER_22_367 ();
 sg13g2_decap_8 FILLER_22_374 ();
 sg13g2_decap_8 FILLER_22_381 ();
 sg13g2_decap_8 FILLER_22_388 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_decap_4 FILLER_23_30 ();
 sg13g2_fill_1 FILLER_23_42 ();
 sg13g2_fill_2 FILLER_23_69 ();
 sg13g2_fill_1 FILLER_23_71 ();
 sg13g2_fill_2 FILLER_23_165 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_fill_2 FILLER_23_200 ();
 sg13g2_fill_1 FILLER_23_214 ();
 sg13g2_fill_1 FILLER_23_224 ();
 sg13g2_decap_4 FILLER_23_254 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_fill_2 FILLER_23_281 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_fill_1 FILLER_23_289 ();
 sg13g2_fill_2 FILLER_23_317 ();
 sg13g2_fill_1 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_359 ();
 sg13g2_decap_8 FILLER_23_366 ();
 sg13g2_decap_8 FILLER_23_373 ();
 sg13g2_decap_8 FILLER_23_380 ();
 sg13g2_decap_8 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_11 ();
 sg13g2_fill_2 FILLER_24_77 ();
 sg13g2_fill_1 FILLER_24_79 ();
 sg13g2_fill_2 FILLER_24_99 ();
 sg13g2_fill_2 FILLER_24_124 ();
 sg13g2_fill_1 FILLER_24_126 ();
 sg13g2_fill_1 FILLER_24_137 ();
 sg13g2_fill_2 FILLER_24_158 ();
 sg13g2_fill_2 FILLER_24_212 ();
 sg13g2_fill_2 FILLER_24_244 ();
 sg13g2_fill_1 FILLER_24_246 ();
 sg13g2_fill_1 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_decap_4 FILLER_24_356 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_fill_1 FILLER_25_78 ();
 sg13g2_fill_2 FILLER_25_101 ();
 sg13g2_fill_1 FILLER_25_133 ();
 sg13g2_fill_2 FILLER_25_173 ();
 sg13g2_fill_1 FILLER_25_195 ();
 sg13g2_fill_1 FILLER_25_221 ();
 sg13g2_fill_1 FILLER_25_249 ();
 sg13g2_fill_2 FILLER_25_291 ();
 sg13g2_fill_2 FILLER_25_319 ();
 sg13g2_fill_1 FILLER_25_321 ();
 sg13g2_fill_2 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_330 ();
 sg13g2_fill_2 FILLER_25_367 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_fill_2 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_67 ();
 sg13g2_fill_2 FILLER_26_138 ();
 sg13g2_fill_1 FILLER_26_140 ();
 sg13g2_fill_2 FILLER_26_159 ();
 sg13g2_fill_1 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_188 ();
 sg13g2_fill_1 FILLER_26_232 ();
 sg13g2_fill_1 FILLER_26_281 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_fill_2 FILLER_26_332 ();
 sg13g2_fill_2 FILLER_26_353 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_4 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_69 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_fill_1 FILLER_27_142 ();
 sg13g2_fill_2 FILLER_27_170 ();
 sg13g2_fill_1 FILLER_27_172 ();
 sg13g2_fill_1 FILLER_27_177 ();
 sg13g2_fill_2 FILLER_27_212 ();
 sg13g2_fill_1 FILLER_27_214 ();
 sg13g2_fill_2 FILLER_27_223 ();
 sg13g2_fill_2 FILLER_27_235 ();
 sg13g2_fill_2 FILLER_27_242 ();
 sg13g2_fill_1 FILLER_27_244 ();
 sg13g2_fill_1 FILLER_27_257 ();
 sg13g2_fill_2 FILLER_27_345 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_4 FILLER_28_49 ();
 sg13g2_fill_2 FILLER_28_61 ();
 sg13g2_fill_2 FILLER_28_316 ();
 sg13g2_fill_2 FILLER_28_323 ();
 sg13g2_fill_1 FILLER_28_330 ();
 sg13g2_fill_2 FILLER_28_345 ();
 sg13g2_fill_1 FILLER_28_393 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_4 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_67 ();
 sg13g2_fill_2 FILLER_29_87 ();
 sg13g2_fill_1 FILLER_29_89 ();
 sg13g2_fill_2 FILLER_29_113 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_fill_2 FILLER_29_180 ();
 sg13g2_fill_1 FILLER_29_182 ();
 sg13g2_decap_4 FILLER_29_209 ();
 sg13g2_fill_2 FILLER_29_213 ();
 sg13g2_fill_2 FILLER_29_250 ();
 sg13g2_fill_2 FILLER_29_290 ();
 sg13g2_decap_8 FILLER_29_296 ();
 sg13g2_decap_4 FILLER_29_303 ();
 sg13g2_fill_2 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_fill_2 FILLER_30_84 ();
 sg13g2_fill_1 FILLER_30_86 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_fill_2 FILLER_30_158 ();
 sg13g2_fill_2 FILLER_30_190 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_fill_1 FILLER_30_219 ();
 sg13g2_fill_1 FILLER_30_232 ();
 sg13g2_fill_2 FILLER_30_242 ();
 sg13g2_fill_1 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_260 ();
 sg13g2_decap_4 FILLER_30_281 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_decap_8 FILLER_30_296 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_4 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_139 ();
 sg13g2_fill_2 FILLER_31_167 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_fill_2 FILLER_31_205 ();
 sg13g2_fill_1 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_fill_1 FILLER_31_243 ();
 sg13g2_fill_2 FILLER_31_270 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_decap_4 FILLER_31_284 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_fill_1 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_fill_1 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_134 ();
 sg13g2_fill_1 FILLER_32_136 ();
 sg13g2_fill_2 FILLER_32_154 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_fill_1 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_4 FILLER_32_210 ();
 sg13g2_fill_2 FILLER_32_214 ();
 sg13g2_decap_4 FILLER_32_220 ();
 sg13g2_fill_2 FILLER_32_282 ();
 sg13g2_fill_1 FILLER_32_284 ();
 sg13g2_decap_4 FILLER_32_304 ();
 sg13g2_fill_1 FILLER_32_318 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_fill_2 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_139 ();
 sg13g2_fill_1 FILLER_33_166 ();
 sg13g2_fill_1 FILLER_33_191 ();
 sg13g2_fill_1 FILLER_33_277 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_307 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_4 FILLER_34_104 ();
 sg13g2_fill_2 FILLER_34_108 ();
 sg13g2_fill_2 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_212 ();
 sg13g2_decap_4 FILLER_34_218 ();
 sg13g2_fill_2 FILLER_34_303 ();
 sg13g2_fill_1 FILLER_34_305 ();
 sg13g2_fill_2 FILLER_34_329 ();
 sg13g2_fill_1 FILLER_34_339 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_4 FILLER_35_98 ();
 sg13g2_fill_2 FILLER_35_102 ();
 sg13g2_fill_2 FILLER_35_114 ();
 sg13g2_fill_2 FILLER_35_132 ();
 sg13g2_fill_1 FILLER_35_169 ();
 sg13g2_fill_1 FILLER_35_193 ();
 sg13g2_fill_2 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_257 ();
 sg13g2_fill_2 FILLER_35_283 ();
 sg13g2_fill_2 FILLER_35_298 ();
 sg13g2_fill_1 FILLER_35_390 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_fill_2 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_135 ();
 sg13g2_fill_2 FILLER_36_181 ();
 sg13g2_decap_8 FILLER_36_223 ();
 sg13g2_fill_2 FILLER_36_230 ();
 sg13g2_fill_1 FILLER_36_232 ();
 sg13g2_fill_1 FILLER_36_237 ();
 sg13g2_fill_2 FILLER_36_273 ();
 sg13g2_fill_2 FILLER_36_306 ();
 sg13g2_fill_1 FILLER_36_308 ();
 sg13g2_fill_2 FILLER_36_346 ();
 sg13g2_fill_1 FILLER_36_348 ();
 sg13g2_fill_2 FILLER_36_377 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_4 FILLER_37_147 ();
 sg13g2_fill_2 FILLER_37_155 ();
 sg13g2_fill_2 FILLER_37_171 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_decap_8 FILLER_37_223 ();
 sg13g2_fill_2 FILLER_37_230 ();
 sg13g2_fill_2 FILLER_37_258 ();
 sg13g2_fill_1 FILLER_37_283 ();
 sg13g2_fill_1 FILLER_37_310 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_202 ();
 sg13g2_decap_4 FILLER_38_211 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_240 ();
 sg13g2_fill_1 FILLER_38_242 ();
 sg13g2_fill_2 FILLER_38_247 ();
 sg13g2_fill_1 FILLER_38_249 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net167;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[2] = net18;
 assign uio_out[3] = net19;
 assign uio_out[4] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
endmodule

module tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire fail;
 wire \i_soc.cnt[0] ;
 wire \i_soc.cnt[1] ;
 wire \i_soc.cnt[2] ;
 wire \i_soc.cnt[3] ;
 wire \i_soc.cnt[4] ;
 wire \i_soc.cnt[5] ;
 wire \i_soc.cnt[6] ;
 wire \i_soc.cnt[7] ;
 wire \i_soc.cpu.pc[2] ;
 wire \i_soc.cpu.pc[3] ;
 wire \i_soc.cpu.pc[4] ;
 wire \i_soc.cpu.pc[5] ;
 wire \i_soc.cpu.rd0[0] ;
 wire \i_soc.cpu.rd0[10] ;
 wire \i_soc.cpu.rd0[11] ;
 wire \i_soc.cpu.rd0[12] ;
 wire \i_soc.cpu.rd0[13] ;
 wire \i_soc.cpu.rd0[14] ;
 wire \i_soc.cpu.rd0[15] ;
 wire \i_soc.cpu.rd0[16] ;
 wire \i_soc.cpu.rd0[17] ;
 wire \i_soc.cpu.rd0[18] ;
 wire \i_soc.cpu.rd0[19] ;
 wire \i_soc.cpu.rd0[1] ;
 wire \i_soc.cpu.rd0[20] ;
 wire \i_soc.cpu.rd0[21] ;
 wire \i_soc.cpu.rd0[22] ;
 wire \i_soc.cpu.rd0[23] ;
 wire \i_soc.cpu.rd0[24] ;
 wire \i_soc.cpu.rd0[25] ;
 wire \i_soc.cpu.rd0[26] ;
 wire \i_soc.cpu.rd0[27] ;
 wire \i_soc.cpu.rd0[28] ;
 wire \i_soc.cpu.rd0[29] ;
 wire \i_soc.cpu.rd0[2] ;
 wire \i_soc.cpu.rd0[30] ;
 wire \i_soc.cpu.rd0[31] ;
 wire \i_soc.cpu.rd0[3] ;
 wire \i_soc.cpu.rd0[4] ;
 wire \i_soc.cpu.rd0[5] ;
 wire \i_soc.cpu.rd0[6] ;
 wire \i_soc.cpu.rd0[7] ;
 wire \i_soc.cpu.rd0[8] ;
 wire \i_soc.cpu.rd0[9] ;
 wire \i_soc.cpu.rf.rf[0][0] ;
 wire \i_soc.cpu.rf.rf[0][1] ;
 wire \i_soc.cpu.rf.rf[0][2] ;
 wire \i_soc.cpu.rf.rf[0][30] ;
 wire \i_soc.cpu.rf.rf[0][3] ;
 wire \i_soc.cpu.rf.rf[11][0] ;
 wire \i_soc.cpu.rf.rf[11][10] ;
 wire \i_soc.cpu.rf.rf[11][11] ;
 wire \i_soc.cpu.rf.rf[11][12] ;
 wire \i_soc.cpu.rf.rf[11][13] ;
 wire \i_soc.cpu.rf.rf[11][14] ;
 wire \i_soc.cpu.rf.rf[11][15] ;
 wire \i_soc.cpu.rf.rf[11][16] ;
 wire \i_soc.cpu.rf.rf[11][17] ;
 wire \i_soc.cpu.rf.rf[11][18] ;
 wire \i_soc.cpu.rf.rf[11][19] ;
 wire \i_soc.cpu.rf.rf[11][1] ;
 wire \i_soc.cpu.rf.rf[11][20] ;
 wire \i_soc.cpu.rf.rf[11][21] ;
 wire \i_soc.cpu.rf.rf[11][22] ;
 wire \i_soc.cpu.rf.rf[11][24] ;
 wire \i_soc.cpu.rf.rf[11][25] ;
 wire \i_soc.cpu.rf.rf[11][26] ;
 wire \i_soc.cpu.rf.rf[11][27] ;
 wire \i_soc.cpu.rf.rf[11][28] ;
 wire \i_soc.cpu.rf.rf[11][29] ;
 wire \i_soc.cpu.rf.rf[11][2] ;
 wire \i_soc.cpu.rf.rf[11][30] ;
 wire \i_soc.cpu.rf.rf[11][31] ;
 wire \i_soc.cpu.rf.rf[11][3] ;
 wire \i_soc.cpu.rf.rf[11][4] ;
 wire \i_soc.cpu.rf.rf[11][5] ;
 wire \i_soc.cpu.rf.rf[11][6] ;
 wire \i_soc.cpu.rf.rf[11][7] ;
 wire \i_soc.cpu.rf.rf[11][8] ;
 wire \i_soc.cpu.rf.rf[11][9] ;
 wire \i_soc.cpu.rf.rf[1][0] ;
 wire \i_soc.cpu.rf.rf[1][10] ;
 wire \i_soc.cpu.rf.rf[1][11] ;
 wire \i_soc.cpu.rf.rf[1][12] ;
 wire \i_soc.cpu.rf.rf[1][13] ;
 wire \i_soc.cpu.rf.rf[1][14] ;
 wire \i_soc.cpu.rf.rf[1][15] ;
 wire \i_soc.cpu.rf.rf[1][16] ;
 wire \i_soc.cpu.rf.rf[1][17] ;
 wire \i_soc.cpu.rf.rf[1][18] ;
 wire \i_soc.cpu.rf.rf[1][19] ;
 wire \i_soc.cpu.rf.rf[1][1] ;
 wire \i_soc.cpu.rf.rf[1][20] ;
 wire \i_soc.cpu.rf.rf[1][21] ;
 wire \i_soc.cpu.rf.rf[1][22] ;
 wire \i_soc.cpu.rf.rf[1][23] ;
 wire \i_soc.cpu.rf.rf[1][24] ;
 wire \i_soc.cpu.rf.rf[1][25] ;
 wire \i_soc.cpu.rf.rf[1][26] ;
 wire \i_soc.cpu.rf.rf[1][27] ;
 wire \i_soc.cpu.rf.rf[1][28] ;
 wire \i_soc.cpu.rf.rf[1][29] ;
 wire \i_soc.cpu.rf.rf[1][2] ;
 wire \i_soc.cpu.rf.rf[1][30] ;
 wire \i_soc.cpu.rf.rf[1][31] ;
 wire \i_soc.cpu.rf.rf[1][3] ;
 wire \i_soc.cpu.rf.rf[1][4] ;
 wire \i_soc.cpu.rf.rf[1][5] ;
 wire \i_soc.cpu.rf.rf[1][6] ;
 wire \i_soc.cpu.rf.rf[1][7] ;
 wire \i_soc.cpu.rf.rf[1][8] ;
 wire \i_soc.cpu.rf.rf[1][9] ;
 wire \i_soc.cpu.rf.rf[27][0] ;
 wire \i_soc.cpu.rf.rf[27][10] ;
 wire \i_soc.cpu.rf.rf[27][11] ;
 wire \i_soc.cpu.rf.rf[27][12] ;
 wire \i_soc.cpu.rf.rf[27][13] ;
 wire \i_soc.cpu.rf.rf[27][14] ;
 wire \i_soc.cpu.rf.rf[27][15] ;
 wire \i_soc.cpu.rf.rf[27][16] ;
 wire \i_soc.cpu.rf.rf[27][17] ;
 wire \i_soc.cpu.rf.rf[27][18] ;
 wire \i_soc.cpu.rf.rf[27][19] ;
 wire \i_soc.cpu.rf.rf[27][1] ;
 wire \i_soc.cpu.rf.rf[27][20] ;
 wire \i_soc.cpu.rf.rf[27][21] ;
 wire \i_soc.cpu.rf.rf[27][22] ;
 wire \i_soc.cpu.rf.rf[27][23] ;
 wire \i_soc.cpu.rf.rf[27][24] ;
 wire \i_soc.cpu.rf.rf[27][25] ;
 wire \i_soc.cpu.rf.rf[27][26] ;
 wire \i_soc.cpu.rf.rf[27][27] ;
 wire \i_soc.cpu.rf.rf[27][28] ;
 wire \i_soc.cpu.rf.rf[27][29] ;
 wire \i_soc.cpu.rf.rf[27][2] ;
 wire \i_soc.cpu.rf.rf[27][30] ;
 wire \i_soc.cpu.rf.rf[27][31] ;
 wire \i_soc.cpu.rf.rf[27][3] ;
 wire \i_soc.cpu.rf.rf[27][4] ;
 wire \i_soc.cpu.rf.rf[27][5] ;
 wire \i_soc.cpu.rf.rf[27][6] ;
 wire \i_soc.cpu.rf.rf[27][7] ;
 wire \i_soc.cpu.rf.rf[27][8] ;
 wire \i_soc.cpu.rf.rf[27][9] ;
 wire \i_soc.cpu.rf.rf[3][0] ;
 wire \i_soc.cpu.rf.rf[3][10] ;
 wire \i_soc.cpu.rf.rf[3][11] ;
 wire \i_soc.cpu.rf.rf[3][12] ;
 wire \i_soc.cpu.rf.rf[3][13] ;
 wire \i_soc.cpu.rf.rf[3][14] ;
 wire \i_soc.cpu.rf.rf[3][15] ;
 wire \i_soc.cpu.rf.rf[3][16] ;
 wire \i_soc.cpu.rf.rf[3][17] ;
 wire \i_soc.cpu.rf.rf[3][18] ;
 wire \i_soc.cpu.rf.rf[3][19] ;
 wire \i_soc.cpu.rf.rf[3][1] ;
 wire \i_soc.cpu.rf.rf[3][20] ;
 wire \i_soc.cpu.rf.rf[3][21] ;
 wire \i_soc.cpu.rf.rf[3][22] ;
 wire \i_soc.cpu.rf.rf[3][23] ;
 wire \i_soc.cpu.rf.rf[3][24] ;
 wire \i_soc.cpu.rf.rf[3][25] ;
 wire \i_soc.cpu.rf.rf[3][26] ;
 wire \i_soc.cpu.rf.rf[3][27] ;
 wire \i_soc.cpu.rf.rf[3][28] ;
 wire \i_soc.cpu.rf.rf[3][29] ;
 wire \i_soc.cpu.rf.rf[3][2] ;
 wire \i_soc.cpu.rf.rf[3][30] ;
 wire \i_soc.cpu.rf.rf[3][31] ;
 wire \i_soc.cpu.rf.rf[3][3] ;
 wire \i_soc.cpu.rf.rf[3][4] ;
 wire \i_soc.cpu.rf.rf[3][5] ;
 wire \i_soc.cpu.rf.rf[3][6] ;
 wire \i_soc.cpu.rf.rf[3][7] ;
 wire \i_soc.cpu.rf.rf[3][8] ;
 wire \i_soc.cpu.rf.rf[3][9] ;
 wire \i_soc.cpu.rf.rf[5][0] ;
 wire \i_soc.cpu.rf.rf[5][10] ;
 wire \i_soc.cpu.rf.rf[5][11] ;
 wire \i_soc.cpu.rf.rf[5][12] ;
 wire \i_soc.cpu.rf.rf[5][13] ;
 wire \i_soc.cpu.rf.rf[5][14] ;
 wire \i_soc.cpu.rf.rf[5][15] ;
 wire \i_soc.cpu.rf.rf[5][16] ;
 wire \i_soc.cpu.rf.rf[5][17] ;
 wire \i_soc.cpu.rf.rf[5][18] ;
 wire \i_soc.cpu.rf.rf[5][19] ;
 wire \i_soc.cpu.rf.rf[5][1] ;
 wire \i_soc.cpu.rf.rf[5][20] ;
 wire \i_soc.cpu.rf.rf[5][21] ;
 wire \i_soc.cpu.rf.rf[5][22] ;
 wire \i_soc.cpu.rf.rf[5][23] ;
 wire \i_soc.cpu.rf.rf[5][24] ;
 wire \i_soc.cpu.rf.rf[5][25] ;
 wire \i_soc.cpu.rf.rf[5][26] ;
 wire \i_soc.cpu.rf.rf[5][27] ;
 wire \i_soc.cpu.rf.rf[5][28] ;
 wire \i_soc.cpu.rf.rf[5][29] ;
 wire \i_soc.cpu.rf.rf[5][2] ;
 wire \i_soc.cpu.rf.rf[5][30] ;
 wire \i_soc.cpu.rf.rf[5][31] ;
 wire \i_soc.cpu.rf.rf[5][3] ;
 wire \i_soc.cpu.rf.rf[5][4] ;
 wire \i_soc.cpu.rf.rf[5][5] ;
 wire \i_soc.cpu.rf.rf[5][6] ;
 wire \i_soc.cpu.rf.rf[5][7] ;
 wire \i_soc.cpu.rf.rf[5][8] ;
 wire \i_soc.cpu.rf.rf[5][9] ;
 wire \i_soc.cpu.rf.rf[6][0] ;
 wire \i_soc.cpu.rf.rf[6][10] ;
 wire \i_soc.cpu.rf.rf[6][11] ;
 wire \i_soc.cpu.rf.rf[6][12] ;
 wire \i_soc.cpu.rf.rf[6][13] ;
 wire \i_soc.cpu.rf.rf[6][14] ;
 wire \i_soc.cpu.rf.rf[6][15] ;
 wire \i_soc.cpu.rf.rf[6][16] ;
 wire \i_soc.cpu.rf.rf[6][17] ;
 wire \i_soc.cpu.rf.rf[6][18] ;
 wire \i_soc.cpu.rf.rf[6][19] ;
 wire \i_soc.cpu.rf.rf[6][1] ;
 wire \i_soc.cpu.rf.rf[6][20] ;
 wire \i_soc.cpu.rf.rf[6][21] ;
 wire \i_soc.cpu.rf.rf[6][22] ;
 wire \i_soc.cpu.rf.rf[6][23] ;
 wire \i_soc.cpu.rf.rf[6][24] ;
 wire \i_soc.cpu.rf.rf[6][25] ;
 wire \i_soc.cpu.rf.rf[6][26] ;
 wire \i_soc.cpu.rf.rf[6][27] ;
 wire \i_soc.cpu.rf.rf[6][28] ;
 wire \i_soc.cpu.rf.rf[6][29] ;
 wire \i_soc.cpu.rf.rf[6][2] ;
 wire \i_soc.cpu.rf.rf[6][30] ;
 wire \i_soc.cpu.rf.rf[6][31] ;
 wire \i_soc.cpu.rf.rf[6][3] ;
 wire \i_soc.cpu.rf.rf[6][4] ;
 wire \i_soc.cpu.rf.rf[6][5] ;
 wire \i_soc.cpu.rf.rf[6][6] ;
 wire \i_soc.cpu.rf.rf[6][7] ;
 wire \i_soc.cpu.rf.rf[6][8] ;
 wire \i_soc.cpu.rf.rf[6][9] ;
 wire \i_soc.cpu.rf.rf[7][0] ;
 wire \i_soc.cpu.rf.rf[7][10] ;
 wire \i_soc.cpu.rf.rf[7][11] ;
 wire \i_soc.cpu.rf.rf[7][12] ;
 wire \i_soc.cpu.rf.rf[7][13] ;
 wire \i_soc.cpu.rf.rf[7][14] ;
 wire \i_soc.cpu.rf.rf[7][15] ;
 wire \i_soc.cpu.rf.rf[7][16] ;
 wire \i_soc.cpu.rf.rf[7][17] ;
 wire \i_soc.cpu.rf.rf[7][18] ;
 wire \i_soc.cpu.rf.rf[7][19] ;
 wire \i_soc.cpu.rf.rf[7][1] ;
 wire \i_soc.cpu.rf.rf[7][20] ;
 wire \i_soc.cpu.rf.rf[7][21] ;
 wire \i_soc.cpu.rf.rf[7][22] ;
 wire \i_soc.cpu.rf.rf[7][23] ;
 wire \i_soc.cpu.rf.rf[7][24] ;
 wire \i_soc.cpu.rf.rf[7][25] ;
 wire \i_soc.cpu.rf.rf[7][26] ;
 wire \i_soc.cpu.rf.rf[7][27] ;
 wire \i_soc.cpu.rf.rf[7][28] ;
 wire \i_soc.cpu.rf.rf[7][29] ;
 wire \i_soc.cpu.rf.rf[7][2] ;
 wire \i_soc.cpu.rf.rf[7][30] ;
 wire \i_soc.cpu.rf.rf[7][31] ;
 wire \i_soc.cpu.rf.rf[7][3] ;
 wire \i_soc.cpu.rf.rf[7][4] ;
 wire \i_soc.cpu.rf.rf[7][5] ;
 wire \i_soc.cpu.rf.rf[7][6] ;
 wire \i_soc.cpu.rf.rf[7][7] ;
 wire \i_soc.cpu.rf.rf[7][8] ;
 wire \i_soc.cpu.rf.rf[7][9] ;
 wire \i_soc.cpu.rf.rf[8][0] ;
 wire \i_soc.cpu.rf.rf[8][10] ;
 wire \i_soc.cpu.rf.rf[8][11] ;
 wire \i_soc.cpu.rf.rf[8][12] ;
 wire \i_soc.cpu.rf.rf[8][13] ;
 wire \i_soc.cpu.rf.rf[8][14] ;
 wire \i_soc.cpu.rf.rf[8][15] ;
 wire \i_soc.cpu.rf.rf[8][16] ;
 wire \i_soc.cpu.rf.rf[8][17] ;
 wire \i_soc.cpu.rf.rf[8][18] ;
 wire \i_soc.cpu.rf.rf[8][19] ;
 wire \i_soc.cpu.rf.rf[8][1] ;
 wire \i_soc.cpu.rf.rf[8][20] ;
 wire \i_soc.cpu.rf.rf[8][21] ;
 wire \i_soc.cpu.rf.rf[8][22] ;
 wire \i_soc.cpu.rf.rf[8][23] ;
 wire \i_soc.cpu.rf.rf[8][24] ;
 wire \i_soc.cpu.rf.rf[8][25] ;
 wire \i_soc.cpu.rf.rf[8][26] ;
 wire \i_soc.cpu.rf.rf[8][27] ;
 wire \i_soc.cpu.rf.rf[8][28] ;
 wire \i_soc.cpu.rf.rf[8][29] ;
 wire \i_soc.cpu.rf.rf[8][2] ;
 wire \i_soc.cpu.rf.rf[8][30] ;
 wire \i_soc.cpu.rf.rf[8][31] ;
 wire \i_soc.cpu.rf.rf[8][3] ;
 wire \i_soc.cpu.rf.rf[8][4] ;
 wire \i_soc.cpu.rf.rf[8][5] ;
 wire \i_soc.cpu.rf.rf[8][6] ;
 wire \i_soc.cpu.rf.rf[8][7] ;
 wire \i_soc.cpu.rf.rf[8][8] ;
 wire \i_soc.cpu.rf.rf[8][9] ;
 wire \i_soc.pass ;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire clknet_leaf_0_clk;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net1;
 wire net2;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;

 sg13g2_inv_1 _1895_ (.Y(_0600_),
    .A(\i_soc.cpu.rf.rf[7][25] ));
 sg13g2_inv_1 _1896_ (.Y(_0601_),
    .A(\i_soc.cpu.rf.rf[7][28] ));
 sg13g2_inv_1 _1897_ (.Y(_0602_),
    .A(net785));
 sg13g2_inv_1 _1898_ (.Y(_0603_),
    .A(net786));
 sg13g2_inv_1 _1899_ (.Y(_0604_),
    .A(\i_soc.cpu.rd0[9] ));
 sg13g2_inv_1 _1900_ (.Y(_0605_),
    .A(\i_soc.cpu.rd0[21] ));
 sg13g2_inv_1 _1901_ (.Y(_0606_),
    .A(_0228_));
 sg13g2_inv_1 _1902_ (.Y(_0607_),
    .A(_0286_));
 sg13g2_inv_1 _1903_ (.Y(_0608_),
    .A(_0083_));
 sg13g2_inv_1 _1904_ (.Y(_0609_),
    .A(_0245_));
 sg13g2_inv_1 _1905_ (.Y(_0610_),
    .A(_0242_));
 sg13g2_inv_1 _1906_ (.Y(_0611_),
    .A(\i_soc.cpu.rf.rf[7][21] ));
 sg13g2_inv_2 _1907_ (.Y(_0612_),
    .A(net611));
 sg13g2_nor2b_2 _1908_ (.A(net603),
    .B_N(net605),
    .Y(_0613_));
 sg13g2_nor2b_2 _1909_ (.A(net608),
    .B_N(net609),
    .Y(_0614_));
 sg13g2_and2_1 _1910_ (.A(_0613_),
    .B(_0614_),
    .X(_0615_));
 sg13g2_nand2_2 _1911_ (.Y(_0616_),
    .A(_0613_),
    .B(_0614_));
 sg13g2_nor2b_2 _1912_ (.A(net609),
    .B_N(net608),
    .Y(_0617_));
 sg13g2_nor2b_2 _1913_ (.A(net606),
    .B_N(net603),
    .Y(_0618_));
 sg13g2_a22oi_1 _1914_ (.Y(_0619_),
    .B1(_0618_),
    .B2(_0614_),
    .A2(_0617_),
    .A1(_0613_));
 sg13g2_nor2b_1 _1915_ (.A(net604),
    .B_N(net610),
    .Y(_0620_));
 sg13g2_nand2b_1 _1916_ (.Y(_0621_),
    .B(net609),
    .A_N(net602));
 sg13g2_nor2_2 _1917_ (.A(net605),
    .B(net602),
    .Y(_0622_));
 sg13g2_nor2_1 _1918_ (.A(net605),
    .B(_0621_),
    .Y(_0623_));
 sg13g2_nand2_1 _1919_ (.Y(_0624_),
    .A(net609),
    .B(_0622_));
 sg13g2_nor2_1 _1920_ (.A(net608),
    .B(net607),
    .Y(_0625_));
 sg13g2_or2_1 _1921_ (.X(_0626_),
    .B(net605),
    .A(net608));
 sg13g2_nor2_2 _1922_ (.A(_0620_),
    .B(_0625_),
    .Y(_0627_));
 sg13g2_a21oi_2 _1923_ (.B1(net602),
    .Y(_0628_),
    .A2(_0617_),
    .A1(net606));
 sg13g2_and2_1 _1924_ (.A(net572),
    .B(_0628_),
    .X(_0629_));
 sg13g2_nand2_1 _1925_ (.Y(_0630_),
    .A(net572),
    .B(_0628_));
 sg13g2_nor2_1 _1926_ (.A(_0627_),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_and2_1 _1927_ (.A(net605),
    .B(net602),
    .X(_0632_));
 sg13g2_nand2_2 _1928_ (.Y(_0633_),
    .A(net605),
    .B(net602));
 sg13g2_a21oi_2 _1929_ (.B1(net601),
    .Y(_0634_),
    .A2(_0622_),
    .A1(net609));
 sg13g2_o21ai_1 _1930_ (.B1(_0633_),
    .Y(_0635_),
    .A1(net605),
    .A2(_0621_));
 sg13g2_nor2_2 _1931_ (.A(net609),
    .B(net608),
    .Y(_0636_));
 sg13g2_nor4_2 _1932_ (.A(net609),
    .B(net608),
    .C(net605),
    .Y(_0637_),
    .D(net602));
 sg13g2_nand2_1 _1933_ (.Y(_0638_),
    .A(_0617_),
    .B(_0618_));
 sg13g2_a21oi_2 _1934_ (.B1(_0637_),
    .Y(_0639_),
    .A2(_0618_),
    .A1(_0617_));
 sg13g2_a21o_1 _1935_ (.A2(_0618_),
    .A1(_0617_),
    .B1(_0637_),
    .X(_0640_));
 sg13g2_nor2_1 _1936_ (.A(_0635_),
    .B(_0640_),
    .Y(_0641_));
 sg13g2_nand2_1 _1937_ (.Y(_0642_),
    .A(_0634_),
    .B(_0639_));
 sg13g2_a21oi_1 _1938_ (.A1(_0621_),
    .A2(_0626_),
    .Y(_0643_),
    .B1(_0160_));
 sg13g2_nor3_2 _1939_ (.A(_0197_),
    .B(_0620_),
    .C(_0625_),
    .Y(_0644_));
 sg13g2_nor4_1 _1940_ (.A(_0635_),
    .B(_0640_),
    .C(_0643_),
    .D(_0644_),
    .Y(_0645_));
 sg13g2_a21oi_2 _1941_ (.B1(net606),
    .Y(_0646_),
    .A2(net608),
    .A1(net610));
 sg13g2_a21oi_1 _1942_ (.A1(net603),
    .A2(_0646_),
    .Y(_0647_),
    .B1(net589));
 sg13g2_a21o_1 _1943_ (.A2(_0646_),
    .A1(net603),
    .B1(net589),
    .X(_0648_));
 sg13g2_o21ai_1 _1944_ (.B1(_0261_),
    .Y(_0649_),
    .A1(_0635_),
    .A2(_0640_));
 sg13g2_nand3b_1 _1945_ (.B(net556),
    .C(_0649_),
    .Y(_0650_),
    .A_N(_0645_));
 sg13g2_nor3_1 _1946_ (.A(net609),
    .B(net606),
    .C(net602),
    .Y(_0651_));
 sg13g2_nand2_1 _1947_ (.Y(_0652_),
    .A(_0617_),
    .B(_0622_));
 sg13g2_a22oi_1 _1948_ (.Y(_0653_),
    .B1(_0617_),
    .B2(_0622_),
    .A2(_0614_),
    .A1(_0613_));
 sg13g2_and2_1 _1949_ (.A(_0633_),
    .B(_0653_),
    .X(_0654_));
 sg13g2_nand2_1 _1950_ (.Y(_0655_),
    .A(_0633_),
    .B(_0653_));
 sg13g2_o21ai_1 _1951_ (.B1(_0031_),
    .Y(_0656_),
    .A1(_0635_),
    .A2(_0640_));
 sg13g2_nand3_1 _1952_ (.B(_0634_),
    .C(_0639_),
    .A(_0128_),
    .Y(_0657_));
 sg13g2_nand3_1 _1953_ (.B(_0656_),
    .C(_0657_),
    .A(net552),
    .Y(_0658_));
 sg13g2_nand3_1 _1954_ (.B(net548),
    .C(_0658_),
    .A(_0650_),
    .Y(_0659_));
 sg13g2_nand4_1 _1955_ (.B(_0634_),
    .C(_0639_),
    .A(_0627_),
    .Y(_0660_),
    .D(_0653_));
 sg13g2_inv_1 _1956_ (.Y(_0661_),
    .A(_0660_));
 sg13g2_nor2_2 _1957_ (.A(_0629_),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_nand2_2 _1958_ (.Y(_0663_),
    .A(_0630_),
    .B(_0660_));
 sg13g2_a21oi_1 _1959_ (.A1(_0229_),
    .A2(net545),
    .Y(_0664_),
    .B1(net499));
 sg13g2_a21oi_2 _1960_ (.B1(_0631_),
    .Y(_0665_),
    .A2(_0664_),
    .A1(_0659_));
 sg13g2_and2_1 _1961_ (.A(_0613_),
    .B(_0636_),
    .X(_0666_));
 sg13g2_nand2_2 _1962_ (.Y(_0667_),
    .A(_0613_),
    .B(_0636_));
 sg13g2_nor2_1 _1963_ (.A(net599),
    .B(net569),
    .Y(_0668_));
 sg13g2_nand2_1 _1964_ (.Y(_0669_),
    .A(_0633_),
    .B(_0667_));
 sg13g2_nand2_2 _1965_ (.Y(_0670_),
    .A(_0618_),
    .B(_0636_));
 sg13g2_and3_1 _1966_ (.X(_0671_),
    .A(_0652_),
    .B(net538),
    .C(_0670_));
 sg13g2_nand3_1 _1967_ (.B(net538),
    .C(_0670_),
    .A(_0652_),
    .Y(_0672_));
 sg13g2_nor2_1 _1968_ (.A(_0229_),
    .B(net528),
    .Y(_0673_));
 sg13g2_o21ai_1 _1969_ (.B1(net484),
    .Y(_0674_),
    .A1(_0094_),
    .A2(net534));
 sg13g2_and2_1 _1970_ (.A(_0634_),
    .B(_0670_),
    .X(_0675_));
 sg13g2_nand2_2 _1971_ (.Y(_0676_),
    .A(_0634_),
    .B(_0670_));
 sg13g2_a21oi_1 _1972_ (.A1(_0192_),
    .A2(net493),
    .Y(_0677_),
    .B1(net518));
 sg13g2_o21ai_1 _1973_ (.B1(_0677_),
    .Y(_0678_),
    .A1(_0673_),
    .A2(_0674_));
 sg13g2_nand2_1 _1974_ (.Y(_0679_),
    .A(_0063_),
    .B(net526));
 sg13g2_a21oi_1 _1975_ (.A1(_0031_),
    .A2(net534),
    .Y(_0680_),
    .B1(net513));
 sg13g2_a21oi_1 _1976_ (.A1(_0679_),
    .A2(_0680_),
    .Y(_0681_),
    .B1(net601));
 sg13g2_nand2b_1 _1977_ (.Y(_0682_),
    .B(_0622_),
    .A_N(_0636_));
 sg13g2_nor2_1 _1978_ (.A(net575),
    .B(_0672_),
    .Y(_0683_));
 sg13g2_nand2_2 _1979_ (.Y(_0684_),
    .A(net572),
    .B(net493));
 sg13g2_a221oi_1 _1980_ (.B2(_0681_),
    .C1(net471),
    .B1(_0678_),
    .A1(_0293_),
    .Y(_0685_),
    .A2(net601));
 sg13g2_or2_1 _1981_ (.X(_0686_),
    .B(_0685_),
    .A(_0665_));
 sg13g2_xnor2_1 _1982_ (.Y(_0687_),
    .A(_0665_),
    .B(_0685_));
 sg13g2_nand2_2 _1983_ (.Y(_0688_),
    .A(net572),
    .B(_0687_));
 sg13g2_nand2_1 _1984_ (.Y(_0689_),
    .A(net782),
    .B(net586));
 sg13g2_o21ai_1 _1985_ (.B1(_0689_),
    .Y(_0358_),
    .A1(net586),
    .A2(_0688_));
 sg13g2_nor2_1 _1986_ (.A(_0606_),
    .B(net525),
    .Y(_0690_));
 sg13g2_a21oi_1 _1987_ (.A1(_0093_),
    .A2(net525),
    .Y(_0691_),
    .B1(_0690_));
 sg13g2_a21oi_1 _1988_ (.A1(_0191_),
    .A2(net491),
    .Y(_0692_),
    .B1(net518));
 sg13g2_o21ai_1 _1989_ (.B1(_0692_),
    .Y(_0693_),
    .A1(net491),
    .A2(_0691_));
 sg13g2_nand2_1 _1990_ (.Y(_0694_),
    .A(_0062_),
    .B(net525));
 sg13g2_a21oi_1 _1991_ (.A1(_0030_),
    .A2(net534),
    .Y(_0695_),
    .B1(net513));
 sg13g2_a21oi_1 _1992_ (.A1(_0694_),
    .A2(_0695_),
    .Y(_0696_),
    .B1(net597));
 sg13g2_a221oi_1 _1993_ (.B2(_0696_),
    .C1(net471),
    .B1(_0693_),
    .A1(_0292_),
    .Y(_0697_),
    .A2(net597));
 sg13g2_mux2_1 _1994_ (.A0(_0159_),
    .A1(_0196_),
    .S(_0627_),
    .X(_0698_));
 sg13g2_mux4_1 _1995_ (.S0(net552),
    .A0(_0260_),
    .A1(_0030_),
    .A2(_0698_),
    .A3(_0127_),
    .S1(net566),
    .X(_0699_));
 sg13g2_o21ai_1 _1996_ (.B1(_0660_),
    .Y(_0700_),
    .A1(_0606_),
    .A2(net548));
 sg13g2_a21oi_1 _1997_ (.A1(net548),
    .A2(_0699_),
    .Y(_0701_),
    .B1(_0700_));
 sg13g2_nand2_1 _1998_ (.Y(_0702_),
    .A(_0628_),
    .B(net566));
 sg13g2_o21ai_1 _1999_ (.B1(_0702_),
    .Y(_0703_),
    .A1(_0629_),
    .A2(_0701_));
 sg13g2_xnor2_1 _2000_ (.Y(_0704_),
    .A(_0665_),
    .B(_0703_));
 sg13g2_and2_1 _2001_ (.A(_0697_),
    .B(_0704_),
    .X(_0705_));
 sg13g2_xor2_1 _2002_ (.B(_0704_),
    .A(_0697_),
    .X(_0706_));
 sg13g2_a21oi_1 _2003_ (.A1(_0686_),
    .A2(_0706_),
    .Y(_0707_),
    .B1(net575));
 sg13g2_o21ai_1 _2004_ (.B1(_0707_),
    .Y(_0708_),
    .A1(_0686_),
    .A2(_0706_));
 sg13g2_nand2_1 _2005_ (.Y(_0709_),
    .A(net777),
    .B(net585));
 sg13g2_o21ai_1 _2006_ (.B1(_0709_),
    .Y(_0359_),
    .A1(net585),
    .A2(_0708_));
 sg13g2_a21oi_1 _2007_ (.A1(_0686_),
    .A2(_0706_),
    .Y(_0710_),
    .B1(_0705_));
 sg13g2_and2_1 _2008_ (.A(_0092_),
    .B(net525),
    .X(_0711_));
 sg13g2_a21oi_1 _2009_ (.A1(_0227_),
    .A2(net534),
    .Y(_0712_),
    .B1(_0711_));
 sg13g2_a21oi_1 _2010_ (.A1(_0190_),
    .A2(net491),
    .Y(_0713_),
    .B1(net518));
 sg13g2_o21ai_1 _2011_ (.B1(_0713_),
    .Y(_0714_),
    .A1(net491),
    .A2(_0712_));
 sg13g2_nand2_1 _2012_ (.Y(_0715_),
    .A(_0061_),
    .B(net525));
 sg13g2_a21oi_1 _2013_ (.A1(_0029_),
    .A2(net534),
    .Y(_0716_),
    .B1(net513));
 sg13g2_a21oi_1 _2014_ (.A1(_0715_),
    .A2(_0716_),
    .Y(_0717_),
    .B1(net597));
 sg13g2_a221oi_1 _2015_ (.B2(_0717_),
    .C1(net471),
    .B1(_0714_),
    .A1(_0291_),
    .Y(_0718_),
    .A2(net597));
 sg13g2_mux2_1 _2016_ (.A0(_0158_),
    .A1(_0195_),
    .S(_0627_),
    .X(_0719_));
 sg13g2_mux4_1 _2017_ (.S0(net552),
    .A0(_0259_),
    .A1(_0029_),
    .A2(_0719_),
    .A3(_0126_),
    .S1(net566),
    .X(_0720_));
 sg13g2_nand2_1 _2018_ (.Y(_0721_),
    .A(net548),
    .B(_0720_));
 sg13g2_a21oi_1 _2019_ (.A1(_0227_),
    .A2(net545),
    .Y(_0722_),
    .B1(net499));
 sg13g2_a21oi_1 _2020_ (.A1(_0721_),
    .A2(_0722_),
    .Y(_0723_),
    .B1(net589));
 sg13g2_a21oi_1 _2021_ (.A1(_0665_),
    .A2(_0703_),
    .Y(_0724_),
    .B1(_0723_));
 sg13g2_nand3_1 _2022_ (.B(_0703_),
    .C(_0723_),
    .A(_0665_),
    .Y(_0725_));
 sg13g2_nor2b_1 _2023_ (.A(_0724_),
    .B_N(_0725_),
    .Y(_0726_));
 sg13g2_nand2b_1 _2024_ (.Y(_0727_),
    .B(_0718_),
    .A_N(_0726_));
 sg13g2_xor2_1 _2025_ (.B(_0726_),
    .A(_0718_),
    .X(_0728_));
 sg13g2_a21oi_1 _2026_ (.A1(_0710_),
    .A2(_0728_),
    .Y(_0729_),
    .B1(net575));
 sg13g2_o21ai_1 _2027_ (.B1(_0729_),
    .Y(_0730_),
    .A1(_0710_),
    .A2(_0728_));
 sg13g2_nand2_1 _2028_ (.Y(_0731_),
    .A(net775),
    .B(net585));
 sg13g2_o21ai_1 _2029_ (.B1(_0731_),
    .Y(_0360_),
    .A1(net585),
    .A2(_0730_));
 sg13g2_o21ai_1 _2030_ (.B1(_0727_),
    .Y(_0732_),
    .A1(_0710_),
    .A2(_0728_));
 sg13g2_nor2_1 _2031_ (.A(_0226_),
    .B(net526),
    .Y(_0733_));
 sg13g2_o21ai_1 _2032_ (.B1(net484),
    .Y(_0734_),
    .A1(_0091_),
    .A2(net535));
 sg13g2_a21oi_1 _2033_ (.A1(_0189_),
    .A2(net491),
    .Y(_0735_),
    .B1(net518));
 sg13g2_o21ai_1 _2034_ (.B1(_0735_),
    .Y(_0736_),
    .A1(_0733_),
    .A2(_0734_));
 sg13g2_nand2_1 _2035_ (.Y(_0737_),
    .A(_0060_),
    .B(net525));
 sg13g2_a21oi_1 _2036_ (.A1(_0028_),
    .A2(net534),
    .Y(_0738_),
    .B1(net513));
 sg13g2_a21oi_1 _2037_ (.A1(_0737_),
    .A2(_0738_),
    .Y(_0739_),
    .B1(net597));
 sg13g2_a22oi_1 _2038_ (.Y(_0740_),
    .B1(_0736_),
    .B2(_0739_),
    .A2(net597),
    .A1(_0290_));
 sg13g2_nand2_1 _2039_ (.Y(_0741_),
    .A(_0684_),
    .B(_0740_));
 sg13g2_mux2_1 _2040_ (.A0(_0157_),
    .A1(_0194_),
    .S(_0627_),
    .X(_0742_));
 sg13g2_mux4_1 _2041_ (.S0(net552),
    .A0(_0258_),
    .A1(_0028_),
    .A2(_0742_),
    .A3(_0125_),
    .S1(net566),
    .X(_0743_));
 sg13g2_o21ai_1 _2042_ (.B1(net548),
    .Y(_0744_),
    .A1(_0629_),
    .A2(_0743_));
 sg13g2_a21oi_1 _2043_ (.A1(_0226_),
    .A2(net545),
    .Y(_0745_),
    .B1(_0661_));
 sg13g2_o21ai_1 _2044_ (.B1(_0744_),
    .Y(_0746_),
    .A1(_0629_),
    .A2(_0745_));
 sg13g2_nand4_1 _2045_ (.B(_0703_),
    .C(_0723_),
    .A(_0665_),
    .Y(_0747_),
    .D(_0746_));
 sg13g2_xor2_1 _2046_ (.B(_0746_),
    .A(_0725_),
    .X(_0748_));
 sg13g2_nor2b_1 _2047_ (.A(_0741_),
    .B_N(_0748_),
    .Y(_0749_));
 sg13g2_nand2b_1 _2048_ (.Y(_0750_),
    .B(_0741_),
    .A_N(_0748_));
 sg13g2_nand2b_1 _2049_ (.Y(_0751_),
    .B(_0750_),
    .A_N(_0749_));
 sg13g2_xnor2_1 _2050_ (.Y(_0752_),
    .A(_0732_),
    .B(_0751_));
 sg13g2_nand2_2 _2051_ (.Y(_0753_),
    .A(net572),
    .B(_0752_));
 sg13g2_nand2_1 _2052_ (.Y(_0754_),
    .A(net767),
    .B(net585));
 sg13g2_o21ai_1 _2053_ (.B1(_0754_),
    .Y(_0361_),
    .A1(net585),
    .A2(_0753_));
 sg13g2_nor2_1 _2054_ (.A(_0090_),
    .B(net534),
    .Y(_0755_));
 sg13g2_nor2_1 _2055_ (.A(_0225_),
    .B(net525),
    .Y(_0756_));
 sg13g2_nor3_1 _2056_ (.A(net491),
    .B(_0755_),
    .C(_0756_),
    .Y(_0757_));
 sg13g2_a21oi_1 _2057_ (.A1(_0188_),
    .A2(net493),
    .Y(_0758_),
    .B1(_0757_));
 sg13g2_nand2_1 _2058_ (.Y(_0759_),
    .A(_0059_),
    .B(net525));
 sg13g2_a21oi_1 _2059_ (.A1(_0027_),
    .A2(net534),
    .Y(_0760_),
    .B1(net513));
 sg13g2_a221oi_1 _2060_ (.B2(_0760_),
    .C1(net597),
    .B1(_0759_),
    .A1(net515),
    .Y(_0761_),
    .A2(_0758_));
 sg13g2_a21oi_1 _2061_ (.A1(_0289_),
    .A2(net597),
    .Y(_0762_),
    .B1(net471));
 sg13g2_nand2b_1 _2062_ (.Y(_0763_),
    .B(_0762_),
    .A_N(_0761_));
 sg13g2_nand2_1 _2063_ (.Y(_0764_),
    .A(_0027_),
    .B(net561));
 sg13g2_a21oi_1 _2064_ (.A1(_0124_),
    .A2(net566),
    .Y(_0765_),
    .B1(net556));
 sg13g2_nand2_1 _2065_ (.Y(_0766_),
    .A(_0257_),
    .B(net561));
 sg13g2_a21oi_1 _2066_ (.A1(_0156_),
    .A2(net566),
    .Y(_0767_),
    .B1(net552));
 sg13g2_a221oi_1 _2067_ (.B2(_0767_),
    .C1(net545),
    .B1(_0766_),
    .A1(_0764_),
    .Y(_0768_),
    .A2(_0765_));
 sg13g2_nand2_1 _2068_ (.Y(_0769_),
    .A(_0653_),
    .B(net497));
 sg13g2_and2_1 _2069_ (.A(_0225_),
    .B(_0630_),
    .X(_0770_));
 sg13g2_a221oi_1 _2070_ (.B2(net545),
    .C1(_0768_),
    .B1(_0770_),
    .A1(_0653_),
    .Y(_0771_),
    .A2(net499));
 sg13g2_nor2_1 _2071_ (.A(_0747_),
    .B(_0771_),
    .Y(_0772_));
 sg13g2_xnor2_1 _2072_ (.Y(_0773_),
    .A(_0747_),
    .B(_0771_));
 sg13g2_nand2b_1 _2073_ (.Y(_0774_),
    .B(_0773_),
    .A_N(_0763_));
 sg13g2_xor2_1 _2074_ (.B(_0773_),
    .A(_0763_),
    .X(_0775_));
 sg13g2_a21oi_2 _2075_ (.B1(_0749_),
    .Y(_0776_),
    .A2(_0750_),
    .A1(_0732_));
 sg13g2_or2_1 _2076_ (.X(_0777_),
    .B(_0776_),
    .A(_0775_));
 sg13g2_a21oi_1 _2077_ (.A1(_0775_),
    .A2(_0776_),
    .Y(_0778_),
    .B1(net575));
 sg13g2_nand2_2 _2078_ (.Y(_0779_),
    .A(_0777_),
    .B(_0778_));
 sg13g2_nand2_1 _2079_ (.Y(_0780_),
    .A(net754),
    .B(net584));
 sg13g2_o21ai_1 _2080_ (.B1(_0780_),
    .Y(_0362_),
    .A1(net584),
    .A2(_0779_));
 sg13g2_nor2_1 _2081_ (.A(_0224_),
    .B(net526),
    .Y(_0781_));
 sg13g2_o21ai_1 _2082_ (.B1(net484),
    .Y(_0782_),
    .A1(_0089_),
    .A2(net535));
 sg13g2_a21oi_1 _2083_ (.A1(_0187_),
    .A2(net491),
    .Y(_0783_),
    .B1(net518));
 sg13g2_o21ai_1 _2084_ (.B1(_0783_),
    .Y(_0784_),
    .A1(_0781_),
    .A2(_0782_));
 sg13g2_nand2_1 _2085_ (.Y(_0785_),
    .A(_0026_),
    .B(net535));
 sg13g2_a21oi_1 _2086_ (.A1(_0058_),
    .A2(net526),
    .Y(_0786_),
    .B1(net513));
 sg13g2_a21oi_1 _2087_ (.A1(_0785_),
    .A2(_0786_),
    .Y(_0787_),
    .B1(net598));
 sg13g2_nand2_1 _2088_ (.Y(_0788_),
    .A(_0288_),
    .B(net598));
 sg13g2_a21oi_1 _2089_ (.A1(_0784_),
    .A2(_0787_),
    .Y(_0789_),
    .B1(net471));
 sg13g2_mux4_1 _2090_ (.S0(net561),
    .A0(_0155_),
    .A1(_0256_),
    .A2(_0123_),
    .A3(_0026_),
    .S1(net553),
    .X(_0790_));
 sg13g2_a21o_1 _2091_ (.A2(net545),
    .A1(_0224_),
    .B1(net498),
    .X(_0791_));
 sg13g2_a21oi_1 _2092_ (.A1(net548),
    .A2(_0790_),
    .Y(_0792_),
    .B1(_0791_));
 sg13g2_nor2_1 _2093_ (.A(_0651_),
    .B(_0792_),
    .Y(_0793_));
 sg13g2_or2_1 _2094_ (.X(_0794_),
    .B(_0792_),
    .A(_0651_));
 sg13g2_nand2_1 _2095_ (.Y(_0795_),
    .A(_0772_),
    .B(_0793_));
 sg13g2_xnor2_1 _2096_ (.Y(_0796_),
    .A(_0772_),
    .B(_0793_));
 sg13g2_a21oi_1 _2097_ (.A1(_0788_),
    .A2(_0789_),
    .Y(_0797_),
    .B1(_0796_));
 sg13g2_inv_1 _2098_ (.Y(_0798_),
    .A(_0797_));
 sg13g2_nand3_1 _2099_ (.B(_0789_),
    .C(_0796_),
    .A(_0788_),
    .Y(_0799_));
 sg13g2_nand2_1 _2100_ (.Y(_0800_),
    .A(_0798_),
    .B(_0799_));
 sg13g2_and2_1 _2101_ (.A(_0774_),
    .B(_0777_),
    .X(_0801_));
 sg13g2_a21oi_1 _2102_ (.A1(_0800_),
    .A2(_0801_),
    .Y(_0802_),
    .B1(net574));
 sg13g2_o21ai_1 _2103_ (.B1(_0802_),
    .Y(_0803_),
    .A1(_0800_),
    .A2(_0801_));
 sg13g2_nand2_1 _2104_ (.Y(_0804_),
    .A(net753),
    .B(net584));
 sg13g2_o21ai_1 _2105_ (.B1(_0804_),
    .Y(_0363_),
    .A1(net584),
    .A2(_0803_));
 sg13g2_nand2_1 _2106_ (.Y(_0805_),
    .A(_0057_),
    .B(net569));
 sg13g2_a21oi_1 _2107_ (.A1(_0025_),
    .A2(net535),
    .Y(_0806_),
    .B1(net513));
 sg13g2_a21oi_1 _2108_ (.A1(_0805_),
    .A2(_0806_),
    .Y(_0807_),
    .B1(net598));
 sg13g2_nor2_1 _2109_ (.A(_0223_),
    .B(net526),
    .Y(_0808_));
 sg13g2_o21ai_1 _2110_ (.B1(net484),
    .Y(_0809_),
    .A1(_0088_),
    .A2(net535));
 sg13g2_a21oi_1 _2111_ (.A1(_0186_),
    .A2(net491),
    .Y(_0810_),
    .B1(net518));
 sg13g2_o21ai_1 _2112_ (.B1(_0810_),
    .Y(_0811_),
    .A1(_0808_),
    .A2(_0809_));
 sg13g2_a221oi_1 _2113_ (.B2(_0811_),
    .C1(net471),
    .B1(_0807_),
    .A1(_0287_),
    .Y(_0812_),
    .A2(net598));
 sg13g2_a21o_1 _2114_ (.A2(net561),
    .A1(_0025_),
    .B1(net556),
    .X(_0813_));
 sg13g2_a21oi_1 _2115_ (.A1(_0122_),
    .A2(net566),
    .Y(_0814_),
    .B1(_0813_));
 sg13g2_a21o_1 _2116_ (.A2(net566),
    .A1(_0154_),
    .B1(net553),
    .X(_0815_));
 sg13g2_a21oi_1 _2117_ (.A1(_0255_),
    .A2(net561),
    .Y(_0816_),
    .B1(_0815_));
 sg13g2_nor3_1 _2118_ (.A(net545),
    .B(_0814_),
    .C(_0816_),
    .Y(_0817_));
 sg13g2_a221oi_1 _2119_ (.B2(net498),
    .C1(_0817_),
    .B1(_0653_),
    .A1(_0223_),
    .Y(_0818_),
    .A2(net598));
 sg13g2_nor4_2 _2120_ (.A(_0747_),
    .B(_0771_),
    .C(_0794_),
    .Y(_0819_),
    .D(_0818_));
 sg13g2_xor2_1 _2121_ (.B(_0818_),
    .A(_0795_),
    .X(_0820_));
 sg13g2_nand2b_1 _2122_ (.Y(_0821_),
    .B(_0812_),
    .A_N(_0820_));
 sg13g2_xor2_1 _2123_ (.B(_0820_),
    .A(_0812_),
    .X(_0822_));
 sg13g2_and2_1 _2124_ (.A(_0774_),
    .B(_0799_),
    .X(_0823_));
 sg13g2_o21ai_1 _2125_ (.B1(_0823_),
    .Y(_0824_),
    .A1(_0775_),
    .A2(_0776_));
 sg13g2_nand2_1 _2126_ (.Y(_0825_),
    .A(_0798_),
    .B(_0824_));
 sg13g2_nand3b_1 _2127_ (.B(_0824_),
    .C(_0798_),
    .Y(_0826_),
    .A_N(_0822_));
 sg13g2_a21oi_1 _2128_ (.A1(_0822_),
    .A2(_0825_),
    .Y(_0827_),
    .B1(net574));
 sg13g2_nand2_2 _2129_ (.Y(_0828_),
    .A(_0826_),
    .B(_0827_));
 sg13g2_nand2_1 _2130_ (.Y(_0829_),
    .A(net750),
    .B(net584));
 sg13g2_o21ai_1 _2131_ (.B1(_0829_),
    .Y(_0364_),
    .A1(net584),
    .A2(_0828_));
 sg13g2_nand2_1 _2132_ (.Y(_0830_),
    .A(_0821_),
    .B(_0826_));
 sg13g2_and2_1 _2133_ (.A(_0087_),
    .B(net526),
    .X(_0831_));
 sg13g2_a21oi_1 _2134_ (.A1(_0222_),
    .A2(net535),
    .Y(_0832_),
    .B1(_0831_));
 sg13g2_a21oi_1 _2135_ (.A1(net484),
    .A2(_0832_),
    .Y(_0833_),
    .B1(net518));
 sg13g2_o21ai_1 _2136_ (.B1(_0833_),
    .Y(_0834_),
    .A1(_0185_),
    .A2(net485));
 sg13g2_a22oi_1 _2137_ (.Y(_0835_),
    .B1(net535),
    .B2(_0024_),
    .A2(net569),
    .A1(_0056_));
 sg13g2_nor2_1 _2138_ (.A(net513),
    .B(_0835_),
    .Y(_0836_));
 sg13g2_nor2_1 _2139_ (.A(net598),
    .B(_0836_),
    .Y(_0837_));
 sg13g2_a22oi_1 _2140_ (.Y(_0838_),
    .B1(_0834_),
    .B2(_0837_),
    .A2(net598),
    .A1(_0607_));
 sg13g2_mux4_1 _2141_ (.S0(net561),
    .A0(_0153_),
    .A1(_0254_),
    .A2(_0121_),
    .A3(_0024_),
    .S1(net553),
    .X(_0839_));
 sg13g2_nand2_1 _2142_ (.Y(_0840_),
    .A(_0222_),
    .B(net545));
 sg13g2_a21oi_1 _2143_ (.A1(net548),
    .A2(_0839_),
    .Y(_0841_),
    .B1(net498));
 sg13g2_a21oi_2 _2144_ (.B1(net590),
    .Y(_0842_),
    .A2(_0841_),
    .A1(_0840_));
 sg13g2_xor2_1 _2145_ (.B(_0842_),
    .A(_0819_),
    .X(_0843_));
 sg13g2_nor3_1 _2146_ (.A(net471),
    .B(_0838_),
    .C(_0843_),
    .Y(_0844_));
 sg13g2_inv_1 _2147_ (.Y(_0845_),
    .A(_0844_));
 sg13g2_o21ai_1 _2148_ (.B1(_0843_),
    .Y(_0846_),
    .A1(net471),
    .A2(_0838_));
 sg13g2_nor2b_1 _2149_ (.A(_0844_),
    .B_N(_0846_),
    .Y(_0847_));
 sg13g2_a21oi_1 _2150_ (.A1(_0830_),
    .A2(_0847_),
    .Y(_0848_),
    .B1(net576));
 sg13g2_o21ai_1 _2151_ (.B1(_0848_),
    .Y(_0849_),
    .A1(_0830_),
    .A2(_0847_));
 sg13g2_nand2_1 _2152_ (.Y(_0850_),
    .A(net765),
    .B(net584));
 sg13g2_o21ai_1 _2153_ (.B1(_0850_),
    .Y(_0365_),
    .A1(net582),
    .A2(_0849_));
 sg13g2_nor2_1 _2154_ (.A(_0221_),
    .B(net522),
    .Y(_0851_));
 sg13g2_o21ai_1 _2155_ (.B1(net485),
    .Y(_0852_),
    .A1(_0086_),
    .A2(net531));
 sg13g2_o21ai_1 _2156_ (.B1(net510),
    .Y(_0853_),
    .A1(_0851_),
    .A2(_0852_));
 sg13g2_a21oi_1 _2157_ (.A1(_0184_),
    .A2(net487),
    .Y(_0854_),
    .B1(_0853_));
 sg13g2_mux2_1 _2158_ (.A0(_0023_),
    .A1(_0055_),
    .S(net522),
    .X(_0855_));
 sg13g2_o21ai_1 _2159_ (.B1(_0633_),
    .Y(_0856_),
    .A1(net510),
    .A2(_0855_));
 sg13g2_a21oi_1 _2160_ (.A1(_0285_),
    .A2(net592),
    .Y(_0857_),
    .B1(net469));
 sg13g2_o21ai_1 _2161_ (.B1(_0857_),
    .Y(_0858_),
    .A1(_0854_),
    .A2(_0856_));
 sg13g2_mux4_1 _2162_ (.S0(net559),
    .A0(_0152_),
    .A1(_0253_),
    .A2(_0120_),
    .A3(_0023_),
    .S1(net554),
    .X(_0859_));
 sg13g2_nand2_1 _2163_ (.Y(_0860_),
    .A(net549),
    .B(_0859_));
 sg13g2_a21oi_1 _2164_ (.A1(_0221_),
    .A2(net542),
    .Y(_0861_),
    .B1(net497));
 sg13g2_a21oi_1 _2165_ (.A1(_0860_),
    .A2(_0861_),
    .Y(_0862_),
    .B1(_0637_));
 sg13g2_a21oi_1 _2166_ (.A1(_0819_),
    .A2(_0842_),
    .Y(_0863_),
    .B1(_0862_));
 sg13g2_nand3_1 _2167_ (.B(_0842_),
    .C(_0862_),
    .A(_0819_),
    .Y(_0864_));
 sg13g2_nor2b_1 _2168_ (.A(_0863_),
    .B_N(_0864_),
    .Y(_0865_));
 sg13g2_or2_1 _2169_ (.X(_0866_),
    .B(_0865_),
    .A(_0858_));
 sg13g2_xor2_1 _2170_ (.B(_0865_),
    .A(_0858_),
    .X(_0867_));
 sg13g2_nand3_1 _2171_ (.B(_0826_),
    .C(_0845_),
    .A(_0821_),
    .Y(_0868_));
 sg13g2_nand2_1 _2172_ (.Y(_0869_),
    .A(_0846_),
    .B(_0868_));
 sg13g2_nand2b_1 _2173_ (.Y(_0870_),
    .B(_0869_),
    .A_N(_0867_));
 sg13g2_nand3_1 _2174_ (.B(_0867_),
    .C(_0868_),
    .A(_0846_),
    .Y(_0871_));
 sg13g2_nand3_1 _2175_ (.B(_0870_),
    .C(_0871_),
    .A(net572),
    .Y(_0872_));
 sg13g2_nand2_1 _2176_ (.Y(_0873_),
    .A(net778),
    .B(net582));
 sg13g2_o21ai_1 _2177_ (.B1(_0873_),
    .Y(_0366_),
    .A1(net582),
    .A2(_0872_));
 sg13g2_nor2_1 _2178_ (.A(_0085_),
    .B(net531),
    .Y(_0874_));
 sg13g2_nor2_1 _2179_ (.A(_0220_),
    .B(net522),
    .Y(_0875_));
 sg13g2_nor3_1 _2180_ (.A(net487),
    .B(_0874_),
    .C(_0875_),
    .Y(_0876_));
 sg13g2_a21oi_1 _2181_ (.A1(_0183_),
    .A2(net487),
    .Y(_0877_),
    .B1(_0876_));
 sg13g2_nand2_1 _2182_ (.Y(_0878_),
    .A(_0054_),
    .B(net522));
 sg13g2_a21oi_1 _2183_ (.A1(_0022_),
    .A2(net531),
    .Y(_0879_),
    .B1(net512));
 sg13g2_a221oi_1 _2184_ (.B2(_0879_),
    .C1(net596),
    .B1(_0878_),
    .A1(net512),
    .Y(_0880_),
    .A2(_0877_));
 sg13g2_a21oi_1 _2185_ (.A1(_0284_),
    .A2(net592),
    .Y(_0881_),
    .B1(net469));
 sg13g2_nand2b_1 _2186_ (.Y(_0882_),
    .B(_0881_),
    .A_N(_0880_));
 sg13g2_mux4_1 _2187_ (.S0(net557),
    .A0(_0151_),
    .A1(_0252_),
    .A2(_0119_),
    .A3(_0022_),
    .S1(net551),
    .X(_0883_));
 sg13g2_a21o_1 _2188_ (.A2(net596),
    .A1(_0220_),
    .B1(net495),
    .X(_0884_));
 sg13g2_a21oi_1 _2189_ (.A1(net549),
    .A2(_0883_),
    .Y(_0885_),
    .B1(_0884_));
 sg13g2_nor2b_1 _2190_ (.A(_0885_),
    .B_N(_0653_),
    .Y(_0886_));
 sg13g2_nand2b_1 _2191_ (.Y(_0887_),
    .B(_0886_),
    .A_N(_0864_));
 sg13g2_xnor2_1 _2192_ (.Y(_0888_),
    .A(_0864_),
    .B(_0886_));
 sg13g2_or2_1 _2193_ (.X(_0889_),
    .B(_0888_),
    .A(_0882_));
 sg13g2_inv_1 _2194_ (.Y(_0890_),
    .A(_0889_));
 sg13g2_xnor2_1 _2195_ (.Y(_0891_),
    .A(_0882_),
    .B(_0888_));
 sg13g2_inv_1 _2196_ (.Y(_0892_),
    .A(_0891_));
 sg13g2_nor2_1 _2197_ (.A(_0866_),
    .B(_0891_),
    .Y(_0893_));
 sg13g2_nand2_1 _2198_ (.Y(_0894_),
    .A(_0867_),
    .B(_0892_));
 sg13g2_nor2_1 _2199_ (.A(_0869_),
    .B(_0894_),
    .Y(_0895_));
 sg13g2_nand3_1 _2200_ (.B(_0871_),
    .C(_0891_),
    .A(_0866_),
    .Y(_0896_));
 sg13g2_nor3_1 _2201_ (.A(net573),
    .B(_0893_),
    .C(_0895_),
    .Y(_0897_));
 sg13g2_nand2_2 _2202_ (.Y(_0898_),
    .A(_0896_),
    .B(_0897_));
 sg13g2_nand2_1 _2203_ (.Y(_0899_),
    .A(net745),
    .B(net578));
 sg13g2_o21ai_1 _2204_ (.B1(_0899_),
    .Y(_0367_),
    .A1(net578),
    .A2(_0898_));
 sg13g2_nor2_1 _2205_ (.A(_0219_),
    .B(net521),
    .Y(_0900_));
 sg13g2_o21ai_1 _2206_ (.B1(net485),
    .Y(_0901_),
    .A1(_0084_),
    .A2(net530));
 sg13g2_a21oi_1 _2207_ (.A1(_0182_),
    .A2(net486),
    .Y(_0902_),
    .B1(net516));
 sg13g2_o21ai_1 _2208_ (.B1(_0902_),
    .Y(_0903_),
    .A1(_0900_),
    .A2(_0901_));
 sg13g2_nand2_1 _2209_ (.Y(_0904_),
    .A(_0021_),
    .B(net530));
 sg13g2_a21oi_1 _2210_ (.A1(_0053_),
    .A2(net521),
    .Y(_0905_),
    .B1(net510));
 sg13g2_a21oi_1 _2211_ (.A1(_0904_),
    .A2(_0905_),
    .Y(_0906_),
    .B1(net591));
 sg13g2_a221oi_1 _2212_ (.B2(_0906_),
    .C1(net469),
    .B1(_0903_),
    .A1(_0283_),
    .Y(_0907_),
    .A2(net591));
 sg13g2_nand2_1 _2213_ (.Y(_0908_),
    .A(_0118_),
    .B(net563));
 sg13g2_a21oi_1 _2214_ (.A1(_0021_),
    .A2(net557),
    .Y(_0909_),
    .B1(net555));
 sg13g2_nand2_1 _2215_ (.Y(_0910_),
    .A(_0251_),
    .B(net557));
 sg13g2_a21oi_1 _2216_ (.A1(_0150_),
    .A2(net563),
    .Y(_0911_),
    .B1(net550));
 sg13g2_a221oi_1 _2217_ (.B2(_0911_),
    .C1(net540),
    .B1(_0910_),
    .A1(_0908_),
    .Y(_0912_),
    .A2(_0909_));
 sg13g2_a21oi_2 _2218_ (.B1(_0912_),
    .Y(_0913_),
    .A2(net591),
    .A1(_0219_));
 sg13g2_nand2_1 _2219_ (.Y(_0914_),
    .A(_0769_),
    .B(_0913_));
 sg13g2_inv_1 _2220_ (.Y(_0915_),
    .A(_0914_));
 sg13g2_and3_1 _2221_ (.X(_0916_),
    .A(_0862_),
    .B(_0886_),
    .C(_0914_));
 sg13g2_and3_1 _2222_ (.X(_0917_),
    .A(_0819_),
    .B(_0842_),
    .C(_0916_));
 sg13g2_a21oi_1 _2223_ (.A1(_0887_),
    .A2(_0915_),
    .Y(_0918_),
    .B1(_0917_));
 sg13g2_nor2b_1 _2224_ (.A(_0918_),
    .B_N(_0907_),
    .Y(_0919_));
 sg13g2_xnor2_1 _2225_ (.Y(_0920_),
    .A(_0907_),
    .B(_0918_));
 sg13g2_nor2_1 _2226_ (.A(_0890_),
    .B(_0893_),
    .Y(_0921_));
 sg13g2_nor2b_1 _2227_ (.A(_0895_),
    .B_N(_0921_),
    .Y(_0922_));
 sg13g2_nor2b_1 _2228_ (.A(_0920_),
    .B_N(_0922_),
    .Y(_0923_));
 sg13g2_nor2b_1 _2229_ (.A(_0922_),
    .B_N(_0920_),
    .Y(_0924_));
 sg13g2_or3_2 _2230_ (.A(net573),
    .B(_0923_),
    .C(_0924_),
    .X(_0925_));
 sg13g2_nand2_1 _2231_ (.Y(_0926_),
    .A(net769),
    .B(net577));
 sg13g2_o21ai_1 _2232_ (.B1(_0926_),
    .Y(_0368_),
    .A1(net577),
    .A2(_0925_));
 sg13g2_a21oi_1 _2233_ (.A1(_0608_),
    .A2(net521),
    .Y(_0927_),
    .B1(net486));
 sg13g2_o21ai_1 _2234_ (.B1(_0927_),
    .Y(_0928_),
    .A1(_0218_),
    .A2(net521));
 sg13g2_a21oi_1 _2235_ (.A1(_0181_),
    .A2(net486),
    .Y(_0929_),
    .B1(net516));
 sg13g2_nand2_1 _2236_ (.Y(_0930_),
    .A(_0052_),
    .B(net521));
 sg13g2_a21oi_1 _2237_ (.A1(_0020_),
    .A2(net530),
    .Y(_0931_),
    .B1(net510));
 sg13g2_a221oi_1 _2238_ (.B2(_0931_),
    .C1(net591),
    .B1(_0930_),
    .A1(_0928_),
    .Y(_0932_),
    .A2(_0929_));
 sg13g2_a21o_1 _2239_ (.A2(net592),
    .A1(_0282_),
    .B1(_0932_),
    .X(_0933_));
 sg13g2_mux4_1 _2240_ (.S0(net557),
    .A0(_0149_),
    .A1(_0250_),
    .A2(_0117_),
    .A3(_0020_),
    .S1(net550),
    .X(_0934_));
 sg13g2_nand2_1 _2241_ (.Y(_0935_),
    .A(_0218_),
    .B(net540));
 sg13g2_a21oi_1 _2242_ (.A1(net547),
    .A2(_0934_),
    .Y(_0936_),
    .B1(net495));
 sg13g2_a21oi_2 _2243_ (.B1(net588),
    .Y(_0937_),
    .A2(_0936_),
    .A1(_0935_));
 sg13g2_nand4_1 _2244_ (.B(_0842_),
    .C(_0916_),
    .A(_0819_),
    .Y(_0938_),
    .D(_0937_));
 sg13g2_xor2_1 _2245_ (.B(_0937_),
    .A(_0917_),
    .X(_0939_));
 sg13g2_nor3_1 _2246_ (.A(net469),
    .B(_0933_),
    .C(_0939_),
    .Y(_0940_));
 sg13g2_o21ai_1 _2247_ (.B1(_0939_),
    .Y(_0941_),
    .A1(net469),
    .A2(_0933_));
 sg13g2_nor2b_1 _2248_ (.A(_0940_),
    .B_N(_0941_),
    .Y(_0942_));
 sg13g2_nor2_1 _2249_ (.A(_0919_),
    .B(_0924_),
    .Y(_0943_));
 sg13g2_xnor2_1 _2250_ (.Y(_0944_),
    .A(_0942_),
    .B(_0943_));
 sg13g2_nand2_2 _2251_ (.Y(_0945_),
    .A(net571),
    .B(_0944_));
 sg13g2_nand2_1 _2252_ (.Y(_0946_),
    .A(net774),
    .B(net577));
 sg13g2_o21ai_1 _2253_ (.B1(_0946_),
    .Y(_0369_),
    .A1(net577),
    .A2(_0945_));
 sg13g2_nor2_1 _2254_ (.A(_0082_),
    .B(net532),
    .Y(_0947_));
 sg13g2_nor2_1 _2255_ (.A(_0217_),
    .B(net524),
    .Y(_0948_));
 sg13g2_nor3_1 _2256_ (.A(net488),
    .B(_0947_),
    .C(_0948_),
    .Y(_0949_));
 sg13g2_a21oi_1 _2257_ (.A1(_0180_),
    .A2(net488),
    .Y(_0950_),
    .B1(_0949_));
 sg13g2_nand2_1 _2258_ (.Y(_0951_),
    .A(_0051_),
    .B(net523));
 sg13g2_a21oi_1 _2259_ (.A1(_0019_),
    .A2(net532),
    .Y(_0952_),
    .B1(net511));
 sg13g2_a221oi_1 _2260_ (.B2(_0952_),
    .C1(net594),
    .B1(_0951_),
    .A1(net511),
    .Y(_0953_),
    .A2(_0950_));
 sg13g2_a21oi_1 _2261_ (.A1(_0281_),
    .A2(net594),
    .Y(_0954_),
    .B1(net470));
 sg13g2_nand2b_1 _2262_ (.Y(_0955_),
    .B(_0954_),
    .A_N(_0953_));
 sg13g2_nand2_1 _2263_ (.Y(_0956_),
    .A(_0019_),
    .B(net559));
 sg13g2_a21oi_1 _2264_ (.A1(_0116_),
    .A2(net564),
    .Y(_0957_),
    .B1(net555));
 sg13g2_nand2_1 _2265_ (.Y(_0958_),
    .A(_0249_),
    .B(net559));
 sg13g2_a21oi_1 _2266_ (.A1(_0148_),
    .A2(net564),
    .Y(_0959_),
    .B1(net551));
 sg13g2_a221oi_1 _2267_ (.B2(_0959_),
    .C1(net542),
    .B1(_0958_),
    .A1(_0956_),
    .Y(_0960_),
    .A2(_0957_));
 sg13g2_a21o_1 _2268_ (.A2(net541),
    .A1(_0217_),
    .B1(net496),
    .X(_0961_));
 sg13g2_o21ai_1 _2269_ (.B1(_0616_),
    .Y(_0962_),
    .A1(_0960_),
    .A2(_0961_));
 sg13g2_xor2_1 _2270_ (.B(_0962_),
    .A(_0938_),
    .X(_0963_));
 sg13g2_nor2_1 _2271_ (.A(_0955_),
    .B(_0963_),
    .Y(_0964_));
 sg13g2_nand2_1 _2272_ (.Y(_0965_),
    .A(_0955_),
    .B(_0963_));
 sg13g2_nand2b_1 _2273_ (.Y(_0966_),
    .B(_0965_),
    .A_N(_0964_));
 sg13g2_a21oi_1 _2274_ (.A1(_0919_),
    .A2(_0941_),
    .Y(_0967_),
    .B1(_0940_));
 sg13g2_nand2_1 _2275_ (.Y(_0968_),
    .A(_0920_),
    .B(_0942_));
 sg13g2_nor2_1 _2276_ (.A(_0894_),
    .B(_0968_),
    .Y(_0969_));
 sg13g2_nand3_1 _2277_ (.B(_0868_),
    .C(_0969_),
    .A(_0846_),
    .Y(_0970_));
 sg13g2_o21ai_1 _2278_ (.B1(_0967_),
    .Y(_0971_),
    .A1(_0921_),
    .A2(_0968_));
 sg13g2_nand2b_1 _2279_ (.Y(_0972_),
    .B(_0970_),
    .A_N(_0971_));
 sg13g2_xnor2_1 _2280_ (.Y(_0973_),
    .A(_0966_),
    .B(_0972_));
 sg13g2_nor2_2 _2281_ (.A(net576),
    .B(_0973_),
    .Y(_0974_));
 sg13g2_nand2_1 _2282_ (.Y(_0975_),
    .A(net752),
    .B(net579));
 sg13g2_o21ai_1 _2283_ (.B1(_0975_),
    .Y(_0370_),
    .A1(net579),
    .A2(_0974_));
 sg13g2_and2_1 _2284_ (.A(_0081_),
    .B(net524),
    .X(_0976_));
 sg13g2_a21oi_1 _2285_ (.A1(_0216_),
    .A2(net533),
    .Y(_0977_),
    .B1(_0976_));
 sg13g2_nand2_1 _2286_ (.Y(_0978_),
    .A(_0050_),
    .B(net570));
 sg13g2_a21oi_1 _2287_ (.A1(_0179_),
    .A2(net489),
    .Y(_0979_),
    .B1(net517));
 sg13g2_o21ai_1 _2288_ (.B1(_0979_),
    .Y(_0980_),
    .A1(net489),
    .A2(_0977_));
 sg13g2_a21oi_1 _2289_ (.A1(_0018_),
    .A2(net533),
    .Y(_0981_),
    .B1(net511));
 sg13g2_a21oi_1 _2290_ (.A1(_0978_),
    .A2(_0981_),
    .Y(_0982_),
    .B1(net594));
 sg13g2_a221oi_1 _2291_ (.B2(_0982_),
    .C1(net470),
    .B1(_0980_),
    .A1(_0280_),
    .Y(_0983_),
    .A2(net594));
 sg13g2_mux4_1 _2292_ (.S0(net558),
    .A0(_0147_),
    .A1(_0248_),
    .A2(_0115_),
    .A3(_0018_),
    .S1(net550),
    .X(_0984_));
 sg13g2_nand2_1 _2293_ (.Y(_0985_),
    .A(_0216_),
    .B(net541));
 sg13g2_a21oi_1 _2294_ (.A1(net547),
    .A2(_0984_),
    .Y(_0986_),
    .B1(net496));
 sg13g2_a21o_1 _2295_ (.A2(_0986_),
    .A1(_0985_),
    .B1(net588),
    .X(_0987_));
 sg13g2_nor3_1 _2296_ (.A(_0938_),
    .B(_0962_),
    .C(_0987_),
    .Y(_0988_));
 sg13g2_o21ai_1 _2297_ (.B1(_0987_),
    .Y(_0989_),
    .A1(_0938_),
    .A2(_0962_));
 sg13g2_nand2b_1 _2298_ (.Y(_0990_),
    .B(_0989_),
    .A_N(_0988_));
 sg13g2_nor2_1 _2299_ (.A(_0983_),
    .B(_0990_),
    .Y(_0991_));
 sg13g2_xor2_1 _2300_ (.B(_0990_),
    .A(_0983_),
    .X(_0992_));
 sg13g2_a21oi_1 _2301_ (.A1(_0965_),
    .A2(_0972_),
    .Y(_0993_),
    .B1(_0964_));
 sg13g2_xnor2_1 _2302_ (.Y(_0994_),
    .A(_0992_),
    .B(_0993_));
 sg13g2_nand2_2 _2303_ (.Y(_0995_),
    .A(net571),
    .B(_0994_));
 sg13g2_nand2_1 _2304_ (.Y(_0996_),
    .A(net756),
    .B(net580));
 sg13g2_o21ai_1 _2305_ (.B1(_0996_),
    .Y(_0371_),
    .A1(net580),
    .A2(_0995_));
 sg13g2_nor2_1 _2306_ (.A(_0215_),
    .B(net524),
    .Y(_0997_));
 sg13g2_nor2_1 _2307_ (.A(_0080_),
    .B(net533),
    .Y(_0998_));
 sg13g2_nor3_1 _2308_ (.A(net490),
    .B(_0997_),
    .C(_0998_),
    .Y(_0999_));
 sg13g2_a21oi_1 _2309_ (.A1(_0178_),
    .A2(net490),
    .Y(_1000_),
    .B1(_0999_));
 sg13g2_nand2_1 _2310_ (.Y(_1001_),
    .A(_0049_),
    .B(net524));
 sg13g2_a21oi_1 _2311_ (.A1(_0017_),
    .A2(_0667_),
    .Y(_1002_),
    .B1(net512));
 sg13g2_a221oi_1 _2312_ (.B2(_1002_),
    .C1(net595),
    .B1(_1001_),
    .A1(net512),
    .Y(_1003_),
    .A2(_1000_));
 sg13g2_a21oi_1 _2313_ (.A1(_0279_),
    .A2(net596),
    .Y(_1004_),
    .B1(net470));
 sg13g2_nand2b_1 _2314_ (.Y(_1005_),
    .B(_1004_),
    .A_N(_1003_));
 sg13g2_nand2_1 _2315_ (.Y(_1006_),
    .A(_0017_),
    .B(net558));
 sg13g2_a21oi_1 _2316_ (.A1(_0114_),
    .A2(net564),
    .Y(_1007_),
    .B1(net555));
 sg13g2_nand2_1 _2317_ (.Y(_1008_),
    .A(_0247_),
    .B(net559));
 sg13g2_a21oi_1 _2318_ (.A1(_0146_),
    .A2(net564),
    .Y(_1009_),
    .B1(net551));
 sg13g2_a221oi_1 _2319_ (.B2(_1009_),
    .C1(net542),
    .B1(_1008_),
    .A1(_1006_),
    .Y(_1010_),
    .A2(_1007_));
 sg13g2_a21o_1 _2320_ (.A2(net541),
    .A1(_0215_),
    .B1(net496),
    .X(_1011_));
 sg13g2_o21ai_1 _2321_ (.B1(_0616_),
    .Y(_1012_),
    .A1(_1010_),
    .A2(_1011_));
 sg13g2_nor4_2 _2322_ (.A(_0938_),
    .B(_0962_),
    .C(_0987_),
    .Y(_1013_),
    .D(_1012_));
 sg13g2_xnor2_1 _2323_ (.Y(_1014_),
    .A(_0988_),
    .B(_1012_));
 sg13g2_or2_1 _2324_ (.X(_1015_),
    .B(_1014_),
    .A(_1005_));
 sg13g2_xnor2_1 _2325_ (.Y(_1016_),
    .A(_1005_),
    .B(_1014_));
 sg13g2_nor2b_1 _2326_ (.A(_0966_),
    .B_N(_0992_),
    .Y(_1017_));
 sg13g2_a21oi_1 _2327_ (.A1(_0983_),
    .A2(_0990_),
    .Y(_1018_),
    .B1(_0964_));
 sg13g2_nor2_1 _2328_ (.A(_0991_),
    .B(_1018_),
    .Y(_1019_));
 sg13g2_a21o_1 _2329_ (.A2(_1017_),
    .A1(_0972_),
    .B1(_1019_),
    .X(_1020_));
 sg13g2_nand2b_1 _2330_ (.Y(_1021_),
    .B(_1020_),
    .A_N(_1016_));
 sg13g2_nand2b_1 _2331_ (.Y(_1022_),
    .B(_1016_),
    .A_N(_1020_));
 sg13g2_a21oi_2 _2332_ (.B1(net573),
    .Y(_1023_),
    .A2(_1022_),
    .A1(_1021_));
 sg13g2_nand2_1 _2333_ (.Y(_1024_),
    .A(net751),
    .B(net581));
 sg13g2_o21ai_1 _2334_ (.B1(_1024_),
    .Y(_0372_),
    .A1(net581),
    .A2(_1023_));
 sg13g2_and2_1 _2335_ (.A(_0079_),
    .B(net523),
    .X(_1025_));
 sg13g2_a21oi_1 _2336_ (.A1(_0214_),
    .A2(net533),
    .Y(_1026_),
    .B1(_1025_));
 sg13g2_nand2_1 _2337_ (.Y(_1027_),
    .A(_0048_),
    .B(net570));
 sg13g2_a21oi_1 _2338_ (.A1(_0177_),
    .A2(net489),
    .Y(_1028_),
    .B1(net517));
 sg13g2_o21ai_1 _2339_ (.B1(_1028_),
    .Y(_1029_),
    .A1(net489),
    .A2(_1026_));
 sg13g2_a21oi_1 _2340_ (.A1(_0016_),
    .A2(net532),
    .Y(_1030_),
    .B1(net511));
 sg13g2_a21oi_1 _2341_ (.A1(_1027_),
    .A2(_1030_),
    .Y(_1031_),
    .B1(net593));
 sg13g2_a221oi_1 _2342_ (.B2(_1031_),
    .C1(net470),
    .B1(_1029_),
    .A1(_0278_),
    .Y(_1032_),
    .A2(net593));
 sg13g2_mux4_1 _2343_ (.S0(net558),
    .A0(_0145_),
    .A1(_0246_),
    .A2(_0113_),
    .A3(_0016_),
    .S1(net550),
    .X(_1033_));
 sg13g2_nand2_1 _2344_ (.Y(_1034_),
    .A(_0214_),
    .B(net541));
 sg13g2_a21oi_1 _2345_ (.A1(net547),
    .A2(_1033_),
    .Y(_1035_),
    .B1(net496));
 sg13g2_a21oi_2 _2346_ (.B1(net588),
    .Y(_1036_),
    .A2(_1035_),
    .A1(_1034_));
 sg13g2_nand2_2 _2347_ (.Y(_1037_),
    .A(_1013_),
    .B(_1036_));
 sg13g2_xnor2_1 _2348_ (.Y(_1038_),
    .A(_1013_),
    .B(_1036_));
 sg13g2_nor2_1 _2349_ (.A(_1032_),
    .B(_1038_),
    .Y(_1039_));
 sg13g2_xnor2_1 _2350_ (.Y(_1040_),
    .A(_1032_),
    .B(_1038_));
 sg13g2_and2_1 _2351_ (.A(_1015_),
    .B(_1021_),
    .X(_1041_));
 sg13g2_a21oi_1 _2352_ (.A1(_1040_),
    .A2(_1041_),
    .Y(_1042_),
    .B1(net573));
 sg13g2_o21ai_1 _2353_ (.B1(_1042_),
    .Y(_1043_),
    .A1(_1040_),
    .A2(_1041_));
 sg13g2_nand2_1 _2354_ (.Y(_1044_),
    .A(net760),
    .B(net580));
 sg13g2_o21ai_1 _2355_ (.B1(_1044_),
    .Y(_0373_),
    .A1(net580),
    .A2(_1043_));
 sg13g2_nor2_1 _2356_ (.A(_1016_),
    .B(_1040_),
    .Y(_1045_));
 sg13g2_and2_1 _2357_ (.A(_1017_),
    .B(_1045_),
    .X(_1046_));
 sg13g2_nand2_1 _2358_ (.Y(_1047_),
    .A(_0971_),
    .B(_1046_));
 sg13g2_nand4_1 _2359_ (.B(_0868_),
    .C(_0969_),
    .A(_0846_),
    .Y(_1048_),
    .D(_1046_));
 sg13g2_nor2_1 _2360_ (.A(_1015_),
    .B(_1039_),
    .Y(_1049_));
 sg13g2_a221oi_1 _2361_ (.B2(_1019_),
    .C1(_1049_),
    .B1(_1045_),
    .A1(_1032_),
    .Y(_1050_),
    .A2(_1038_));
 sg13g2_nand3_1 _2362_ (.B(_1048_),
    .C(_1050_),
    .A(_1047_),
    .Y(_1051_));
 sg13g2_nand2_1 _2363_ (.Y(_1052_),
    .A(_0047_),
    .B(net569));
 sg13g2_a21oi_1 _2364_ (.A1(_0015_),
    .A2(net537),
    .Y(_1053_),
    .B1(net515));
 sg13g2_a21oi_1 _2365_ (.A1(_1052_),
    .A2(_1053_),
    .Y(_1054_),
    .B1(net599));
 sg13g2_nor2_1 _2366_ (.A(_0213_),
    .B(net528),
    .Y(_1055_));
 sg13g2_o21ai_1 _2367_ (.B1(net484),
    .Y(_1056_),
    .A1(_0078_),
    .A2(net537));
 sg13g2_a21oi_1 _2368_ (.A1(_0176_),
    .A2(net492),
    .Y(_1057_),
    .B1(net519));
 sg13g2_o21ai_1 _2369_ (.B1(_1057_),
    .Y(_1058_),
    .A1(_1055_),
    .A2(_1056_));
 sg13g2_a221oi_1 _2370_ (.B2(_1058_),
    .C1(net472),
    .B1(_1054_),
    .A1(_0277_),
    .Y(_1059_),
    .A2(net599));
 sg13g2_nand2_1 _2371_ (.Y(_1060_),
    .A(_0015_),
    .B(net560));
 sg13g2_a21oi_1 _2372_ (.A1(_0112_),
    .A2(net567),
    .Y(_1061_),
    .B1(net555));
 sg13g2_a21oi_1 _2373_ (.A1(_0144_),
    .A2(net567),
    .Y(_1062_),
    .B1(net552));
 sg13g2_o21ai_1 _2374_ (.B1(_1062_),
    .Y(_1063_),
    .A1(_0609_),
    .A2(net567));
 sg13g2_a21oi_1 _2375_ (.A1(_1060_),
    .A2(_1061_),
    .Y(_1064_),
    .B1(net544));
 sg13g2_a221oi_1 _2376_ (.B2(_1064_),
    .C1(net499),
    .B1(_1063_),
    .A1(_0213_),
    .Y(_1065_),
    .A2(net544));
 sg13g2_nor2_1 _2377_ (.A(net589),
    .B(_1065_),
    .Y(_1066_));
 sg13g2_nand3_1 _2378_ (.B(_1036_),
    .C(_1066_),
    .A(_1013_),
    .Y(_1067_));
 sg13g2_xnor2_1 _2379_ (.Y(_1068_),
    .A(_1037_),
    .B(_1066_));
 sg13g2_nand2b_1 _2380_ (.Y(_1069_),
    .B(_1059_),
    .A_N(_1068_));
 sg13g2_xnor2_1 _2381_ (.Y(_1070_),
    .A(_1059_),
    .B(_1068_));
 sg13g2_nand2_1 _2382_ (.Y(_1071_),
    .A(_1051_),
    .B(_1070_));
 sg13g2_inv_1 _2383_ (.Y(_1072_),
    .A(_1071_));
 sg13g2_nor2_1 _2384_ (.A(net574),
    .B(_1072_),
    .Y(_1073_));
 sg13g2_o21ai_1 _2385_ (.B1(_1073_),
    .Y(_1074_),
    .A1(_1051_),
    .A2(_1070_));
 sg13g2_nand2_1 _2386_ (.Y(_1075_),
    .A(net738),
    .B(net587));
 sg13g2_o21ai_1 _2387_ (.B1(_1075_),
    .Y(_0374_),
    .A1(net586),
    .A2(_1074_));
 sg13g2_nand2_1 _2388_ (.Y(_1076_),
    .A(_0046_),
    .B(net569));
 sg13g2_nand2_1 _2389_ (.Y(_1077_),
    .A(_0276_),
    .B(net600));
 sg13g2_a21oi_1 _2390_ (.A1(_0014_),
    .A2(net537),
    .Y(_1078_),
    .B1(net515));
 sg13g2_a21oi_1 _2391_ (.A1(_1076_),
    .A2(_1078_),
    .Y(_1079_),
    .B1(net599));
 sg13g2_nor2_1 _2392_ (.A(_0212_),
    .B(net527),
    .Y(_1080_));
 sg13g2_o21ai_1 _2393_ (.B1(net484),
    .Y(_1081_),
    .A1(_0077_),
    .A2(net537));
 sg13g2_a21oi_1 _2394_ (.A1(_0175_),
    .A2(net492),
    .Y(_1082_),
    .B1(net519));
 sg13g2_o21ai_1 _2395_ (.B1(_1082_),
    .Y(_1083_),
    .A1(_1080_),
    .A2(_1081_));
 sg13g2_a21oi_1 _2396_ (.A1(_1079_),
    .A2(_1083_),
    .Y(_1084_),
    .B1(net472));
 sg13g2_nand2_1 _2397_ (.Y(_1085_),
    .A(_0014_),
    .B(net562));
 sg13g2_a21oi_1 _2398_ (.A1(_0111_),
    .A2(net565),
    .Y(_1086_),
    .B1(net556));
 sg13g2_nand2_1 _2399_ (.Y(_1087_),
    .A(_0244_),
    .B(net562));
 sg13g2_a21oi_1 _2400_ (.A1(_0143_),
    .A2(net565),
    .Y(_1088_),
    .B1(net554));
 sg13g2_a221oi_1 _2401_ (.B2(_1088_),
    .C1(net544),
    .B1(_1087_),
    .A1(_1085_),
    .Y(_1089_),
    .A2(_1086_));
 sg13g2_a21o_1 _2402_ (.A2(net543),
    .A1(_0212_),
    .B1(net498),
    .X(_1090_));
 sg13g2_o21ai_1 _2403_ (.B1(_0616_),
    .Y(_1091_),
    .A1(_1089_),
    .A2(_1090_));
 sg13g2_inv_1 _2404_ (.Y(_1092_),
    .A(_1091_));
 sg13g2_nand4_1 _2405_ (.B(_1036_),
    .C(_1066_),
    .A(_1013_),
    .Y(_1093_),
    .D(_1092_));
 sg13g2_xnor2_1 _2406_ (.Y(_1094_),
    .A(_1067_),
    .B(_1091_));
 sg13g2_a21oi_1 _2407_ (.A1(_1077_),
    .A2(_1084_),
    .Y(_1095_),
    .B1(_1094_));
 sg13g2_nand3_1 _2408_ (.B(_1084_),
    .C(_1094_),
    .A(_1077_),
    .Y(_1096_));
 sg13g2_nor2b_1 _2409_ (.A(_1095_),
    .B_N(_1096_),
    .Y(_1097_));
 sg13g2_nand2_1 _2410_ (.Y(_1098_),
    .A(_1069_),
    .B(_1071_));
 sg13g2_a21oi_1 _2411_ (.A1(_1097_),
    .A2(_1098_),
    .Y(_1099_),
    .B1(net574));
 sg13g2_o21ai_1 _2412_ (.B1(_1099_),
    .Y(_1100_),
    .A1(_1097_),
    .A2(_1098_));
 sg13g2_nand2_1 _2413_ (.Y(_1101_),
    .A(net739),
    .B(net586));
 sg13g2_o21ai_1 _2414_ (.B1(_1101_),
    .Y(_0375_),
    .A1(net586),
    .A2(_1100_));
 sg13g2_nand2_1 _2415_ (.Y(_1102_),
    .A(_0013_),
    .B(_0667_));
 sg13g2_a21oi_1 _2416_ (.A1(_0045_),
    .A2(net527),
    .Y(_1103_),
    .B1(net514));
 sg13g2_a21oi_1 _2417_ (.A1(_1102_),
    .A2(_1103_),
    .Y(_1104_),
    .B1(net599));
 sg13g2_nor2_1 _2418_ (.A(_0211_),
    .B(net527),
    .Y(_1105_));
 sg13g2_o21ai_1 _2419_ (.B1(_0672_),
    .Y(_1106_),
    .A1(_0076_),
    .A2(net536));
 sg13g2_a21oi_1 _2420_ (.A1(_0174_),
    .A2(net492),
    .Y(_1107_),
    .B1(net519));
 sg13g2_o21ai_1 _2421_ (.B1(_1107_),
    .Y(_1108_),
    .A1(_1105_),
    .A2(_1106_));
 sg13g2_a221oi_1 _2422_ (.B2(_1108_),
    .C1(net472),
    .B1(_1104_),
    .A1(_0275_),
    .Y(_1109_),
    .A2(net599));
 sg13g2_mux4_1 _2423_ (.S0(net562),
    .A0(_0142_),
    .A1(_0243_),
    .A2(_0110_),
    .A3(_0013_),
    .S1(net552),
    .X(_1110_));
 sg13g2_a21o_1 _2424_ (.A2(_1110_),
    .A1(net549),
    .B1(net498),
    .X(_1111_));
 sg13g2_a21oi_1 _2425_ (.A1(_0211_),
    .A2(net544),
    .Y(_1112_),
    .B1(_1111_));
 sg13g2_nor2_1 _2426_ (.A(_1093_),
    .B(_1112_),
    .Y(_1113_));
 sg13g2_o21ai_1 _2427_ (.B1(_1093_),
    .Y(_1114_),
    .A1(net589),
    .A2(_1112_));
 sg13g2_nor2b_1 _2428_ (.A(_1113_),
    .B_N(_1114_),
    .Y(_1115_));
 sg13g2_nor2b_1 _2429_ (.A(_1115_),
    .B_N(_1109_),
    .Y(_1116_));
 sg13g2_xnor2_1 _2430_ (.Y(_1117_),
    .A(_1109_),
    .B(_1115_));
 sg13g2_o21ai_1 _2431_ (.B1(_1096_),
    .Y(_1118_),
    .A1(_1069_),
    .A2(_1095_));
 sg13g2_a21oi_1 _2432_ (.A1(_1072_),
    .A2(_1097_),
    .Y(_1119_),
    .B1(_1118_));
 sg13g2_nor2b_1 _2433_ (.A(_1119_),
    .B_N(_1117_),
    .Y(_1120_));
 sg13g2_xnor2_1 _2434_ (.Y(_1121_),
    .A(_1117_),
    .B(_1119_));
 sg13g2_nor2_2 _2435_ (.A(net574),
    .B(_1121_),
    .Y(_1122_));
 sg13g2_nand2_1 _2436_ (.Y(_1123_),
    .A(net724),
    .B(net587));
 sg13g2_o21ai_1 _2437_ (.B1(_1123_),
    .Y(_0376_),
    .A1(net587),
    .A2(_1122_));
 sg13g2_and2_1 _2438_ (.A(_0075_),
    .B(net527),
    .X(_1124_));
 sg13g2_a21oi_1 _2439_ (.A1(_0210_),
    .A2(net536),
    .Y(_1125_),
    .B1(_1124_));
 sg13g2_nand2_1 _2440_ (.Y(_1126_),
    .A(_0012_),
    .B(_0667_));
 sg13g2_a21oi_1 _2441_ (.A1(_0173_),
    .A2(net492),
    .Y(_1127_),
    .B1(net518));
 sg13g2_o21ai_1 _2442_ (.B1(_1127_),
    .Y(_1128_),
    .A1(net492),
    .A2(_1125_));
 sg13g2_a21oi_1 _2443_ (.A1(_0044_),
    .A2(net528),
    .Y(_1129_),
    .B1(net514));
 sg13g2_a21oi_1 _2444_ (.A1(_1126_),
    .A2(_1129_),
    .Y(_1130_),
    .B1(net599));
 sg13g2_a221oi_1 _2445_ (.B2(_1130_),
    .C1(net472),
    .B1(_1128_),
    .A1(_0274_),
    .Y(_1131_),
    .A2(net599));
 sg13g2_nand2_1 _2446_ (.Y(_1132_),
    .A(_0012_),
    .B(net560));
 sg13g2_a21oi_1 _2447_ (.A1(_0109_),
    .A2(net565),
    .Y(_1133_),
    .B1(net556));
 sg13g2_a21oi_1 _2448_ (.A1(_0141_),
    .A2(net565),
    .Y(_1134_),
    .B1(net552));
 sg13g2_o21ai_1 _2449_ (.B1(_1134_),
    .Y(_1135_),
    .A1(_0610_),
    .A2(net565));
 sg13g2_a21oi_1 _2450_ (.A1(_1132_),
    .A2(_1133_),
    .Y(_1136_),
    .B1(net544));
 sg13g2_a221oi_1 _2451_ (.B2(_1136_),
    .C1(net498),
    .B1(_1135_),
    .A1(_0210_),
    .Y(_1137_),
    .A2(net543));
 sg13g2_nor2_1 _2452_ (.A(net590),
    .B(_1137_),
    .Y(_1138_));
 sg13g2_or4_2 _2453_ (.A(_1065_),
    .B(_1091_),
    .C(_1112_),
    .D(_1137_),
    .X(_1139_));
 sg13g2_xor2_1 _2454_ (.B(_1138_),
    .A(_1113_),
    .X(_1140_));
 sg13g2_nor2b_1 _2455_ (.A(_1140_),
    .B_N(_1131_),
    .Y(_1141_));
 sg13g2_nand2b_1 _2456_ (.Y(_1142_),
    .B(_1140_),
    .A_N(_1131_));
 sg13g2_xnor2_1 _2457_ (.Y(_1143_),
    .A(_1131_),
    .B(_1140_));
 sg13g2_nor2_1 _2458_ (.A(_1116_),
    .B(_1120_),
    .Y(_1144_));
 sg13g2_xnor2_1 _2459_ (.Y(_1145_),
    .A(_1143_),
    .B(_1144_));
 sg13g2_nand2_2 _2460_ (.Y(_1146_),
    .A(net572),
    .B(_1145_));
 sg13g2_nand2_1 _2461_ (.Y(_1147_),
    .A(net746),
    .B(net586));
 sg13g2_o21ai_1 _2462_ (.B1(_1147_),
    .Y(_0377_),
    .A1(net586),
    .A2(_1146_));
 sg13g2_nor2_1 _2463_ (.A(_0074_),
    .B(net536),
    .Y(_1148_));
 sg13g2_nor2_1 _2464_ (.A(_0209_),
    .B(net527),
    .Y(_1149_));
 sg13g2_nor3_1 _2465_ (.A(net492),
    .B(_1148_),
    .C(_1149_),
    .Y(_1150_));
 sg13g2_a21oi_1 _2466_ (.A1(_0172_),
    .A2(net492),
    .Y(_1151_),
    .B1(_1150_));
 sg13g2_nand2_1 _2467_ (.Y(_1152_),
    .A(_0043_),
    .B(net527));
 sg13g2_a21oi_1 _2468_ (.A1(_0011_),
    .A2(net536),
    .Y(_1153_),
    .B1(net514));
 sg13g2_a221oi_1 _2469_ (.B2(_1153_),
    .C1(net600),
    .B1(_1152_),
    .A1(net514),
    .Y(_1154_),
    .A2(_1151_));
 sg13g2_a21oi_1 _2470_ (.A1(_0273_),
    .A2(net600),
    .Y(_1155_),
    .B1(net472));
 sg13g2_nand2b_1 _2471_ (.Y(_1156_),
    .B(_1155_),
    .A_N(_1154_));
 sg13g2_mux4_1 _2472_ (.S0(net560),
    .A0(_0140_),
    .A1(_0241_),
    .A2(_0108_),
    .A3(_0011_),
    .S1(net553),
    .X(_1157_));
 sg13g2_nand2_1 _2473_ (.Y(_1158_),
    .A(net548),
    .B(_1157_));
 sg13g2_a21oi_1 _2474_ (.A1(_0209_),
    .A2(net543),
    .Y(_1159_),
    .B1(net498));
 sg13g2_a21oi_1 _2475_ (.A1(_1158_),
    .A2(_1159_),
    .Y(_1160_),
    .B1(net589));
 sg13g2_inv_1 _2476_ (.Y(_1161_),
    .A(_1160_));
 sg13g2_nor3_1 _2477_ (.A(_1037_),
    .B(_1139_),
    .C(_1161_),
    .Y(_1162_));
 sg13g2_o21ai_1 _2478_ (.B1(_1161_),
    .Y(_1163_),
    .A1(_1037_),
    .A2(_1139_));
 sg13g2_nand2b_1 _2479_ (.Y(_1164_),
    .B(_1163_),
    .A_N(_1162_));
 sg13g2_nor2b_1 _2480_ (.A(_1156_),
    .B_N(_1164_),
    .Y(_1165_));
 sg13g2_xnor2_1 _2481_ (.Y(_1166_),
    .A(_1156_),
    .B(_1164_));
 sg13g2_and2_1 _2482_ (.A(_1117_),
    .B(_1143_),
    .X(_1167_));
 sg13g2_and3_1 _2483_ (.X(_1168_),
    .A(_1070_),
    .B(_1097_),
    .C(_1167_));
 sg13g2_a21o_1 _2484_ (.A2(_1142_),
    .A1(_1116_),
    .B1(_1141_),
    .X(_1169_));
 sg13g2_a221oi_1 _2485_ (.B2(_1051_),
    .C1(_1169_),
    .B1(_1168_),
    .A1(_1118_),
    .Y(_1170_),
    .A2(_1167_));
 sg13g2_nand2b_1 _2486_ (.Y(_1171_),
    .B(_1166_),
    .A_N(_1170_));
 sg13g2_nand2b_1 _2487_ (.Y(_1172_),
    .B(_1170_),
    .A_N(_1166_));
 sg13g2_a21oi_2 _2488_ (.B1(net574),
    .Y(_1173_),
    .A2(_1172_),
    .A1(_1171_));
 sg13g2_nand2_1 _2489_ (.Y(_1174_),
    .A(net768),
    .B(net587));
 sg13g2_o21ai_1 _2490_ (.B1(_1174_),
    .Y(_0378_),
    .A1(net587),
    .A2(_1173_));
 sg13g2_nor2_1 _2491_ (.A(_0208_),
    .B(net527),
    .Y(_1175_));
 sg13g2_o21ai_1 _2492_ (.B1(net484),
    .Y(_1176_),
    .A1(_0073_),
    .A2(net536));
 sg13g2_a21oi_1 _2493_ (.A1(_0171_),
    .A2(net492),
    .Y(_1177_),
    .B1(net519));
 sg13g2_o21ai_1 _2494_ (.B1(_1177_),
    .Y(_1178_),
    .A1(_1175_),
    .A2(_1176_));
 sg13g2_nand2_1 _2495_ (.Y(_1179_),
    .A(_0010_),
    .B(net536));
 sg13g2_a21oi_1 _2496_ (.A1(_0042_),
    .A2(net569),
    .Y(_1180_),
    .B1(net514));
 sg13g2_a21oi_1 _2497_ (.A1(_1179_),
    .A2(_1180_),
    .Y(_1181_),
    .B1(net600));
 sg13g2_a221oi_1 _2498_ (.B2(_1181_),
    .C1(net472),
    .B1(_1178_),
    .A1(_0272_),
    .Y(_1182_),
    .A2(net600));
 sg13g2_nand2_1 _2499_ (.Y(_1183_),
    .A(_0010_),
    .B(net560));
 sg13g2_a21oi_1 _2500_ (.A1(_0107_),
    .A2(net565),
    .Y(_1184_),
    .B1(net556));
 sg13g2_nand2_1 _2501_ (.Y(_1185_),
    .A(_0240_),
    .B(net560));
 sg13g2_a21oi_1 _2502_ (.A1(_0139_),
    .A2(net565),
    .Y(_1186_),
    .B1(net553));
 sg13g2_a221oi_1 _2503_ (.B2(_1186_),
    .C1(net543),
    .B1(_1185_),
    .A1(_1183_),
    .Y(_1187_),
    .A2(_1184_));
 sg13g2_a21oi_1 _2504_ (.A1(_0208_),
    .A2(net543),
    .Y(_1188_),
    .B1(_1187_));
 sg13g2_nand2_1 _2505_ (.Y(_1189_),
    .A(_0662_),
    .B(_1188_));
 sg13g2_nand2_1 _2506_ (.Y(_1190_),
    .A(_0616_),
    .B(_1189_));
 sg13g2_nand2_1 _2507_ (.Y(_1191_),
    .A(_1160_),
    .B(_1189_));
 sg13g2_nor3_1 _2508_ (.A(_1037_),
    .B(_1139_),
    .C(_1191_),
    .Y(_1192_));
 sg13g2_xnor2_1 _2509_ (.Y(_1193_),
    .A(_1162_),
    .B(_1190_));
 sg13g2_nand2b_1 _2510_ (.Y(_1194_),
    .B(_1193_),
    .A_N(_1182_));
 sg13g2_nor2b_1 _2511_ (.A(_1193_),
    .B_N(_1182_),
    .Y(_1195_));
 sg13g2_xnor2_1 _2512_ (.Y(_1196_),
    .A(_1182_),
    .B(_1193_));
 sg13g2_nand2b_1 _2513_ (.Y(_1197_),
    .B(_1171_),
    .A_N(_1165_));
 sg13g2_xor2_1 _2514_ (.B(_1197_),
    .A(_1196_),
    .X(_1198_));
 sg13g2_nor2_2 _2515_ (.A(net574),
    .B(_1198_),
    .Y(_1199_));
 sg13g2_nand2_1 _2516_ (.Y(_1200_),
    .A(net733),
    .B(net587));
 sg13g2_o21ai_1 _2517_ (.B1(_1200_),
    .Y(_0379_),
    .A1(net584),
    .A2(_1199_));
 sg13g2_nand2_1 _2518_ (.Y(_1201_),
    .A(_0041_),
    .B(net569));
 sg13g2_a21oi_1 _2519_ (.A1(_0009_),
    .A2(net536),
    .Y(_1202_),
    .B1(net514));
 sg13g2_a21oi_1 _2520_ (.A1(_1201_),
    .A2(_1202_),
    .Y(_1203_),
    .B1(net595));
 sg13g2_nor2_1 _2521_ (.A(_0207_),
    .B(net527),
    .Y(_1204_));
 sg13g2_o21ai_1 _2522_ (.B1(net485),
    .Y(_1205_),
    .A1(_0072_),
    .A2(net536));
 sg13g2_a21oi_1 _2523_ (.A1(_0170_),
    .A2(net490),
    .Y(_1206_),
    .B1(net517));
 sg13g2_o21ai_1 _2524_ (.B1(_1206_),
    .Y(_1207_),
    .A1(_1204_),
    .A2(_1205_));
 sg13g2_a22oi_1 _2525_ (.Y(_1208_),
    .B1(_1203_),
    .B2(_1207_),
    .A2(net595),
    .A1(_0271_));
 sg13g2_nand2_1 _2526_ (.Y(_1209_),
    .A(_0684_),
    .B(_1208_));
 sg13g2_mux4_1 _2527_ (.S0(net560),
    .A0(_0138_),
    .A1(_0239_),
    .A2(_0106_),
    .A3(_0009_),
    .S1(net553),
    .X(_1210_));
 sg13g2_nand2_1 _2528_ (.Y(_1211_),
    .A(net549),
    .B(_1210_));
 sg13g2_a21oi_1 _2529_ (.A1(_0207_),
    .A2(net543),
    .Y(_1212_),
    .B1(net498));
 sg13g2_a21oi_1 _2530_ (.A1(_1211_),
    .A2(_1212_),
    .Y(_1213_),
    .B1(net589));
 sg13g2_inv_1 _2531_ (.Y(_1214_),
    .A(_1213_));
 sg13g2_nor4_2 _2532_ (.A(_1037_),
    .B(_1139_),
    .C(_1191_),
    .Y(_1215_),
    .D(_1214_));
 sg13g2_xnor2_1 _2533_ (.Y(_1216_),
    .A(_1192_),
    .B(_1213_));
 sg13g2_nand2b_1 _2534_ (.Y(_1217_),
    .B(_1216_),
    .A_N(_1209_));
 sg13g2_xnor2_1 _2535_ (.Y(_1218_),
    .A(_1209_),
    .B(_1216_));
 sg13g2_a21oi_1 _2536_ (.A1(_1165_),
    .A2(_1194_),
    .Y(_1219_),
    .B1(_1195_));
 sg13g2_nand2_1 _2537_ (.Y(_1220_),
    .A(_1166_),
    .B(_1196_));
 sg13g2_o21ai_1 _2538_ (.B1(_1219_),
    .Y(_1221_),
    .A1(_1170_),
    .A2(_1220_));
 sg13g2_nand2_1 _2539_ (.Y(_1222_),
    .A(_1218_),
    .B(_1221_));
 sg13g2_o21ai_1 _2540_ (.B1(net571),
    .Y(_1223_),
    .A1(_1218_),
    .A2(_1221_));
 sg13g2_nand2b_2 _2541_ (.Y(_1224_),
    .B(_1222_),
    .A_N(_1223_));
 sg13g2_nand2_1 _2542_ (.Y(_1225_),
    .A(net773),
    .B(net582));
 sg13g2_o21ai_1 _2543_ (.B1(_1225_),
    .Y(_0380_),
    .A1(net582),
    .A2(_1224_));
 sg13g2_nand2b_1 _2544_ (.Y(_1226_),
    .B(net485),
    .A_N(_0206_));
 sg13g2_o21ai_1 _2545_ (.B1(_1226_),
    .Y(_1227_),
    .A1(_0169_),
    .A2(net485));
 sg13g2_nand2_1 _2546_ (.Y(_1228_),
    .A(_0040_),
    .B(net524));
 sg13g2_a21oi_1 _2547_ (.A1(_0008_),
    .A2(_0667_),
    .Y(_1229_),
    .B1(net514));
 sg13g2_a221oi_1 _2548_ (.B2(_1229_),
    .C1(net600),
    .B1(_1228_),
    .A1(net514),
    .Y(_1230_),
    .A2(_1227_));
 sg13g2_a21oi_1 _2549_ (.A1(_0270_),
    .A2(net595),
    .Y(_1231_),
    .B1(_1230_));
 sg13g2_nand2_1 _2550_ (.Y(_1232_),
    .A(_0684_),
    .B(_1231_));
 sg13g2_nand2_1 _2551_ (.Y(_1233_),
    .A(_0008_),
    .B(net560));
 sg13g2_a21oi_1 _2552_ (.A1(_0105_),
    .A2(net563),
    .Y(_1234_),
    .B1(net555));
 sg13g2_nand2_1 _2553_ (.Y(_1235_),
    .A(_0238_),
    .B(net560));
 sg13g2_a21oi_1 _2554_ (.A1(_0137_),
    .A2(net565),
    .Y(_1236_),
    .B1(net553));
 sg13g2_a221oi_1 _2555_ (.B2(_1236_),
    .C1(net543),
    .B1(_1235_),
    .A1(_1233_),
    .Y(_1237_),
    .A2(_1234_));
 sg13g2_a21oi_1 _2556_ (.A1(_0206_),
    .A2(net543),
    .Y(_1238_),
    .B1(_1237_));
 sg13g2_nand2_2 _2557_ (.Y(_1239_),
    .A(_0662_),
    .B(_1238_));
 sg13g2_inv_1 _2558_ (.Y(_1240_),
    .A(_1239_));
 sg13g2_nor2_1 _2559_ (.A(net590),
    .B(_1240_),
    .Y(_1241_));
 sg13g2_mux2_1 _2560_ (.A0(_1241_),
    .A1(_1240_),
    .S(_1215_),
    .X(_1242_));
 sg13g2_nand2_1 _2561_ (.Y(_1243_),
    .A(_1232_),
    .B(_1242_));
 sg13g2_nor2_1 _2562_ (.A(_1232_),
    .B(_1242_),
    .Y(_1244_));
 sg13g2_xnor2_1 _2563_ (.Y(_1245_),
    .A(_1232_),
    .B(_1242_));
 sg13g2_nand2_1 _2564_ (.Y(_1246_),
    .A(_1217_),
    .B(_1222_));
 sg13g2_xnor2_1 _2565_ (.Y(_1247_),
    .A(_1245_),
    .B(_1246_));
 sg13g2_nand2_2 _2566_ (.Y(_1248_),
    .A(net571),
    .B(_1247_));
 sg13g2_nand2_1 _2567_ (.Y(_1249_),
    .A(net772),
    .B(net583));
 sg13g2_o21ai_1 _2568_ (.B1(_1249_),
    .Y(_0381_),
    .A1(net582),
    .A2(_1248_));
 sg13g2_nand3b_1 _2569_ (.B(_1218_),
    .C(_1243_),
    .Y(_1250_),
    .A_N(_1244_));
 sg13g2_or2_1 _2570_ (.X(_1251_),
    .B(_1250_),
    .A(_1220_));
 sg13g2_nor2_1 _2571_ (.A(_1170_),
    .B(_1251_),
    .Y(_1252_));
 sg13g2_nor2_1 _2572_ (.A(_1219_),
    .B(_1250_),
    .Y(_1253_));
 sg13g2_nor2b_1 _2573_ (.A(_1217_),
    .B_N(_1243_),
    .Y(_1254_));
 sg13g2_nor3_1 _2574_ (.A(_1244_),
    .B(_1253_),
    .C(_1254_),
    .Y(_1255_));
 sg13g2_nor2b_2 _2575_ (.A(_1252_),
    .B_N(_1255_),
    .Y(_1256_));
 sg13g2_o21ai_1 _2576_ (.B1(_1255_),
    .Y(_1257_),
    .A1(_1170_),
    .A2(_1251_));
 sg13g2_and2_1 _2577_ (.A(_0071_),
    .B(net523),
    .X(_1258_));
 sg13g2_a21oi_1 _2578_ (.A1(_0205_),
    .A2(net532),
    .Y(_1259_),
    .B1(_1258_));
 sg13g2_a21oi_1 _2579_ (.A1(_0168_),
    .A2(net488),
    .Y(_1260_),
    .B1(net516));
 sg13g2_o21ai_1 _2580_ (.B1(_1260_),
    .Y(_1261_),
    .A1(net488),
    .A2(_1259_));
 sg13g2_nand2_1 _2581_ (.Y(_1262_),
    .A(_0007_),
    .B(net532));
 sg13g2_a21oi_1 _2582_ (.A1(_0039_),
    .A2(net523),
    .Y(_1263_),
    .B1(net511));
 sg13g2_a21oi_1 _2583_ (.A1(_1262_),
    .A2(_1263_),
    .Y(_1264_),
    .B1(net593));
 sg13g2_a221oi_1 _2584_ (.B2(_1264_),
    .C1(net470),
    .B1(_1261_),
    .A1(_0269_),
    .Y(_1265_),
    .A2(net593));
 sg13g2_mux4_1 _2585_ (.S0(net558),
    .A0(_0136_),
    .A1(_0237_),
    .A2(_0104_),
    .A3(_0007_),
    .S1(net551),
    .X(_1266_));
 sg13g2_nand2_1 _2586_ (.Y(_1267_),
    .A(net547),
    .B(_1266_));
 sg13g2_a21oi_1 _2587_ (.A1(_0205_),
    .A2(net541),
    .Y(_1268_),
    .B1(net495));
 sg13g2_a21oi_2 _2588_ (.B1(net588),
    .Y(_1269_),
    .A2(_1268_),
    .A1(_1267_));
 sg13g2_nand3_1 _2589_ (.B(_1239_),
    .C(_1269_),
    .A(_1215_),
    .Y(_1270_));
 sg13g2_a21o_1 _2590_ (.A2(_1239_),
    .A1(_1215_),
    .B1(_1269_),
    .X(_1271_));
 sg13g2_and2_1 _2591_ (.A(_1270_),
    .B(_1271_),
    .X(_1272_));
 sg13g2_nor2b_1 _2592_ (.A(_1272_),
    .B_N(_1265_),
    .Y(_1273_));
 sg13g2_xnor2_1 _2593_ (.Y(_1274_),
    .A(_1265_),
    .B(_1272_));
 sg13g2_a21oi_1 _2594_ (.A1(_1257_),
    .A2(_1274_),
    .Y(_1275_),
    .B1(net573));
 sg13g2_o21ai_1 _2595_ (.B1(_1275_),
    .Y(_1276_),
    .A1(_1257_),
    .A2(_1274_));
 sg13g2_nand2_1 _2596_ (.Y(_1277_),
    .A(net761),
    .B(net579));
 sg13g2_o21ai_1 _2597_ (.B1(_1277_),
    .Y(_0382_),
    .A1(net579),
    .A2(_1276_));
 sg13g2_nand2b_1 _2598_ (.Y(_1278_),
    .B(net523),
    .A_N(_0070_));
 sg13g2_o21ai_1 _2599_ (.B1(_1278_),
    .Y(_1279_),
    .A1(_0204_),
    .A2(net523));
 sg13g2_a21oi_1 _2600_ (.A1(_0167_),
    .A2(net488),
    .Y(_1280_),
    .B1(net517));
 sg13g2_o21ai_1 _2601_ (.B1(_1280_),
    .Y(_1281_),
    .A1(net488),
    .A2(_1279_));
 sg13g2_nand2_1 _2602_ (.Y(_1282_),
    .A(_0006_),
    .B(net532));
 sg13g2_a21oi_1 _2603_ (.A1(_0038_),
    .A2(net570),
    .Y(_1283_),
    .B1(net511));
 sg13g2_a21oi_1 _2604_ (.A1(_1282_),
    .A2(_1283_),
    .Y(_1284_),
    .B1(net593));
 sg13g2_a221oi_1 _2605_ (.B2(_1284_),
    .C1(net470),
    .B1(_1281_),
    .A1(_0268_),
    .Y(_1285_),
    .A2(net593));
 sg13g2_nand2_1 _2606_ (.Y(_1286_),
    .A(_0006_),
    .B(net558));
 sg13g2_a21oi_1 _2607_ (.A1(_0103_),
    .A2(net564),
    .Y(_1287_),
    .B1(net555));
 sg13g2_nand2_1 _2608_ (.Y(_1288_),
    .A(_0236_),
    .B(net558));
 sg13g2_a21oi_1 _2609_ (.A1(_0135_),
    .A2(net564),
    .Y(_1289_),
    .B1(net550));
 sg13g2_a221oi_1 _2610_ (.B2(_1289_),
    .C1(net541),
    .B1(_1288_),
    .A1(_1286_),
    .Y(_1290_),
    .A2(_1287_));
 sg13g2_a21o_1 _2611_ (.A2(net541),
    .A1(_0204_),
    .B1(net495),
    .X(_1291_));
 sg13g2_o21ai_1 _2612_ (.B1(_0616_),
    .Y(_1292_),
    .A1(_1290_),
    .A2(_1291_));
 sg13g2_inv_1 _2613_ (.Y(_1293_),
    .A(_1292_));
 sg13g2_nand4_1 _2614_ (.B(_1239_),
    .C(_1269_),
    .A(_1215_),
    .Y(_1294_),
    .D(_1293_));
 sg13g2_xnor2_1 _2615_ (.Y(_1295_),
    .A(_1270_),
    .B(_1293_));
 sg13g2_nand2b_1 _2616_ (.Y(_1296_),
    .B(_1295_),
    .A_N(_1285_));
 sg13g2_nor2b_1 _2617_ (.A(_1295_),
    .B_N(_1285_),
    .Y(_1297_));
 sg13g2_xnor2_1 _2618_ (.Y(_1298_),
    .A(_1285_),
    .B(_1295_));
 sg13g2_a21oi_1 _2619_ (.A1(_1257_),
    .A2(_1274_),
    .Y(_1299_),
    .B1(_1273_));
 sg13g2_o21ai_1 _2620_ (.B1(net571),
    .Y(_1300_),
    .A1(_1298_),
    .A2(_1299_));
 sg13g2_a21oi_2 _2621_ (.B1(_1300_),
    .Y(_1301_),
    .A2(_1299_),
    .A1(_1298_));
 sg13g2_nand2_1 _2622_ (.Y(_1302_),
    .A(net735),
    .B(net579));
 sg13g2_o21ai_1 _2623_ (.B1(_1302_),
    .Y(_0383_),
    .A1(net579),
    .A2(_1301_));
 sg13g2_nor2_1 _2624_ (.A(_0069_),
    .B(net532),
    .Y(_1303_));
 sg13g2_nor2_1 _2625_ (.A(_0203_),
    .B(net523),
    .Y(_1304_));
 sg13g2_nor3_1 _2626_ (.A(net488),
    .B(_1303_),
    .C(_1304_),
    .Y(_1305_));
 sg13g2_a21oi_1 _2627_ (.A1(_0166_),
    .A2(net488),
    .Y(_1306_),
    .B1(_1305_));
 sg13g2_nand2_1 _2628_ (.Y(_1307_),
    .A(_0037_),
    .B(net523));
 sg13g2_a21oi_1 _2629_ (.A1(_0005_),
    .A2(net532),
    .Y(_1308_),
    .B1(net511));
 sg13g2_a221oi_1 _2630_ (.B2(_1308_),
    .C1(net593),
    .B1(_1307_),
    .A1(net511),
    .Y(_1309_),
    .A2(_1306_));
 sg13g2_a21oi_1 _2631_ (.A1(_0267_),
    .A2(net593),
    .Y(_1310_),
    .B1(net470));
 sg13g2_nand2b_1 _2632_ (.Y(_1311_),
    .B(_1310_),
    .A_N(_1309_));
 sg13g2_mux4_1 _2633_ (.S0(net558),
    .A0(_0134_),
    .A1(_0235_),
    .A2(_0102_),
    .A3(_0005_),
    .S1(net550),
    .X(_1312_));
 sg13g2_nand2_1 _2634_ (.Y(_1313_),
    .A(net547),
    .B(_1312_));
 sg13g2_a21oi_1 _2635_ (.A1(_0203_),
    .A2(net541),
    .Y(_1314_),
    .B1(net496));
 sg13g2_a21oi_1 _2636_ (.A1(_1313_),
    .A2(_1314_),
    .Y(_1315_),
    .B1(net588));
 sg13g2_nor2b_1 _2637_ (.A(_1294_),
    .B_N(_1315_),
    .Y(_1316_));
 sg13g2_xnor2_1 _2638_ (.Y(_1317_),
    .A(_1294_),
    .B(_1315_));
 sg13g2_nor2_1 _2639_ (.A(_1311_),
    .B(_1317_),
    .Y(_1318_));
 sg13g2_inv_1 _2640_ (.Y(_1319_),
    .A(_1318_));
 sg13g2_xnor2_1 _2641_ (.Y(_1320_),
    .A(_1311_),
    .B(_1317_));
 sg13g2_a21oi_1 _2642_ (.A1(_1273_),
    .A2(_1296_),
    .Y(_1321_),
    .B1(_1297_));
 sg13g2_nand2_1 _2643_ (.Y(_1322_),
    .A(_1274_),
    .B(_1298_));
 sg13g2_o21ai_1 _2644_ (.B1(_1321_),
    .Y(_1323_),
    .A1(_1256_),
    .A2(_1322_));
 sg13g2_nand2b_1 _2645_ (.Y(_1324_),
    .B(_1320_),
    .A_N(_1323_));
 sg13g2_nand2b_1 _2646_ (.Y(_1325_),
    .B(_1323_),
    .A_N(_1320_));
 sg13g2_nand3_1 _2647_ (.B(_1324_),
    .C(_1325_),
    .A(net571),
    .Y(_1326_));
 sg13g2_nand2_1 _2648_ (.Y(_1327_),
    .A(net762),
    .B(net579));
 sg13g2_o21ai_1 _2649_ (.B1(_1327_),
    .Y(_0384_),
    .A1(net579),
    .A2(_1326_));
 sg13g2_nand2b_1 _2650_ (.Y(_1328_),
    .B(net526),
    .A_N(_0068_));
 sg13g2_o21ai_1 _2651_ (.B1(_1328_),
    .Y(_1329_),
    .A1(_0202_),
    .A2(net524));
 sg13g2_a21oi_1 _2652_ (.A1(_0165_),
    .A2(net490),
    .Y(_1330_),
    .B1(net516));
 sg13g2_o21ai_1 _2653_ (.B1(_1330_),
    .Y(_1331_),
    .A1(net486),
    .A2(_1329_));
 sg13g2_nand2_1 _2654_ (.Y(_1332_),
    .A(_0004_),
    .B(net531));
 sg13g2_a21oi_1 _2655_ (.A1(_0036_),
    .A2(net524),
    .Y(_1333_),
    .B1(net512));
 sg13g2_a21oi_1 _2656_ (.A1(_1332_),
    .A2(_1333_),
    .Y(_1334_),
    .B1(net595));
 sg13g2_a221oi_1 _2657_ (.B2(_1334_),
    .C1(net470),
    .B1(_1331_),
    .A1(_0266_),
    .Y(_1335_),
    .A2(net595));
 sg13g2_nand2_1 _2658_ (.Y(_1336_),
    .A(_0004_),
    .B(net558));
 sg13g2_a21oi_1 _2659_ (.A1(_0101_),
    .A2(net563),
    .Y(_1337_),
    .B1(net555));
 sg13g2_nand2_1 _2660_ (.Y(_1338_),
    .A(_0234_),
    .B(net561));
 sg13g2_a21oi_1 _2661_ (.A1(_0133_),
    .A2(net563),
    .Y(_1339_),
    .B1(net551));
 sg13g2_a221oi_1 _2662_ (.B2(_1339_),
    .C1(net540),
    .B1(_1338_),
    .A1(_1336_),
    .Y(_1340_),
    .A2(_1337_));
 sg13g2_a21o_1 _2663_ (.A2(net542),
    .A1(_0202_),
    .B1(net497),
    .X(_1341_));
 sg13g2_o21ai_1 _2664_ (.B1(_0616_),
    .Y(_1342_),
    .A1(_1340_),
    .A2(_1341_));
 sg13g2_inv_1 _2665_ (.Y(_1343_),
    .A(_1342_));
 sg13g2_nand2_1 _2666_ (.Y(_1344_),
    .A(_1316_),
    .B(_1343_));
 sg13g2_xnor2_1 _2667_ (.Y(_1345_),
    .A(_1316_),
    .B(_1343_));
 sg13g2_nand2_1 _2668_ (.Y(_1346_),
    .A(_1335_),
    .B(_1345_));
 sg13g2_xnor2_1 _2669_ (.Y(_1347_),
    .A(_1335_),
    .B(_1345_));
 sg13g2_nand3_1 _2670_ (.B(_1325_),
    .C(_1347_),
    .A(_1319_),
    .Y(_1348_));
 sg13g2_a21o_1 _2671_ (.A2(_1325_),
    .A1(_1319_),
    .B1(_1347_),
    .X(_1349_));
 sg13g2_nand3_1 _2672_ (.B(_1348_),
    .C(_1349_),
    .A(net571),
    .Y(_1350_));
 sg13g2_nand2_1 _2673_ (.Y(_1351_),
    .A(net764),
    .B(net582));
 sg13g2_o21ai_1 _2674_ (.B1(_1351_),
    .Y(_0385_),
    .A1(net582),
    .A2(_1350_));
 sg13g2_nor2_1 _2675_ (.A(_0201_),
    .B(net521),
    .Y(_1352_));
 sg13g2_o21ai_1 _2676_ (.B1(net485),
    .Y(_1353_),
    .A1(_0067_),
    .A2(net530));
 sg13g2_a21oi_1 _2677_ (.A1(_0164_),
    .A2(net486),
    .Y(_1354_),
    .B1(net516));
 sg13g2_o21ai_1 _2678_ (.B1(_1354_),
    .Y(_1355_),
    .A1(_1352_),
    .A2(_1353_));
 sg13g2_nand2_1 _2679_ (.Y(_1356_),
    .A(_0003_),
    .B(net530));
 sg13g2_a21oi_1 _2680_ (.A1(_0035_),
    .A2(net570),
    .Y(_1357_),
    .B1(net510));
 sg13g2_a21oi_1 _2681_ (.A1(_1356_),
    .A2(_1357_),
    .Y(_1358_),
    .B1(net592));
 sg13g2_a221oi_1 _2682_ (.B2(_1358_),
    .C1(net469),
    .B1(_1355_),
    .A1(_0265_),
    .Y(_1359_),
    .A2(net592));
 sg13g2_mux4_1 _2683_ (.S0(net557),
    .A0(_0132_),
    .A1(_0233_),
    .A2(_0100_),
    .A3(_0003_),
    .S1(net550),
    .X(_1360_));
 sg13g2_nand2_1 _2684_ (.Y(_1361_),
    .A(net547),
    .B(_1360_));
 sg13g2_a21oi_1 _2685_ (.A1(_0201_),
    .A2(net540),
    .Y(_1362_),
    .B1(net495));
 sg13g2_a21oi_1 _2686_ (.A1(_1361_),
    .A2(_1362_),
    .Y(_1363_),
    .B1(net588));
 sg13g2_nand3_1 _2687_ (.B(_1343_),
    .C(_1363_),
    .A(_1316_),
    .Y(_1364_));
 sg13g2_xor2_1 _2688_ (.B(_1363_),
    .A(_1344_),
    .X(_1365_));
 sg13g2_and2_1 _2689_ (.A(_1359_),
    .B(_1365_),
    .X(_1366_));
 sg13g2_xor2_1 _2690_ (.B(_1365_),
    .A(_1359_),
    .X(_1367_));
 sg13g2_nor3_1 _2691_ (.A(_1320_),
    .B(_1322_),
    .C(_1347_),
    .Y(_1368_));
 sg13g2_or3_1 _2692_ (.A(_1320_),
    .B(_1321_),
    .C(_1347_),
    .X(_1369_));
 sg13g2_o21ai_1 _2693_ (.B1(_1318_),
    .Y(_1370_),
    .A1(_1335_),
    .A2(_1345_));
 sg13g2_nand3_1 _2694_ (.B(_1369_),
    .C(_1370_),
    .A(_1346_),
    .Y(_1371_));
 sg13g2_a21oi_1 _2695_ (.A1(_1257_),
    .A2(_1368_),
    .Y(_1372_),
    .B1(_1371_));
 sg13g2_nand2b_2 _2696_ (.Y(_1373_),
    .B(_1367_),
    .A_N(_1372_));
 sg13g2_nand2b_1 _2697_ (.Y(_1374_),
    .B(_1372_),
    .A_N(_1367_));
 sg13g2_a21oi_2 _2698_ (.B1(net573),
    .Y(_1375_),
    .A2(_1374_),
    .A1(_1373_));
 sg13g2_nand2_1 _2699_ (.Y(_1376_),
    .A(net770),
    .B(net577));
 sg13g2_o21ai_1 _2700_ (.B1(_1376_),
    .Y(_0386_),
    .A1(net578),
    .A2(_1375_));
 sg13g2_nand2b_1 _2701_ (.Y(_1377_),
    .B(_1373_),
    .A_N(_1366_));
 sg13g2_nand2b_1 _2702_ (.Y(_1378_),
    .B(net522),
    .A_N(_0066_));
 sg13g2_o21ai_1 _2703_ (.B1(_1378_),
    .Y(_1379_),
    .A1(_0200_),
    .A2(net522));
 sg13g2_a21oi_1 _2704_ (.A1(_0163_),
    .A2(net487),
    .Y(_1380_),
    .B1(net516));
 sg13g2_o21ai_1 _2705_ (.B1(_1380_),
    .Y(_1381_),
    .A1(net487),
    .A2(_1379_));
 sg13g2_nand2_1 _2706_ (.Y(_1382_),
    .A(_0002_),
    .B(net531));
 sg13g2_a21oi_1 _2707_ (.A1(_0034_),
    .A2(net522),
    .Y(_1383_),
    .B1(net510));
 sg13g2_a21oi_1 _2708_ (.A1(_1382_),
    .A2(_1383_),
    .Y(_1384_),
    .B1(net592));
 sg13g2_a22oi_1 _2709_ (.Y(_1385_),
    .B1(_1381_),
    .B2(_1384_),
    .A2(net592),
    .A1(_0264_));
 sg13g2_nand2_1 _2710_ (.Y(_1386_),
    .A(_0684_),
    .B(_1385_));
 sg13g2_nand2_1 _2711_ (.Y(_1387_),
    .A(_0002_),
    .B(net557));
 sg13g2_a21oi_1 _2712_ (.A1(_0099_),
    .A2(net563),
    .Y(_1388_),
    .B1(net555));
 sg13g2_nand2_1 _2713_ (.Y(_1389_),
    .A(_0232_),
    .B(net557));
 sg13g2_a21oi_1 _2714_ (.A1(_0131_),
    .A2(net563),
    .Y(_1390_),
    .B1(net551));
 sg13g2_a221oi_1 _2715_ (.B2(_1390_),
    .C1(net540),
    .B1(_1389_),
    .A1(_1387_),
    .Y(_1391_),
    .A2(_1388_));
 sg13g2_a21o_1 _2716_ (.A2(net540),
    .A1(_0200_),
    .B1(net495),
    .X(_1392_));
 sg13g2_o21ai_1 _2717_ (.B1(_0616_),
    .Y(_1393_),
    .A1(_1391_),
    .A2(_1392_));
 sg13g2_nor2_1 _2718_ (.A(_1364_),
    .B(_1393_),
    .Y(_1394_));
 sg13g2_xor2_1 _2719_ (.B(_1393_),
    .A(_1364_),
    .X(_1395_));
 sg13g2_and2_1 _2720_ (.A(_1386_),
    .B(_1395_),
    .X(_1396_));
 sg13g2_nor2_1 _2721_ (.A(_1386_),
    .B(_1395_),
    .Y(_1397_));
 sg13g2_nor2_1 _2722_ (.A(_1396_),
    .B(_1397_),
    .Y(_1398_));
 sg13g2_a21oi_1 _2723_ (.A1(_1377_),
    .A2(_1398_),
    .Y(_1399_),
    .B1(net573));
 sg13g2_o21ai_1 _2724_ (.B1(_1399_),
    .Y(_1400_),
    .A1(_1377_),
    .A2(_1398_));
 sg13g2_nand2_1 _2725_ (.Y(_1401_),
    .A(net763),
    .B(net578));
 sg13g2_o21ai_1 _2726_ (.B1(_1401_),
    .Y(_0387_),
    .A1(net578),
    .A2(_1400_));
 sg13g2_nor2_1 _2727_ (.A(_0199_),
    .B(net521),
    .Y(_1402_));
 sg13g2_o21ai_1 _2728_ (.B1(net485),
    .Y(_1403_),
    .A1(_0065_),
    .A2(net530));
 sg13g2_a21oi_1 _2729_ (.A1(_0162_),
    .A2(net486),
    .Y(_1404_),
    .B1(net516));
 sg13g2_o21ai_1 _2730_ (.B1(_1404_),
    .Y(_1405_),
    .A1(_1402_),
    .A2(_1403_));
 sg13g2_nand2_1 _2731_ (.Y(_1406_),
    .A(_0001_),
    .B(net531));
 sg13g2_a21oi_1 _2732_ (.A1(_0033_),
    .A2(net522),
    .Y(_1407_),
    .B1(net510));
 sg13g2_a21oi_1 _2733_ (.A1(_1406_),
    .A2(_1407_),
    .Y(_1408_),
    .B1(net591));
 sg13g2_a221oi_1 _2734_ (.B2(_1408_),
    .C1(net469),
    .B1(_1405_),
    .A1(_0263_),
    .Y(_1409_),
    .A2(net591));
 sg13g2_mux2_1 _2735_ (.A0(_0130_),
    .A1(_0193_),
    .S(_0627_),
    .X(_1410_));
 sg13g2_mux4_1 _2736_ (.S0(net551),
    .A0(_0231_),
    .A1(_0001_),
    .A2(_1410_),
    .A3(_0098_),
    .S1(net563),
    .X(_1411_));
 sg13g2_nand2_1 _2737_ (.Y(_1412_),
    .A(_0199_),
    .B(net540));
 sg13g2_a21oi_1 _2738_ (.A1(net547),
    .A2(_1411_),
    .Y(_1413_),
    .B1(net495));
 sg13g2_a21oi_1 _2739_ (.A1(_1412_),
    .A2(_1413_),
    .Y(_1414_),
    .B1(net588));
 sg13g2_nand2_1 _2740_ (.Y(_1415_),
    .A(_1394_),
    .B(_1414_));
 sg13g2_xnor2_1 _2741_ (.Y(_1416_),
    .A(_1394_),
    .B(_1414_));
 sg13g2_and2_1 _2742_ (.A(_1409_),
    .B(_1416_),
    .X(_1417_));
 sg13g2_xnor2_1 _2743_ (.Y(_1418_),
    .A(_1409_),
    .B(_1416_));
 sg13g2_inv_1 _2744_ (.Y(_1419_),
    .A(_1418_));
 sg13g2_nor2_1 _2745_ (.A(_1366_),
    .B(_1397_),
    .Y(_1420_));
 sg13g2_a21oi_1 _2746_ (.A1(_1373_),
    .A2(_1420_),
    .Y(_1421_),
    .B1(_1396_));
 sg13g2_a221oi_1 _2747_ (.B2(_1373_),
    .C1(_1418_),
    .B1(_1420_),
    .A1(_1386_),
    .Y(_1422_),
    .A2(_1395_));
 sg13g2_nor2_1 _2748_ (.A(net573),
    .B(_1422_),
    .Y(_1423_));
 sg13g2_o21ai_1 _2749_ (.B1(_1423_),
    .Y(_1424_),
    .A1(_1419_),
    .A2(_1421_));
 sg13g2_nand2_1 _2750_ (.Y(_1425_),
    .A(net771),
    .B(net578));
 sg13g2_o21ai_1 _2751_ (.B1(_1425_),
    .Y(_0388_),
    .A1(net577),
    .A2(_1424_));
 sg13g2_and2_1 _2752_ (.A(_0064_),
    .B(net521),
    .X(_1426_));
 sg13g2_a21oi_1 _2753_ (.A1(_0198_),
    .A2(net530),
    .Y(_1427_),
    .B1(_1426_));
 sg13g2_nand2_1 _2754_ (.Y(_1428_),
    .A(_0032_),
    .B(net570));
 sg13g2_a21oi_1 _2755_ (.A1(_0161_),
    .A2(net486),
    .Y(_1429_),
    .B1(net516));
 sg13g2_o21ai_1 _2756_ (.B1(_1429_),
    .Y(_1430_),
    .A1(net486),
    .A2(_1427_));
 sg13g2_a21oi_1 _2757_ (.A1(_0000_),
    .A2(net530),
    .Y(_1431_),
    .B1(net510));
 sg13g2_a21oi_1 _2758_ (.A1(_1428_),
    .A2(_1431_),
    .Y(_1432_),
    .B1(net591));
 sg13g2_a221oi_1 _2759_ (.B2(_1432_),
    .C1(net469),
    .B1(_1430_),
    .A1(_0262_),
    .Y(_1433_),
    .A2(net591));
 sg13g2_mux4_1 _2760_ (.S0(net557),
    .A0(_0129_),
    .A1(_0230_),
    .A2(_0097_),
    .A3(_0000_),
    .S1(net550),
    .X(_1434_));
 sg13g2_nand2_1 _2761_ (.Y(_1435_),
    .A(net547),
    .B(_1434_));
 sg13g2_a21oi_1 _2762_ (.A1(_0198_),
    .A2(net540),
    .Y(_1436_),
    .B1(net495));
 sg13g2_a21oi_1 _2763_ (.A1(_1435_),
    .A2(_1436_),
    .Y(_1437_),
    .B1(net588));
 sg13g2_xnor2_1 _2764_ (.Y(_1438_),
    .A(_1433_),
    .B(_1437_));
 sg13g2_xnor2_1 _2765_ (.Y(_1439_),
    .A(_1415_),
    .B(_1438_));
 sg13g2_or3_1 _2766_ (.A(_1417_),
    .B(_1422_),
    .C(_1439_),
    .X(_1440_));
 sg13g2_o21ai_1 _2767_ (.B1(_1439_),
    .Y(_1441_),
    .A1(_1417_),
    .A2(_1422_));
 sg13g2_nand3_1 _2768_ (.B(_1440_),
    .C(_1441_),
    .A(net571),
    .Y(_1442_));
 sg13g2_nand2_1 _2769_ (.Y(_1443_),
    .A(net766),
    .B(net577));
 sg13g2_o21ai_1 _2770_ (.B1(_1443_),
    .Y(_0389_),
    .A1(net577),
    .A2(_1442_));
 sg13g2_and4_1 _2771_ (.A(net585),
    .B(_0667_),
    .C(_0670_),
    .D(_0682_),
    .X(_1444_));
 sg13g2_or2_1 _2772_ (.X(_1445_),
    .B(_0617_),
    .A(_0614_));
 sg13g2_or2_1 _2773_ (.X(_1446_),
    .B(_1445_),
    .A(net603));
 sg13g2_nand2_1 _2774_ (.Y(_1447_),
    .A(_0638_),
    .B(_1446_));
 sg13g2_nand2_2 _2775_ (.Y(_1448_),
    .A(_1444_),
    .B(_1447_));
 sg13g2_nand2_1 _2776_ (.Y(_1449_),
    .A(net674),
    .B(net466));
 sg13g2_o21ai_1 _2777_ (.B1(_1449_),
    .Y(_0459_),
    .A1(_0688_),
    .A2(net466));
 sg13g2_nand2_1 _2778_ (.Y(_1450_),
    .A(net709),
    .B(net467));
 sg13g2_o21ai_1 _2779_ (.B1(_1450_),
    .Y(_0460_),
    .A1(_0708_),
    .A2(net467));
 sg13g2_nand2_1 _2780_ (.Y(_1451_),
    .A(net690),
    .B(net466));
 sg13g2_o21ai_1 _2781_ (.B1(_1451_),
    .Y(_0461_),
    .A1(_0730_),
    .A2(net466));
 sg13g2_nand2_1 _2782_ (.Y(_1452_),
    .A(net742),
    .B(net466));
 sg13g2_o21ai_1 _2783_ (.B1(_1452_),
    .Y(_0462_),
    .A1(_0753_),
    .A2(net466));
 sg13g2_nand2_1 _2784_ (.Y(_1453_),
    .A(net726),
    .B(net466));
 sg13g2_o21ai_1 _2785_ (.B1(_1453_),
    .Y(_0463_),
    .A1(_0779_),
    .A2(net466));
 sg13g2_nand2_1 _2786_ (.Y(_1454_),
    .A(net696),
    .B(net465));
 sg13g2_o21ai_1 _2787_ (.B1(_1454_),
    .Y(_0464_),
    .A1(_0803_),
    .A2(net465));
 sg13g2_nand2_1 _2788_ (.Y(_1455_),
    .A(net658),
    .B(net465));
 sg13g2_o21ai_1 _2789_ (.B1(_1455_),
    .Y(_0465_),
    .A1(_0828_),
    .A2(net465));
 sg13g2_nand2_1 _2790_ (.Y(_1456_),
    .A(net652),
    .B(net465));
 sg13g2_o21ai_1 _2791_ (.B1(_1456_),
    .Y(_0466_),
    .A1(_0849_),
    .A2(net465));
 sg13g2_nand2_1 _2792_ (.Y(_1457_),
    .A(net719),
    .B(net461));
 sg13g2_o21ai_1 _2793_ (.B1(_1457_),
    .Y(_0467_),
    .A1(_0872_),
    .A2(net461));
 sg13g2_nand2_1 _2794_ (.Y(_1458_),
    .A(net749),
    .B(net461));
 sg13g2_o21ai_1 _2795_ (.B1(_1458_),
    .Y(_0468_),
    .A1(_0898_),
    .A2(net461));
 sg13g2_nand2_1 _2796_ (.Y(_1459_),
    .A(net692),
    .B(net460));
 sg13g2_o21ai_1 _2797_ (.B1(_1459_),
    .Y(_0469_),
    .A1(_0925_),
    .A2(net460));
 sg13g2_nand2_1 _2798_ (.Y(_1460_),
    .A(net740),
    .B(net460));
 sg13g2_o21ai_1 _2799_ (.B1(_1460_),
    .Y(_0470_),
    .A1(_0945_),
    .A2(net460));
 sg13g2_nand2_1 _2800_ (.Y(_1461_),
    .A(net734),
    .B(net462));
 sg13g2_o21ai_1 _2801_ (.B1(_1461_),
    .Y(_0471_),
    .A1(_0974_),
    .A2(net462));
 sg13g2_nand2_1 _2802_ (.Y(_1462_),
    .A(net684),
    .B(net459));
 sg13g2_o21ai_1 _2803_ (.B1(_1462_),
    .Y(_0472_),
    .A1(_0995_),
    .A2(net459));
 sg13g2_nand2_1 _2804_ (.Y(_1463_),
    .A(net649),
    .B(net462));
 sg13g2_o21ai_1 _2805_ (.B1(_1463_),
    .Y(_0473_),
    .A1(_1023_),
    .A2(net461));
 sg13g2_nand2_1 _2806_ (.Y(_1464_),
    .A(net682),
    .B(net459));
 sg13g2_o21ai_1 _2807_ (.B1(_1464_),
    .Y(_0474_),
    .A1(_1043_),
    .A2(net459));
 sg13g2_nand2_1 _2808_ (.Y(_1465_),
    .A(net675),
    .B(net468));
 sg13g2_o21ai_1 _2809_ (.B1(_1465_),
    .Y(_0475_),
    .A1(_1074_),
    .A2(net468));
 sg13g2_nand2_1 _2810_ (.Y(_1466_),
    .A(net729),
    .B(net468));
 sg13g2_o21ai_1 _2811_ (.B1(_1466_),
    .Y(_0476_),
    .A1(_1100_),
    .A2(net467));
 sg13g2_nand2_1 _2812_ (.Y(_1467_),
    .A(net715),
    .B(net467));
 sg13g2_o21ai_1 _2813_ (.B1(_1467_),
    .Y(_0477_),
    .A1(_1122_),
    .A2(net467));
 sg13g2_nand2_1 _2814_ (.Y(_1468_),
    .A(net728),
    .B(net467));
 sg13g2_o21ai_1 _2815_ (.B1(_1468_),
    .Y(_0478_),
    .A1(_1146_),
    .A2(net467));
 sg13g2_nand2_1 _2816_ (.Y(_1469_),
    .A(net659),
    .B(net464));
 sg13g2_o21ai_1 _2817_ (.B1(_1469_),
    .Y(_0479_),
    .A1(_1173_),
    .A2(net464));
 sg13g2_nand2_1 _2818_ (.Y(_1470_),
    .A(net723),
    .B(net465));
 sg13g2_o21ai_1 _2819_ (.B1(_1470_),
    .Y(_0480_),
    .A1(_1199_),
    .A2(net468));
 sg13g2_nand2_1 _2820_ (.Y(_1471_),
    .A(net660),
    .B(net464));
 sg13g2_o21ai_1 _2821_ (.B1(_1471_),
    .Y(_0481_),
    .A1(_1224_),
    .A2(net464));
 sg13g2_nand2_1 _2822_ (.Y(_1472_),
    .A(net712),
    .B(net464));
 sg13g2_o21ai_1 _2823_ (.B1(_1472_),
    .Y(_0482_),
    .A1(_1248_),
    .A2(net464));
 sg13g2_nand2_1 _2824_ (.Y(_1473_),
    .A(net699),
    .B(net459));
 sg13g2_o21ai_1 _2825_ (.B1(_1473_),
    .Y(_0483_),
    .A1(_1276_),
    .A2(net459));
 sg13g2_nand2_1 _2826_ (.Y(_1474_),
    .A(net718),
    .B(net463));
 sg13g2_o21ai_1 _2827_ (.B1(_1474_),
    .Y(_0484_),
    .A1(_1301_),
    .A2(net463));
 sg13g2_nand2_1 _2828_ (.Y(_1475_),
    .A(net702),
    .B(net459));
 sg13g2_o21ai_1 _2829_ (.B1(_1475_),
    .Y(_0485_),
    .A1(_1326_),
    .A2(net459));
 sg13g2_nand2_1 _2830_ (.Y(_1476_),
    .A(net685),
    .B(net464));
 sg13g2_o21ai_1 _2831_ (.B1(_1476_),
    .Y(_0486_),
    .A1(_1350_),
    .A2(net464));
 sg13g2_nand2_1 _2832_ (.Y(_1477_),
    .A(net731),
    .B(net460));
 sg13g2_o21ai_1 _2833_ (.B1(_1477_),
    .Y(_0487_),
    .A1(_1375_),
    .A2(net460));
 sg13g2_nand2_1 _2834_ (.Y(_1478_),
    .A(net666),
    .B(net462));
 sg13g2_o21ai_1 _2835_ (.B1(_1478_),
    .Y(_0488_),
    .A1(_1400_),
    .A2(net461));
 sg13g2_nand2_1 _2836_ (.Y(_1479_),
    .A(net706),
    .B(net461));
 sg13g2_o21ai_1 _2837_ (.B1(_1479_),
    .Y(_0489_),
    .A1(_1424_),
    .A2(net461));
 sg13g2_nand2_1 _2838_ (.Y(_1480_),
    .A(net683),
    .B(net460));
 sg13g2_o21ai_1 _2839_ (.B1(_1480_),
    .Y(_0490_),
    .A1(_1442_),
    .A2(net460));
 sg13g2_and2_1 _2840_ (.A(net322),
    .B(net1),
    .X(_0491_));
 sg13g2_o21ai_1 _2841_ (.B1(net611),
    .Y(_1481_),
    .A1(net743),
    .A2(\i_soc.cnt[1] ));
 sg13g2_a21oi_1 _2842_ (.A1(net743),
    .A2(\i_soc.cnt[1] ),
    .Y(_0492_),
    .B1(_1481_));
 sg13g2_a21oi_1 _2843_ (.A1(net743),
    .A2(\i_soc.cnt[1] ),
    .Y(_1482_),
    .B1(net747));
 sg13g2_nand3_1 _2844_ (.B(net747),
    .C(\i_soc.cnt[1] ),
    .A(net743),
    .Y(_1483_));
 sg13g2_nand2_1 _2845_ (.Y(_1484_),
    .A(net611),
    .B(_1483_));
 sg13g2_nor2_1 _2846_ (.A(net748),
    .B(_1484_),
    .Y(_0493_));
 sg13g2_and2_1 _2847_ (.A(_0603_),
    .B(_1483_),
    .X(_1485_));
 sg13g2_nor2_1 _2848_ (.A(_0603_),
    .B(_1483_),
    .Y(_1486_));
 sg13g2_nor3_1 _2849_ (.A(_0612_),
    .B(net787),
    .C(_1486_),
    .Y(_0494_));
 sg13g2_and2_1 _2850_ (.A(net779),
    .B(_1486_),
    .X(_1487_));
 sg13g2_o21ai_1 _2851_ (.B1(net611),
    .Y(_1488_),
    .A1(net779),
    .A2(_1486_));
 sg13g2_nor2_1 _2852_ (.A(_1487_),
    .B(net780),
    .Y(_0495_));
 sg13g2_xnor2_1 _2853_ (.Y(_1489_),
    .A(net781),
    .B(_1487_));
 sg13g2_nor2_1 _2854_ (.A(_0612_),
    .B(_1489_),
    .Y(_0496_));
 sg13g2_a21oi_1 _2855_ (.A1(\i_soc.cnt[5] ),
    .A2(_1487_),
    .Y(_1490_),
    .B1(net757));
 sg13g2_nand3_1 _2856_ (.B(net781),
    .C(_1487_),
    .A(net757),
    .Y(_1491_));
 sg13g2_nand2_1 _2857_ (.Y(_1492_),
    .A(net611),
    .B(_1491_));
 sg13g2_nor2_1 _2858_ (.A(net758),
    .B(_1492_),
    .Y(_0497_));
 sg13g2_xnor2_1 _2859_ (.Y(_1493_),
    .A(_0602_),
    .B(_1491_));
 sg13g2_nor2_1 _2860_ (.A(_0612_),
    .B(_1493_),
    .Y(_0498_));
 sg13g2_and2_1 _2861_ (.A(net323),
    .B(net611),
    .X(_0499_));
 sg13g2_and2_1 _2862_ (.A(net611),
    .B(_1445_),
    .X(_0500_));
 sg13g2_nand3_1 _2863_ (.B(net790),
    .C(net607),
    .A(net610),
    .Y(_1494_));
 sg13g2_nor3_1 _2864_ (.A(_0612_),
    .B(_0618_),
    .C(_0646_),
    .Y(_1495_));
 sg13g2_and2_1 _2865_ (.A(_1494_),
    .B(_1495_),
    .X(_0501_));
 sg13g2_xor2_1 _2866_ (.B(_1494_),
    .A(net604),
    .X(_1496_));
 sg13g2_nor2_1 _2867_ (.A(_0612_),
    .B(net789),
    .Y(_0502_));
 sg13g2_a21oi_1 _2868_ (.A1(net608),
    .A2(net574),
    .Y(_1497_),
    .B1(net569));
 sg13g2_nand2_1 _2869_ (.Y(_1498_),
    .A(net648),
    .B(net507));
 sg13g2_o21ai_1 _2870_ (.B1(_1498_),
    .Y(_0534_),
    .A1(_0688_),
    .A2(net507));
 sg13g2_nand2_1 _2871_ (.Y(_1499_),
    .A(net755),
    .B(net508));
 sg13g2_o21ai_1 _2872_ (.B1(_1499_),
    .Y(_0535_),
    .A1(_0708_),
    .A2(net508));
 sg13g2_nand2_1 _2873_ (.Y(_1500_),
    .A(net700),
    .B(net507));
 sg13g2_o21ai_1 _2874_ (.B1(_1500_),
    .Y(_0536_),
    .A1(_0730_),
    .A2(net507));
 sg13g2_nand2_1 _2875_ (.Y(_1501_),
    .A(net687),
    .B(net507));
 sg13g2_o21ai_1 _2876_ (.B1(_1501_),
    .Y(_0537_),
    .A1(_0753_),
    .A2(net507));
 sg13g2_nand2_1 _2877_ (.Y(_1502_),
    .A(net695),
    .B(net507));
 sg13g2_o21ai_1 _2878_ (.B1(_1502_),
    .Y(_0538_),
    .A1(_0779_),
    .A2(net507));
 sg13g2_nand2_1 _2879_ (.Y(_1503_),
    .A(net697),
    .B(net505));
 sg13g2_o21ai_1 _2880_ (.B1(_1503_),
    .Y(_0539_),
    .A1(_0803_),
    .A2(net505));
 sg13g2_nand2_1 _2881_ (.Y(_1504_),
    .A(net711),
    .B(net505));
 sg13g2_o21ai_1 _2882_ (.B1(_1504_),
    .Y(_0540_),
    .A1(_0828_),
    .A2(net505));
 sg13g2_nand2_1 _2883_ (.Y(_1505_),
    .A(net701),
    .B(net505));
 sg13g2_o21ai_1 _2884_ (.B1(_1505_),
    .Y(_0541_),
    .A1(_0849_),
    .A2(net505));
 sg13g2_nand2_1 _2885_ (.Y(_1506_),
    .A(net681),
    .B(net502));
 sg13g2_o21ai_1 _2886_ (.B1(_1506_),
    .Y(_0542_),
    .A1(_0872_),
    .A2(net502));
 sg13g2_nand2_1 _2887_ (.Y(_1507_),
    .A(net707),
    .B(net502));
 sg13g2_o21ai_1 _2888_ (.B1(_1507_),
    .Y(_0543_),
    .A1(_0898_),
    .A2(net502));
 sg13g2_nand2_1 _2889_ (.Y(_1508_),
    .A(net720),
    .B(net501));
 sg13g2_o21ai_1 _2890_ (.B1(_1508_),
    .Y(_0544_),
    .A1(_0925_),
    .A2(net501));
 sg13g2_nand2_1 _2891_ (.Y(_1509_),
    .A(net686),
    .B(net501));
 sg13g2_o21ai_1 _2892_ (.B1(_1509_),
    .Y(_0545_),
    .A1(_0945_),
    .A2(net501));
 sg13g2_nand2_1 _2893_ (.Y(_1510_),
    .A(net691),
    .B(net504));
 sg13g2_o21ai_1 _2894_ (.B1(_1510_),
    .Y(_0546_),
    .A1(_0974_),
    .A2(net504));
 sg13g2_nand2_1 _2895_ (.Y(_1511_),
    .A(net651),
    .B(net500));
 sg13g2_o21ai_1 _2896_ (.B1(_1511_),
    .Y(_0547_),
    .A1(_0995_),
    .A2(net500));
 sg13g2_nand2_1 _2897_ (.Y(_1512_),
    .A(net705),
    .B(net503));
 sg13g2_o21ai_1 _2898_ (.B1(_1512_),
    .Y(_0548_),
    .A1(_1023_),
    .A2(net503));
 sg13g2_nand2_1 _2899_ (.Y(_1513_),
    .A(net730),
    .B(net500));
 sg13g2_o21ai_1 _2900_ (.B1(_1513_),
    .Y(_0549_),
    .A1(_1043_),
    .A2(net500));
 sg13g2_nand2_1 _2901_ (.Y(_1514_),
    .A(net656),
    .B(net509));
 sg13g2_o21ai_1 _2902_ (.B1(_1514_),
    .Y(_0550_),
    .A1(_1074_),
    .A2(net509));
 sg13g2_nand2_1 _2903_ (.Y(_1515_),
    .A(net725),
    .B(net508));
 sg13g2_o21ai_1 _2904_ (.B1(_1515_),
    .Y(_0551_),
    .A1(_1100_),
    .A2(net508));
 sg13g2_nand2_1 _2905_ (.Y(_1516_),
    .A(net673),
    .B(net508));
 sg13g2_o21ai_1 _2906_ (.B1(_1516_),
    .Y(_0552_),
    .A1(_1122_),
    .A2(net508));
 sg13g2_nand2_1 _2907_ (.Y(_1517_),
    .A(net657),
    .B(net508));
 sg13g2_o21ai_1 _2908_ (.B1(_1517_),
    .Y(_0553_),
    .A1(_1146_),
    .A2(net509));
 sg13g2_nand2_1 _2909_ (.Y(_1518_),
    .A(net676),
    .B(net506));
 sg13g2_o21ai_1 _2910_ (.B1(_1518_),
    .Y(_0554_),
    .A1(_1173_),
    .A2(net506));
 sg13g2_a22oi_1 _2911_ (.Y(_0555_),
    .B1(net506),
    .B2(_0611_),
    .A2(_0666_),
    .A1(net328));
 sg13g2_nand2_1 _2912_ (.Y(_1519_),
    .A(net721),
    .B(net506));
 sg13g2_o21ai_1 _2913_ (.B1(_1519_),
    .Y(_0556_),
    .A1(_1224_),
    .A2(net506));
 sg13g2_nand2_1 _2914_ (.Y(_1520_),
    .A(net727),
    .B(net505));
 sg13g2_o21ai_1 _2915_ (.B1(_1520_),
    .Y(_0557_),
    .A1(_1248_),
    .A2(net505));
 sg13g2_nand2_1 _2916_ (.Y(_1521_),
    .A(net668),
    .B(net500));
 sg13g2_o21ai_1 _2917_ (.B1(_1521_),
    .Y(_0558_),
    .A1(_1276_),
    .A2(net500));
 sg13g2_a22oi_1 _2918_ (.Y(_0559_),
    .B1(net504),
    .B2(_0600_),
    .A2(net570),
    .A1(net381));
 sg13g2_nand2_1 _2919_ (.Y(_1522_),
    .A(net703),
    .B(net500));
 sg13g2_o21ai_1 _2920_ (.B1(_1522_),
    .Y(_0560_),
    .A1(_1326_),
    .A2(net500));
 sg13g2_nand2_1 _2921_ (.Y(_1523_),
    .A(net736),
    .B(net503));
 sg13g2_o21ai_1 _2922_ (.B1(_1523_),
    .Y(_0561_),
    .A1(_1350_),
    .A2(net503));
 sg13g2_a22oi_1 _2923_ (.Y(_0562_),
    .B1(net501),
    .B2(_0601_),
    .A2(net570),
    .A1(net339));
 sg13g2_nand2_1 _2924_ (.Y(_1524_),
    .A(net741),
    .B(net502));
 sg13g2_o21ai_1 _2925_ (.B1(_1524_),
    .Y(_0563_),
    .A1(_1400_),
    .A2(net502));
 sg13g2_nand2_1 _2926_ (.Y(_1525_),
    .A(net688),
    .B(net502));
 sg13g2_o21ai_1 _2927_ (.B1(_1525_),
    .Y(_0564_),
    .A1(_1424_),
    .A2(net502));
 sg13g2_nand2_1 _2928_ (.Y(_1526_),
    .A(net713),
    .B(net501));
 sg13g2_o21ai_1 _2929_ (.B1(_1526_),
    .Y(_0565_),
    .A1(_1442_),
    .A2(net501));
 sg13g2_nand2_1 _2930_ (.Y(_1527_),
    .A(\i_soc.cpu.rd0[13] ),
    .B(\i_soc.cpu.rd0[12] ));
 sg13g2_nand4_1 _2931_ (.B(\i_soc.cpu.rd0[8] ),
    .C(\i_soc.cpu.rd0[11] ),
    .A(_0604_),
    .Y(_1528_),
    .D(\i_soc.cpu.rd0[10] ));
 sg13g2_nor4_1 _2932_ (.A(\i_soc.cpu.rd0[15] ),
    .B(\i_soc.cpu.rd0[14] ),
    .C(_1527_),
    .D(_1528_),
    .Y(_1529_));
 sg13g2_nor4_2 _2933_ (.A(\i_soc.cpu.rd0[20] ),
    .B(_0605_),
    .C(\i_soc.cpu.rd0[23] ),
    .Y(_1530_),
    .D(\i_soc.cpu.rd0[22] ));
 sg13g2_nor4_2 _2934_ (.A(\i_soc.cpu.rd0[28] ),
    .B(\i_soc.cpu.rd0[29] ),
    .C(\i_soc.cpu.rd0[30] ),
    .Y(_1531_),
    .D(\i_soc.cpu.rd0[31] ));
 sg13g2_nor3_1 _2935_ (.A(\i_soc.cpu.rd0[24] ),
    .B(\i_soc.cpu.rd0[25] ),
    .C(\i_soc.cpu.rd0[26] ),
    .Y(_1532_));
 sg13g2_nor4_1 _2936_ (.A(\i_soc.cpu.rd0[5] ),
    .B(\i_soc.cpu.rd0[4] ),
    .C(\i_soc.cpu.rd0[7] ),
    .D(\i_soc.cpu.rd0[6] ),
    .Y(_1533_));
 sg13g2_nand3b_1 _2937_ (.B(_1530_),
    .C(net738),
    .Y(_1534_),
    .A_N(net724));
 sg13g2_nor3_1 _2938_ (.A(net739),
    .B(net746),
    .C(_1534_),
    .Y(_1535_));
 sg13g2_nand3_1 _2939_ (.B(\i_soc.cpu.rd0[2] ),
    .C(_1533_),
    .A(\i_soc.cpu.rd0[0] ),
    .Y(_1536_));
 sg13g2_nor2_2 _2940_ (.A(\i_soc.cpu.rd0[1] ),
    .B(\i_soc.cpu.rd0[3] ),
    .Y(_1537_));
 sg13g2_nand4_1 _2941_ (.B(_1531_),
    .C(_1532_),
    .A(_1529_),
    .Y(_1538_),
    .D(_1537_));
 sg13g2_nor3_2 _2942_ (.A(net764),
    .B(_1536_),
    .C(_1538_),
    .Y(_1539_));
 sg13g2_a21oi_1 _2943_ (.A1(_1535_),
    .A2(_1539_),
    .Y(_1540_),
    .B1(net776));
 sg13g2_nor2_1 _2944_ (.A(_0612_),
    .B(_1540_),
    .Y(_0566_));
 sg13g2_nor3_1 _2945_ (.A(net776),
    .B(_0602_),
    .C(_1491_),
    .Y(_1541_));
 sg13g2_o21ai_1 _2946_ (.B1(net611),
    .Y(_1542_),
    .A1(net783),
    .A2(_1541_));
 sg13g2_inv_1 _2947_ (.Y(_0567_),
    .A(net784));
 sg13g2_a21oi_1 _2948_ (.A1(net602),
    .A2(_0626_),
    .Y(_1543_),
    .B1(net589));
 sg13g2_nand3_1 _2949_ (.B(_1446_),
    .C(_1543_),
    .A(net585),
    .Y(_1544_));
 sg13g2_nand2_1 _2950_ (.Y(_1545_),
    .A(net654),
    .B(net481));
 sg13g2_o21ai_1 _2951_ (.B1(_1545_),
    .Y(_0568_),
    .A1(_0688_),
    .A2(net481));
 sg13g2_nand2_1 _2952_ (.Y(_1546_),
    .A(net677),
    .B(net482));
 sg13g2_o21ai_1 _2953_ (.B1(_1546_),
    .Y(_0569_),
    .A1(_0708_),
    .A2(net482));
 sg13g2_nand2_1 _2954_ (.Y(_1547_),
    .A(net665),
    .B(net481));
 sg13g2_o21ai_1 _2955_ (.B1(_1547_),
    .Y(_0570_),
    .A1(_0730_),
    .A2(net481));
 sg13g2_nand2_1 _2956_ (.Y(_1548_),
    .A(net680),
    .B(net481));
 sg13g2_o21ai_1 _2957_ (.B1(_1548_),
    .Y(_0571_),
    .A1(_0753_),
    .A2(net481));
 sg13g2_nand2_1 _2958_ (.Y(_1549_),
    .A(net655),
    .B(net481));
 sg13g2_o21ai_1 _2959_ (.B1(_1549_),
    .Y(_0572_),
    .A1(_0779_),
    .A2(net481));
 sg13g2_nand2_1 _2960_ (.Y(_1550_),
    .A(net708),
    .B(net479));
 sg13g2_o21ai_1 _2961_ (.B1(_1550_),
    .Y(_0573_),
    .A1(_0803_),
    .A2(net479));
 sg13g2_nand2_1 _2962_ (.Y(_1551_),
    .A(net704),
    .B(net479));
 sg13g2_o21ai_1 _2963_ (.B1(_1551_),
    .Y(_0574_),
    .A1(_0828_),
    .A2(net479));
 sg13g2_nand2_1 _2964_ (.Y(_1552_),
    .A(net671),
    .B(net479));
 sg13g2_o21ai_1 _2965_ (.B1(_1552_),
    .Y(_0575_),
    .A1(_0849_),
    .A2(net479));
 sg13g2_nand2_1 _2966_ (.Y(_1553_),
    .A(net710),
    .B(net476));
 sg13g2_o21ai_1 _2967_ (.B1(_1553_),
    .Y(_0576_),
    .A1(_0872_),
    .A2(net476));
 sg13g2_nand2_1 _2968_ (.Y(_1554_),
    .A(net737),
    .B(net476));
 sg13g2_o21ai_1 _2969_ (.B1(_1554_),
    .Y(_0577_),
    .A1(_0898_),
    .A2(net476));
 sg13g2_nand2_1 _2970_ (.Y(_1555_),
    .A(net689),
    .B(net475));
 sg13g2_o21ai_1 _2971_ (.B1(_1555_),
    .Y(_0578_),
    .A1(_0925_),
    .A2(net475));
 sg13g2_nand2_1 _2972_ (.Y(_1556_),
    .A(net653),
    .B(net475));
 sg13g2_o21ai_1 _2973_ (.B1(_1556_),
    .Y(_0579_),
    .A1(_0945_),
    .A2(net475));
 sg13g2_nand2_1 _2974_ (.Y(_1557_),
    .A(net716),
    .B(net477));
 sg13g2_o21ai_1 _2975_ (.B1(_1557_),
    .Y(_0580_),
    .A1(_0974_),
    .A2(net477));
 sg13g2_nand2_1 _2976_ (.Y(_1558_),
    .A(net670),
    .B(net474));
 sg13g2_o21ai_1 _2977_ (.B1(_1558_),
    .Y(_0581_),
    .A1(_0995_),
    .A2(net474));
 sg13g2_nand2_1 _2978_ (.Y(_1559_),
    .A(net714),
    .B(net477));
 sg13g2_o21ai_1 _2979_ (.B1(_1559_),
    .Y(_0582_),
    .A1(_1023_),
    .A2(net477));
 sg13g2_nand2_1 _2980_ (.Y(_1560_),
    .A(net647),
    .B(net474));
 sg13g2_o21ai_1 _2981_ (.B1(_1560_),
    .Y(_0583_),
    .A1(_1043_),
    .A2(net474));
 sg13g2_nand2_1 _2982_ (.Y(_1561_),
    .A(net664),
    .B(net483));
 sg13g2_o21ai_1 _2983_ (.B1(_1561_),
    .Y(_0584_),
    .A1(_1074_),
    .A2(net483));
 sg13g2_nand2_1 _2984_ (.Y(_1562_),
    .A(net698),
    .B(net482));
 sg13g2_o21ai_1 _2985_ (.B1(_1562_),
    .Y(_0585_),
    .A1(_1100_),
    .A2(net482));
 sg13g2_nand2_1 _2986_ (.Y(_1563_),
    .A(net693),
    .B(net483));
 sg13g2_o21ai_1 _2987_ (.B1(_1563_),
    .Y(_0586_),
    .A1(_1122_),
    .A2(net482));
 sg13g2_nand2_1 _2988_ (.Y(_1564_),
    .A(net650),
    .B(net482));
 sg13g2_o21ai_1 _2989_ (.B1(_1564_),
    .Y(_0587_),
    .A1(_1146_),
    .A2(net482));
 sg13g2_nand2_1 _2990_ (.Y(_1565_),
    .A(net661),
    .B(net480));
 sg13g2_o21ai_1 _2991_ (.B1(_1565_),
    .Y(_0588_),
    .A1(_1173_),
    .A2(net480));
 sg13g2_nand2_1 _2992_ (.Y(_1566_),
    .A(net669),
    .B(net480));
 sg13g2_o21ai_1 _2993_ (.B1(_1566_),
    .Y(_0589_),
    .A1(_1199_),
    .A2(net480));
 sg13g2_nand2_1 _2994_ (.Y(_1567_),
    .A(net678),
    .B(net480));
 sg13g2_o21ai_1 _2995_ (.B1(_1567_),
    .Y(_0590_),
    .A1(_1224_),
    .A2(net480));
 sg13g2_nand2_1 _2996_ (.Y(_1568_),
    .A(net667),
    .B(net479));
 sg13g2_o21ai_1 _2997_ (.B1(_1568_),
    .Y(_0591_),
    .A1(_1248_),
    .A2(net479));
 sg13g2_nand2_1 _2998_ (.Y(_1569_),
    .A(net722),
    .B(net474));
 sg13g2_o21ai_1 _2999_ (.B1(_1569_),
    .Y(_0592_),
    .A1(_1276_),
    .A2(net474));
 sg13g2_nand2_1 _3000_ (.Y(_1570_),
    .A(net717),
    .B(net478));
 sg13g2_o21ai_1 _3001_ (.B1(_1570_),
    .Y(_0593_),
    .A1(_1301_),
    .A2(net478));
 sg13g2_nand2_1 _3002_ (.Y(_1571_),
    .A(net672),
    .B(net474));
 sg13g2_o21ai_1 _3003_ (.B1(_1571_),
    .Y(_0594_),
    .A1(_1326_),
    .A2(net474));
 sg13g2_nand2_1 _3004_ (.Y(_1572_),
    .A(net694),
    .B(net477));
 sg13g2_o21ai_1 _3005_ (.B1(_1572_),
    .Y(_0595_),
    .A1(_1350_),
    .A2(net477));
 sg13g2_nand2_1 _3006_ (.Y(_1573_),
    .A(net679),
    .B(net475));
 sg13g2_o21ai_1 _3007_ (.B1(_1573_),
    .Y(_0596_),
    .A1(_1375_),
    .A2(net475));
 sg13g2_nand2_1 _3008_ (.Y(_1574_),
    .A(net662),
    .B(net476));
 sg13g2_o21ai_1 _3009_ (.B1(_1574_),
    .Y(_0597_),
    .A1(_1400_),
    .A2(net476));
 sg13g2_nand2_1 _3010_ (.Y(_1575_),
    .A(net732),
    .B(net476));
 sg13g2_o21ai_1 _3011_ (.B1(_1575_),
    .Y(_0598_),
    .A1(_1424_),
    .A2(net476));
 sg13g2_nand2_1 _3012_ (.Y(_1576_),
    .A(net663),
    .B(net475));
 sg13g2_o21ai_1 _3013_ (.B1(_1576_),
    .Y(_0599_),
    .A1(_1442_),
    .A2(net475));
 sg13g2_buf_1 _3014_ (.A(net391),
    .X(_0294_));
 sg13g2_buf_1 _3015_ (.A(net352),
    .X(_0295_));
 sg13g2_buf_1 _3016_ (.A(net351),
    .X(_0296_));
 sg13g2_buf_1 _3017_ (.A(net350),
    .X(_0297_));
 sg13g2_buf_1 _3018_ (.A(net386),
    .X(_0298_));
 sg13g2_buf_1 _3019_ (.A(net620),
    .X(_0299_));
 sg13g2_buf_1 _3020_ (.A(net385),
    .X(_0300_));
 sg13g2_buf_1 _3021_ (.A(net358),
    .X(_0301_));
 sg13g2_buf_1 _3022_ (.A(net331),
    .X(_0302_));
 sg13g2_buf_1 _3023_ (.A(net400),
    .X(_0303_));
 sg13g2_buf_1 _3024_ (.A(net440),
    .X(_0304_));
 sg13g2_buf_1 _3025_ (.A(net324),
    .X(_0305_));
 sg13g2_buf_1 _3026_ (.A(net449),
    .X(_0306_));
 sg13g2_buf_1 _3027_ (.A(net442),
    .X(_0307_));
 sg13g2_buf_1 _3028_ (.A(net444),
    .X(_0308_));
 sg13g2_buf_1 _3029_ (.A(net417),
    .X(_0309_));
 sg13g2_buf_1 _3030_ (.A(net428),
    .X(_0310_));
 sg13g2_buf_1 _3031_ (.A(net375),
    .X(_0311_));
 sg13g2_buf_1 _3032_ (.A(net635),
    .X(_0312_));
 sg13g2_buf_1 _3033_ (.A(net380),
    .X(_0313_));
 sg13g2_buf_1 _3034_ (.A(net621),
    .X(_0314_));
 sg13g2_buf_1 _3035_ (.A(net633),
    .X(_0315_));
 sg13g2_buf_1 _3036_ (.A(net342),
    .X(_0316_));
 sg13g2_buf_1 _3037_ (.A(net458),
    .X(_0317_));
 sg13g2_buf_1 _3038_ (.A(net456),
    .X(_0318_));
 sg13g2_buf_1 _3039_ (.A(net379),
    .X(_0319_));
 sg13g2_buf_1 _3040_ (.A(net455),
    .X(_0320_));
 sg13g2_buf_1 _3041_ (.A(net644),
    .X(_0321_));
 sg13g2_buf_1 _3042_ (.A(net618),
    .X(_0322_));
 sg13g2_buf_1 _3043_ (.A(net617),
    .X(_0323_));
 sg13g2_buf_1 _3044_ (.A(net441),
    .X(_0324_));
 sg13g2_buf_1 _3045_ (.A(net346),
    .X(_0325_));
 sg13g2_buf_1 _3046_ (.A(net636),
    .X(_0326_));
 sg13g2_buf_1 _3047_ (.A(net396),
    .X(_0327_));
 sg13g2_buf_1 _3048_ (.A(net387),
    .X(_0328_));
 sg13g2_buf_1 _3049_ (.A(net348),
    .X(_0329_));
 sg13g2_buf_1 _3050_ (.A(net619),
    .X(_0330_));
 sg13g2_buf_1 _3051_ (.A(net405),
    .X(_0331_));
 sg13g2_buf_1 _3052_ (.A(net622),
    .X(_0332_));
 sg13g2_buf_1 _3053_ (.A(net407),
    .X(_0333_));
 sg13g2_buf_1 _3054_ (.A(net390),
    .X(_0334_));
 sg13g2_buf_1 _3055_ (.A(net645),
    .X(_0335_));
 sg13g2_buf_1 _3056_ (.A(net336),
    .X(_0336_));
 sg13g2_buf_1 _3057_ (.A(net625),
    .X(_0337_));
 sg13g2_buf_1 _3058_ (.A(net435),
    .X(_0338_));
 sg13g2_buf_1 _3059_ (.A(net425),
    .X(_0339_));
 sg13g2_buf_1 _3060_ (.A(net452),
    .X(_0340_));
 sg13g2_buf_1 _3061_ (.A(net416),
    .X(_0341_));
 sg13g2_buf_1 _3062_ (.A(net374),
    .X(_0342_));
 sg13g2_buf_1 _3063_ (.A(net434),
    .X(_0343_));
 sg13g2_buf_1 _3064_ (.A(net368),
    .X(_0344_));
 sg13g2_buf_1 _3065_ (.A(net367),
    .X(_0345_));
 sg13g2_buf_1 _3066_ (.A(net640),
    .X(_0346_));
 sg13g2_buf_1 _3067_ (.A(net626),
    .X(_0347_));
 sg13g2_buf_1 _3068_ (.A(net641),
    .X(_0348_));
 sg13g2_buf_1 _3069_ (.A(net432),
    .X(_0349_));
 sg13g2_buf_1 _3070_ (.A(net392),
    .X(_0350_));
 sg13g2_buf_1 _3071_ (.A(net438),
    .X(_0351_));
 sg13g2_buf_1 _3072_ (.A(net393),
    .X(_0352_));
 sg13g2_buf_1 _3073_ (.A(net623),
    .X(_0353_));
 sg13g2_buf_1 _3074_ (.A(net401),
    .X(_0354_));
 sg13g2_buf_1 _3075_ (.A(net436),
    .X(_0355_));
 sg13g2_buf_1 _3076_ (.A(net427),
    .X(_0356_));
 sg13g2_buf_1 _3077_ (.A(net612),
    .X(_0357_));
 sg13g2_buf_1 _3078_ (.A(net395),
    .X(_0390_));
 sg13g2_buf_1 _3079_ (.A(net349),
    .X(_0391_));
 sg13g2_buf_1 _3080_ (.A(net421),
    .X(_0392_));
 sg13g2_buf_1 _3081_ (.A(net353),
    .X(_0393_));
 sg13g2_buf_1 _3082_ (.A(net402),
    .X(_0394_));
 sg13g2_buf_1 _3083_ (.A(net345),
    .X(_0395_));
 sg13g2_buf_1 _3084_ (.A(net624),
    .X(_0396_));
 sg13g2_buf_1 _3085_ (.A(net327),
    .X(_0397_));
 sg13g2_buf_1 _3086_ (.A(net347),
    .X(_0398_));
 sg13g2_buf_1 _3087_ (.A(net388),
    .X(_0399_));
 sg13g2_buf_1 _3088_ (.A(net412),
    .X(_0400_));
 sg13g2_buf_1 _3089_ (.A(net355),
    .X(_0401_));
 sg13g2_buf_1 _3090_ (.A(net359),
    .X(_0402_));
 sg13g2_buf_1 _3091_ (.A(net639),
    .X(_0403_));
 sg13g2_buf_1 _3092_ (.A(net398),
    .X(_0404_));
 sg13g2_buf_1 _3093_ (.A(net338),
    .X(_0405_));
 sg13g2_buf_1 _3094_ (.A(net614),
    .X(_0406_));
 sg13g2_buf_1 _3095_ (.A(net423),
    .X(_0407_));
 sg13g2_buf_1 _3096_ (.A(net419),
    .X(_0408_));
 sg13g2_buf_1 _3097_ (.A(net410),
    .X(_0409_));
 sg13g2_buf_1 _3098_ (.A(net335),
    .X(_0410_));
 sg13g2_buf_1 _3099_ (.A(net376),
    .X(_0411_));
 sg13g2_buf_1 _3100_ (.A(net373),
    .X(_0412_));
 sg13g2_buf_1 _3101_ (.A(net361),
    .X(_0413_));
 sg13g2_buf_1 _3102_ (.A(net646),
    .X(_0414_));
 sg13g2_buf_1 _3103_ (.A(net360),
    .X(_0415_));
 sg13g2_buf_1 _3104_ (.A(net371),
    .X(_0416_));
 sg13g2_buf_1 _3105_ (.A(net448),
    .X(_0417_));
 sg13g2_buf_1 _3106_ (.A(net439),
    .X(_0418_));
 sg13g2_buf_1 _3107_ (.A(net437),
    .X(_0419_));
 sg13g2_buf_1 _3108_ (.A(net362),
    .X(_0420_));
 sg13g2_buf_1 _3109_ (.A(net377),
    .X(_0421_));
 sg13g2_buf_1 _3110_ (.A(net642),
    .X(_0422_));
 sg13g2_buf_1 _3111_ (.A(net632),
    .X(_0423_));
 sg13g2_buf_1 _3112_ (.A(net445),
    .X(_0424_));
 sg13g2_buf_1 _3113_ (.A(net334),
    .X(_0425_));
 sg13g2_buf_1 _3114_ (.A(net326),
    .X(_0426_));
 sg13g2_buf_1 _3115_ (.A(net330),
    .X(_0427_));
 sg13g2_buf_1 _3116_ (.A(net631),
    .X(_0428_));
 sg13g2_buf_1 _3117_ (.A(net637),
    .X(_0429_));
 sg13g2_buf_1 _3118_ (.A(net627),
    .X(_0430_));
 sg13g2_buf_1 _3119_ (.A(net424),
    .X(_0431_));
 sg13g2_buf_1 _3120_ (.A(net422),
    .X(_0432_));
 sg13g2_buf_1 _3121_ (.A(net332),
    .X(_0433_));
 sg13g2_buf_1 _3122_ (.A(net357),
    .X(_0434_));
 sg13g2_buf_1 _3123_ (.A(net406),
    .X(_0435_));
 sg13g2_buf_1 _3124_ (.A(net643),
    .X(_0436_));
 sg13g2_buf_1 _3125_ (.A(net613),
    .X(_0437_));
 sg13g2_buf_1 _3126_ (.A(net418),
    .X(_0438_));
 sg13g2_buf_1 _3127_ (.A(net457),
    .X(_0439_));
 sg13g2_buf_1 _3128_ (.A(net426),
    .X(_0440_));
 sg13g2_buf_1 _3129_ (.A(net411),
    .X(_0441_));
 sg13g2_buf_1 _3130_ (.A(net630),
    .X(_0442_));
 sg13g2_buf_1 _3131_ (.A(net433),
    .X(_0443_));
 sg13g2_buf_1 _3132_ (.A(net450),
    .X(_0444_));
 sg13g2_buf_1 _3133_ (.A(net369),
    .X(_0445_));
 sg13g2_buf_1 _3134_ (.A(net366),
    .X(_0446_));
 sg13g2_buf_1 _3135_ (.A(net447),
    .X(_0447_));
 sg13g2_buf_1 _3136_ (.A(net408),
    .X(_0448_));
 sg13g2_buf_1 _3137_ (.A(net446),
    .X(_0449_));
 sg13g2_buf_1 _3138_ (.A(net431),
    .X(_0450_));
 sg13g2_buf_1 _3139_ (.A(net394),
    .X(_0451_));
 sg13g2_buf_1 _3140_ (.A(net378),
    .X(_0452_));
 sg13g2_buf_1 _3141_ (.A(net397),
    .X(_0453_));
 sg13g2_buf_1 _3142_ (.A(net443),
    .X(_0454_));
 sg13g2_buf_1 _3143_ (.A(net414),
    .X(_0455_));
 sg13g2_buf_1 _3144_ (.A(net453),
    .X(_0456_));
 sg13g2_buf_1 _3145_ (.A(net399),
    .X(_0457_));
 sg13g2_buf_1 _3146_ (.A(net615),
    .X(_0458_));
 sg13g2_buf_1 _3147_ (.A(net354),
    .X(_0503_));
 sg13g2_buf_1 _3148_ (.A(net343),
    .X(_0504_));
 sg13g2_buf_1 _3149_ (.A(net384),
    .X(_0505_));
 sg13g2_buf_1 _3150_ (.A(net344),
    .X(_0506_));
 sg13g2_buf_1 _3151_ (.A(net413),
    .X(_0507_));
 sg13g2_buf_1 _3152_ (.A(net356),
    .X(_0508_));
 sg13g2_buf_1 _3153_ (.A(net629),
    .X(_0509_));
 sg13g2_buf_1 _3154_ (.A(net389),
    .X(_0510_));
 sg13g2_buf_1 _3155_ (.A(net451),
    .X(_0511_));
 sg13g2_buf_1 _3156_ (.A(net370),
    .X(_0512_));
 sg13g2_buf_1 _3157_ (.A(net429),
    .X(_0513_));
 sg13g2_buf_1 _3158_ (.A(net337),
    .X(_0514_));
 sg13g2_buf_1 _3159_ (.A(net409),
    .X(_0515_));
 sg13g2_buf_1 _3160_ (.A(net333),
    .X(_0516_));
 sg13g2_buf_1 _3161_ (.A(net420),
    .X(_0517_));
 sg13g2_buf_1 _3162_ (.A(net415),
    .X(_0518_));
 sg13g2_buf_1 _3163_ (.A(net383),
    .X(_0519_));
 sg13g2_buf_1 _3164_ (.A(net638),
    .X(_0520_));
 sg13g2_buf_1 _3165_ (.A(net634),
    .X(_0521_));
 sg13g2_buf_1 _3166_ (.A(net404),
    .X(_0522_));
 sg13g2_buf_1 _3167_ (.A(net372),
    .X(_0523_));
 sg13g2_buf_1 _3168_ (.A(net341),
    .X(_0524_));
 sg13g2_buf_1 _3169_ (.A(net454),
    .X(_0525_));
 sg13g2_buf_1 _3170_ (.A(net363),
    .X(_0526_));
 sg13g2_buf_1 _3171_ (.A(net364),
    .X(_0527_));
 sg13g2_buf_1 _3172_ (.A(net365),
    .X(_0528_));
 sg13g2_buf_1 _3173_ (.A(net628),
    .X(_0529_));
 sg13g2_buf_1 _3174_ (.A(net403),
    .X(_0530_));
 sg13g2_buf_1 _3175_ (.A(net616),
    .X(_0531_));
 sg13g2_buf_1 _3176_ (.A(net430),
    .X(_0532_));
 sg13g2_buf_1 _3177_ (.A(net325),
    .X(_0533_));
 sg13g2_dfrbp_1 _3178_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net39),
    .D(_0294_),
    .Q_N(_0293_),
    .Q(\i_soc.cpu.rf.rf[27][0] ));
 sg13g2_dfrbp_1 _3179_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net38),
    .D(_0295_),
    .Q_N(_0292_),
    .Q(\i_soc.cpu.rf.rf[27][1] ));
 sg13g2_dfrbp_1 _3180_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net37),
    .D(_0296_),
    .Q_N(_0291_),
    .Q(\i_soc.cpu.rf.rf[27][2] ));
 sg13g2_dfrbp_1 _3181_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net36),
    .D(_0297_),
    .Q_N(_0290_),
    .Q(\i_soc.cpu.rf.rf[27][3] ));
 sg13g2_dfrbp_1 _3182_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net35),
    .D(_0298_),
    .Q_N(_0289_),
    .Q(\i_soc.cpu.rf.rf[27][4] ));
 sg13g2_dfrbp_1 _3183_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net34),
    .D(_0299_),
    .Q_N(_0288_),
    .Q(\i_soc.cpu.rf.rf[27][5] ));
 sg13g2_dfrbp_1 _3184_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net33),
    .D(_0300_),
    .Q_N(_0287_),
    .Q(\i_soc.cpu.rf.rf[27][6] ));
 sg13g2_dfrbp_1 _3185_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net32),
    .D(_0301_),
    .Q_N(_0286_),
    .Q(\i_soc.cpu.rf.rf[27][7] ));
 sg13g2_dfrbp_1 _3186_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net31),
    .D(_0302_),
    .Q_N(_0285_),
    .Q(\i_soc.cpu.rf.rf[27][8] ));
 sg13g2_dfrbp_1 _3187_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net30),
    .D(_0303_),
    .Q_N(_0284_),
    .Q(\i_soc.cpu.rf.rf[27][9] ));
 sg13g2_dfrbp_1 _3188_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net29),
    .D(_0304_),
    .Q_N(_0283_),
    .Q(\i_soc.cpu.rf.rf[27][10] ));
 sg13g2_dfrbp_1 _3189_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net28),
    .D(_0305_),
    .Q_N(_0282_),
    .Q(\i_soc.cpu.rf.rf[27][11] ));
 sg13g2_dfrbp_1 _3190_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net27),
    .D(_0306_),
    .Q_N(_0281_),
    .Q(\i_soc.cpu.rf.rf[27][12] ));
 sg13g2_dfrbp_1 _3191_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net26),
    .D(_0307_),
    .Q_N(_0280_),
    .Q(\i_soc.cpu.rf.rf[27][13] ));
 sg13g2_dfrbp_1 _3192_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net25),
    .D(_0308_),
    .Q_N(_0279_),
    .Q(\i_soc.cpu.rf.rf[27][14] ));
 sg13g2_dfrbp_1 _3193_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net24),
    .D(_0309_),
    .Q_N(_0278_),
    .Q(\i_soc.cpu.rf.rf[27][15] ));
 sg13g2_dfrbp_1 _3194_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net23),
    .D(_0310_),
    .Q_N(_0277_),
    .Q(\i_soc.cpu.rf.rf[27][16] ));
 sg13g2_dfrbp_1 _3195_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net22),
    .D(_0311_),
    .Q_N(_0276_),
    .Q(\i_soc.cpu.rf.rf[27][17] ));
 sg13g2_dfrbp_1 _3196_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net21),
    .D(_0312_),
    .Q_N(_0275_),
    .Q(\i_soc.cpu.rf.rf[27][18] ));
 sg13g2_dfrbp_1 _3197_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net20),
    .D(_0313_),
    .Q_N(_0274_),
    .Q(\i_soc.cpu.rf.rf[27][19] ));
 sg13g2_dfrbp_1 _3198_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net19),
    .D(_0314_),
    .Q_N(_0273_),
    .Q(\i_soc.cpu.rf.rf[27][20] ));
 sg13g2_dfrbp_1 _3199_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net18),
    .D(_0315_),
    .Q_N(_0272_),
    .Q(\i_soc.cpu.rf.rf[27][21] ));
 sg13g2_dfrbp_1 _3200_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net17),
    .D(_0316_),
    .Q_N(_0271_),
    .Q(\i_soc.cpu.rf.rf[27][22] ));
 sg13g2_dfrbp_1 _3201_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net16),
    .D(_0317_),
    .Q_N(_0270_),
    .Q(\i_soc.cpu.rf.rf[27][23] ));
 sg13g2_dfrbp_1 _3202_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net15),
    .D(_0318_),
    .Q_N(_0269_),
    .Q(\i_soc.cpu.rf.rf[27][24] ));
 sg13g2_dfrbp_1 _3203_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net14),
    .D(_0319_),
    .Q_N(_0268_),
    .Q(\i_soc.cpu.rf.rf[27][25] ));
 sg13g2_dfrbp_1 _3204_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net13),
    .D(_0320_),
    .Q_N(_0267_),
    .Q(\i_soc.cpu.rf.rf[27][26] ));
 sg13g2_dfrbp_1 _3205_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net12),
    .D(_0321_),
    .Q_N(_0266_),
    .Q(\i_soc.cpu.rf.rf[27][27] ));
 sg13g2_dfrbp_1 _3206_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net11),
    .D(_0322_),
    .Q_N(_0265_),
    .Q(\i_soc.cpu.rf.rf[27][28] ));
 sg13g2_dfrbp_1 _3207_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net10),
    .D(_0323_),
    .Q_N(_0264_),
    .Q(\i_soc.cpu.rf.rf[27][29] ));
 sg13g2_dfrbp_1 _3208_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net9),
    .D(_0324_),
    .Q_N(_0263_),
    .Q(\i_soc.cpu.rf.rf[27][30] ));
 sg13g2_dfrbp_1 _3209_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net8),
    .D(_0325_),
    .Q_N(_0262_),
    .Q(\i_soc.cpu.rf.rf[27][31] ));
 sg13g2_dfrbp_1 _3210_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net313),
    .D(_0326_),
    .Q_N(_0261_),
    .Q(\i_soc.cpu.rf.rf[3][0] ));
 sg13g2_dfrbp_1 _3211_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net312),
    .D(_0327_),
    .Q_N(_0260_),
    .Q(\i_soc.cpu.rf.rf[3][1] ));
 sg13g2_dfrbp_1 _3212_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net311),
    .D(_0328_),
    .Q_N(_0259_),
    .Q(\i_soc.cpu.rf.rf[3][2] ));
 sg13g2_dfrbp_1 _3213_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net310),
    .D(_0329_),
    .Q_N(_0258_),
    .Q(\i_soc.cpu.rf.rf[3][3] ));
 sg13g2_dfrbp_1 _3214_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net309),
    .D(_0330_),
    .Q_N(_0257_),
    .Q(\i_soc.cpu.rf.rf[3][4] ));
 sg13g2_dfrbp_1 _3215_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net308),
    .D(_0331_),
    .Q_N(_0256_),
    .Q(\i_soc.cpu.rf.rf[3][5] ));
 sg13g2_dfrbp_1 _3216_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net307),
    .D(_0332_),
    .Q_N(_0255_),
    .Q(\i_soc.cpu.rf.rf[3][6] ));
 sg13g2_dfrbp_1 _3217_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net306),
    .D(_0333_),
    .Q_N(_0254_),
    .Q(\i_soc.cpu.rf.rf[3][7] ));
 sg13g2_dfrbp_1 _3218_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net305),
    .D(_0334_),
    .Q_N(_0253_),
    .Q(\i_soc.cpu.rf.rf[3][8] ));
 sg13g2_dfrbp_1 _3219_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net304),
    .D(_0335_),
    .Q_N(_0252_),
    .Q(\i_soc.cpu.rf.rf[3][9] ));
 sg13g2_dfrbp_1 _3220_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net303),
    .D(_0336_),
    .Q_N(_0251_),
    .Q(\i_soc.cpu.rf.rf[3][10] ));
 sg13g2_dfrbp_1 _3221_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net302),
    .D(_0337_),
    .Q_N(_0250_),
    .Q(\i_soc.cpu.rf.rf[3][11] ));
 sg13g2_dfrbp_1 _3222_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net301),
    .D(_0338_),
    .Q_N(_0249_),
    .Q(\i_soc.cpu.rf.rf[3][12] ));
 sg13g2_dfrbp_1 _3223_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net300),
    .D(_0339_),
    .Q_N(_0248_),
    .Q(\i_soc.cpu.rf.rf[3][13] ));
 sg13g2_dfrbp_1 _3224_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net299),
    .D(_0340_),
    .Q_N(_0247_),
    .Q(\i_soc.cpu.rf.rf[3][14] ));
 sg13g2_dfrbp_1 _3225_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net298),
    .D(_0341_),
    .Q_N(_0246_),
    .Q(\i_soc.cpu.rf.rf[3][15] ));
 sg13g2_dfrbp_1 _3226_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net297),
    .D(_0342_),
    .Q_N(_0245_),
    .Q(\i_soc.cpu.rf.rf[3][16] ));
 sg13g2_dfrbp_1 _3227_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net296),
    .D(_0343_),
    .Q_N(_0244_),
    .Q(\i_soc.cpu.rf.rf[3][17] ));
 sg13g2_dfrbp_1 _3228_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net295),
    .D(_0344_),
    .Q_N(_0243_),
    .Q(\i_soc.cpu.rf.rf[3][18] ));
 sg13g2_dfrbp_1 _3229_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net294),
    .D(_0345_),
    .Q_N(_0242_),
    .Q(\i_soc.cpu.rf.rf[3][19] ));
 sg13g2_dfrbp_1 _3230_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net293),
    .D(_0346_),
    .Q_N(_0241_),
    .Q(\i_soc.cpu.rf.rf[3][20] ));
 sg13g2_dfrbp_1 _3231_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net292),
    .D(_0347_),
    .Q_N(_0240_),
    .Q(\i_soc.cpu.rf.rf[3][21] ));
 sg13g2_dfrbp_1 _3232_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net291),
    .D(_0348_),
    .Q_N(_0239_),
    .Q(\i_soc.cpu.rf.rf[3][22] ));
 sg13g2_dfrbp_1 _3233_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net290),
    .D(_0349_),
    .Q_N(_0238_),
    .Q(\i_soc.cpu.rf.rf[3][23] ));
 sg13g2_dfrbp_1 _3234_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net289),
    .D(_0350_),
    .Q_N(_0237_),
    .Q(\i_soc.cpu.rf.rf[3][24] ));
 sg13g2_dfrbp_1 _3235_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net288),
    .D(_0351_),
    .Q_N(_0236_),
    .Q(\i_soc.cpu.rf.rf[3][25] ));
 sg13g2_dfrbp_1 _3236_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net287),
    .D(_0352_),
    .Q_N(_0235_),
    .Q(\i_soc.cpu.rf.rf[3][26] ));
 sg13g2_dfrbp_1 _3237_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net286),
    .D(_0353_),
    .Q_N(_0234_),
    .Q(\i_soc.cpu.rf.rf[3][27] ));
 sg13g2_dfrbp_1 _3238_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net285),
    .D(_0354_),
    .Q_N(_0233_),
    .Q(\i_soc.cpu.rf.rf[3][28] ));
 sg13g2_dfrbp_1 _3239_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net284),
    .D(_0355_),
    .Q_N(_0232_),
    .Q(\i_soc.cpu.rf.rf[3][29] ));
 sg13g2_dfrbp_1 _3240_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net283),
    .D(_0356_),
    .Q_N(_0231_),
    .Q(\i_soc.cpu.rf.rf[3][30] ));
 sg13g2_dfrbp_1 _3241_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net282),
    .D(_0357_),
    .Q_N(_0230_),
    .Q(\i_soc.cpu.rf.rf[3][31] ));
 sg13g2_dfrbp_1 _3242_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net281),
    .D(_0358_),
    .Q_N(_0229_),
    .Q(\i_soc.cpu.rd0[0] ));
 sg13g2_dfrbp_1 _3243_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net280),
    .D(_0359_),
    .Q_N(_0228_),
    .Q(\i_soc.cpu.rd0[1] ));
 sg13g2_dfrbp_1 _3244_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net279),
    .D(_0360_),
    .Q_N(_0227_),
    .Q(\i_soc.cpu.rd0[2] ));
 sg13g2_dfrbp_1 _3245_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net278),
    .D(_0361_),
    .Q_N(_0226_),
    .Q(\i_soc.cpu.rd0[3] ));
 sg13g2_dfrbp_1 _3246_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net277),
    .D(_0362_),
    .Q_N(_0225_),
    .Q(\i_soc.cpu.rd0[4] ));
 sg13g2_dfrbp_1 _3247_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net276),
    .D(_0363_),
    .Q_N(_0224_),
    .Q(\i_soc.cpu.rd0[5] ));
 sg13g2_dfrbp_1 _3248_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net275),
    .D(_0364_),
    .Q_N(_0223_),
    .Q(\i_soc.cpu.rd0[6] ));
 sg13g2_dfrbp_1 _3249_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net274),
    .D(_0365_),
    .Q_N(_0222_),
    .Q(\i_soc.cpu.rd0[7] ));
 sg13g2_dfrbp_1 _3250_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net273),
    .D(_0366_),
    .Q_N(_0221_),
    .Q(\i_soc.cpu.rd0[8] ));
 sg13g2_dfrbp_1 _3251_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net272),
    .D(_0367_),
    .Q_N(_0220_),
    .Q(\i_soc.cpu.rd0[9] ));
 sg13g2_dfrbp_1 _3252_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net271),
    .D(_0368_),
    .Q_N(_0219_),
    .Q(\i_soc.cpu.rd0[10] ));
 sg13g2_dfrbp_1 _3253_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net270),
    .D(_0369_),
    .Q_N(_0218_),
    .Q(\i_soc.cpu.rd0[11] ));
 sg13g2_dfrbp_1 _3254_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net269),
    .D(_0370_),
    .Q_N(_0217_),
    .Q(\i_soc.cpu.rd0[12] ));
 sg13g2_dfrbp_1 _3255_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net268),
    .D(_0371_),
    .Q_N(_0216_),
    .Q(\i_soc.cpu.rd0[13] ));
 sg13g2_dfrbp_1 _3256_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net267),
    .D(_0372_),
    .Q_N(_0215_),
    .Q(\i_soc.cpu.rd0[14] ));
 sg13g2_dfrbp_1 _3257_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net266),
    .D(_0373_),
    .Q_N(_0214_),
    .Q(\i_soc.cpu.rd0[15] ));
 sg13g2_dfrbp_1 _3258_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net265),
    .D(_0374_),
    .Q_N(_0213_),
    .Q(\i_soc.cpu.rd0[16] ));
 sg13g2_dfrbp_1 _3259_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net264),
    .D(_0375_),
    .Q_N(_0212_),
    .Q(\i_soc.cpu.rd0[17] ));
 sg13g2_dfrbp_1 _3260_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net263),
    .D(_0376_),
    .Q_N(_0211_),
    .Q(\i_soc.cpu.rd0[18] ));
 sg13g2_dfrbp_1 _3261_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net262),
    .D(_0377_),
    .Q_N(_0210_),
    .Q(\i_soc.cpu.rd0[19] ));
 sg13g2_dfrbp_1 _3262_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net261),
    .D(_0378_),
    .Q_N(_0209_),
    .Q(\i_soc.cpu.rd0[20] ));
 sg13g2_dfrbp_1 _3263_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net260),
    .D(_0379_),
    .Q_N(_0208_),
    .Q(\i_soc.cpu.rd0[21] ));
 sg13g2_dfrbp_1 _3264_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net259),
    .D(_0380_),
    .Q_N(_0207_),
    .Q(\i_soc.cpu.rd0[22] ));
 sg13g2_dfrbp_1 _3265_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net258),
    .D(_0381_),
    .Q_N(_0206_),
    .Q(\i_soc.cpu.rd0[23] ));
 sg13g2_dfrbp_1 _3266_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net257),
    .D(_0382_),
    .Q_N(_0205_),
    .Q(\i_soc.cpu.rd0[24] ));
 sg13g2_dfrbp_1 _3267_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net256),
    .D(_0383_),
    .Q_N(_0204_),
    .Q(\i_soc.cpu.rd0[25] ));
 sg13g2_dfrbp_1 _3268_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net255),
    .D(_0384_),
    .Q_N(_0203_),
    .Q(\i_soc.cpu.rd0[26] ));
 sg13g2_dfrbp_1 _3269_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net254),
    .D(_0385_),
    .Q_N(_0202_),
    .Q(\i_soc.cpu.rd0[27] ));
 sg13g2_dfrbp_1 _3270_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net253),
    .D(_0386_),
    .Q_N(_0201_),
    .Q(\i_soc.cpu.rd0[28] ));
 sg13g2_dfrbp_1 _3271_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net252),
    .D(_0387_),
    .Q_N(_0200_),
    .Q(\i_soc.cpu.rd0[29] ));
 sg13g2_dfrbp_1 _3272_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net251),
    .D(_0388_),
    .Q_N(_0199_),
    .Q(\i_soc.cpu.rd0[30] ));
 sg13g2_dfrbp_1 _3273_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net250),
    .D(_0389_),
    .Q_N(_0198_),
    .Q(\i_soc.cpu.rd0[31] ));
 sg13g2_dfrbp_1 _3274_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net249),
    .D(_0390_),
    .Q_N(_0197_),
    .Q(\i_soc.cpu.rf.rf[0][0] ));
 sg13g2_dfrbp_1 _3275_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net248),
    .D(_0391_),
    .Q_N(_0196_),
    .Q(\i_soc.cpu.rf.rf[0][1] ));
 sg13g2_dfrbp_1 _3276_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net247),
    .D(_0392_),
    .Q_N(_0195_),
    .Q(\i_soc.cpu.rf.rf[0][2] ));
 sg13g2_dfrbp_1 _3277_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net246),
    .D(_0393_),
    .Q_N(_0194_),
    .Q(\i_soc.cpu.rf.rf[0][3] ));
 sg13g2_dfrbp_1 _3278_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net245),
    .D(_0394_),
    .Q_N(_0193_),
    .Q(\i_soc.cpu.rf.rf[0][30] ));
 sg13g2_dfrbp_1 _3279_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net244),
    .D(_0395_),
    .Q_N(_0192_),
    .Q(\i_soc.cpu.rf.rf[8][0] ));
 sg13g2_dfrbp_1 _3280_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net243),
    .D(_0396_),
    .Q_N(_0191_),
    .Q(\i_soc.cpu.rf.rf[8][1] ));
 sg13g2_dfrbp_1 _3281_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net242),
    .D(_0397_),
    .Q_N(_0190_),
    .Q(\i_soc.cpu.rf.rf[8][2] ));
 sg13g2_dfrbp_1 _3282_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net241),
    .D(_0398_),
    .Q_N(_0189_),
    .Q(\i_soc.cpu.rf.rf[8][3] ));
 sg13g2_dfrbp_1 _3283_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net240),
    .D(_0399_),
    .Q_N(_0188_),
    .Q(\i_soc.cpu.rf.rf[8][4] ));
 sg13g2_dfrbp_1 _3284_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net239),
    .D(_0400_),
    .Q_N(_0187_),
    .Q(\i_soc.cpu.rf.rf[8][5] ));
 sg13g2_dfrbp_1 _3285_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net238),
    .D(_0401_),
    .Q_N(_0186_),
    .Q(\i_soc.cpu.rf.rf[8][6] ));
 sg13g2_dfrbp_1 _3286_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net237),
    .D(_0402_),
    .Q_N(_0185_),
    .Q(\i_soc.cpu.rf.rf[8][7] ));
 sg13g2_dfrbp_1 _3287_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net236),
    .D(_0403_),
    .Q_N(_0184_),
    .Q(\i_soc.cpu.rf.rf[8][8] ));
 sg13g2_dfrbp_1 _3288_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net235),
    .D(_0404_),
    .Q_N(_0183_),
    .Q(\i_soc.cpu.rf.rf[8][9] ));
 sg13g2_dfrbp_1 _3289_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net234),
    .D(_0405_),
    .Q_N(_0182_),
    .Q(\i_soc.cpu.rf.rf[8][10] ));
 sg13g2_dfrbp_1 _3290_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net233),
    .D(_0406_),
    .Q_N(_0181_),
    .Q(\i_soc.cpu.rf.rf[8][11] ));
 sg13g2_dfrbp_1 _3291_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net232),
    .D(_0407_),
    .Q_N(_0180_),
    .Q(\i_soc.cpu.rf.rf[8][12] ));
 sg13g2_dfrbp_1 _3292_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net231),
    .D(_0408_),
    .Q_N(_0179_),
    .Q(\i_soc.cpu.rf.rf[8][13] ));
 sg13g2_dfrbp_1 _3293_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net230),
    .D(_0409_),
    .Q_N(_0178_),
    .Q(\i_soc.cpu.rf.rf[8][14] ));
 sg13g2_dfrbp_1 _3294_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net229),
    .D(_0410_),
    .Q_N(_0177_),
    .Q(\i_soc.cpu.rf.rf[8][15] ));
 sg13g2_dfrbp_1 _3295_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net228),
    .D(_0411_),
    .Q_N(_0176_),
    .Q(\i_soc.cpu.rf.rf[8][16] ));
 sg13g2_dfrbp_1 _3296_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net227),
    .D(_0412_),
    .Q_N(_0175_),
    .Q(\i_soc.cpu.rf.rf[8][17] ));
 sg13g2_dfrbp_1 _3297_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net226),
    .D(_0413_),
    .Q_N(_0174_),
    .Q(\i_soc.cpu.rf.rf[8][18] ));
 sg13g2_dfrbp_1 _3298_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net225),
    .D(_0414_),
    .Q_N(_0173_),
    .Q(\i_soc.cpu.rf.rf[8][19] ));
 sg13g2_dfrbp_1 _3299_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net224),
    .D(_0415_),
    .Q_N(_0172_),
    .Q(\i_soc.cpu.rf.rf[8][20] ));
 sg13g2_dfrbp_1 _3300_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net223),
    .D(_0416_),
    .Q_N(_0171_),
    .Q(\i_soc.cpu.rf.rf[8][21] ));
 sg13g2_dfrbp_1 _3301_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net222),
    .D(_0417_),
    .Q_N(_0170_),
    .Q(\i_soc.cpu.rf.rf[8][22] ));
 sg13g2_dfrbp_1 _3302_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net221),
    .D(_0418_),
    .Q_N(_0169_),
    .Q(\i_soc.cpu.rf.rf[8][23] ));
 sg13g2_dfrbp_1 _3303_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net220),
    .D(_0419_),
    .Q_N(_0168_),
    .Q(\i_soc.cpu.rf.rf[8][24] ));
 sg13g2_dfrbp_1 _3304_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net219),
    .D(_0420_),
    .Q_N(_0167_),
    .Q(\i_soc.cpu.rf.rf[8][25] ));
 sg13g2_dfrbp_1 _3305_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net218),
    .D(_0421_),
    .Q_N(_0166_),
    .Q(\i_soc.cpu.rf.rf[8][26] ));
 sg13g2_dfrbp_1 _3306_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net217),
    .D(_0422_),
    .Q_N(_0165_),
    .Q(\i_soc.cpu.rf.rf[8][27] ));
 sg13g2_dfrbp_1 _3307_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net216),
    .D(_0423_),
    .Q_N(_0164_),
    .Q(\i_soc.cpu.rf.rf[8][28] ));
 sg13g2_dfrbp_1 _3308_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net215),
    .D(_0424_),
    .Q_N(_0163_),
    .Q(\i_soc.cpu.rf.rf[8][29] ));
 sg13g2_dfrbp_1 _3309_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net214),
    .D(_0425_),
    .Q_N(_0162_),
    .Q(\i_soc.cpu.rf.rf[8][30] ));
 sg13g2_dfrbp_1 _3310_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net213),
    .D(_0426_),
    .Q_N(_0161_),
    .Q(\i_soc.cpu.rf.rf[8][31] ));
 sg13g2_dfrbp_1 _3311_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net212),
    .D(_0427_),
    .Q_N(_0160_),
    .Q(\i_soc.cpu.rf.rf[1][0] ));
 sg13g2_dfrbp_1 _3312_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net211),
    .D(_0428_),
    .Q_N(_0159_),
    .Q(\i_soc.cpu.rf.rf[1][1] ));
 sg13g2_dfrbp_1 _3313_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net210),
    .D(_0429_),
    .Q_N(_0158_),
    .Q(\i_soc.cpu.rf.rf[1][2] ));
 sg13g2_dfrbp_1 _3314_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net209),
    .D(_0430_),
    .Q_N(_0157_),
    .Q(\i_soc.cpu.rf.rf[1][3] ));
 sg13g2_dfrbp_1 _3315_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net208),
    .D(_0431_),
    .Q_N(_0156_),
    .Q(\i_soc.cpu.rf.rf[1][4] ));
 sg13g2_dfrbp_1 _3316_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net207),
    .D(_0432_),
    .Q_N(_0155_),
    .Q(\i_soc.cpu.rf.rf[1][5] ));
 sg13g2_dfrbp_1 _3317_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net206),
    .D(_0433_),
    .Q_N(_0154_),
    .Q(\i_soc.cpu.rf.rf[1][6] ));
 sg13g2_dfrbp_1 _3318_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net205),
    .D(_0434_),
    .Q_N(_0153_),
    .Q(\i_soc.cpu.rf.rf[1][7] ));
 sg13g2_dfrbp_1 _3319_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net204),
    .D(_0435_),
    .Q_N(_0152_),
    .Q(\i_soc.cpu.rf.rf[1][8] ));
 sg13g2_dfrbp_1 _3320_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net203),
    .D(_0436_),
    .Q_N(_0151_),
    .Q(\i_soc.cpu.rf.rf[1][9] ));
 sg13g2_dfrbp_1 _3321_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net202),
    .D(_0437_),
    .Q_N(_0150_),
    .Q(\i_soc.cpu.rf.rf[1][10] ));
 sg13g2_dfrbp_1 _3322_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net201),
    .D(_0438_),
    .Q_N(_0149_),
    .Q(\i_soc.cpu.rf.rf[1][11] ));
 sg13g2_dfrbp_1 _3323_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net200),
    .D(_0439_),
    .Q_N(_0148_),
    .Q(\i_soc.cpu.rf.rf[1][12] ));
 sg13g2_dfrbp_1 _3324_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net199),
    .D(_0440_),
    .Q_N(_0147_),
    .Q(\i_soc.cpu.rf.rf[1][13] ));
 sg13g2_dfrbp_1 _3325_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net198),
    .D(_0441_),
    .Q_N(_0146_),
    .Q(\i_soc.cpu.rf.rf[1][14] ));
 sg13g2_dfrbp_1 _3326_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net197),
    .D(_0442_),
    .Q_N(_0145_),
    .Q(\i_soc.cpu.rf.rf[1][15] ));
 sg13g2_dfrbp_1 _3327_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net196),
    .D(_0443_),
    .Q_N(_0144_),
    .Q(\i_soc.cpu.rf.rf[1][16] ));
 sg13g2_dfrbp_1 _3328_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net195),
    .D(_0444_),
    .Q_N(_0143_),
    .Q(\i_soc.cpu.rf.rf[1][17] ));
 sg13g2_dfrbp_1 _3329_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net194),
    .D(_0445_),
    .Q_N(_0142_),
    .Q(\i_soc.cpu.rf.rf[1][18] ));
 sg13g2_dfrbp_1 _3330_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net193),
    .D(_0446_),
    .Q_N(_0141_),
    .Q(\i_soc.cpu.rf.rf[1][19] ));
 sg13g2_dfrbp_1 _3331_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net192),
    .D(_0447_),
    .Q_N(_0140_),
    .Q(\i_soc.cpu.rf.rf[1][20] ));
 sg13g2_dfrbp_1 _3332_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net191),
    .D(_0448_),
    .Q_N(_0139_),
    .Q(\i_soc.cpu.rf.rf[1][21] ));
 sg13g2_dfrbp_1 _3333_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net190),
    .D(_0449_),
    .Q_N(_0138_),
    .Q(\i_soc.cpu.rf.rf[1][22] ));
 sg13g2_dfrbp_1 _3334_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net189),
    .D(_0450_),
    .Q_N(_0137_),
    .Q(\i_soc.cpu.rf.rf[1][23] ));
 sg13g2_dfrbp_1 _3335_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net188),
    .D(_0451_),
    .Q_N(_0136_),
    .Q(\i_soc.cpu.rf.rf[1][24] ));
 sg13g2_dfrbp_1 _3336_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net187),
    .D(_0452_),
    .Q_N(_0135_),
    .Q(\i_soc.cpu.rf.rf[1][25] ));
 sg13g2_dfrbp_1 _3337_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net186),
    .D(_0453_),
    .Q_N(_0134_),
    .Q(\i_soc.cpu.rf.rf[1][26] ));
 sg13g2_dfrbp_1 _3338_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net185),
    .D(_0454_),
    .Q_N(_0133_),
    .Q(\i_soc.cpu.rf.rf[1][27] ));
 sg13g2_dfrbp_1 _3339_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net184),
    .D(_0455_),
    .Q_N(_0132_),
    .Q(\i_soc.cpu.rf.rf[1][28] ));
 sg13g2_dfrbp_1 _3340_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net183),
    .D(_0456_),
    .Q_N(_0131_),
    .Q(\i_soc.cpu.rf.rf[1][29] ));
 sg13g2_dfrbp_1 _3341_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net182),
    .D(_0457_),
    .Q_N(_0130_),
    .Q(\i_soc.cpu.rf.rf[1][30] ));
 sg13g2_dfrbp_1 _3342_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net181),
    .D(_0458_),
    .Q_N(_0129_),
    .Q(\i_soc.cpu.rf.rf[1][31] ));
 sg13g2_dfrbp_1 _3343_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net180),
    .D(_0459_),
    .Q_N(_0128_),
    .Q(\i_soc.cpu.rf.rf[5][0] ));
 sg13g2_dfrbp_1 _3344_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net179),
    .D(_0460_),
    .Q_N(_0127_),
    .Q(\i_soc.cpu.rf.rf[5][1] ));
 sg13g2_dfrbp_1 _3345_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net178),
    .D(_0461_),
    .Q_N(_0126_),
    .Q(\i_soc.cpu.rf.rf[5][2] ));
 sg13g2_dfrbp_1 _3346_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net177),
    .D(_0462_),
    .Q_N(_0125_),
    .Q(\i_soc.cpu.rf.rf[5][3] ));
 sg13g2_dfrbp_1 _3347_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net176),
    .D(_0463_),
    .Q_N(_0124_),
    .Q(\i_soc.cpu.rf.rf[5][4] ));
 sg13g2_dfrbp_1 _3348_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net175),
    .D(_0464_),
    .Q_N(_0123_),
    .Q(\i_soc.cpu.rf.rf[5][5] ));
 sg13g2_dfrbp_1 _3349_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net174),
    .D(_0465_),
    .Q_N(_0122_),
    .Q(\i_soc.cpu.rf.rf[5][6] ));
 sg13g2_dfrbp_1 _3350_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net173),
    .D(_0466_),
    .Q_N(_0121_),
    .Q(\i_soc.cpu.rf.rf[5][7] ));
 sg13g2_dfrbp_1 _3351_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net172),
    .D(_0467_),
    .Q_N(_0120_),
    .Q(\i_soc.cpu.rf.rf[5][8] ));
 sg13g2_dfrbp_1 _3352_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net171),
    .D(_0468_),
    .Q_N(_0119_),
    .Q(\i_soc.cpu.rf.rf[5][9] ));
 sg13g2_dfrbp_1 _3353_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net170),
    .D(_0469_),
    .Q_N(_0118_),
    .Q(\i_soc.cpu.rf.rf[5][10] ));
 sg13g2_dfrbp_1 _3354_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net169),
    .D(_0470_),
    .Q_N(_0117_),
    .Q(\i_soc.cpu.rf.rf[5][11] ));
 sg13g2_dfrbp_1 _3355_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net168),
    .D(_0471_),
    .Q_N(_0116_),
    .Q(\i_soc.cpu.rf.rf[5][12] ));
 sg13g2_dfrbp_1 _3356_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net167),
    .D(_0472_),
    .Q_N(_0115_),
    .Q(\i_soc.cpu.rf.rf[5][13] ));
 sg13g2_dfrbp_1 _3357_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net166),
    .D(_0473_),
    .Q_N(_0114_),
    .Q(\i_soc.cpu.rf.rf[5][14] ));
 sg13g2_dfrbp_1 _3358_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net165),
    .D(_0474_),
    .Q_N(_0113_),
    .Q(\i_soc.cpu.rf.rf[5][15] ));
 sg13g2_dfrbp_1 _3359_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net164),
    .D(_0475_),
    .Q_N(_0112_),
    .Q(\i_soc.cpu.rf.rf[5][16] ));
 sg13g2_dfrbp_1 _3360_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net163),
    .D(_0476_),
    .Q_N(_0111_),
    .Q(\i_soc.cpu.rf.rf[5][17] ));
 sg13g2_dfrbp_1 _3361_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net162),
    .D(_0477_),
    .Q_N(_0110_),
    .Q(\i_soc.cpu.rf.rf[5][18] ));
 sg13g2_dfrbp_1 _3362_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net161),
    .D(_0478_),
    .Q_N(_0109_),
    .Q(\i_soc.cpu.rf.rf[5][19] ));
 sg13g2_dfrbp_1 _3363_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net160),
    .D(_0479_),
    .Q_N(_0108_),
    .Q(\i_soc.cpu.rf.rf[5][20] ));
 sg13g2_dfrbp_1 _3364_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net159),
    .D(_0480_),
    .Q_N(_0107_),
    .Q(\i_soc.cpu.rf.rf[5][21] ));
 sg13g2_dfrbp_1 _3365_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net158),
    .D(_0481_),
    .Q_N(_0106_),
    .Q(\i_soc.cpu.rf.rf[5][22] ));
 sg13g2_dfrbp_1 _3366_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net157),
    .D(_0482_),
    .Q_N(_0105_),
    .Q(\i_soc.cpu.rf.rf[5][23] ));
 sg13g2_dfrbp_1 _3367_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net156),
    .D(_0483_),
    .Q_N(_0104_),
    .Q(\i_soc.cpu.rf.rf[5][24] ));
 sg13g2_dfrbp_1 _3368_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net155),
    .D(_0484_),
    .Q_N(_0103_),
    .Q(\i_soc.cpu.rf.rf[5][25] ));
 sg13g2_dfrbp_1 _3369_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net154),
    .D(_0485_),
    .Q_N(_0102_),
    .Q(\i_soc.cpu.rf.rf[5][26] ));
 sg13g2_dfrbp_1 _3370_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net153),
    .D(_0486_),
    .Q_N(_0101_),
    .Q(\i_soc.cpu.rf.rf[5][27] ));
 sg13g2_dfrbp_1 _3371_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net152),
    .D(_0487_),
    .Q_N(_0100_),
    .Q(\i_soc.cpu.rf.rf[5][28] ));
 sg13g2_dfrbp_1 _3372_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net151),
    .D(_0488_),
    .Q_N(_0099_),
    .Q(\i_soc.cpu.rf.rf[5][29] ));
 sg13g2_dfrbp_1 _3373_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net150),
    .D(_0489_),
    .Q_N(_0098_),
    .Q(\i_soc.cpu.rf.rf[5][30] ));
 sg13g2_dfrbp_1 _3374_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net149),
    .D(_0490_),
    .Q_N(_0097_),
    .Q(\i_soc.cpu.rf.rf[5][31] ));
 sg13g2_dfrbp_1 _3375_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net148),
    .D(_0491_),
    .Q_N(_0096_),
    .Q(\i_soc.cnt[0] ));
 sg13g2_dfrbp_1 _3376_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net147),
    .D(net744),
    .Q_N(_1588_),
    .Q(\i_soc.cnt[1] ));
 sg13g2_dfrbp_1 _3377_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net146),
    .D(_0493_),
    .Q_N(_1587_),
    .Q(\i_soc.cnt[2] ));
 sg13g2_dfrbp_1 _3378_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net145),
    .D(_0494_),
    .Q_N(_1586_),
    .Q(\i_soc.cnt[3] ));
 sg13g2_dfrbp_1 _3379_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net144),
    .D(_0495_),
    .Q_N(_1585_),
    .Q(\i_soc.cnt[4] ));
 sg13g2_dfrbp_1 _3380_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net143),
    .D(_0496_),
    .Q_N(_1584_),
    .Q(\i_soc.cnt[5] ));
 sg13g2_dfrbp_1 _3381_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net142),
    .D(net759),
    .Q_N(_1583_),
    .Q(\i_soc.cnt[6] ));
 sg13g2_dfrbp_1 _3382_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net141),
    .D(_0498_),
    .Q_N(_1582_),
    .Q(\i_soc.cnt[7] ));
 sg13g2_dfrbp_1 _3383_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net139),
    .D(_0499_),
    .Q_N(_0095_),
    .Q(\i_soc.cpu.pc[2] ));
 sg13g2_dfrbp_1 _3384_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net138),
    .D(_0500_),
    .Q_N(_1581_),
    .Q(\i_soc.cpu.pc[3] ));
 sg13g2_dfrbp_1 _3385_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net137),
    .D(_0501_),
    .Q_N(_1580_),
    .Q(\i_soc.cpu.pc[4] ));
 sg13g2_dfrbp_1 _3386_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net136),
    .D(_0502_),
    .Q_N(_1579_),
    .Q(\i_soc.cpu.pc[5] ));
 sg13g2_dfrbp_1 _3387_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net135),
    .D(_0503_),
    .Q_N(_0094_),
    .Q(\i_soc.cpu.rf.rf[11][0] ));
 sg13g2_dfrbp_1 _3388_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net134),
    .D(_0504_),
    .Q_N(_0093_),
    .Q(\i_soc.cpu.rf.rf[11][1] ));
 sg13g2_dfrbp_1 _3389_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net133),
    .D(_0505_),
    .Q_N(_0092_),
    .Q(\i_soc.cpu.rf.rf[11][2] ));
 sg13g2_dfrbp_1 _3390_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net132),
    .D(_0506_),
    .Q_N(_0091_),
    .Q(\i_soc.cpu.rf.rf[11][3] ));
 sg13g2_dfrbp_1 _3391_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net131),
    .D(_0507_),
    .Q_N(_0090_),
    .Q(\i_soc.cpu.rf.rf[11][4] ));
 sg13g2_dfrbp_1 _3392_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net130),
    .D(_0508_),
    .Q_N(_0089_),
    .Q(\i_soc.cpu.rf.rf[11][5] ));
 sg13g2_dfrbp_1 _3393_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net129),
    .D(_0509_),
    .Q_N(_0088_),
    .Q(\i_soc.cpu.rf.rf[11][6] ));
 sg13g2_dfrbp_1 _3394_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net128),
    .D(_0510_),
    .Q_N(_0087_),
    .Q(\i_soc.cpu.rf.rf[11][7] ));
 sg13g2_dfrbp_1 _3395_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net127),
    .D(_0511_),
    .Q_N(_0086_),
    .Q(\i_soc.cpu.rf.rf[11][8] ));
 sg13g2_dfrbp_1 _3396_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net126),
    .D(_0512_),
    .Q_N(_0085_),
    .Q(\i_soc.cpu.rf.rf[11][9] ));
 sg13g2_dfrbp_1 _3397_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net125),
    .D(_0513_),
    .Q_N(_0084_),
    .Q(\i_soc.cpu.rf.rf[11][10] ));
 sg13g2_dfrbp_1 _3398_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net124),
    .D(_0514_),
    .Q_N(_0083_),
    .Q(\i_soc.cpu.rf.rf[11][11] ));
 sg13g2_dfrbp_1 _3399_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net123),
    .D(_0515_),
    .Q_N(_0082_),
    .Q(\i_soc.cpu.rf.rf[11][12] ));
 sg13g2_dfrbp_1 _3400_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net122),
    .D(_0516_),
    .Q_N(_0081_),
    .Q(\i_soc.cpu.rf.rf[11][13] ));
 sg13g2_dfrbp_1 _3401_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net121),
    .D(_0517_),
    .Q_N(_0080_),
    .Q(\i_soc.cpu.rf.rf[11][14] ));
 sg13g2_dfrbp_1 _3402_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net120),
    .D(_0518_),
    .Q_N(_0079_),
    .Q(\i_soc.cpu.rf.rf[11][15] ));
 sg13g2_dfrbp_1 _3403_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net119),
    .D(_0519_),
    .Q_N(_0078_),
    .Q(\i_soc.cpu.rf.rf[11][16] ));
 sg13g2_dfrbp_1 _3404_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net118),
    .D(_0520_),
    .Q_N(_0077_),
    .Q(\i_soc.cpu.rf.rf[11][17] ));
 sg13g2_dfrbp_1 _3405_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net117),
    .D(_0521_),
    .Q_N(_0076_),
    .Q(\i_soc.cpu.rf.rf[11][18] ));
 sg13g2_dfrbp_1 _3406_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net116),
    .D(_0522_),
    .Q_N(_0075_),
    .Q(\i_soc.cpu.rf.rf[11][19] ));
 sg13g2_dfrbp_1 _3407_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net115),
    .D(_0523_),
    .Q_N(_0074_),
    .Q(\i_soc.cpu.rf.rf[11][20] ));
 sg13g2_dfrbp_1 _3408_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net114),
    .D(_0524_),
    .Q_N(_0073_),
    .Q(\i_soc.cpu.rf.rf[11][21] ));
 sg13g2_dfrbp_1 _3409_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net113),
    .D(_0525_),
    .Q_N(_0072_),
    .Q(\i_soc.cpu.rf.rf[11][22] ));
 sg13g2_dfrbp_1 _3410_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net112),
    .D(_0526_),
    .Q_N(_0071_),
    .Q(\i_soc.cpu.rf.rf[11][24] ));
 sg13g2_dfrbp_1 _3411_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net111),
    .D(_0527_),
    .Q_N(_0070_),
    .Q(\i_soc.cpu.rf.rf[11][25] ));
 sg13g2_dfrbp_1 _3412_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net110),
    .D(_0528_),
    .Q_N(_0069_),
    .Q(\i_soc.cpu.rf.rf[11][26] ));
 sg13g2_dfrbp_1 _3413_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net109),
    .D(_0529_),
    .Q_N(_0068_),
    .Q(\i_soc.cpu.rf.rf[11][27] ));
 sg13g2_dfrbp_1 _3414_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net108),
    .D(_0530_),
    .Q_N(_0067_),
    .Q(\i_soc.cpu.rf.rf[11][28] ));
 sg13g2_dfrbp_1 _3415_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net107),
    .D(_0531_),
    .Q_N(_0066_),
    .Q(\i_soc.cpu.rf.rf[11][29] ));
 sg13g2_dfrbp_1 _3416_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net106),
    .D(_0532_),
    .Q_N(_0065_),
    .Q(\i_soc.cpu.rf.rf[11][30] ));
 sg13g2_dfrbp_1 _3417_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net105),
    .D(_0533_),
    .Q_N(_0064_),
    .Q(\i_soc.cpu.rf.rf[11][31] ));
 sg13g2_dfrbp_1 _3418_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net104),
    .D(_0534_),
    .Q_N(_0063_),
    .Q(\i_soc.cpu.rf.rf[7][0] ));
 sg13g2_dfrbp_1 _3419_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net103),
    .D(_0535_),
    .Q_N(_0062_),
    .Q(\i_soc.cpu.rf.rf[7][1] ));
 sg13g2_dfrbp_1 _3420_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net102),
    .D(_0536_),
    .Q_N(_0061_),
    .Q(\i_soc.cpu.rf.rf[7][2] ));
 sg13g2_dfrbp_1 _3421_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net101),
    .D(_0537_),
    .Q_N(_0060_),
    .Q(\i_soc.cpu.rf.rf[7][3] ));
 sg13g2_dfrbp_1 _3422_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net100),
    .D(_0538_),
    .Q_N(_0059_),
    .Q(\i_soc.cpu.rf.rf[7][4] ));
 sg13g2_dfrbp_1 _3423_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net99),
    .D(_0539_),
    .Q_N(_0058_),
    .Q(\i_soc.cpu.rf.rf[7][5] ));
 sg13g2_dfrbp_1 _3424_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net98),
    .D(_0540_),
    .Q_N(_0057_),
    .Q(\i_soc.cpu.rf.rf[7][6] ));
 sg13g2_dfrbp_1 _3425_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net97),
    .D(_0541_),
    .Q_N(_0056_),
    .Q(\i_soc.cpu.rf.rf[7][7] ));
 sg13g2_dfrbp_1 _3426_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net96),
    .D(_0542_),
    .Q_N(_0055_),
    .Q(\i_soc.cpu.rf.rf[7][8] ));
 sg13g2_dfrbp_1 _3427_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net95),
    .D(_0543_),
    .Q_N(_0054_),
    .Q(\i_soc.cpu.rf.rf[7][9] ));
 sg13g2_dfrbp_1 _3428_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net94),
    .D(_0544_),
    .Q_N(_0053_),
    .Q(\i_soc.cpu.rf.rf[7][10] ));
 sg13g2_dfrbp_1 _3429_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net93),
    .D(_0545_),
    .Q_N(_0052_),
    .Q(\i_soc.cpu.rf.rf[7][11] ));
 sg13g2_dfrbp_1 _3430_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net92),
    .D(_0546_),
    .Q_N(_0051_),
    .Q(\i_soc.cpu.rf.rf[7][12] ));
 sg13g2_dfrbp_1 _3431_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net91),
    .D(_0547_),
    .Q_N(_0050_),
    .Q(\i_soc.cpu.rf.rf[7][13] ));
 sg13g2_dfrbp_1 _3432_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net90),
    .D(_0548_),
    .Q_N(_0049_),
    .Q(\i_soc.cpu.rf.rf[7][14] ));
 sg13g2_dfrbp_1 _3433_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net89),
    .D(_0549_),
    .Q_N(_0048_),
    .Q(\i_soc.cpu.rf.rf[7][15] ));
 sg13g2_dfrbp_1 _3434_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net88),
    .D(_0550_),
    .Q_N(_0047_),
    .Q(\i_soc.cpu.rf.rf[7][16] ));
 sg13g2_dfrbp_1 _3435_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net87),
    .D(_0551_),
    .Q_N(_0046_),
    .Q(\i_soc.cpu.rf.rf[7][17] ));
 sg13g2_dfrbp_1 _3436_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net86),
    .D(_0552_),
    .Q_N(_0045_),
    .Q(\i_soc.cpu.rf.rf[7][18] ));
 sg13g2_dfrbp_1 _3437_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net85),
    .D(_0553_),
    .Q_N(_0044_),
    .Q(\i_soc.cpu.rf.rf[7][19] ));
 sg13g2_dfrbp_1 _3438_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net84),
    .D(_0554_),
    .Q_N(_0043_),
    .Q(\i_soc.cpu.rf.rf[7][20] ));
 sg13g2_dfrbp_1 _3439_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net83),
    .D(net329),
    .Q_N(_0042_),
    .Q(\i_soc.cpu.rf.rf[7][21] ));
 sg13g2_dfrbp_1 _3440_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net82),
    .D(_0556_),
    .Q_N(_0041_),
    .Q(\i_soc.cpu.rf.rf[7][22] ));
 sg13g2_dfrbp_1 _3441_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net81),
    .D(_0557_),
    .Q_N(_0040_),
    .Q(\i_soc.cpu.rf.rf[7][23] ));
 sg13g2_dfrbp_1 _3442_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net80),
    .D(_0558_),
    .Q_N(_0039_),
    .Q(\i_soc.cpu.rf.rf[7][24] ));
 sg13g2_dfrbp_1 _3443_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net79),
    .D(net382),
    .Q_N(_0038_),
    .Q(\i_soc.cpu.rf.rf[7][25] ));
 sg13g2_dfrbp_1 _3444_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net78),
    .D(_0560_),
    .Q_N(_0037_),
    .Q(\i_soc.cpu.rf.rf[7][26] ));
 sg13g2_dfrbp_1 _3445_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net77),
    .D(_0561_),
    .Q_N(_0036_),
    .Q(\i_soc.cpu.rf.rf[7][27] ));
 sg13g2_dfrbp_1 _3446_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net76),
    .D(net340),
    .Q_N(_0035_),
    .Q(\i_soc.cpu.rf.rf[7][28] ));
 sg13g2_dfrbp_1 _3447_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net75),
    .D(_0563_),
    .Q_N(_0034_),
    .Q(\i_soc.cpu.rf.rf[7][29] ));
 sg13g2_dfrbp_1 _3448_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net74),
    .D(_0564_),
    .Q_N(_0033_),
    .Q(\i_soc.cpu.rf.rf[7][30] ));
 sg13g2_dfrbp_1 _3449_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net73),
    .D(_0565_),
    .Q_N(_0032_),
    .Q(\i_soc.cpu.rf.rf[7][31] ));
 sg13g2_dfrbp_1 _3450_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net72),
    .D(_0566_),
    .Q_N(_1578_),
    .Q(\i_soc.pass ));
 sg13g2_dfrbp_1 _3451_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net70),
    .D(_0567_),
    .Q_N(_1577_),
    .Q(fail));
 sg13g2_dfrbp_1 _3452_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net69),
    .D(_0568_),
    .Q_N(_0031_),
    .Q(\i_soc.cpu.rf.rf[6][0] ));
 sg13g2_dfrbp_1 _3453_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net68),
    .D(_0569_),
    .Q_N(_0030_),
    .Q(\i_soc.cpu.rf.rf[6][1] ));
 sg13g2_dfrbp_1 _3454_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net67),
    .D(_0570_),
    .Q_N(_0029_),
    .Q(\i_soc.cpu.rf.rf[6][2] ));
 sg13g2_dfrbp_1 _3455_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net66),
    .D(_0571_),
    .Q_N(_0028_),
    .Q(\i_soc.cpu.rf.rf[6][3] ));
 sg13g2_dfrbp_1 _3456_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net65),
    .D(_0572_),
    .Q_N(_0027_),
    .Q(\i_soc.cpu.rf.rf[6][4] ));
 sg13g2_dfrbp_1 _3457_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net64),
    .D(_0573_),
    .Q_N(_0026_),
    .Q(\i_soc.cpu.rf.rf[6][5] ));
 sg13g2_dfrbp_1 _3458_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net63),
    .D(_0574_),
    .Q_N(_0025_),
    .Q(\i_soc.cpu.rf.rf[6][6] ));
 sg13g2_dfrbp_1 _3459_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net62),
    .D(_0575_),
    .Q_N(_0024_),
    .Q(\i_soc.cpu.rf.rf[6][7] ));
 sg13g2_dfrbp_1 _3460_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net61),
    .D(_0576_),
    .Q_N(_0023_),
    .Q(\i_soc.cpu.rf.rf[6][8] ));
 sg13g2_dfrbp_1 _3461_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net60),
    .D(_0577_),
    .Q_N(_0022_),
    .Q(\i_soc.cpu.rf.rf[6][9] ));
 sg13g2_dfrbp_1 _3462_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net59),
    .D(_0578_),
    .Q_N(_0021_),
    .Q(\i_soc.cpu.rf.rf[6][10] ));
 sg13g2_dfrbp_1 _3463_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net58),
    .D(_0579_),
    .Q_N(_0020_),
    .Q(\i_soc.cpu.rf.rf[6][11] ));
 sg13g2_dfrbp_1 _3464_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net57),
    .D(_0580_),
    .Q_N(_0019_),
    .Q(\i_soc.cpu.rf.rf[6][12] ));
 sg13g2_dfrbp_1 _3465_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net56),
    .D(_0581_),
    .Q_N(_0018_),
    .Q(\i_soc.cpu.rf.rf[6][13] ));
 sg13g2_dfrbp_1 _3466_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net55),
    .D(_0582_),
    .Q_N(_0017_),
    .Q(\i_soc.cpu.rf.rf[6][14] ));
 sg13g2_dfrbp_1 _3467_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net54),
    .D(_0583_),
    .Q_N(_0016_),
    .Q(\i_soc.cpu.rf.rf[6][15] ));
 sg13g2_dfrbp_1 _3468_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net53),
    .D(_0584_),
    .Q_N(_0015_),
    .Q(\i_soc.cpu.rf.rf[6][16] ));
 sg13g2_dfrbp_1 _3469_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net52),
    .D(_0585_),
    .Q_N(_0014_),
    .Q(\i_soc.cpu.rf.rf[6][17] ));
 sg13g2_dfrbp_1 _3470_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net51),
    .D(_0586_),
    .Q_N(_0013_),
    .Q(\i_soc.cpu.rf.rf[6][18] ));
 sg13g2_dfrbp_1 _3471_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net50),
    .D(_0587_),
    .Q_N(_0012_),
    .Q(\i_soc.cpu.rf.rf[6][19] ));
 sg13g2_dfrbp_1 _3472_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net49),
    .D(_0588_),
    .Q_N(_0011_),
    .Q(\i_soc.cpu.rf.rf[6][20] ));
 sg13g2_dfrbp_1 _3473_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net48),
    .D(_0589_),
    .Q_N(_0010_),
    .Q(\i_soc.cpu.rf.rf[6][21] ));
 sg13g2_dfrbp_1 _3474_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net47),
    .D(_0590_),
    .Q_N(_0009_),
    .Q(\i_soc.cpu.rf.rf[6][22] ));
 sg13g2_dfrbp_1 _3475_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net46),
    .D(_0591_),
    .Q_N(_0008_),
    .Q(\i_soc.cpu.rf.rf[6][23] ));
 sg13g2_dfrbp_1 _3476_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net45),
    .D(_0592_),
    .Q_N(_0007_),
    .Q(\i_soc.cpu.rf.rf[6][24] ));
 sg13g2_dfrbp_1 _3477_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net44),
    .D(_0593_),
    .Q_N(_0006_),
    .Q(\i_soc.cpu.rf.rf[6][25] ));
 sg13g2_dfrbp_1 _3478_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net43),
    .D(_0594_),
    .Q_N(_0005_),
    .Q(\i_soc.cpu.rf.rf[6][26] ));
 sg13g2_dfrbp_1 _3479_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net42),
    .D(_0595_),
    .Q_N(_0004_),
    .Q(\i_soc.cpu.rf.rf[6][27] ));
 sg13g2_dfrbp_1 _3480_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net41),
    .D(_0596_),
    .Q_N(_0003_),
    .Q(\i_soc.cpu.rf.rf[6][28] ));
 sg13g2_dfrbp_1 _3481_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net40),
    .D(_0597_),
    .Q_N(_0002_),
    .Q(\i_soc.cpu.rf.rf[6][29] ));
 sg13g2_dfrbp_1 _3482_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net140),
    .D(_0598_),
    .Q_N(_0001_),
    .Q(\i_soc.cpu.rf.rf[6][30] ));
 sg13g2_dfrbp_1 _3483_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net71),
    .D(_0599_),
    .Q_N(_0000_),
    .Q(\i_soc.cpu.rf.rf[6][31] ));
 sg13g2_tiehi _3208__9 (.L_HI(net9));
 sg13g2_tiehi _3207__10 (.L_HI(net10));
 sg13g2_tiehi _3206__11 (.L_HI(net11));
 sg13g2_tiehi _3205__12 (.L_HI(net12));
 sg13g2_tiehi _3204__13 (.L_HI(net13));
 sg13g2_tiehi _3203__14 (.L_HI(net14));
 sg13g2_tiehi _3202__15 (.L_HI(net15));
 sg13g2_tiehi _3201__16 (.L_HI(net16));
 sg13g2_tiehi _3200__17 (.L_HI(net17));
 sg13g2_tiehi _3199__18 (.L_HI(net18));
 sg13g2_tiehi _3198__19 (.L_HI(net19));
 sg13g2_tiehi _3197__20 (.L_HI(net20));
 sg13g2_tiehi _3196__21 (.L_HI(net21));
 sg13g2_tiehi _3195__22 (.L_HI(net22));
 sg13g2_tiehi _3194__23 (.L_HI(net23));
 sg13g2_tiehi _3193__24 (.L_HI(net24));
 sg13g2_tiehi _3192__25 (.L_HI(net25));
 sg13g2_tiehi _3191__26 (.L_HI(net26));
 sg13g2_tiehi _3190__27 (.L_HI(net27));
 sg13g2_tiehi _3189__28 (.L_HI(net28));
 sg13g2_tiehi _3188__29 (.L_HI(net29));
 sg13g2_tiehi _3187__30 (.L_HI(net30));
 sg13g2_tiehi _3186__31 (.L_HI(net31));
 sg13g2_tiehi _3185__32 (.L_HI(net32));
 sg13g2_tiehi _3184__33 (.L_HI(net33));
 sg13g2_tiehi _3183__34 (.L_HI(net34));
 sg13g2_tiehi _3182__35 (.L_HI(net35));
 sg13g2_tiehi _3181__36 (.L_HI(net36));
 sg13g2_tiehi _3180__37 (.L_HI(net37));
 sg13g2_tiehi _3179__38 (.L_HI(net38));
 sg13g2_tiehi _3178__39 (.L_HI(net39));
 sg13g2_tiehi _3481__40 (.L_HI(net40));
 sg13g2_tiehi _3480__41 (.L_HI(net41));
 sg13g2_tiehi _3479__42 (.L_HI(net42));
 sg13g2_tiehi _3478__43 (.L_HI(net43));
 sg13g2_tiehi _3477__44 (.L_HI(net44));
 sg13g2_tiehi _3476__45 (.L_HI(net45));
 sg13g2_tiehi _3475__46 (.L_HI(net46));
 sg13g2_tiehi _3474__47 (.L_HI(net47));
 sg13g2_tiehi _3473__48 (.L_HI(net48));
 sg13g2_tiehi _3472__49 (.L_HI(net49));
 sg13g2_tiehi _3471__50 (.L_HI(net50));
 sg13g2_tiehi _3470__51 (.L_HI(net51));
 sg13g2_tiehi _3469__52 (.L_HI(net52));
 sg13g2_tiehi _3468__53 (.L_HI(net53));
 sg13g2_tiehi _3467__54 (.L_HI(net54));
 sg13g2_tiehi _3466__55 (.L_HI(net55));
 sg13g2_tiehi _3465__56 (.L_HI(net56));
 sg13g2_tiehi _3464__57 (.L_HI(net57));
 sg13g2_tiehi _3463__58 (.L_HI(net58));
 sg13g2_tiehi _3462__59 (.L_HI(net59));
 sg13g2_tiehi _3461__60 (.L_HI(net60));
 sg13g2_tiehi _3460__61 (.L_HI(net61));
 sg13g2_tiehi _3459__62 (.L_HI(net62));
 sg13g2_tiehi _3458__63 (.L_HI(net63));
 sg13g2_tiehi _3457__64 (.L_HI(net64));
 sg13g2_tiehi _3456__65 (.L_HI(net65));
 sg13g2_tiehi _3455__66 (.L_HI(net66));
 sg13g2_tiehi _3454__67 (.L_HI(net67));
 sg13g2_tiehi _3453__68 (.L_HI(net68));
 sg13g2_tiehi _3452__69 (.L_HI(net69));
 sg13g2_tiehi _3451__70 (.L_HI(net70));
 sg13g2_tiehi _3483__71 (.L_HI(net71));
 sg13g2_tiehi _3450__72 (.L_HI(net72));
 sg13g2_tiehi _3449__73 (.L_HI(net73));
 sg13g2_tiehi _3448__74 (.L_HI(net74));
 sg13g2_tiehi _3447__75 (.L_HI(net75));
 sg13g2_tiehi _3446__76 (.L_HI(net76));
 sg13g2_tiehi _3445__77 (.L_HI(net77));
 sg13g2_tiehi _3444__78 (.L_HI(net78));
 sg13g2_tiehi _3443__79 (.L_HI(net79));
 sg13g2_tiehi _3442__80 (.L_HI(net80));
 sg13g2_tiehi _3441__81 (.L_HI(net81));
 sg13g2_tiehi _3440__82 (.L_HI(net82));
 sg13g2_tiehi _3439__83 (.L_HI(net83));
 sg13g2_tiehi _3438__84 (.L_HI(net84));
 sg13g2_tiehi _3437__85 (.L_HI(net85));
 sg13g2_tiehi _3436__86 (.L_HI(net86));
 sg13g2_tiehi _3435__87 (.L_HI(net87));
 sg13g2_tiehi _3434__88 (.L_HI(net88));
 sg13g2_tiehi _3433__89 (.L_HI(net89));
 sg13g2_tiehi _3432__90 (.L_HI(net90));
 sg13g2_tiehi _3431__91 (.L_HI(net91));
 sg13g2_tiehi _3430__92 (.L_HI(net92));
 sg13g2_tiehi _3429__93 (.L_HI(net93));
 sg13g2_tiehi _3428__94 (.L_HI(net94));
 sg13g2_tiehi _3427__95 (.L_HI(net95));
 sg13g2_tiehi _3426__96 (.L_HI(net96));
 sg13g2_tiehi _3425__97 (.L_HI(net97));
 sg13g2_tiehi _3424__98 (.L_HI(net98));
 sg13g2_tiehi _3423__99 (.L_HI(net99));
 sg13g2_tiehi _3422__100 (.L_HI(net100));
 sg13g2_tiehi _3421__101 (.L_HI(net101));
 sg13g2_tiehi _3420__102 (.L_HI(net102));
 sg13g2_tiehi _3419__103 (.L_HI(net103));
 sg13g2_tiehi _3418__104 (.L_HI(net104));
 sg13g2_tiehi _3417__105 (.L_HI(net105));
 sg13g2_tiehi _3416__106 (.L_HI(net106));
 sg13g2_tiehi _3415__107 (.L_HI(net107));
 sg13g2_tiehi _3414__108 (.L_HI(net108));
 sg13g2_tiehi _3413__109 (.L_HI(net109));
 sg13g2_tiehi _3412__110 (.L_HI(net110));
 sg13g2_tiehi _3411__111 (.L_HI(net111));
 sg13g2_tiehi _3410__112 (.L_HI(net112));
 sg13g2_tiehi _3409__113 (.L_HI(net113));
 sg13g2_tiehi _3408__114 (.L_HI(net114));
 sg13g2_tiehi _3407__115 (.L_HI(net115));
 sg13g2_tiehi _3406__116 (.L_HI(net116));
 sg13g2_tiehi _3405__117 (.L_HI(net117));
 sg13g2_tiehi _3404__118 (.L_HI(net118));
 sg13g2_tiehi _3403__119 (.L_HI(net119));
 sg13g2_tiehi _3402__120 (.L_HI(net120));
 sg13g2_tiehi _3401__121 (.L_HI(net121));
 sg13g2_tiehi _3400__122 (.L_HI(net122));
 sg13g2_tiehi _3399__123 (.L_HI(net123));
 sg13g2_tiehi _3398__124 (.L_HI(net124));
 sg13g2_tiehi _3397__125 (.L_HI(net125));
 sg13g2_tiehi _3396__126 (.L_HI(net126));
 sg13g2_tiehi _3395__127 (.L_HI(net127));
 sg13g2_tiehi _3394__128 (.L_HI(net128));
 sg13g2_tiehi _3393__129 (.L_HI(net129));
 sg13g2_tiehi _3392__130 (.L_HI(net130));
 sg13g2_tiehi _3391__131 (.L_HI(net131));
 sg13g2_tiehi _3390__132 (.L_HI(net132));
 sg13g2_tiehi _3389__133 (.L_HI(net133));
 sg13g2_tiehi _3388__134 (.L_HI(net134));
 sg13g2_tiehi _3387__135 (.L_HI(net135));
 sg13g2_tiehi _3386__136 (.L_HI(net136));
 sg13g2_tiehi _3385__137 (.L_HI(net137));
 sg13g2_tiehi _3384__138 (.L_HI(net138));
 sg13g2_tiehi _3383__139 (.L_HI(net139));
 sg13g2_tiehi _3482__140 (.L_HI(net140));
 sg13g2_tiehi _3382__141 (.L_HI(net141));
 sg13g2_tiehi _3381__142 (.L_HI(net142));
 sg13g2_tiehi _3380__143 (.L_HI(net143));
 sg13g2_tiehi _3379__144 (.L_HI(net144));
 sg13g2_tiehi _3378__145 (.L_HI(net145));
 sg13g2_tiehi _3377__146 (.L_HI(net146));
 sg13g2_tiehi _3376__147 (.L_HI(net147));
 sg13g2_tiehi _3375__148 (.L_HI(net148));
 sg13g2_tiehi _3374__149 (.L_HI(net149));
 sg13g2_tiehi _3373__150 (.L_HI(net150));
 sg13g2_tiehi _3372__151 (.L_HI(net151));
 sg13g2_tiehi _3371__152 (.L_HI(net152));
 sg13g2_tiehi _3370__153 (.L_HI(net153));
 sg13g2_tiehi _3369__154 (.L_HI(net154));
 sg13g2_tiehi _3368__155 (.L_HI(net155));
 sg13g2_tiehi _3367__156 (.L_HI(net156));
 sg13g2_tiehi _3366__157 (.L_HI(net157));
 sg13g2_tiehi _3365__158 (.L_HI(net158));
 sg13g2_tiehi _3364__159 (.L_HI(net159));
 sg13g2_tiehi _3363__160 (.L_HI(net160));
 sg13g2_tiehi _3362__161 (.L_HI(net161));
 sg13g2_tiehi _3361__162 (.L_HI(net162));
 sg13g2_tiehi _3360__163 (.L_HI(net163));
 sg13g2_tiehi _3359__164 (.L_HI(net164));
 sg13g2_tiehi _3358__165 (.L_HI(net165));
 sg13g2_tiehi _3357__166 (.L_HI(net166));
 sg13g2_tiehi _3356__167 (.L_HI(net167));
 sg13g2_tiehi _3355__168 (.L_HI(net168));
 sg13g2_tiehi _3354__169 (.L_HI(net169));
 sg13g2_tiehi _3353__170 (.L_HI(net170));
 sg13g2_tiehi _3352__171 (.L_HI(net171));
 sg13g2_tiehi _3351__172 (.L_HI(net172));
 sg13g2_tiehi _3350__173 (.L_HI(net173));
 sg13g2_tiehi _3349__174 (.L_HI(net174));
 sg13g2_tiehi _3348__175 (.L_HI(net175));
 sg13g2_tiehi _3347__176 (.L_HI(net176));
 sg13g2_tiehi _3346__177 (.L_HI(net177));
 sg13g2_tiehi _3345__178 (.L_HI(net178));
 sg13g2_tiehi _3344__179 (.L_HI(net179));
 sg13g2_tiehi _3343__180 (.L_HI(net180));
 sg13g2_tiehi _3342__181 (.L_HI(net181));
 sg13g2_tiehi _3341__182 (.L_HI(net182));
 sg13g2_tiehi _3340__183 (.L_HI(net183));
 sg13g2_tiehi _3339__184 (.L_HI(net184));
 sg13g2_tiehi _3338__185 (.L_HI(net185));
 sg13g2_tiehi _3337__186 (.L_HI(net186));
 sg13g2_tiehi _3336__187 (.L_HI(net187));
 sg13g2_tiehi _3335__188 (.L_HI(net188));
 sg13g2_tiehi _3334__189 (.L_HI(net189));
 sg13g2_tiehi _3333__190 (.L_HI(net190));
 sg13g2_tiehi _3332__191 (.L_HI(net191));
 sg13g2_tiehi _3331__192 (.L_HI(net192));
 sg13g2_tiehi _3330__193 (.L_HI(net193));
 sg13g2_tiehi _3329__194 (.L_HI(net194));
 sg13g2_tiehi _3328__195 (.L_HI(net195));
 sg13g2_tiehi _3327__196 (.L_HI(net196));
 sg13g2_tiehi _3326__197 (.L_HI(net197));
 sg13g2_tiehi _3325__198 (.L_HI(net198));
 sg13g2_tiehi _3324__199 (.L_HI(net199));
 sg13g2_tiehi _3323__200 (.L_HI(net200));
 sg13g2_tiehi _3322__201 (.L_HI(net201));
 sg13g2_tiehi _3321__202 (.L_HI(net202));
 sg13g2_tiehi _3320__203 (.L_HI(net203));
 sg13g2_tiehi _3319__204 (.L_HI(net204));
 sg13g2_tiehi _3318__205 (.L_HI(net205));
 sg13g2_tiehi _3317__206 (.L_HI(net206));
 sg13g2_tiehi _3316__207 (.L_HI(net207));
 sg13g2_tiehi _3315__208 (.L_HI(net208));
 sg13g2_tiehi _3314__209 (.L_HI(net209));
 sg13g2_tiehi _3313__210 (.L_HI(net210));
 sg13g2_tiehi _3312__211 (.L_HI(net211));
 sg13g2_tiehi _3311__212 (.L_HI(net212));
 sg13g2_tiehi _3310__213 (.L_HI(net213));
 sg13g2_tiehi _3309__214 (.L_HI(net214));
 sg13g2_tiehi _3308__215 (.L_HI(net215));
 sg13g2_tiehi _3307__216 (.L_HI(net216));
 sg13g2_tiehi _3306__217 (.L_HI(net217));
 sg13g2_tiehi _3305__218 (.L_HI(net218));
 sg13g2_tiehi _3304__219 (.L_HI(net219));
 sg13g2_tiehi _3303__220 (.L_HI(net220));
 sg13g2_tiehi _3302__221 (.L_HI(net221));
 sg13g2_tiehi _3301__222 (.L_HI(net222));
 sg13g2_tiehi _3300__223 (.L_HI(net223));
 sg13g2_tiehi _3299__224 (.L_HI(net224));
 sg13g2_tiehi _3298__225 (.L_HI(net225));
 sg13g2_tiehi _3297__226 (.L_HI(net226));
 sg13g2_tiehi _3296__227 (.L_HI(net227));
 sg13g2_tiehi _3295__228 (.L_HI(net228));
 sg13g2_tiehi _3294__229 (.L_HI(net229));
 sg13g2_tiehi _3293__230 (.L_HI(net230));
 sg13g2_tiehi _3292__231 (.L_HI(net231));
 sg13g2_tiehi _3291__232 (.L_HI(net232));
 sg13g2_tiehi _3290__233 (.L_HI(net233));
 sg13g2_tiehi _3289__234 (.L_HI(net234));
 sg13g2_tiehi _3288__235 (.L_HI(net235));
 sg13g2_tiehi _3287__236 (.L_HI(net236));
 sg13g2_tiehi _3286__237 (.L_HI(net237));
 sg13g2_tiehi _3285__238 (.L_HI(net238));
 sg13g2_tiehi _3284__239 (.L_HI(net239));
 sg13g2_tiehi _3283__240 (.L_HI(net240));
 sg13g2_tiehi _3282__241 (.L_HI(net241));
 sg13g2_tiehi _3281__242 (.L_HI(net242));
 sg13g2_tiehi _3280__243 (.L_HI(net243));
 sg13g2_tiehi _3279__244 (.L_HI(net244));
 sg13g2_tiehi _3278__245 (.L_HI(net245));
 sg13g2_tiehi _3277__246 (.L_HI(net246));
 sg13g2_tiehi _3276__247 (.L_HI(net247));
 sg13g2_tiehi _3275__248 (.L_HI(net248));
 sg13g2_tiehi _3274__249 (.L_HI(net249));
 sg13g2_tiehi _3273__250 (.L_HI(net250));
 sg13g2_tiehi _3272__251 (.L_HI(net251));
 sg13g2_tiehi _3271__252 (.L_HI(net252));
 sg13g2_tiehi _3270__253 (.L_HI(net253));
 sg13g2_tiehi _3269__254 (.L_HI(net254));
 sg13g2_tiehi _3268__255 (.L_HI(net255));
 sg13g2_tiehi _3267__256 (.L_HI(net256));
 sg13g2_tiehi _3266__257 (.L_HI(net257));
 sg13g2_tiehi _3265__258 (.L_HI(net258));
 sg13g2_tiehi _3264__259 (.L_HI(net259));
 sg13g2_tiehi _3263__260 (.L_HI(net260));
 sg13g2_tiehi _3262__261 (.L_HI(net261));
 sg13g2_tiehi _3261__262 (.L_HI(net262));
 sg13g2_tiehi _3260__263 (.L_HI(net263));
 sg13g2_tiehi _3259__264 (.L_HI(net264));
 sg13g2_tiehi _3258__265 (.L_HI(net265));
 sg13g2_tiehi _3257__266 (.L_HI(net266));
 sg13g2_tiehi _3256__267 (.L_HI(net267));
 sg13g2_tiehi _3255__268 (.L_HI(net268));
 sg13g2_tiehi _3254__269 (.L_HI(net269));
 sg13g2_tiehi _3253__270 (.L_HI(net270));
 sg13g2_tiehi _3252__271 (.L_HI(net271));
 sg13g2_tiehi _3251__272 (.L_HI(net272));
 sg13g2_tiehi _3250__273 (.L_HI(net273));
 sg13g2_tiehi _3249__274 (.L_HI(net274));
 sg13g2_tiehi _3248__275 (.L_HI(net275));
 sg13g2_tiehi _3247__276 (.L_HI(net276));
 sg13g2_tiehi _3246__277 (.L_HI(net277));
 sg13g2_tiehi _3245__278 (.L_HI(net278));
 sg13g2_tiehi _3244__279 (.L_HI(net279));
 sg13g2_tiehi _3243__280 (.L_HI(net280));
 sg13g2_tiehi _3242__281 (.L_HI(net281));
 sg13g2_tiehi _3241__282 (.L_HI(net282));
 sg13g2_tiehi _3240__283 (.L_HI(net283));
 sg13g2_tiehi _3239__284 (.L_HI(net284));
 sg13g2_tiehi _3238__285 (.L_HI(net285));
 sg13g2_tiehi _3237__286 (.L_HI(net286));
 sg13g2_tiehi _3236__287 (.L_HI(net287));
 sg13g2_tiehi _3235__288 (.L_HI(net288));
 sg13g2_tiehi _3234__289 (.L_HI(net289));
 sg13g2_tiehi _3233__290 (.L_HI(net290));
 sg13g2_tiehi _3232__291 (.L_HI(net291));
 sg13g2_tiehi _3231__292 (.L_HI(net292));
 sg13g2_tiehi _3230__293 (.L_HI(net293));
 sg13g2_tiehi _3229__294 (.L_HI(net294));
 sg13g2_tiehi _3228__295 (.L_HI(net295));
 sg13g2_tiehi _3227__296 (.L_HI(net296));
 sg13g2_tiehi _3226__297 (.L_HI(net297));
 sg13g2_tiehi _3225__298 (.L_HI(net298));
 sg13g2_tiehi _3224__299 (.L_HI(net299));
 sg13g2_tiehi _3223__300 (.L_HI(net300));
 sg13g2_tiehi _3222__301 (.L_HI(net301));
 sg13g2_tiehi _3221__302 (.L_HI(net302));
 sg13g2_tiehi _3220__303 (.L_HI(net303));
 sg13g2_tiehi _3219__304 (.L_HI(net304));
 sg13g2_tiehi _3218__305 (.L_HI(net305));
 sg13g2_tiehi _3217__306 (.L_HI(net306));
 sg13g2_tiehi _3216__307 (.L_HI(net307));
 sg13g2_tiehi _3215__308 (.L_HI(net308));
 sg13g2_tiehi _3214__309 (.L_HI(net309));
 sg13g2_tiehi _3213__310 (.L_HI(net310));
 sg13g2_tiehi _3212__311 (.L_HI(net311));
 sg13g2_tiehi _3211__312 (.L_HI(net312));
 sg13g2_tiehi _3210__313 (.L_HI(net313));
 sg13g2_tiehi tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_314 (.L_HI(net314));
 sg13g2_tiehi tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_315 (.L_HI(net315));
 sg13g2_tiehi tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_316 (.L_HI(net316));
 sg13g2_tiehi tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_317 (.L_HI(net317));
 sg13g2_tiehi tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_318 (.L_HI(net318));
 sg13g2_tiehi tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_319 (.L_HI(net319));
 sg13g2_tiehi tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_320 (.L_HI(net320));
 sg13g2_tiehi tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_321 (.L_HI(net321));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_3 (.L_LO(net3));
 sg13g2_tielo tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_4 (.L_LO(net4));
 sg13g2_tielo tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_5 (.L_LO(net5));
 sg13g2_tielo tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_6 (.L_LO(net6));
 sg13g2_tielo tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_7 (.L_LO(net7));
 sg13g2_tiehi _3209__8 (.L_HI(net8));
 sg13g2_buf_2 _3804_ (.A(\i_soc.cpu.rd0[0] ),
    .X(uio_out[0]));
 sg13g2_buf_1 _3805_ (.A(\i_soc.cpu.rd0[1] ),
    .X(uio_out[1]));
 sg13g2_buf_2 _3806_ (.A(\i_soc.cpu.rd0[2] ),
    .X(uio_out[2]));
 sg13g2_buf_1 _3807_ (.A(\i_soc.cpu.rd0[3] ),
    .X(uio_out[3]));
 sg13g2_buf_1 _3808_ (.A(net610),
    .X(uio_out[4]));
 sg13g2_buf_1 _3809_ (.A(\i_soc.cpu.pc[3] ),
    .X(uio_out[5]));
 sg13g2_buf_1 _3810_ (.A(net607),
    .X(uio_out[6]));
 sg13g2_buf_1 _3811_ (.A(net604),
    .X(uio_out[7]));
 sg13g2_buf_1 _3812_ (.A(\i_soc.pass ),
    .X(uo_out[0]));
 sg13g2_buf_1 _3813_ (.A(fail),
    .X(uo_out[1]));
 sg13g2_buf_2 fanout459 (.A(net463),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(net463),
    .X(net460));
 sg13g2_buf_4 fanout461 (.X(net461),
    .A(net463));
 sg13g2_buf_2 fanout462 (.A(net463),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_1448_),
    .X(net463));
 sg13g2_buf_4 fanout464 (.X(net464),
    .A(net465));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(net468));
 sg13g2_buf_4 fanout466 (.X(net466),
    .A(net467));
 sg13g2_buf_2 fanout467 (.A(net468),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_1448_),
    .X(net468));
 sg13g2_buf_4 fanout469 (.X(net469),
    .A(net473));
 sg13g2_buf_4 fanout470 (.X(net470),
    .A(net473));
 sg13g2_buf_4 fanout471 (.X(net471),
    .A(net473));
 sg13g2_buf_2 fanout472 (.A(net473),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(_0683_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net478),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(net478),
    .X(net475));
 sg13g2_buf_4 fanout476 (.X(net476),
    .A(net478));
 sg13g2_buf_2 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_4 fanout478 (.X(net478),
    .A(_1544_));
 sg13g2_buf_4 fanout479 (.X(net479),
    .A(net483));
 sg13g2_buf_2 fanout480 (.A(net483),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(net482),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(net483),
    .X(net482));
 sg13g2_buf_4 fanout483 (.X(net483),
    .A(_1544_));
 sg13g2_buf_4 fanout484 (.X(net484),
    .A(_0672_));
 sg13g2_buf_4 fanout485 (.X(net485),
    .A(_0672_));
 sg13g2_buf_4 fanout486 (.X(net486),
    .A(net494));
 sg13g2_buf_2 fanout487 (.A(net494),
    .X(net487));
 sg13g2_buf_4 fanout488 (.X(net488),
    .A(net490));
 sg13g2_buf_1 fanout489 (.A(net490),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(net494),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(net493),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(net493),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(net494),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_0671_),
    .X(net494));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(net497));
 sg13g2_buf_2 fanout496 (.A(net497),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_0663_),
    .X(net497));
 sg13g2_buf_4 fanout498 (.X(net498),
    .A(_0663_));
 sg13g2_buf_2 fanout499 (.A(_0663_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(net501),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(net504),
    .X(net501));
 sg13g2_buf_4 fanout502 (.X(net502),
    .A(net504));
 sg13g2_buf_1 fanout503 (.A(net504),
    .X(net503));
 sg13g2_buf_4 fanout504 (.X(net504),
    .A(_1497_));
 sg13g2_buf_2 fanout505 (.A(net509),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(net509),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(net508),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_1497_),
    .X(net509));
 sg13g2_buf_4 fanout510 (.X(net510),
    .A(net512));
 sg13g2_buf_2 fanout511 (.A(net512),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_0676_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(net515),
    .X(net513));
 sg13g2_buf_4 fanout514 (.X(net514),
    .A(net515));
 sg13g2_buf_2 fanout515 (.A(_0676_),
    .X(net515));
 sg13g2_buf_4 fanout516 (.X(net516),
    .A(net520));
 sg13g2_buf_2 fanout517 (.A(net520),
    .X(net517));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(net520));
 sg13g2_buf_2 fanout519 (.A(net520),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_0675_),
    .X(net520));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(net529));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(net529));
 sg13g2_buf_2 fanout523 (.A(net524),
    .X(net523));
 sg13g2_buf_4 fanout524 (.X(net524),
    .A(net529));
 sg13g2_buf_2 fanout525 (.A(net526),
    .X(net525));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(net528));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(net529),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_0669_),
    .X(net529));
 sg13g2_buf_4 fanout530 (.X(net530),
    .A(net539));
 sg13g2_buf_2 fanout531 (.A(net539),
    .X(net531));
 sg13g2_buf_4 fanout532 (.X(net532),
    .A(net533));
 sg13g2_buf_2 fanout533 (.A(net539),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net535),
    .X(net534));
 sg13g2_buf_4 fanout535 (.X(net535),
    .A(net538));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(net538));
 sg13g2_buf_1 fanout537 (.A(net538),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(net539),
    .X(net538));
 sg13g2_buf_4 fanout539 (.X(net539),
    .A(_0668_));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(net542));
 sg13g2_buf_2 fanout541 (.A(net542),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(net546),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(net546),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(net546),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net546),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_0655_),
    .X(net546));
 sg13g2_buf_4 fanout547 (.X(net547),
    .A(net549));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(net549));
 sg13g2_buf_4 fanout549 (.X(net549),
    .A(_0654_));
 sg13g2_buf_4 fanout550 (.X(net550),
    .A(net551));
 sg13g2_buf_8 fanout551 (.A(net554),
    .X(net551));
 sg13g2_buf_8 fanout552 (.A(net553),
    .X(net552));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(net554));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(_0648_));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(_0647_));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(_0647_));
 sg13g2_buf_8 fanout557 (.A(net559),
    .X(net557));
 sg13g2_buf_8 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_4 fanout559 (.X(net559),
    .A(net562));
 sg13g2_buf_4 fanout560 (.X(net560),
    .A(net561));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(net562));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(_0642_));
 sg13g2_buf_4 fanout563 (.X(net563),
    .A(net568));
 sg13g2_buf_2 fanout564 (.A(net568),
    .X(net564));
 sg13g2_buf_4 fanout565 (.X(net565),
    .A(net567));
 sg13g2_buf_4 fanout566 (.X(net566),
    .A(net568));
 sg13g2_buf_1 fanout567 (.A(net568),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_0641_),
    .X(net568));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(net570));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(_0666_));
 sg13g2_buf_4 fanout571 (.X(net571),
    .A(net572));
 sg13g2_buf_4 fanout572 (.X(net572),
    .A(_0624_));
 sg13g2_buf_4 fanout573 (.X(net573),
    .A(net576));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(net576));
 sg13g2_buf_2 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_0623_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(net583),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(net581),
    .X(net579));
 sg13g2_buf_1 fanout580 (.A(net581),
    .X(net580));
 sg13g2_buf_1 fanout581 (.A(net583),
    .X(net581));
 sg13g2_buf_4 fanout582 (.X(net582),
    .A(net583));
 sg13g2_buf_2 fanout583 (.A(_0619_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(net587),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(net586),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(net587),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_0619_),
    .X(net587));
 sg13g2_buf_4 fanout588 (.X(net588),
    .A(net590));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(net590));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(_0615_));
 sg13g2_buf_2 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_4 fanout592 (.X(net592),
    .A(net596));
 sg13g2_buf_2 fanout593 (.A(net595),
    .X(net593));
 sg13g2_buf_1 fanout594 (.A(net595),
    .X(net594));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(net596));
 sg13g2_buf_2 fanout596 (.A(_0632_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(net598),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(net601),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(net600),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(net601),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_0632_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(net604),
    .X(net603));
 sg13g2_buf_1 fanout604 (.A(net788),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(net606),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_1 fanout607 (.A(\i_soc.cpu.pc[4] ),
    .X(net607));
 sg13g2_buf_4 fanout608 (.X(net608),
    .A(\i_soc.cpu.pc[3] ));
 sg13g2_buf_4 fanout609 (.X(net609),
    .A(net610));
 sg13g2_buf_2 fanout610 (.A(\i_soc.cpu.pc[2] ),
    .X(net610));
 sg13g2_buf_4 fanout611 (.X(net611),
    .A(net1));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_tielo tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload0 (.A(clknet_leaf_39_clk));
 sg13g2_inv_4 clkload1 (.A(clknet_leaf_24_clk));
 sg13g2_inv_4 clkload2 (.A(clknet_leaf_14_clk));
 sg13g2_inv_2 clkload3 (.A(clknet_leaf_23_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0096_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0095_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold3 (.A(\i_soc.cpu.rf.rf[27][11] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold4 (.A(\i_soc.cpu.rf.rf[11][31] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold5 (.A(\i_soc.cpu.rf.rf[8][31] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold6 (.A(\i_soc.cpu.rf.rf[8][2] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0042_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0555_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold9 (.A(\i_soc.cpu.rf.rf[1][0] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold10 (.A(\i_soc.cpu.rf.rf[27][8] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold11 (.A(\i_soc.cpu.rf.rf[1][6] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold12 (.A(\i_soc.cpu.rf.rf[11][13] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold13 (.A(\i_soc.cpu.rf.rf[8][30] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_soc.cpu.rf.rf[8][15] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold15 (.A(\i_soc.cpu.rf.rf[3][10] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold16 (.A(\i_soc.cpu.rf.rf[11][11] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold17 (.A(\i_soc.cpu.rf.rf[8][10] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0035_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0562_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_soc.cpu.rf.rf[11][21] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold21 (.A(\i_soc.cpu.rf.rf[27][22] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold22 (.A(\i_soc.cpu.rf.rf[11][1] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold23 (.A(\i_soc.cpu.rf.rf[11][3] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold24 (.A(\i_soc.cpu.rf.rf[8][0] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold25 (.A(\i_soc.cpu.rf.rf[27][31] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold26 (.A(\i_soc.cpu.rf.rf[8][3] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold27 (.A(\i_soc.cpu.rf.rf[3][3] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold28 (.A(\i_soc.cpu.rf.rf[0][1] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold29 (.A(\i_soc.cpu.rf.rf[27][3] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i_soc.cpu.rf.rf[27][2] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold31 (.A(\i_soc.cpu.rf.rf[27][1] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_soc.cpu.rf.rf[0][3] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold33 (.A(\i_soc.cpu.rf.rf[11][0] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold34 (.A(\i_soc.cpu.rf.rf[8][6] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold35 (.A(\i_soc.cpu.rf.rf[11][5] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold36 (.A(\i_soc.cpu.rf.rf[1][7] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold37 (.A(\i_soc.cpu.rf.rf[27][7] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold38 (.A(\i_soc.cpu.rf.rf[8][7] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold39 (.A(\i_soc.cpu.rf.rf[8][20] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold40 (.A(\i_soc.cpu.rf.rf[8][18] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold41 (.A(\i_soc.cpu.rf.rf[8][25] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold42 (.A(\i_soc.cpu.rf.rf[11][24] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold43 (.A(\i_soc.cpu.rf.rf[11][25] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold44 (.A(\i_soc.cpu.rf.rf[11][26] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold45 (.A(\i_soc.cpu.rf.rf[1][19] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold46 (.A(\i_soc.cpu.rf.rf[3][19] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold47 (.A(\i_soc.cpu.rf.rf[3][18] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold48 (.A(\i_soc.cpu.rf.rf[1][18] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold49 (.A(\i_soc.cpu.rf.rf[11][9] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold50 (.A(\i_soc.cpu.rf.rf[8][21] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold51 (.A(\i_soc.cpu.rf.rf[11][20] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold52 (.A(\i_soc.cpu.rf.rf[8][17] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold53 (.A(\i_soc.cpu.rf.rf[3][16] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold54 (.A(\i_soc.cpu.rf.rf[27][17] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold55 (.A(\i_soc.cpu.rf.rf[8][16] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold56 (.A(\i_soc.cpu.rf.rf[8][26] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold57 (.A(\i_soc.cpu.rf.rf[1][25] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold58 (.A(\i_soc.cpu.rf.rf[27][25] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold59 (.A(\i_soc.cpu.rf.rf[27][19] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0038_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0559_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold62 (.A(\i_soc.cpu.rf.rf[11][16] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold63 (.A(\i_soc.cpu.rf.rf[11][2] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold64 (.A(\i_soc.cpu.rf.rf[27][6] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold65 (.A(\i_soc.cpu.rf.rf[27][4] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold66 (.A(\i_soc.cpu.rf.rf[3][2] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold67 (.A(\i_soc.cpu.rf.rf[8][4] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold68 (.A(\i_soc.cpu.rf.rf[11][7] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold69 (.A(\i_soc.cpu.rf.rf[3][8] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_soc.cpu.rf.rf[27][0] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold71 (.A(\i_soc.cpu.rf.rf[3][24] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold72 (.A(\i_soc.cpu.rf.rf[3][26] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold73 (.A(\i_soc.cpu.rf.rf[1][24] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold74 (.A(\i_soc.cpu.rf.rf[0][0] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold75 (.A(\i_soc.cpu.rf.rf[3][1] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold76 (.A(\i_soc.cpu.rf.rf[1][26] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold77 (.A(\i_soc.cpu.rf.rf[8][9] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold78 (.A(\i_soc.cpu.rf.rf[1][30] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold79 (.A(\i_soc.cpu.rf.rf[27][9] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold80 (.A(\i_soc.cpu.rf.rf[3][28] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold81 (.A(\i_soc.cpu.rf.rf[0][30] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_soc.cpu.rf.rf[11][28] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold83 (.A(\i_soc.cpu.rf.rf[11][19] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold84 (.A(\i_soc.cpu.rf.rf[3][5] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold85 (.A(\i_soc.cpu.rf.rf[1][8] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold86 (.A(\i_soc.cpu.rf.rf[3][7] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold87 (.A(\i_soc.cpu.rf.rf[1][21] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold88 (.A(\i_soc.cpu.rf.rf[11][12] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold89 (.A(\i_soc.cpu.rf.rf[8][14] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold90 (.A(\i_soc.cpu.rf.rf[1][14] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold91 (.A(\i_soc.cpu.rf.rf[8][5] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold92 (.A(\i_soc.cpu.rf.rf[11][4] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold93 (.A(\i_soc.cpu.rf.rf[1][28] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold94 (.A(\i_soc.cpu.rf.rf[11][15] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold95 (.A(\i_soc.cpu.rf.rf[3][15] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold96 (.A(\i_soc.cpu.rf.rf[27][15] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold97 (.A(\i_soc.cpu.rf.rf[1][11] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold98 (.A(\i_soc.cpu.rf.rf[8][13] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_soc.cpu.rf.rf[11][14] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold100 (.A(\i_soc.cpu.rf.rf[0][2] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold101 (.A(\i_soc.cpu.rf.rf[1][5] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold102 (.A(\i_soc.cpu.rf.rf[8][12] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold103 (.A(\i_soc.cpu.rf.rf[1][4] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold104 (.A(\i_soc.cpu.rf.rf[3][13] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold105 (.A(\i_soc.cpu.rf.rf[1][13] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold106 (.A(\i_soc.cpu.rf.rf[3][30] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold107 (.A(\i_soc.cpu.rf.rf[27][16] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold108 (.A(\i_soc.cpu.rf.rf[11][10] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold109 (.A(\i_soc.cpu.rf.rf[11][30] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold110 (.A(\i_soc.cpu.rf.rf[1][23] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold111 (.A(\i_soc.cpu.rf.rf[3][23] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold112 (.A(\i_soc.cpu.rf.rf[1][16] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold113 (.A(\i_soc.cpu.rf.rf[3][17] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold114 (.A(\i_soc.cpu.rf.rf[3][12] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold115 (.A(\i_soc.cpu.rf.rf[3][29] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold116 (.A(\i_soc.cpu.rf.rf[8][24] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold117 (.A(\i_soc.cpu.rf.rf[3][25] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_soc.cpu.rf.rf[8][23] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold119 (.A(\i_soc.cpu.rf.rf[27][10] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold120 (.A(\i_soc.cpu.rf.rf[27][30] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold121 (.A(\i_soc.cpu.rf.rf[27][13] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold122 (.A(\i_soc.cpu.rf.rf[1][27] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold123 (.A(\i_soc.cpu.rf.rf[27][14] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold124 (.A(\i_soc.cpu.rf.rf[8][29] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold125 (.A(\i_soc.cpu.rf.rf[1][22] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold126 (.A(\i_soc.cpu.rf.rf[1][20] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold127 (.A(\i_soc.cpu.rf.rf[8][22] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold128 (.A(\i_soc.cpu.rf.rf[27][12] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold129 (.A(\i_soc.cpu.rf.rf[1][17] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold130 (.A(\i_soc.cpu.rf.rf[11][8] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold131 (.A(\i_soc.cpu.rf.rf[3][14] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold132 (.A(\i_soc.cpu.rf.rf[1][29] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold133 (.A(\i_soc.cpu.rf.rf[11][22] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold134 (.A(\i_soc.cpu.rf.rf[27][26] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold135 (.A(\i_soc.cpu.rf.rf[27][24] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold136 (.A(\i_soc.cpu.rf.rf[1][12] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold137 (.A(\i_soc.cpu.rf.rf[27][23] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold138 (.A(\i_soc.cpu.rf.rf[3][31] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold139 (.A(\i_soc.cpu.rf.rf[1][10] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold140 (.A(\i_soc.cpu.rf.rf[8][11] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold141 (.A(\i_soc.cpu.rf.rf[1][31] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold142 (.A(\i_soc.cpu.rf.rf[11][29] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold143 (.A(\i_soc.cpu.rf.rf[27][29] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold144 (.A(\i_soc.cpu.rf.rf[27][28] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold145 (.A(\i_soc.cpu.rf.rf[3][4] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold146 (.A(\i_soc.cpu.rf.rf[27][5] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold147 (.A(\i_soc.cpu.rf.rf[27][20] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold148 (.A(\i_soc.cpu.rf.rf[3][6] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold149 (.A(\i_soc.cpu.rf.rf[3][27] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold150 (.A(\i_soc.cpu.rf.rf[8][1] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_soc.cpu.rf.rf[3][11] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold152 (.A(\i_soc.cpu.rf.rf[3][21] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold153 (.A(\i_soc.cpu.rf.rf[1][3] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold154 (.A(\i_soc.cpu.rf.rf[11][27] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold155 (.A(\i_soc.cpu.rf.rf[11][6] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold156 (.A(\i_soc.cpu.rf.rf[1][15] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold157 (.A(\i_soc.cpu.rf.rf[1][1] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold158 (.A(\i_soc.cpu.rf.rf[8][28] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold159 (.A(\i_soc.cpu.rf.rf[27][21] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold160 (.A(\i_soc.cpu.rf.rf[11][18] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold161 (.A(\i_soc.cpu.rf.rf[27][18] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold162 (.A(\i_soc.cpu.rf.rf[3][0] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold163 (.A(\i_soc.cpu.rf.rf[1][2] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold164 (.A(\i_soc.cpu.rf.rf[11][17] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold165 (.A(\i_soc.cpu.rf.rf[8][8] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold166 (.A(\i_soc.cpu.rf.rf[3][20] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold167 (.A(\i_soc.cpu.rf.rf[3][22] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold168 (.A(\i_soc.cpu.rf.rf[8][27] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold169 (.A(\i_soc.cpu.rf.rf[1][9] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold170 (.A(\i_soc.cpu.rf.rf[27][27] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold171 (.A(\i_soc.cpu.rf.rf[3][9] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold172 (.A(\i_soc.cpu.rf.rf[8][19] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold173 (.A(\i_soc.cpu.rf.rf[6][15] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold174 (.A(\i_soc.cpu.rf.rf[7][0] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold175 (.A(\i_soc.cpu.rf.rf[5][14] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold176 (.A(\i_soc.cpu.rf.rf[6][19] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold177 (.A(\i_soc.cpu.rf.rf[7][13] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold178 (.A(\i_soc.cpu.rf.rf[5][7] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold179 (.A(\i_soc.cpu.rf.rf[6][11] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold180 (.A(\i_soc.cpu.rf.rf[6][0] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold181 (.A(\i_soc.cpu.rf.rf[6][4] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold182 (.A(\i_soc.cpu.rf.rf[7][16] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold183 (.A(\i_soc.cpu.rf.rf[7][19] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold184 (.A(\i_soc.cpu.rf.rf[5][6] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold185 (.A(\i_soc.cpu.rf.rf[5][20] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold186 (.A(\i_soc.cpu.rf.rf[5][22] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold187 (.A(\i_soc.cpu.rf.rf[6][20] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold188 (.A(\i_soc.cpu.rf.rf[6][29] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold189 (.A(\i_soc.cpu.rf.rf[6][31] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold190 (.A(\i_soc.cpu.rf.rf[6][16] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold191 (.A(\i_soc.cpu.rf.rf[6][2] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold192 (.A(\i_soc.cpu.rf.rf[5][29] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold193 (.A(\i_soc.cpu.rf.rf[6][23] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold194 (.A(\i_soc.cpu.rf.rf[7][24] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold195 (.A(\i_soc.cpu.rf.rf[6][21] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold196 (.A(\i_soc.cpu.rf.rf[6][13] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold197 (.A(\i_soc.cpu.rf.rf[6][7] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold198 (.A(\i_soc.cpu.rf.rf[6][26] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold199 (.A(\i_soc.cpu.rf.rf[7][18] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold200 (.A(\i_soc.cpu.rf.rf[5][0] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold201 (.A(\i_soc.cpu.rf.rf[5][16] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold202 (.A(\i_soc.cpu.rf.rf[7][20] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold203 (.A(\i_soc.cpu.rf.rf[6][1] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold204 (.A(\i_soc.cpu.rf.rf[6][22] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold205 (.A(\i_soc.cpu.rf.rf[6][28] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold206 (.A(\i_soc.cpu.rf.rf[6][3] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold207 (.A(\i_soc.cpu.rf.rf[7][8] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold208 (.A(\i_soc.cpu.rf.rf[5][15] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold209 (.A(\i_soc.cpu.rf.rf[5][31] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold210 (.A(\i_soc.cpu.rf.rf[5][13] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold211 (.A(\i_soc.cpu.rf.rf[5][27] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold212 (.A(\i_soc.cpu.rf.rf[7][11] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold213 (.A(\i_soc.cpu.rf.rf[7][3] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold214 (.A(\i_soc.cpu.rf.rf[7][30] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold215 (.A(\i_soc.cpu.rf.rf[6][10] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold216 (.A(\i_soc.cpu.rf.rf[5][2] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold217 (.A(\i_soc.cpu.rf.rf[7][12] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold218 (.A(\i_soc.cpu.rf.rf[5][10] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold219 (.A(\i_soc.cpu.rf.rf[6][18] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold220 (.A(\i_soc.cpu.rf.rf[6][27] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold221 (.A(\i_soc.cpu.rf.rf[7][4] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold222 (.A(\i_soc.cpu.rf.rf[5][5] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold223 (.A(\i_soc.cpu.rf.rf[7][5] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold224 (.A(\i_soc.cpu.rf.rf[6][17] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold225 (.A(\i_soc.cpu.rf.rf[5][24] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold226 (.A(\i_soc.cpu.rf.rf[7][2] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold227 (.A(\i_soc.cpu.rf.rf[7][7] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold228 (.A(\i_soc.cpu.rf.rf[5][26] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold229 (.A(\i_soc.cpu.rf.rf[7][26] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold230 (.A(\i_soc.cpu.rf.rf[6][6] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold231 (.A(\i_soc.cpu.rf.rf[7][14] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold232 (.A(\i_soc.cpu.rf.rf[5][30] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold233 (.A(\i_soc.cpu.rf.rf[7][9] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold234 (.A(\i_soc.cpu.rf.rf[6][5] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold235 (.A(\i_soc.cpu.rf.rf[5][1] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold236 (.A(\i_soc.cpu.rf.rf[6][8] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold237 (.A(\i_soc.cpu.rf.rf[7][6] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold238 (.A(\i_soc.cpu.rf.rf[5][23] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold239 (.A(\i_soc.cpu.rf.rf[7][31] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold240 (.A(\i_soc.cpu.rf.rf[6][14] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold241 (.A(\i_soc.cpu.rf.rf[5][18] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold242 (.A(\i_soc.cpu.rf.rf[6][12] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold243 (.A(\i_soc.cpu.rf.rf[6][25] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold244 (.A(\i_soc.cpu.rf.rf[5][25] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold245 (.A(\i_soc.cpu.rf.rf[5][8] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold246 (.A(\i_soc.cpu.rf.rf[7][10] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold247 (.A(\i_soc.cpu.rf.rf[7][22] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold248 (.A(\i_soc.cpu.rf.rf[6][24] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold249 (.A(\i_soc.cpu.rf.rf[5][21] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold250 (.A(\i_soc.cpu.rd0[18] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold251 (.A(\i_soc.cpu.rf.rf[7][17] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold252 (.A(\i_soc.cpu.rf.rf[5][4] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold253 (.A(\i_soc.cpu.rf.rf[7][23] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold254 (.A(\i_soc.cpu.rf.rf[5][19] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold255 (.A(\i_soc.cpu.rf.rf[5][17] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold256 (.A(\i_soc.cpu.rf.rf[7][15] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold257 (.A(\i_soc.cpu.rf.rf[5][28] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold258 (.A(\i_soc.cpu.rf.rf[6][30] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold259 (.A(\i_soc.cpu.rd0[21] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold260 (.A(\i_soc.cpu.rf.rf[5][12] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold261 (.A(\i_soc.cpu.rd0[25] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold262 (.A(\i_soc.cpu.rf.rf[7][27] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold263 (.A(\i_soc.cpu.rf.rf[6][9] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold264 (.A(\i_soc.cpu.rd0[16] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold265 (.A(\i_soc.cpu.rd0[17] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold266 (.A(\i_soc.cpu.rf.rf[5][11] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold267 (.A(\i_soc.cpu.rf.rf[7][29] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold268 (.A(\i_soc.cpu.rf.rf[5][3] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold269 (.A(\i_soc.cnt[0] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0492_),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold271 (.A(\i_soc.cpu.rd0[9] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold272 (.A(\i_soc.cpu.rd0[19] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold273 (.A(\i_soc.cnt[2] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold274 (.A(_1482_),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold275 (.A(\i_soc.cpu.rf.rf[5][9] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold276 (.A(\i_soc.cpu.rd0[6] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold277 (.A(\i_soc.cpu.rd0[14] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold278 (.A(\i_soc.cpu.rd0[12] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold279 (.A(\i_soc.cpu.rd0[5] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold280 (.A(\i_soc.cpu.rd0[4] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold281 (.A(\i_soc.cpu.rf.rf[7][1] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold282 (.A(\i_soc.cpu.rd0[13] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold283 (.A(\i_soc.cnt[6] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold284 (.A(_1490_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0497_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold286 (.A(\i_soc.cpu.rd0[15] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold287 (.A(\i_soc.cpu.rd0[24] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold288 (.A(\i_soc.cpu.rd0[26] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold289 (.A(\i_soc.cpu.rd0[29] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold290 (.A(\i_soc.cpu.rd0[27] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold291 (.A(\i_soc.cpu.rd0[7] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold292 (.A(\i_soc.cpu.rd0[31] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold293 (.A(\i_soc.cpu.rd0[3] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold294 (.A(\i_soc.cpu.rd0[20] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold295 (.A(\i_soc.cpu.rd0[10] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold296 (.A(\i_soc.cpu.rd0[28] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold297 (.A(\i_soc.cpu.rd0[30] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold298 (.A(\i_soc.cpu.rd0[23] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold299 (.A(\i_soc.cpu.rd0[22] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold300 (.A(\i_soc.cpu.rd0[11] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold301 (.A(\i_soc.cpu.rd0[2] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold302 (.A(\i_soc.pass ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold303 (.A(\i_soc.cpu.rd0[1] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold304 (.A(\i_soc.cpu.rd0[8] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold305 (.A(\i_soc.cnt[4] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold306 (.A(_1488_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold307 (.A(\i_soc.cnt[5] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold308 (.A(\i_soc.cpu.rd0[0] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold309 (.A(fail),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold310 (.A(_1542_),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold311 (.A(\i_soc.cnt[7] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold312 (.A(\i_soc.cnt[3] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold313 (.A(_1485_),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold314 (.A(\i_soc.cpu.pc[5] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold315 (.A(_1496_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold316 (.A(\i_soc.cpu.pc[3] ),
    .X(net790));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_fill_2 FILLER_0_91 ();
 sg13g2_decap_4 FILLER_0_106 ();
 sg13g2_fill_1 FILLER_0_110 ();
 sg13g2_decap_8 FILLER_0_115 ();
 sg13g2_fill_2 FILLER_0_122 ();
 sg13g2_fill_2 FILLER_0_150 ();
 sg13g2_decap_8 FILLER_0_156 ();
 sg13g2_fill_2 FILLER_0_163 ();
 sg13g2_decap_8 FILLER_0_191 ();
 sg13g2_decap_8 FILLER_0_198 ();
 sg13g2_decap_8 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_212 ();
 sg13g2_decap_8 FILLER_0_219 ();
 sg13g2_decap_8 FILLER_0_226 ();
 sg13g2_decap_8 FILLER_0_233 ();
 sg13g2_decap_8 FILLER_0_240 ();
 sg13g2_decap_8 FILLER_0_247 ();
 sg13g2_fill_2 FILLER_0_254 ();
 sg13g2_fill_2 FILLER_0_260 ();
 sg13g2_fill_1 FILLER_0_262 ();
 sg13g2_decap_8 FILLER_0_272 ();
 sg13g2_decap_4 FILLER_0_279 ();
 sg13g2_fill_2 FILLER_0_283 ();
 sg13g2_decap_4 FILLER_0_289 ();
 sg13g2_fill_1 FILLER_0_293 ();
 sg13g2_decap_4 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_decap_8 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_0_334 ();
 sg13g2_decap_8 FILLER_0_341 ();
 sg13g2_decap_8 FILLER_0_348 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_4 FILLER_0_404 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_fill_2 FILLER_1_84 ();
 sg13g2_decap_4 FILLER_1_121 ();
 sg13g2_fill_1 FILLER_1_125 ();
 sg13g2_fill_2 FILLER_1_134 ();
 sg13g2_fill_1 FILLER_1_136 ();
 sg13g2_fill_2 FILLER_1_172 ();
 sg13g2_fill_1 FILLER_1_174 ();
 sg13g2_decap_8 FILLER_1_201 ();
 sg13g2_decap_8 FILLER_1_208 ();
 sg13g2_decap_8 FILLER_1_215 ();
 sg13g2_decap_8 FILLER_1_222 ();
 sg13g2_decap_8 FILLER_1_229 ();
 sg13g2_decap_8 FILLER_1_236 ();
 sg13g2_decap_4 FILLER_1_269 ();
 sg13g2_fill_2 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_327 ();
 sg13g2_decap_8 FILLER_1_334 ();
 sg13g2_decap_8 FILLER_1_341 ();
 sg13g2_decap_8 FILLER_1_348 ();
 sg13g2_decap_8 FILLER_1_355 ();
 sg13g2_decap_8 FILLER_1_362 ();
 sg13g2_decap_8 FILLER_1_369 ();
 sg13g2_decap_8 FILLER_1_376 ();
 sg13g2_decap_8 FILLER_1_383 ();
 sg13g2_decap_8 FILLER_1_390 ();
 sg13g2_decap_8 FILLER_1_397 ();
 sg13g2_decap_4 FILLER_1_404 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_4 FILLER_2_77 ();
 sg13g2_fill_1 FILLER_2_111 ();
 sg13g2_fill_2 FILLER_2_125 ();
 sg13g2_fill_1 FILLER_2_136 ();
 sg13g2_decap_4 FILLER_2_158 ();
 sg13g2_fill_1 FILLER_2_162 ();
 sg13g2_fill_2 FILLER_2_171 ();
 sg13g2_fill_1 FILLER_2_173 ();
 sg13g2_fill_1 FILLER_2_195 ();
 sg13g2_decap_8 FILLER_2_205 ();
 sg13g2_decap_8 FILLER_2_212 ();
 sg13g2_decap_8 FILLER_2_219 ();
 sg13g2_decap_8 FILLER_2_226 ();
 sg13g2_fill_2 FILLER_2_233 ();
 sg13g2_fill_1 FILLER_2_235 ();
 sg13g2_fill_2 FILLER_2_270 ();
 sg13g2_fill_1 FILLER_2_272 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_4 FILLER_3_84 ();
 sg13g2_fill_1 FILLER_3_88 ();
 sg13g2_fill_1 FILLER_3_146 ();
 sg13g2_decap_8 FILLER_3_177 ();
 sg13g2_fill_1 FILLER_3_184 ();
 sg13g2_decap_8 FILLER_3_206 ();
 sg13g2_decap_8 FILLER_3_213 ();
 sg13g2_decap_8 FILLER_3_220 ();
 sg13g2_decap_8 FILLER_3_227 ();
 sg13g2_decap_4 FILLER_3_234 ();
 sg13g2_fill_2 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_4 FILLER_4_92 ();
 sg13g2_fill_1 FILLER_4_100 ();
 sg13g2_decap_8 FILLER_4_131 ();
 sg13g2_fill_2 FILLER_4_138 ();
 sg13g2_fill_1 FILLER_4_140 ();
 sg13g2_fill_2 FILLER_4_171 ();
 sg13g2_decap_8 FILLER_4_212 ();
 sg13g2_decap_4 FILLER_4_219 ();
 sg13g2_fill_2 FILLER_4_223 ();
 sg13g2_decap_8 FILLER_4_234 ();
 sg13g2_fill_1 FILLER_4_241 ();
 sg13g2_fill_2 FILLER_4_268 ();
 sg13g2_fill_1 FILLER_4_270 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_318 ();
 sg13g2_decap_8 FILLER_4_325 ();
 sg13g2_decap_8 FILLER_4_332 ();
 sg13g2_decap_8 FILLER_4_339 ();
 sg13g2_decap_8 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_367 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_fill_1 FILLER_5_112 ();
 sg13g2_fill_2 FILLER_5_170 ();
 sg13g2_fill_1 FILLER_5_172 ();
 sg13g2_fill_2 FILLER_5_207 ();
 sg13g2_fill_1 FILLER_5_209 ();
 sg13g2_fill_1 FILLER_5_253 ();
 sg13g2_fill_2 FILLER_5_275 ();
 sg13g2_fill_2 FILLER_5_299 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_354 ();
 sg13g2_decap_8 FILLER_5_361 ();
 sg13g2_decap_8 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_decap_8 FILLER_5_382 ();
 sg13g2_decap_8 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_4 FILLER_5_403 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_fill_2 FILLER_6_96 ();
 sg13g2_fill_1 FILLER_6_98 ();
 sg13g2_fill_2 FILLER_6_112 ();
 sg13g2_fill_2 FILLER_6_122 ();
 sg13g2_fill_2 FILLER_6_129 ();
 sg13g2_fill_2 FILLER_6_153 ();
 sg13g2_fill_2 FILLER_6_183 ();
 sg13g2_fill_1 FILLER_6_190 ();
 sg13g2_decap_8 FILLER_6_200 ();
 sg13g2_fill_2 FILLER_6_207 ();
 sg13g2_fill_1 FILLER_6_209 ();
 sg13g2_decap_4 FILLER_6_263 ();
 sg13g2_fill_1 FILLER_6_267 ();
 sg13g2_fill_2 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_fill_2 FILLER_7_134 ();
 sg13g2_fill_2 FILLER_7_141 ();
 sg13g2_fill_2 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_4 FILLER_7_210 ();
 sg13g2_fill_2 FILLER_7_214 ();
 sg13g2_decap_4 FILLER_7_258 ();
 sg13g2_fill_1 FILLER_7_262 ();
 sg13g2_decap_8 FILLER_7_354 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_4 FILLER_8_84 ();
 sg13g2_fill_2 FILLER_8_205 ();
 sg13g2_decap_8 FILLER_8_214 ();
 sg13g2_decap_8 FILLER_8_221 ();
 sg13g2_decap_8 FILLER_8_228 ();
 sg13g2_decap_4 FILLER_8_278 ();
 sg13g2_fill_1 FILLER_8_282 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_4 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_fill_2 FILLER_9_77 ();
 sg13g2_fill_2 FILLER_9_142 ();
 sg13g2_fill_1 FILLER_9_144 ();
 sg13g2_fill_1 FILLER_9_219 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_4 FILLER_9_240 ();
 sg13g2_fill_2 FILLER_9_244 ();
 sg13g2_decap_4 FILLER_9_289 ();
 sg13g2_fill_1 FILLER_9_297 ();
 sg13g2_decap_8 FILLER_9_331 ();
 sg13g2_decap_8 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_345 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_decap_8 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_4 FILLER_10_63 ();
 sg13g2_fill_1 FILLER_10_114 ();
 sg13g2_fill_1 FILLER_10_130 ();
 sg13g2_decap_8 FILLER_10_295 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_4 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_339 ();
 sg13g2_decap_8 FILLER_10_346 ();
 sg13g2_decap_8 FILLER_10_353 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_4 FILLER_11_56 ();
 sg13g2_fill_2 FILLER_11_60 ();
 sg13g2_decap_4 FILLER_11_142 ();
 sg13g2_fill_1 FILLER_11_146 ();
 sg13g2_fill_2 FILLER_11_152 ();
 sg13g2_decap_8 FILLER_11_159 ();
 sg13g2_fill_2 FILLER_11_166 ();
 sg13g2_fill_1 FILLER_11_168 ();
 sg13g2_fill_1 FILLER_11_212 ();
 sg13g2_fill_1 FILLER_11_218 ();
 sg13g2_fill_2 FILLER_11_245 ();
 sg13g2_fill_1 FILLER_11_317 ();
 sg13g2_decap_8 FILLER_11_344 ();
 sg13g2_decap_8 FILLER_11_351 ();
 sg13g2_decap_8 FILLER_11_358 ();
 sg13g2_decap_8 FILLER_11_365 ();
 sg13g2_decap_8 FILLER_11_372 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_8 FILLER_11_393 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_4 FILLER_12_56 ();
 sg13g2_fill_1 FILLER_12_60 ();
 sg13g2_fill_1 FILLER_12_96 ();
 sg13g2_fill_1 FILLER_12_109 ();
 sg13g2_fill_2 FILLER_12_153 ();
 sg13g2_decap_8 FILLER_12_164 ();
 sg13g2_decap_4 FILLER_12_171 ();
 sg13g2_fill_2 FILLER_12_175 ();
 sg13g2_fill_2 FILLER_12_185 ();
 sg13g2_fill_1 FILLER_12_187 ();
 sg13g2_fill_2 FILLER_12_223 ();
 sg13g2_fill_2 FILLER_12_233 ();
 sg13g2_fill_1 FILLER_12_235 ();
 sg13g2_fill_2 FILLER_12_258 ();
 sg13g2_fill_2 FILLER_12_278 ();
 sg13g2_fill_1 FILLER_12_280 ();
 sg13g2_fill_2 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_decap_8 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_fill_2 FILLER_13_63 ();
 sg13g2_fill_1 FILLER_13_65 ();
 sg13g2_fill_1 FILLER_13_123 ();
 sg13g2_fill_2 FILLER_13_134 ();
 sg13g2_fill_1 FILLER_13_136 ();
 sg13g2_fill_2 FILLER_13_171 ();
 sg13g2_fill_1 FILLER_13_173 ();
 sg13g2_fill_2 FILLER_13_178 ();
 sg13g2_fill_1 FILLER_13_180 ();
 sg13g2_decap_8 FILLER_13_190 ();
 sg13g2_fill_1 FILLER_13_205 ();
 sg13g2_decap_4 FILLER_13_214 ();
 sg13g2_fill_2 FILLER_13_218 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_fill_2 FILLER_13_260 ();
 sg13g2_fill_1 FILLER_13_262 ();
 sg13g2_fill_1 FILLER_13_318 ();
 sg13g2_fill_1 FILLER_13_337 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_decap_8 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_4 FILLER_14_56 ();
 sg13g2_fill_2 FILLER_14_70 ();
 sg13g2_fill_2 FILLER_14_112 ();
 sg13g2_fill_1 FILLER_14_114 ();
 sg13g2_fill_2 FILLER_14_128 ();
 sg13g2_fill_1 FILLER_14_138 ();
 sg13g2_fill_1 FILLER_14_147 ();
 sg13g2_fill_1 FILLER_14_162 ();
 sg13g2_fill_2 FILLER_14_194 ();
 sg13g2_fill_2 FILLER_14_201 ();
 sg13g2_fill_1 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_fill_2 FILLER_14_224 ();
 sg13g2_fill_1 FILLER_14_226 ();
 sg13g2_fill_2 FILLER_14_236 ();
 sg13g2_fill_2 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_fill_2 FILLER_15_86 ();
 sg13g2_fill_1 FILLER_15_100 ();
 sg13g2_fill_2 FILLER_15_136 ();
 sg13g2_decap_4 FILLER_15_148 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_decap_4 FILLER_15_189 ();
 sg13g2_fill_2 FILLER_15_193 ();
 sg13g2_decap_4 FILLER_15_221 ();
 sg13g2_fill_2 FILLER_15_225 ();
 sg13g2_fill_2 FILLER_15_232 ();
 sg13g2_fill_2 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_240 ();
 sg13g2_fill_1 FILLER_15_258 ();
 sg13g2_fill_1 FILLER_15_264 ();
 sg13g2_decap_4 FILLER_15_270 ();
 sg13g2_fill_2 FILLER_15_274 ();
 sg13g2_fill_1 FILLER_15_311 ();
 sg13g2_fill_2 FILLER_15_338 ();
 sg13g2_decap_8 FILLER_15_344 ();
 sg13g2_decap_8 FILLER_15_351 ();
 sg13g2_decap_8 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_fill_1 FILLER_16_63 ();
 sg13g2_fill_1 FILLER_16_103 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_142 ();
 sg13g2_fill_2 FILLER_16_154 ();
 sg13g2_fill_1 FILLER_16_156 ();
 sg13g2_fill_2 FILLER_16_167 ();
 sg13g2_fill_2 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_fill_2 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_4 FILLER_16_233 ();
 sg13g2_decap_8 FILLER_16_246 ();
 sg13g2_fill_1 FILLER_16_253 ();
 sg13g2_decap_8 FILLER_16_264 ();
 sg13g2_decap_8 FILLER_16_271 ();
 sg13g2_decap_8 FILLER_16_278 ();
 sg13g2_decap_8 FILLER_16_285 ();
 sg13g2_fill_2 FILLER_16_300 ();
 sg13g2_fill_1 FILLER_16_320 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_fill_2 FILLER_17_63 ();
 sg13g2_fill_1 FILLER_17_65 ();
 sg13g2_fill_1 FILLER_17_87 ();
 sg13g2_decap_8 FILLER_17_131 ();
 sg13g2_fill_2 FILLER_17_138 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_fill_2 FILLER_17_161 ();
 sg13g2_fill_2 FILLER_17_211 ();
 sg13g2_fill_1 FILLER_17_223 ();
 sg13g2_fill_1 FILLER_17_231 ();
 sg13g2_fill_2 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_282 ();
 sg13g2_decap_4 FILLER_17_289 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_fill_1 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_358 ();
 sg13g2_decap_8 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_56 ();
 sg13g2_fill_1 FILLER_18_83 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_fill_1 FILLER_18_112 ();
 sg13g2_fill_2 FILLER_18_130 ();
 sg13g2_fill_1 FILLER_18_132 ();
 sg13g2_fill_1 FILLER_18_180 ();
 sg13g2_fill_1 FILLER_18_202 ();
 sg13g2_fill_1 FILLER_18_219 ();
 sg13g2_fill_1 FILLER_18_257 ();
 sg13g2_fill_2 FILLER_18_284 ();
 sg13g2_fill_1 FILLER_18_286 ();
 sg13g2_fill_1 FILLER_18_313 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_fill_1 FILLER_19_63 ();
 sg13g2_fill_2 FILLER_19_90 ();
 sg13g2_fill_1 FILLER_19_92 ();
 sg13g2_fill_2 FILLER_19_110 ();
 sg13g2_fill_2 FILLER_19_152 ();
 sg13g2_fill_1 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_decap_4 FILLER_19_199 ();
 sg13g2_fill_2 FILLER_19_228 ();
 sg13g2_fill_1 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_360 ();
 sg13g2_decap_8 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_374 ();
 sg13g2_decap_8 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_19_395 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_4 FILLER_20_70 ();
 sg13g2_fill_2 FILLER_20_82 ();
 sg13g2_fill_1 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_fill_2 FILLER_20_110 ();
 sg13g2_fill_1 FILLER_20_152 ();
 sg13g2_fill_1 FILLER_20_166 ();
 sg13g2_fill_2 FILLER_20_192 ();
 sg13g2_fill_1 FILLER_20_194 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_fill_2 FILLER_20_217 ();
 sg13g2_fill_2 FILLER_20_254 ();
 sg13g2_fill_1 FILLER_20_256 ();
 sg13g2_fill_2 FILLER_20_266 ();
 sg13g2_fill_1 FILLER_20_295 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_fill_2 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_107 ();
 sg13g2_fill_1 FILLER_21_113 ();
 sg13g2_fill_2 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_121 ();
 sg13g2_fill_2 FILLER_21_143 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_fill_2 FILLER_21_159 ();
 sg13g2_fill_1 FILLER_21_161 ();
 sg13g2_fill_2 FILLER_21_167 ();
 sg13g2_decap_4 FILLER_21_173 ();
 sg13g2_fill_1 FILLER_21_191 ();
 sg13g2_fill_2 FILLER_21_196 ();
 sg13g2_fill_2 FILLER_21_210 ();
 sg13g2_fill_1 FILLER_21_212 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_4 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_235 ();
 sg13g2_decap_8 FILLER_21_251 ();
 sg13g2_decap_4 FILLER_21_258 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_292 ();
 sg13g2_fill_2 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_317 ();
 sg13g2_fill_2 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_21_338 ();
 sg13g2_decap_8 FILLER_21_345 ();
 sg13g2_decap_8 FILLER_21_352 ();
 sg13g2_decap_8 FILLER_21_359 ();
 sg13g2_decap_8 FILLER_21_366 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_140 ();
 sg13g2_decap_4 FILLER_22_152 ();
 sg13g2_fill_2 FILLER_22_156 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_186 ();
 sg13g2_decap_4 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_237 ();
 sg13g2_fill_1 FILLER_22_253 ();
 sg13g2_decap_4 FILLER_22_258 ();
 sg13g2_fill_1 FILLER_22_262 ();
 sg13g2_fill_2 FILLER_22_299 ();
 sg13g2_fill_1 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_4 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_53 ();
 sg13g2_fill_1 FILLER_23_80 ();
 sg13g2_fill_1 FILLER_23_166 ();
 sg13g2_fill_1 FILLER_23_198 ();
 sg13g2_fill_2 FILLER_23_217 ();
 sg13g2_fill_1 FILLER_23_254 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_117 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_2 FILLER_24_134 ();
 sg13g2_fill_1 FILLER_24_143 ();
 sg13g2_fill_1 FILLER_24_321 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_4 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_90 ();
 sg13g2_fill_1 FILLER_25_92 ();
 sg13g2_decap_8 FILLER_25_101 ();
 sg13g2_fill_1 FILLER_25_108 ();
 sg13g2_fill_2 FILLER_25_143 ();
 sg13g2_fill_2 FILLER_25_185 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_decap_8 FILLER_25_192 ();
 sg13g2_decap_4 FILLER_25_199 ();
 sg13g2_fill_2 FILLER_25_203 ();
 sg13g2_fill_1 FILLER_25_229 ();
 sg13g2_fill_1 FILLER_25_249 ();
 sg13g2_fill_2 FILLER_25_259 ();
 sg13g2_fill_1 FILLER_25_267 ();
 sg13g2_fill_2 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_279 ();
 sg13g2_fill_2 FILLER_25_311 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_decap_4 FILLER_25_324 ();
 sg13g2_fill_2 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_55 ();
 sg13g2_fill_1 FILLER_26_57 ();
 sg13g2_fill_1 FILLER_26_84 ();
 sg13g2_fill_1 FILLER_26_94 ();
 sg13g2_fill_2 FILLER_26_113 ();
 sg13g2_fill_2 FILLER_26_125 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_2 FILLER_26_148 ();
 sg13g2_fill_2 FILLER_26_167 ();
 sg13g2_decap_8 FILLER_26_184 ();
 sg13g2_decap_4 FILLER_26_191 ();
 sg13g2_decap_8 FILLER_26_199 ();
 sg13g2_fill_1 FILLER_26_216 ();
 sg13g2_fill_1 FILLER_26_234 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_fill_1 FILLER_26_259 ();
 sg13g2_fill_2 FILLER_26_267 ();
 sg13g2_decap_4 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_295 ();
 sg13g2_decap_4 FILLER_26_302 ();
 sg13g2_fill_1 FILLER_26_319 ();
 sg13g2_decap_8 FILLER_26_354 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_128 ();
 sg13g2_decap_4 FILLER_27_153 ();
 sg13g2_fill_1 FILLER_27_157 ();
 sg13g2_decap_8 FILLER_27_166 ();
 sg13g2_decap_8 FILLER_27_173 ();
 sg13g2_decap_4 FILLER_27_180 ();
 sg13g2_fill_1 FILLER_27_184 ();
 sg13g2_fill_2 FILLER_27_211 ();
 sg13g2_fill_1 FILLER_27_213 ();
 sg13g2_fill_2 FILLER_27_223 ();
 sg13g2_fill_2 FILLER_27_251 ();
 sg13g2_fill_1 FILLER_27_253 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_285 ();
 sg13g2_decap_4 FILLER_27_292 ();
 sg13g2_decap_8 FILLER_27_362 ();
 sg13g2_decap_8 FILLER_27_369 ();
 sg13g2_decap_8 FILLER_27_376 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_decap_8 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_65 ();
 sg13g2_decap_4 FILLER_28_164 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_fill_2 FILLER_28_244 ();
 sg13g2_fill_1 FILLER_28_246 ();
 sg13g2_fill_2 FILLER_28_276 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_319 ();
 sg13g2_fill_1 FILLER_28_321 ();
 sg13g2_decap_8 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_28_359 ();
 sg13g2_decap_8 FILLER_28_366 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_4 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_39 ();
 sg13g2_fill_2 FILLER_29_48 ();
 sg13g2_decap_4 FILLER_29_59 ();
 sg13g2_fill_2 FILLER_29_127 ();
 sg13g2_fill_1 FILLER_29_129 ();
 sg13g2_fill_2 FILLER_29_243 ();
 sg13g2_fill_1 FILLER_29_245 ();
 sg13g2_fill_2 FILLER_29_255 ();
 sg13g2_fill_1 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_decap_8 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_29_370 ();
 sg13g2_decap_8 FILLER_29_377 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_4 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_53 ();
 sg13g2_decap_4 FILLER_30_59 ();
 sg13g2_fill_1 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_73 ();
 sg13g2_decap_4 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_88 ();
 sg13g2_fill_1 FILLER_30_103 ();
 sg13g2_fill_2 FILLER_30_131 ();
 sg13g2_fill_1 FILLER_30_133 ();
 sg13g2_fill_2 FILLER_30_139 ();
 sg13g2_decap_8 FILLER_30_145 ();
 sg13g2_fill_1 FILLER_30_173 ();
 sg13g2_fill_2 FILLER_30_187 ();
 sg13g2_fill_1 FILLER_30_189 ();
 sg13g2_fill_2 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_202 ();
 sg13g2_fill_2 FILLER_30_207 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_fill_2 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_226 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_277 ();
 sg13g2_fill_2 FILLER_30_311 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_decap_8 FILLER_30_344 ();
 sg13g2_decap_8 FILLER_30_351 ();
 sg13g2_decap_8 FILLER_30_358 ();
 sg13g2_decap_8 FILLER_30_365 ();
 sg13g2_decap_8 FILLER_30_372 ();
 sg13g2_decap_8 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_30_386 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_fill_2 FILLER_31_42 ();
 sg13g2_fill_1 FILLER_31_44 ();
 sg13g2_fill_2 FILLER_31_97 ();
 sg13g2_fill_1 FILLER_31_99 ();
 sg13g2_fill_1 FILLER_31_141 ();
 sg13g2_decap_8 FILLER_31_146 ();
 sg13g2_decap_4 FILLER_31_153 ();
 sg13g2_fill_1 FILLER_31_157 ();
 sg13g2_fill_2 FILLER_31_166 ();
 sg13g2_decap_4 FILLER_31_181 ();
 sg13g2_fill_2 FILLER_31_185 ();
 sg13g2_decap_8 FILLER_31_201 ();
 sg13g2_decap_8 FILLER_31_212 ();
 sg13g2_decap_8 FILLER_31_219 ();
 sg13g2_fill_1 FILLER_31_226 ();
 sg13g2_fill_2 FILLER_31_271 ();
 sg13g2_fill_1 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_278 ();
 sg13g2_decap_8 FILLER_31_285 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_decap_4 FILLER_31_312 ();
 sg13g2_fill_2 FILLER_31_316 ();
 sg13g2_decap_8 FILLER_31_348 ();
 sg13g2_decap_8 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_362 ();
 sg13g2_decap_8 FILLER_31_369 ();
 sg13g2_decap_8 FILLER_31_376 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_4 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_81 ();
 sg13g2_fill_2 FILLER_32_118 ();
 sg13g2_fill_2 FILLER_32_153 ();
 sg13g2_fill_1 FILLER_32_192 ();
 sg13g2_decap_4 FILLER_32_243 ();
 sg13g2_decap_4 FILLER_32_292 ();
 sg13g2_fill_1 FILLER_32_296 ();
 sg13g2_fill_2 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_309 ();
 sg13g2_decap_8 FILLER_32_354 ();
 sg13g2_decap_8 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_375 ();
 sg13g2_decap_8 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_32_389 ();
 sg13g2_decap_8 FILLER_32_396 ();
 sg13g2_decap_4 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_fill_1 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_78 ();
 sg13g2_fill_2 FILLER_33_128 ();
 sg13g2_fill_2 FILLER_33_138 ();
 sg13g2_decap_8 FILLER_33_164 ();
 sg13g2_fill_2 FILLER_33_210 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_349 ();
 sg13g2_decap_8 FILLER_33_356 ();
 sg13g2_decap_8 FILLER_33_363 ();
 sg13g2_decap_8 FILLER_33_370 ();
 sg13g2_decap_8 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_384 ();
 sg13g2_decap_8 FILLER_33_391 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_4 FILLER_34_49 ();
 sg13g2_fill_1 FILLER_34_53 ();
 sg13g2_decap_4 FILLER_34_63 ();
 sg13g2_fill_2 FILLER_34_67 ();
 sg13g2_decap_4 FILLER_34_73 ();
 sg13g2_fill_1 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_82 ();
 sg13g2_fill_2 FILLER_34_92 ();
 sg13g2_fill_2 FILLER_34_107 ();
 sg13g2_fill_2 FILLER_34_123 ();
 sg13g2_fill_1 FILLER_34_125 ();
 sg13g2_decap_4 FILLER_34_153 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_decap_8 FILLER_34_166 ();
 sg13g2_fill_1 FILLER_34_181 ();
 sg13g2_fill_2 FILLER_34_190 ();
 sg13g2_fill_2 FILLER_34_217 ();
 sg13g2_fill_1 FILLER_34_252 ();
 sg13g2_fill_2 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_277 ();
 sg13g2_decap_8 FILLER_34_338 ();
 sg13g2_decap_8 FILLER_34_345 ();
 sg13g2_decap_8 FILLER_34_352 ();
 sg13g2_decap_8 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_34_366 ();
 sg13g2_decap_8 FILLER_34_373 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_fill_2 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_81 ();
 sg13g2_fill_2 FILLER_35_88 ();
 sg13g2_fill_1 FILLER_35_90 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_157 ();
 sg13g2_fill_1 FILLER_35_159 ();
 sg13g2_fill_2 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_174 ();
 sg13g2_decap_8 FILLER_35_181 ();
 sg13g2_fill_1 FILLER_35_188 ();
 sg13g2_fill_1 FILLER_35_194 ();
 sg13g2_fill_1 FILLER_35_221 ();
 sg13g2_fill_2 FILLER_35_290 ();
 sg13g2_fill_1 FILLER_35_292 ();
 sg13g2_decap_8 FILLER_35_328 ();
 sg13g2_decap_8 FILLER_35_335 ();
 sg13g2_decap_8 FILLER_35_342 ();
 sg13g2_decap_8 FILLER_35_349 ();
 sg13g2_decap_8 FILLER_35_356 ();
 sg13g2_decap_8 FILLER_35_363 ();
 sg13g2_decap_8 FILLER_35_370 ();
 sg13g2_decap_8 FILLER_35_377 ();
 sg13g2_decap_8 FILLER_35_384 ();
 sg13g2_decap_8 FILLER_35_391 ();
 sg13g2_decap_8 FILLER_35_398 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_133 ();
 sg13g2_fill_2 FILLER_36_149 ();
 sg13g2_fill_1 FILLER_36_151 ();
 sg13g2_decap_8 FILLER_36_183 ();
 sg13g2_decap_4 FILLER_36_190 ();
 sg13g2_fill_2 FILLER_36_194 ();
 sg13g2_fill_2 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_203 ();
 sg13g2_fill_2 FILLER_36_209 ();
 sg13g2_fill_2 FILLER_36_215 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_decap_4 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_250 ();
 sg13g2_decap_8 FILLER_36_265 ();
 sg13g2_fill_2 FILLER_36_302 ();
 sg13g2_fill_1 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_fill_2 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_44 ();
 sg13g2_decap_4 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_53 ();
 sg13g2_decap_4 FILLER_37_93 ();
 sg13g2_fill_2 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_116 ();
 sg13g2_fill_2 FILLER_37_123 ();
 sg13g2_fill_2 FILLER_37_130 ();
 sg13g2_fill_1 FILLER_37_132 ();
 sg13g2_fill_1 FILLER_37_142 ();
 sg13g2_fill_2 FILLER_37_148 ();
 sg13g2_fill_1 FILLER_37_150 ();
 sg13g2_fill_1 FILLER_37_181 ();
 sg13g2_fill_2 FILLER_37_212 ();
 sg13g2_decap_8 FILLER_37_226 ();
 sg13g2_decap_8 FILLER_37_233 ();
 sg13g2_decap_8 FILLER_37_240 ();
 sg13g2_decap_8 FILLER_37_247 ();
 sg13g2_decap_8 FILLER_37_254 ();
 sg13g2_decap_4 FILLER_37_261 ();
 sg13g2_decap_8 FILLER_37_270 ();
 sg13g2_decap_4 FILLER_37_277 ();
 sg13g2_fill_2 FILLER_37_281 ();
 sg13g2_decap_8 FILLER_37_291 ();
 sg13g2_fill_2 FILLER_37_298 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_decap_8 FILLER_37_327 ();
 sg13g2_decap_8 FILLER_37_334 ();
 sg13g2_decap_8 FILLER_37_341 ();
 sg13g2_decap_8 FILLER_37_348 ();
 sg13g2_decap_8 FILLER_37_355 ();
 sg13g2_decap_8 FILLER_37_362 ();
 sg13g2_decap_8 FILLER_37_369 ();
 sg13g2_decap_8 FILLER_37_376 ();
 sg13g2_decap_8 FILLER_37_383 ();
 sg13g2_decap_8 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_4 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_32 ();
 sg13g2_decap_8 FILLER_38_100 ();
 sg13g2_decap_8 FILLER_38_107 ();
 sg13g2_fill_2 FILLER_38_114 ();
 sg13g2_fill_2 FILLER_38_142 ();
 sg13g2_fill_1 FILLER_38_162 ();
 sg13g2_fill_2 FILLER_38_193 ();
 sg13g2_decap_4 FILLER_38_217 ();
 sg13g2_fill_2 FILLER_38_221 ();
 sg13g2_decap_8 FILLER_38_227 ();
 sg13g2_decap_4 FILLER_38_247 ();
 sg13g2_decap_8 FILLER_38_277 ();
 sg13g2_decap_8 FILLER_38_284 ();
 sg13g2_fill_2 FILLER_38_291 ();
 sg13g2_decap_4 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_decap_8 FILLER_38_316 ();
 sg13g2_decap_8 FILLER_38_323 ();
 sg13g2_decap_8 FILLER_38_330 ();
 sg13g2_decap_8 FILLER_38_337 ();
 sg13g2_decap_8 FILLER_38_344 ();
 sg13g2_decap_8 FILLER_38_351 ();
 sg13g2_decap_8 FILLER_38_358 ();
 sg13g2_decap_8 FILLER_38_365 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_fill_1 FILLER_39_61 ();
 sg13g2_fill_2 FILLER_39_71 ();
 sg13g2_decap_4 FILLER_39_99 ();
 sg13g2_fill_1 FILLER_39_103 ();
 sg13g2_fill_2 FILLER_39_109 ();
 sg13g2_fill_2 FILLER_39_119 ();
 sg13g2_fill_1 FILLER_39_121 ();
 sg13g2_fill_1 FILLER_39_126 ();
 sg13g2_fill_2 FILLER_39_135 ();
 sg13g2_fill_2 FILLER_39_146 ();
 sg13g2_fill_2 FILLER_39_191 ();
 sg13g2_fill_2 FILLER_39_197 ();
 sg13g2_decap_8 FILLER_39_240 ();
 sg13g2_decap_8 FILLER_39_247 ();
 sg13g2_decap_8 FILLER_39_254 ();
 sg13g2_fill_1 FILLER_39_261 ();
 sg13g2_fill_2 FILLER_39_270 ();
 sg13g2_decap_4 FILLER_39_281 ();
 sg13g2_decap_8 FILLER_39_320 ();
 sg13g2_decap_8 FILLER_39_327 ();
 sg13g2_decap_8 FILLER_39_334 ();
 sg13g2_decap_8 FILLER_39_341 ();
 sg13g2_decap_8 FILLER_39_348 ();
 sg13g2_decap_8 FILLER_39_355 ();
 sg13g2_decap_8 FILLER_39_362 ();
 sg13g2_decap_8 FILLER_39_369 ();
 sg13g2_decap_8 FILLER_39_376 ();
 sg13g2_decap_8 FILLER_39_383 ();
 sg13g2_decap_8 FILLER_39_390 ();
 sg13g2_decap_8 FILLER_39_397 ();
 sg13g2_decap_4 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_4 FILLER_40_28 ();
 sg13g2_fill_2 FILLER_40_66 ();
 sg13g2_fill_1 FILLER_40_68 ();
 sg13g2_fill_2 FILLER_40_78 ();
 sg13g2_decap_8 FILLER_40_142 ();
 sg13g2_decap_8 FILLER_40_149 ();
 sg13g2_fill_2 FILLER_40_156 ();
 sg13g2_fill_1 FILLER_40_158 ();
 sg13g2_fill_2 FILLER_40_168 ();
 sg13g2_fill_1 FILLER_40_170 ();
 sg13g2_fill_2 FILLER_40_180 ();
 sg13g2_decap_8 FILLER_40_190 ();
 sg13g2_fill_1 FILLER_40_223 ();
 sg13g2_fill_1 FILLER_40_243 ();
 sg13g2_fill_2 FILLER_40_264 ();
 sg13g2_fill_1 FILLER_40_266 ();
 sg13g2_fill_1 FILLER_40_271 ();
 sg13g2_fill_2 FILLER_40_315 ();
 sg13g2_fill_1 FILLER_40_317 ();
 sg13g2_decap_8 FILLER_40_326 ();
 sg13g2_decap_8 FILLER_40_333 ();
 sg13g2_decap_8 FILLER_40_340 ();
 sg13g2_decap_8 FILLER_40_347 ();
 sg13g2_decap_8 FILLER_40_354 ();
 sg13g2_decap_8 FILLER_40_361 ();
 sg13g2_decap_8 FILLER_40_368 ();
 sg13g2_decap_8 FILLER_40_375 ();
 sg13g2_decap_8 FILLER_40_382 ();
 sg13g2_decap_8 FILLER_40_389 ();
 sg13g2_decap_8 FILLER_40_396 ();
 sg13g2_decap_4 FILLER_40_403 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_4 FILLER_41_21 ();
 sg13g2_fill_1 FILLER_41_25 ();
 sg13g2_decap_8 FILLER_41_87 ();
 sg13g2_fill_2 FILLER_41_94 ();
 sg13g2_decap_8 FILLER_41_152 ();
 sg13g2_decap_8 FILLER_41_159 ();
 sg13g2_decap_8 FILLER_41_166 ();
 sg13g2_fill_2 FILLER_41_173 ();
 sg13g2_fill_1 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_195 ();
 sg13g2_fill_2 FILLER_41_216 ();
 sg13g2_fill_1 FILLER_41_218 ();
 sg13g2_fill_2 FILLER_41_234 ();
 sg13g2_decap_4 FILLER_41_302 ();
 sg13g2_fill_1 FILLER_41_306 ();
 sg13g2_decap_8 FILLER_41_342 ();
 sg13g2_decap_8 FILLER_41_349 ();
 sg13g2_decap_8 FILLER_41_356 ();
 sg13g2_decap_8 FILLER_41_363 ();
 sg13g2_decap_8 FILLER_41_370 ();
 sg13g2_decap_8 FILLER_41_377 ();
 sg13g2_decap_8 FILLER_41_384 ();
 sg13g2_decap_8 FILLER_41_391 ();
 sg13g2_decap_8 FILLER_41_398 ();
 sg13g2_decap_4 FILLER_41_405 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_fill_2 FILLER_42_21 ();
 sg13g2_fill_2 FILLER_42_101 ();
 sg13g2_fill_1 FILLER_42_103 ();
 sg13g2_fill_2 FILLER_42_145 ();
 sg13g2_fill_2 FILLER_42_155 ();
 sg13g2_decap_4 FILLER_42_203 ();
 sg13g2_fill_2 FILLER_42_207 ();
 sg13g2_fill_2 FILLER_42_217 ();
 sg13g2_fill_2 FILLER_42_272 ();
 sg13g2_fill_1 FILLER_42_279 ();
 sg13g2_fill_1 FILLER_42_285 ();
 sg13g2_fill_1 FILLER_42_296 ();
 sg13g2_fill_2 FILLER_42_302 ();
 sg13g2_fill_1 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_335 ();
 sg13g2_decap_8 FILLER_42_342 ();
 sg13g2_decap_8 FILLER_42_349 ();
 sg13g2_decap_8 FILLER_42_356 ();
 sg13g2_decap_8 FILLER_42_363 ();
 sg13g2_decap_8 FILLER_42_370 ();
 sg13g2_decap_8 FILLER_42_377 ();
 sg13g2_decap_8 FILLER_42_384 ();
 sg13g2_decap_8 FILLER_42_391 ();
 sg13g2_decap_8 FILLER_42_398 ();
 sg13g2_decap_4 FILLER_42_405 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_fill_2 FILLER_43_28 ();
 sg13g2_fill_2 FILLER_43_38 ();
 sg13g2_fill_2 FILLER_43_49 ();
 sg13g2_fill_1 FILLER_43_76 ();
 sg13g2_fill_2 FILLER_43_113 ();
 sg13g2_fill_1 FILLER_43_115 ();
 sg13g2_fill_2 FILLER_43_161 ();
 sg13g2_fill_1 FILLER_43_163 ();
 sg13g2_fill_2 FILLER_43_172 ();
 sg13g2_fill_1 FILLER_43_174 ();
 sg13g2_fill_2 FILLER_43_180 ();
 sg13g2_fill_2 FILLER_43_213 ();
 sg13g2_decap_4 FILLER_43_220 ();
 sg13g2_fill_2 FILLER_43_224 ();
 sg13g2_decap_4 FILLER_43_231 ();
 sg13g2_fill_1 FILLER_43_239 ();
 sg13g2_fill_2 FILLER_43_253 ();
 sg13g2_fill_2 FILLER_43_265 ();
 sg13g2_fill_1 FILLER_43_271 ();
 sg13g2_decap_8 FILLER_43_345 ();
 sg13g2_decap_8 FILLER_43_352 ();
 sg13g2_decap_8 FILLER_43_359 ();
 sg13g2_decap_8 FILLER_43_366 ();
 sg13g2_decap_8 FILLER_43_373 ();
 sg13g2_decap_8 FILLER_43_380 ();
 sg13g2_decap_8 FILLER_43_387 ();
 sg13g2_decap_8 FILLER_43_394 ();
 sg13g2_decap_8 FILLER_43_401 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_fill_2 FILLER_44_21 ();
 sg13g2_fill_1 FILLER_44_23 ();
 sg13g2_decap_8 FILLER_44_50 ();
 sg13g2_fill_2 FILLER_44_57 ();
 sg13g2_decap_8 FILLER_44_67 ();
 sg13g2_fill_2 FILLER_44_74 ();
 sg13g2_fill_2 FILLER_44_129 ();
 sg13g2_fill_1 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_153 ();
 sg13g2_decap_4 FILLER_44_160 ();
 sg13g2_fill_2 FILLER_44_219 ();
 sg13g2_fill_1 FILLER_44_221 ();
 sg13g2_decap_8 FILLER_44_256 ();
 sg13g2_decap_8 FILLER_44_263 ();
 sg13g2_fill_1 FILLER_44_274 ();
 sg13g2_fill_2 FILLER_44_328 ();
 sg13g2_decap_8 FILLER_44_343 ();
 sg13g2_decap_8 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_fill_2 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_14 ();
 sg13g2_fill_2 FILLER_45_64 ();
 sg13g2_fill_1 FILLER_45_66 ();
 sg13g2_fill_1 FILLER_45_71 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_fill_1 FILLER_45_84 ();
 sg13g2_fill_1 FILLER_45_106 ();
 sg13g2_fill_2 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_165 ();
 sg13g2_decap_4 FILLER_45_172 ();
 sg13g2_fill_2 FILLER_45_176 ();
 sg13g2_fill_1 FILLER_45_234 ();
 sg13g2_decap_8 FILLER_45_257 ();
 sg13g2_decap_8 FILLER_45_264 ();
 sg13g2_decap_8 FILLER_45_271 ();
 sg13g2_decap_4 FILLER_45_278 ();
 sg13g2_fill_1 FILLER_45_290 ();
 sg13g2_fill_2 FILLER_45_308 ();
 sg13g2_fill_1 FILLER_45_310 ();
 sg13g2_decap_8 FILLER_45_333 ();
 sg13g2_decap_8 FILLER_45_340 ();
 sg13g2_decap_8 FILLER_45_347 ();
 sg13g2_decap_8 FILLER_45_354 ();
 sg13g2_decap_8 FILLER_45_361 ();
 sg13g2_decap_8 FILLER_45_368 ();
 sg13g2_decap_8 FILLER_45_375 ();
 sg13g2_decap_8 FILLER_45_382 ();
 sg13g2_decap_8 FILLER_45_389 ();
 sg13g2_decap_8 FILLER_45_396 ();
 sg13g2_decap_4 FILLER_45_403 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_fill_1 FILLER_46_73 ();
 sg13g2_fill_2 FILLER_46_79 ();
 sg13g2_fill_1 FILLER_46_81 ();
 sg13g2_fill_2 FILLER_46_87 ();
 sg13g2_fill_1 FILLER_46_89 ();
 sg13g2_decap_8 FILLER_46_94 ();
 sg13g2_decap_4 FILLER_46_106 ();
 sg13g2_fill_2 FILLER_46_124 ();
 sg13g2_fill_2 FILLER_46_186 ();
 sg13g2_fill_1 FILLER_46_188 ();
 sg13g2_fill_1 FILLER_46_201 ();
 sg13g2_fill_1 FILLER_46_224 ();
 sg13g2_fill_1 FILLER_46_231 ();
 sg13g2_fill_2 FILLER_46_253 ();
 sg13g2_decap_4 FILLER_46_300 ();
 sg13g2_decap_8 FILLER_46_333 ();
 sg13g2_decap_8 FILLER_46_340 ();
 sg13g2_decap_8 FILLER_46_347 ();
 sg13g2_decap_8 FILLER_46_354 ();
 sg13g2_decap_8 FILLER_46_361 ();
 sg13g2_decap_8 FILLER_46_368 ();
 sg13g2_decap_8 FILLER_46_375 ();
 sg13g2_decap_8 FILLER_46_382 ();
 sg13g2_decap_8 FILLER_46_389 ();
 sg13g2_decap_8 FILLER_46_396 ();
 sg13g2_decap_4 FILLER_46_403 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_4 FILLER_47_14 ();
 sg13g2_fill_1 FILLER_47_18 ();
 sg13g2_fill_2 FILLER_47_48 ();
 sg13g2_fill_1 FILLER_47_64 ();
 sg13g2_decap_8 FILLER_47_92 ();
 sg13g2_fill_2 FILLER_47_99 ();
 sg13g2_fill_1 FILLER_47_101 ();
 sg13g2_fill_1 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_128 ();
 sg13g2_decap_8 FILLER_47_135 ();
 sg13g2_fill_2 FILLER_47_176 ();
 sg13g2_fill_1 FILLER_47_178 ();
 sg13g2_decap_4 FILLER_47_213 ();
 sg13g2_fill_1 FILLER_47_217 ();
 sg13g2_fill_2 FILLER_47_227 ();
 sg13g2_fill_1 FILLER_47_229 ();
 sg13g2_fill_2 FILLER_47_275 ();
 sg13g2_fill_1 FILLER_47_277 ();
 sg13g2_fill_2 FILLER_47_283 ();
 sg13g2_fill_1 FILLER_47_285 ();
 sg13g2_fill_1 FILLER_47_317 ();
 sg13g2_decap_8 FILLER_47_344 ();
 sg13g2_decap_8 FILLER_47_351 ();
 sg13g2_decap_8 FILLER_47_358 ();
 sg13g2_decap_8 FILLER_47_365 ();
 sg13g2_decap_8 FILLER_47_372 ();
 sg13g2_decap_8 FILLER_47_379 ();
 sg13g2_decap_8 FILLER_47_386 ();
 sg13g2_decap_8 FILLER_47_393 ();
 sg13g2_decap_8 FILLER_47_400 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_fill_2 FILLER_48_67 ();
 sg13g2_fill_2 FILLER_48_109 ();
 sg13g2_fill_1 FILLER_48_127 ();
 sg13g2_decap_8 FILLER_48_136 ();
 sg13g2_decap_4 FILLER_48_143 ();
 sg13g2_fill_1 FILLER_48_147 ();
 sg13g2_fill_2 FILLER_48_186 ();
 sg13g2_fill_1 FILLER_48_205 ();
 sg13g2_fill_2 FILLER_48_219 ();
 sg13g2_decap_4 FILLER_48_226 ();
 sg13g2_fill_2 FILLER_48_230 ();
 sg13g2_fill_1 FILLER_48_282 ();
 sg13g2_fill_2 FILLER_48_296 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_fill_2 FILLER_48_406 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_4 FILLER_49_14 ();
 sg13g2_fill_2 FILLER_49_18 ();
 sg13g2_fill_2 FILLER_49_46 ();
 sg13g2_fill_1 FILLER_49_48 ();
 sg13g2_fill_2 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_150 ();
 sg13g2_fill_1 FILLER_49_157 ();
 sg13g2_fill_2 FILLER_49_163 ();
 sg13g2_fill_1 FILLER_49_165 ();
 sg13g2_fill_1 FILLER_49_193 ();
 sg13g2_decap_8 FILLER_49_212 ();
 sg13g2_fill_1 FILLER_49_219 ();
 sg13g2_fill_2 FILLER_49_225 ();
 sg13g2_fill_2 FILLER_49_244 ();
 sg13g2_fill_2 FILLER_49_256 ();
 sg13g2_fill_1 FILLER_49_271 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_decap_8 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_fill_2 FILLER_50_14 ();
 sg13g2_fill_1 FILLER_50_16 ();
 sg13g2_fill_2 FILLER_50_47 ();
 sg13g2_fill_1 FILLER_50_49 ();
 sg13g2_fill_2 FILLER_50_75 ();
 sg13g2_fill_1 FILLER_50_118 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_fill_2 FILLER_50_152 ();
 sg13g2_decap_8 FILLER_50_159 ();
 sg13g2_decap_4 FILLER_50_166 ();
 sg13g2_fill_1 FILLER_50_170 ();
 sg13g2_decap_4 FILLER_50_210 ();
 sg13g2_fill_1 FILLER_50_214 ();
 sg13g2_decap_8 FILLER_50_250 ();
 sg13g2_fill_2 FILLER_50_257 ();
 sg13g2_fill_1 FILLER_50_259 ();
 sg13g2_decap_8 FILLER_50_265 ();
 sg13g2_fill_2 FILLER_50_272 ();
 sg13g2_fill_1 FILLER_50_323 ();
 sg13g2_fill_1 FILLER_50_328 ();
 sg13g2_decap_8 FILLER_50_342 ();
 sg13g2_decap_8 FILLER_50_349 ();
 sg13g2_decap_8 FILLER_50_356 ();
 sg13g2_decap_8 FILLER_50_363 ();
 sg13g2_decap_8 FILLER_50_370 ();
 sg13g2_decap_8 FILLER_50_377 ();
 sg13g2_decap_8 FILLER_50_384 ();
 sg13g2_decap_8 FILLER_50_391 ();
 sg13g2_decap_8 FILLER_50_398 ();
 sg13g2_decap_4 FILLER_50_405 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_4 FILLER_51_14 ();
 sg13g2_fill_1 FILLER_51_18 ();
 sg13g2_fill_2 FILLER_51_85 ();
 sg13g2_fill_1 FILLER_51_87 ();
 sg13g2_fill_2 FILLER_51_102 ();
 sg13g2_fill_1 FILLER_51_104 ();
 sg13g2_decap_4 FILLER_51_119 ();
 sg13g2_fill_2 FILLER_51_123 ();
 sg13g2_fill_2 FILLER_51_133 ();
 sg13g2_fill_2 FILLER_51_151 ();
 sg13g2_fill_1 FILLER_51_153 ();
 sg13g2_decap_8 FILLER_51_164 ();
 sg13g2_decap_8 FILLER_51_171 ();
 sg13g2_decap_4 FILLER_51_178 ();
 sg13g2_decap_4 FILLER_51_187 ();
 sg13g2_fill_1 FILLER_51_191 ();
 sg13g2_fill_1 FILLER_51_209 ();
 sg13g2_fill_2 FILLER_51_215 ();
 sg13g2_fill_2 FILLER_51_221 ();
 sg13g2_fill_2 FILLER_51_231 ();
 sg13g2_decap_4 FILLER_51_251 ();
 sg13g2_fill_2 FILLER_51_255 ();
 sg13g2_fill_1 FILLER_51_268 ();
 sg13g2_fill_1 FILLER_51_289 ();
 sg13g2_decap_8 FILLER_51_293 ();
 sg13g2_decap_8 FILLER_51_300 ();
 sg13g2_decap_8 FILLER_51_307 ();
 sg13g2_decap_8 FILLER_51_314 ();
 sg13g2_decap_8 FILLER_51_321 ();
 sg13g2_decap_8 FILLER_51_328 ();
 sg13g2_decap_8 FILLER_51_335 ();
 sg13g2_decap_8 FILLER_51_342 ();
 sg13g2_decap_8 FILLER_51_349 ();
 sg13g2_decap_8 FILLER_51_356 ();
 sg13g2_decap_8 FILLER_51_363 ();
 sg13g2_decap_8 FILLER_51_370 ();
 sg13g2_decap_8 FILLER_51_377 ();
 sg13g2_decap_8 FILLER_51_384 ();
 sg13g2_decap_8 FILLER_51_391 ();
 sg13g2_decap_8 FILLER_51_398 ();
 sg13g2_decap_4 FILLER_51_405 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_4 FILLER_52_28 ();
 sg13g2_fill_2 FILLER_52_36 ();
 sg13g2_decap_4 FILLER_52_47 ();
 sg13g2_decap_4 FILLER_52_55 ();
 sg13g2_fill_1 FILLER_52_59 ();
 sg13g2_fill_2 FILLER_52_73 ();
 sg13g2_fill_2 FILLER_52_92 ();
 sg13g2_fill_1 FILLER_52_94 ();
 sg13g2_fill_2 FILLER_52_127 ();
 sg13g2_decap_8 FILLER_52_174 ();
 sg13g2_decap_8 FILLER_52_181 ();
 sg13g2_fill_1 FILLER_52_197 ();
 sg13g2_fill_2 FILLER_52_207 ();
 sg13g2_fill_1 FILLER_52_244 ();
 sg13g2_fill_2 FILLER_52_255 ();
 sg13g2_fill_1 FILLER_52_257 ();
 sg13g2_fill_1 FILLER_52_286 ();
 sg13g2_fill_2 FILLER_52_317 ();
 sg13g2_fill_1 FILLER_52_319 ();
 sg13g2_decap_8 FILLER_52_350 ();
 sg13g2_decap_8 FILLER_52_357 ();
 sg13g2_decap_8 FILLER_52_364 ();
 sg13g2_decap_8 FILLER_52_371 ();
 sg13g2_decap_8 FILLER_52_378 ();
 sg13g2_decap_8 FILLER_52_385 ();
 sg13g2_decap_8 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_fill_2 FILLER_52_406 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_40 ();
 sg13g2_decap_4 FILLER_53_47 ();
 sg13g2_fill_1 FILLER_53_51 ();
 sg13g2_decap_4 FILLER_53_124 ();
 sg13g2_decap_8 FILLER_53_136 ();
 sg13g2_decap_4 FILLER_53_143 ();
 sg13g2_decap_4 FILLER_53_167 ();
 sg13g2_fill_1 FILLER_53_171 ();
 sg13g2_decap_8 FILLER_53_188 ();
 sg13g2_fill_2 FILLER_53_195 ();
 sg13g2_fill_2 FILLER_53_228 ();
 sg13g2_fill_1 FILLER_53_230 ();
 sg13g2_fill_2 FILLER_53_234 ();
 sg13g2_fill_1 FILLER_53_236 ();
 sg13g2_fill_2 FILLER_53_250 ();
 sg13g2_fill_1 FILLER_53_252 ();
 sg13g2_decap_8 FILLER_53_357 ();
 sg13g2_decap_8 FILLER_53_364 ();
 sg13g2_decap_8 FILLER_53_371 ();
 sg13g2_decap_8 FILLER_53_378 ();
 sg13g2_decap_8 FILLER_53_385 ();
 sg13g2_decap_8 FILLER_53_392 ();
 sg13g2_decap_8 FILLER_53_399 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_4 FILLER_54_21 ();
 sg13g2_fill_1 FILLER_54_25 ();
 sg13g2_fill_2 FILLER_54_52 ();
 sg13g2_fill_1 FILLER_54_54 ();
 sg13g2_fill_2 FILLER_54_80 ();
 sg13g2_fill_1 FILLER_54_82 ();
 sg13g2_fill_2 FILLER_54_88 ();
 sg13g2_fill_2 FILLER_54_99 ();
 sg13g2_fill_2 FILLER_54_110 ();
 sg13g2_decap_4 FILLER_54_152 ();
 sg13g2_decap_4 FILLER_54_192 ();
 sg13g2_fill_1 FILLER_54_196 ();
 sg13g2_fill_2 FILLER_54_202 ();
 sg13g2_fill_1 FILLER_54_204 ();
 sg13g2_decap_8 FILLER_54_219 ();
 sg13g2_decap_8 FILLER_54_226 ();
 sg13g2_decap_4 FILLER_54_233 ();
 sg13g2_fill_2 FILLER_54_237 ();
 sg13g2_fill_2 FILLER_54_258 ();
 sg13g2_fill_1 FILLER_54_264 ();
 sg13g2_fill_2 FILLER_54_274 ();
 sg13g2_fill_1 FILLER_54_276 ();
 sg13g2_fill_2 FILLER_54_292 ();
 sg13g2_fill_1 FILLER_54_294 ();
 sg13g2_fill_1 FILLER_54_304 ();
 sg13g2_decap_8 FILLER_54_348 ();
 sg13g2_decap_8 FILLER_54_355 ();
 sg13g2_decap_8 FILLER_54_362 ();
 sg13g2_decap_8 FILLER_54_369 ();
 sg13g2_decap_8 FILLER_54_376 ();
 sg13g2_decap_8 FILLER_54_383 ();
 sg13g2_decap_8 FILLER_54_390 ();
 sg13g2_decap_8 FILLER_54_397 ();
 sg13g2_decap_4 FILLER_54_404 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_fill_2 FILLER_55_85 ();
 sg13g2_decap_4 FILLER_55_100 ();
 sg13g2_fill_1 FILLER_55_104 ();
 sg13g2_decap_4 FILLER_55_122 ();
 sg13g2_fill_2 FILLER_55_126 ();
 sg13g2_decap_4 FILLER_55_132 ();
 sg13g2_fill_1 FILLER_55_136 ();
 sg13g2_fill_2 FILLER_55_142 ();
 sg13g2_fill_1 FILLER_55_144 ();
 sg13g2_fill_2 FILLER_55_174 ();
 sg13g2_decap_8 FILLER_55_215 ();
 sg13g2_decap_8 FILLER_55_222 ();
 sg13g2_fill_2 FILLER_55_229 ();
 sg13g2_fill_2 FILLER_55_247 ();
 sg13g2_decap_8 FILLER_55_257 ();
 sg13g2_decap_4 FILLER_55_268 ();
 sg13g2_fill_2 FILLER_55_272 ();
 sg13g2_fill_1 FILLER_55_279 ();
 sg13g2_fill_2 FILLER_55_290 ();
 sg13g2_fill_1 FILLER_55_292 ();
 sg13g2_fill_2 FILLER_55_310 ();
 sg13g2_fill_1 FILLER_55_312 ();
 sg13g2_decap_8 FILLER_55_339 ();
 sg13g2_decap_8 FILLER_55_346 ();
 sg13g2_decap_8 FILLER_55_353 ();
 sg13g2_decap_8 FILLER_55_360 ();
 sg13g2_decap_8 FILLER_55_367 ();
 sg13g2_decap_8 FILLER_55_374 ();
 sg13g2_decap_8 FILLER_55_381 ();
 sg13g2_decap_8 FILLER_55_388 ();
 sg13g2_decap_8 FILLER_55_395 ();
 sg13g2_decap_8 FILLER_55_402 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_fill_2 FILLER_56_75 ();
 sg13g2_fill_1 FILLER_56_77 ();
 sg13g2_decap_4 FILLER_56_109 ();
 sg13g2_fill_2 FILLER_56_113 ();
 sg13g2_fill_1 FILLER_56_119 ();
 sg13g2_decap_4 FILLER_56_125 ();
 sg13g2_fill_2 FILLER_56_141 ();
 sg13g2_decap_4 FILLER_56_151 ();
 sg13g2_fill_2 FILLER_56_163 ();
 sg13g2_fill_1 FILLER_56_165 ();
 sg13g2_decap_8 FILLER_56_192 ();
 sg13g2_decap_4 FILLER_56_199 ();
 sg13g2_fill_2 FILLER_56_203 ();
 sg13g2_decap_8 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_217 ();
 sg13g2_fill_2 FILLER_56_224 ();
 sg13g2_decap_4 FILLER_56_244 ();
 sg13g2_fill_2 FILLER_56_248 ();
 sg13g2_decap_8 FILLER_56_278 ();
 sg13g2_fill_2 FILLER_56_285 ();
 sg13g2_fill_1 FILLER_56_287 ();
 sg13g2_fill_1 FILLER_56_301 ();
 sg13g2_fill_1 FILLER_56_315 ();
 sg13g2_decap_8 FILLER_56_338 ();
 sg13g2_decap_8 FILLER_56_345 ();
 sg13g2_decap_8 FILLER_56_352 ();
 sg13g2_decap_8 FILLER_56_359 ();
 sg13g2_decap_8 FILLER_56_366 ();
 sg13g2_decap_8 FILLER_56_373 ();
 sg13g2_decap_8 FILLER_56_380 ();
 sg13g2_decap_8 FILLER_56_387 ();
 sg13g2_decap_8 FILLER_56_394 ();
 sg13g2_decap_8 FILLER_56_401 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_4 FILLER_57_28 ();
 sg13g2_fill_1 FILLER_57_32 ();
 sg13g2_fill_1 FILLER_57_59 ();
 sg13g2_fill_1 FILLER_57_90 ();
 sg13g2_fill_1 FILLER_57_96 ();
 sg13g2_fill_1 FILLER_57_136 ();
 sg13g2_decap_4 FILLER_57_168 ();
 sg13g2_fill_2 FILLER_57_182 ();
 sg13g2_decap_8 FILLER_57_194 ();
 sg13g2_fill_1 FILLER_57_201 ();
 sg13g2_fill_2 FILLER_57_218 ();
 sg13g2_fill_1 FILLER_57_220 ();
 sg13g2_fill_1 FILLER_57_233 ();
 sg13g2_fill_1 FILLER_57_252 ();
 sg13g2_decap_4 FILLER_57_288 ();
 sg13g2_fill_1 FILLER_57_292 ();
 sg13g2_decap_8 FILLER_57_323 ();
 sg13g2_decap_8 FILLER_57_330 ();
 sg13g2_decap_8 FILLER_57_337 ();
 sg13g2_decap_8 FILLER_57_344 ();
 sg13g2_decap_8 FILLER_57_351 ();
 sg13g2_decap_8 FILLER_57_358 ();
 sg13g2_decap_8 FILLER_57_365 ();
 sg13g2_decap_8 FILLER_57_372 ();
 sg13g2_decap_8 FILLER_57_379 ();
 sg13g2_decap_8 FILLER_57_386 ();
 sg13g2_decap_8 FILLER_57_393 ();
 sg13g2_decap_8 FILLER_57_400 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_4 FILLER_58_28 ();
 sg13g2_fill_1 FILLER_58_32 ();
 sg13g2_decap_8 FILLER_58_50 ();
 sg13g2_decap_8 FILLER_58_57 ();
 sg13g2_fill_1 FILLER_58_64 ();
 sg13g2_fill_2 FILLER_58_79 ();
 sg13g2_fill_2 FILLER_58_163 ();
 sg13g2_fill_2 FILLER_58_173 ();
 sg13g2_fill_1 FILLER_58_175 ();
 sg13g2_fill_2 FILLER_58_274 ();
 sg13g2_fill_2 FILLER_58_297 ();
 sg13g2_decap_8 FILLER_58_320 ();
 sg13g2_decap_8 FILLER_58_327 ();
 sg13g2_decap_8 FILLER_58_334 ();
 sg13g2_decap_8 FILLER_58_341 ();
 sg13g2_decap_8 FILLER_58_348 ();
 sg13g2_decap_8 FILLER_58_355 ();
 sg13g2_decap_8 FILLER_58_362 ();
 sg13g2_decap_8 FILLER_58_369 ();
 sg13g2_decap_8 FILLER_58_376 ();
 sg13g2_decap_8 FILLER_58_383 ();
 sg13g2_decap_8 FILLER_58_390 ();
 sg13g2_decap_8 FILLER_58_397 ();
 sg13g2_decap_4 FILLER_58_404 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_61 ();
 sg13g2_decap_8 FILLER_59_68 ();
 sg13g2_fill_1 FILLER_59_75 ();
 sg13g2_decap_4 FILLER_59_85 ();
 sg13g2_decap_4 FILLER_59_93 ();
 sg13g2_fill_1 FILLER_59_97 ();
 sg13g2_decap_8 FILLER_59_123 ();
 sg13g2_fill_2 FILLER_59_130 ();
 sg13g2_fill_1 FILLER_59_132 ();
 sg13g2_decap_8 FILLER_59_137 ();
 sg13g2_decap_4 FILLER_59_144 ();
 sg13g2_fill_2 FILLER_59_148 ();
 sg13g2_decap_4 FILLER_59_159 ();
 sg13g2_fill_2 FILLER_59_182 ();
 sg13g2_decap_8 FILLER_59_194 ();
 sg13g2_decap_4 FILLER_59_201 ();
 sg13g2_fill_2 FILLER_59_205 ();
 sg13g2_fill_2 FILLER_59_212 ();
 sg13g2_fill_1 FILLER_59_214 ();
 sg13g2_decap_4 FILLER_59_232 ();
 sg13g2_decap_8 FILLER_59_337 ();
 sg13g2_decap_8 FILLER_59_344 ();
 sg13g2_decap_8 FILLER_59_351 ();
 sg13g2_decap_8 FILLER_59_358 ();
 sg13g2_decap_8 FILLER_59_365 ();
 sg13g2_decap_8 FILLER_59_372 ();
 sg13g2_decap_8 FILLER_59_379 ();
 sg13g2_decap_8 FILLER_59_386 ();
 sg13g2_decap_8 FILLER_59_393 ();
 sg13g2_decap_8 FILLER_59_400 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_4 FILLER_60_87 ();
 sg13g2_fill_1 FILLER_60_126 ();
 sg13g2_decap_8 FILLER_60_131 ();
 sg13g2_decap_8 FILLER_60_150 ();
 sg13g2_fill_2 FILLER_60_157 ();
 sg13g2_fill_1 FILLER_60_159 ();
 sg13g2_fill_2 FILLER_60_176 ();
 sg13g2_fill_1 FILLER_60_178 ();
 sg13g2_decap_8 FILLER_60_187 ();
 sg13g2_decap_4 FILLER_60_194 ();
 sg13g2_decap_8 FILLER_60_203 ();
 sg13g2_fill_2 FILLER_60_210 ();
 sg13g2_fill_1 FILLER_60_217 ();
 sg13g2_fill_2 FILLER_60_237 ();
 sg13g2_fill_2 FILLER_60_284 ();
 sg13g2_fill_1 FILLER_60_286 ();
 sg13g2_fill_2 FILLER_60_296 ();
 sg13g2_decap_8 FILLER_60_332 ();
 sg13g2_decap_8 FILLER_60_339 ();
 sg13g2_decap_8 FILLER_60_346 ();
 sg13g2_decap_8 FILLER_60_353 ();
 sg13g2_decap_8 FILLER_60_360 ();
 sg13g2_decap_8 FILLER_60_367 ();
 sg13g2_decap_8 FILLER_60_374 ();
 sg13g2_decap_8 FILLER_60_381 ();
 sg13g2_decap_8 FILLER_60_388 ();
 sg13g2_decap_8 FILLER_60_395 ();
 sg13g2_decap_8 FILLER_60_402 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_fill_1 FILLER_61_21 ();
 sg13g2_fill_2 FILLER_61_65 ();
 sg13g2_fill_1 FILLER_61_67 ();
 sg13g2_fill_1 FILLER_61_114 ();
 sg13g2_fill_2 FILLER_61_120 ();
 sg13g2_fill_2 FILLER_61_156 ();
 sg13g2_decap_4 FILLER_61_178 ();
 sg13g2_decap_8 FILLER_61_243 ();
 sg13g2_decap_8 FILLER_61_250 ();
 sg13g2_decap_8 FILLER_61_257 ();
 sg13g2_decap_4 FILLER_61_264 ();
 sg13g2_fill_1 FILLER_61_286 ();
 sg13g2_decap_8 FILLER_61_339 ();
 sg13g2_decap_8 FILLER_61_346 ();
 sg13g2_decap_8 FILLER_61_353 ();
 sg13g2_decap_8 FILLER_61_360 ();
 sg13g2_decap_8 FILLER_61_367 ();
 sg13g2_decap_8 FILLER_61_374 ();
 sg13g2_decap_8 FILLER_61_381 ();
 sg13g2_decap_8 FILLER_61_388 ();
 sg13g2_decap_8 FILLER_61_395 ();
 sg13g2_decap_8 FILLER_61_402 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_4 FILLER_62_21 ();
 sg13g2_fill_2 FILLER_62_25 ();
 sg13g2_fill_2 FILLER_62_48 ();
 sg13g2_fill_1 FILLER_62_50 ();
 sg13g2_fill_2 FILLER_62_77 ();
 sg13g2_fill_1 FILLER_62_79 ();
 sg13g2_fill_2 FILLER_62_111 ();
 sg13g2_fill_1 FILLER_62_147 ();
 sg13g2_decap_4 FILLER_62_170 ();
 sg13g2_decap_4 FILLER_62_180 ();
 sg13g2_fill_1 FILLER_62_184 ();
 sg13g2_decap_4 FILLER_62_190 ();
 sg13g2_fill_1 FILLER_62_224 ();
 sg13g2_decap_8 FILLER_62_238 ();
 sg13g2_fill_2 FILLER_62_249 ();
 sg13g2_decap_8 FILLER_62_255 ();
 sg13g2_decap_8 FILLER_62_266 ();
 sg13g2_fill_2 FILLER_62_273 ();
 sg13g2_fill_2 FILLER_62_293 ();
 sg13g2_decap_8 FILLER_62_308 ();
 sg13g2_fill_1 FILLER_62_315 ();
 sg13g2_decap_8 FILLER_62_329 ();
 sg13g2_decap_8 FILLER_62_336 ();
 sg13g2_decap_8 FILLER_62_343 ();
 sg13g2_decap_8 FILLER_62_350 ();
 sg13g2_decap_8 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_364 ();
 sg13g2_decap_8 FILLER_62_371 ();
 sg13g2_decap_8 FILLER_62_378 ();
 sg13g2_decap_8 FILLER_62_385 ();
 sg13g2_decap_8 FILLER_62_392 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_4 FILLER_63_42 ();
 sg13g2_fill_2 FILLER_63_59 ();
 sg13g2_fill_1 FILLER_63_61 ();
 sg13g2_fill_2 FILLER_63_93 ();
 sg13g2_fill_1 FILLER_63_95 ();
 sg13g2_fill_2 FILLER_63_118 ();
 sg13g2_fill_1 FILLER_63_128 ();
 sg13g2_decap_4 FILLER_63_137 ();
 sg13g2_decap_8 FILLER_63_156 ();
 sg13g2_decap_8 FILLER_63_163 ();
 sg13g2_fill_2 FILLER_63_196 ();
 sg13g2_fill_1 FILLER_63_198 ();
 sg13g2_decap_4 FILLER_63_204 ();
 sg13g2_decap_4 FILLER_63_217 ();
 sg13g2_fill_2 FILLER_63_221 ();
 sg13g2_fill_2 FILLER_63_228 ();
 sg13g2_fill_1 FILLER_63_245 ();
 sg13g2_fill_1 FILLER_63_254 ();
 sg13g2_decap_4 FILLER_63_300 ();
 sg13g2_decap_8 FILLER_63_316 ();
 sg13g2_decap_8 FILLER_63_323 ();
 sg13g2_decap_8 FILLER_63_330 ();
 sg13g2_decap_8 FILLER_63_337 ();
 sg13g2_decap_8 FILLER_63_344 ();
 sg13g2_decap_8 FILLER_63_351 ();
 sg13g2_decap_8 FILLER_63_358 ();
 sg13g2_decap_8 FILLER_63_365 ();
 sg13g2_decap_8 FILLER_63_372 ();
 sg13g2_decap_8 FILLER_63_379 ();
 sg13g2_decap_8 FILLER_63_386 ();
 sg13g2_decap_8 FILLER_63_393 ();
 sg13g2_decap_8 FILLER_63_400 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_4 FILLER_64_49 ();
 sg13g2_fill_1 FILLER_64_61 ();
 sg13g2_decap_4 FILLER_64_79 ();
 sg13g2_fill_2 FILLER_64_88 ();
 sg13g2_fill_2 FILLER_64_108 ();
 sg13g2_fill_1 FILLER_64_110 ();
 sg13g2_fill_2 FILLER_64_134 ();
 sg13g2_fill_1 FILLER_64_136 ();
 sg13g2_decap_8 FILLER_64_146 ();
 sg13g2_decap_4 FILLER_64_153 ();
 sg13g2_fill_2 FILLER_64_157 ();
 sg13g2_fill_1 FILLER_64_259 ();
 sg13g2_fill_2 FILLER_64_283 ();
 sg13g2_decap_8 FILLER_64_330 ();
 sg13g2_decap_8 FILLER_64_337 ();
 sg13g2_decap_8 FILLER_64_344 ();
 sg13g2_decap_8 FILLER_64_351 ();
 sg13g2_decap_8 FILLER_64_358 ();
 sg13g2_decap_8 FILLER_64_365 ();
 sg13g2_decap_8 FILLER_64_372 ();
 sg13g2_decap_8 FILLER_64_379 ();
 sg13g2_decap_8 FILLER_64_386 ();
 sg13g2_decap_8 FILLER_64_393 ();
 sg13g2_decap_8 FILLER_64_400 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_fill_2 FILLER_65_28 ();
 sg13g2_fill_1 FILLER_65_30 ();
 sg13g2_fill_2 FILLER_65_61 ();
 sg13g2_fill_1 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_69 ();
 sg13g2_decap_4 FILLER_65_76 ();
 sg13g2_fill_1 FILLER_65_92 ();
 sg13g2_decap_4 FILLER_65_101 ();
 sg13g2_fill_2 FILLER_65_105 ();
 sg13g2_decap_4 FILLER_65_125 ();
 sg13g2_fill_2 FILLER_65_135 ();
 sg13g2_fill_1 FILLER_65_137 ();
 sg13g2_fill_2 FILLER_65_149 ();
 sg13g2_fill_1 FILLER_65_151 ();
 sg13g2_fill_2 FILLER_65_179 ();
 sg13g2_decap_4 FILLER_65_224 ();
 sg13g2_fill_2 FILLER_65_237 ();
 sg13g2_fill_1 FILLER_65_253 ();
 sg13g2_fill_2 FILLER_65_304 ();
 sg13g2_decap_8 FILLER_65_310 ();
 sg13g2_decap_8 FILLER_65_317 ();
 sg13g2_decap_8 FILLER_65_324 ();
 sg13g2_decap_8 FILLER_65_331 ();
 sg13g2_decap_8 FILLER_65_338 ();
 sg13g2_decap_8 FILLER_65_345 ();
 sg13g2_decap_8 FILLER_65_352 ();
 sg13g2_decap_8 FILLER_65_359 ();
 sg13g2_decap_8 FILLER_65_366 ();
 sg13g2_decap_8 FILLER_65_373 ();
 sg13g2_decap_8 FILLER_65_380 ();
 sg13g2_decap_8 FILLER_65_387 ();
 sg13g2_decap_8 FILLER_65_394 ();
 sg13g2_decap_8 FILLER_65_401 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_fill_1 FILLER_66_35 ();
 sg13g2_fill_1 FILLER_66_66 ();
 sg13g2_fill_2 FILLER_66_95 ();
 sg13g2_fill_2 FILLER_66_102 ();
 sg13g2_fill_1 FILLER_66_104 ();
 sg13g2_fill_2 FILLER_66_128 ();
 sg13g2_fill_1 FILLER_66_130 ();
 sg13g2_fill_1 FILLER_66_139 ();
 sg13g2_decap_8 FILLER_66_171 ();
 sg13g2_fill_2 FILLER_66_195 ();
 sg13g2_fill_1 FILLER_66_197 ();
 sg13g2_fill_1 FILLER_66_207 ();
 sg13g2_decap_8 FILLER_66_214 ();
 sg13g2_decap_8 FILLER_66_221 ();
 sg13g2_decap_8 FILLER_66_228 ();
 sg13g2_fill_2 FILLER_66_235 ();
 sg13g2_fill_1 FILLER_66_245 ();
 sg13g2_fill_2 FILLER_66_251 ();
 sg13g2_decap_4 FILLER_66_257 ();
 sg13g2_fill_2 FILLER_66_261 ();
 sg13g2_fill_2 FILLER_66_268 ();
 sg13g2_fill_1 FILLER_66_270 ();
 sg13g2_decap_4 FILLER_66_280 ();
 sg13g2_fill_2 FILLER_66_284 ();
 sg13g2_decap_8 FILLER_66_303 ();
 sg13g2_decap_8 FILLER_66_310 ();
 sg13g2_decap_8 FILLER_66_317 ();
 sg13g2_decap_8 FILLER_66_324 ();
 sg13g2_decap_8 FILLER_66_331 ();
 sg13g2_decap_8 FILLER_66_338 ();
 sg13g2_decap_8 FILLER_66_345 ();
 sg13g2_decap_8 FILLER_66_352 ();
 sg13g2_decap_8 FILLER_66_359 ();
 sg13g2_decap_8 FILLER_66_366 ();
 sg13g2_decap_8 FILLER_66_373 ();
 sg13g2_decap_8 FILLER_66_380 ();
 sg13g2_decap_8 FILLER_66_387 ();
 sg13g2_decap_8 FILLER_66_394 ();
 sg13g2_decap_8 FILLER_66_401 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_fill_2 FILLER_67_28 ();
 sg13g2_fill_1 FILLER_67_79 ();
 sg13g2_fill_2 FILLER_67_86 ();
 sg13g2_fill_2 FILLER_67_98 ();
 sg13g2_fill_2 FILLER_67_105 ();
 sg13g2_fill_1 FILLER_67_107 ();
 sg13g2_fill_1 FILLER_67_113 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_fill_2 FILLER_67_147 ();
 sg13g2_fill_1 FILLER_67_157 ();
 sg13g2_decap_8 FILLER_67_167 ();
 sg13g2_fill_2 FILLER_67_174 ();
 sg13g2_decap_8 FILLER_67_202 ();
 sg13g2_decap_4 FILLER_67_209 ();
 sg13g2_fill_2 FILLER_67_213 ();
 sg13g2_decap_4 FILLER_67_280 ();
 sg13g2_decap_8 FILLER_67_323 ();
 sg13g2_decap_8 FILLER_67_330 ();
 sg13g2_decap_8 FILLER_67_337 ();
 sg13g2_decap_8 FILLER_67_344 ();
 sg13g2_decap_8 FILLER_67_351 ();
 sg13g2_decap_8 FILLER_67_358 ();
 sg13g2_decap_8 FILLER_67_365 ();
 sg13g2_decap_8 FILLER_67_372 ();
 sg13g2_decap_8 FILLER_67_379 ();
 sg13g2_decap_8 FILLER_67_386 ();
 sg13g2_decap_8 FILLER_67_393 ();
 sg13g2_decap_8 FILLER_67_400 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_4 FILLER_68_42 ();
 sg13g2_fill_1 FILLER_68_46 ();
 sg13g2_fill_2 FILLER_68_82 ();
 sg13g2_fill_2 FILLER_68_133 ();
 sg13g2_fill_1 FILLER_68_135 ();
 sg13g2_decap_4 FILLER_68_140 ();
 sg13g2_fill_1 FILLER_68_144 ();
 sg13g2_decap_4 FILLER_68_149 ();
 sg13g2_decap_4 FILLER_68_178 ();
 sg13g2_fill_2 FILLER_68_182 ();
 sg13g2_fill_2 FILLER_68_192 ();
 sg13g2_fill_1 FILLER_68_208 ();
 sg13g2_fill_1 FILLER_68_249 ();
 sg13g2_decap_8 FILLER_68_333 ();
 sg13g2_decap_8 FILLER_68_340 ();
 sg13g2_decap_8 FILLER_68_347 ();
 sg13g2_decap_8 FILLER_68_354 ();
 sg13g2_decap_8 FILLER_68_361 ();
 sg13g2_decap_8 FILLER_68_368 ();
 sg13g2_decap_8 FILLER_68_375 ();
 sg13g2_decap_8 FILLER_68_382 ();
 sg13g2_decap_8 FILLER_68_389 ();
 sg13g2_decap_8 FILLER_68_396 ();
 sg13g2_decap_4 FILLER_68_403 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_4 FILLER_69_35 ();
 sg13g2_fill_2 FILLER_69_39 ();
 sg13g2_fill_2 FILLER_69_67 ();
 sg13g2_fill_1 FILLER_69_69 ();
 sg13g2_fill_1 FILLER_69_119 ();
 sg13g2_fill_2 FILLER_69_124 ();
 sg13g2_fill_1 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_180 ();
 sg13g2_fill_2 FILLER_69_213 ();
 sg13g2_fill_1 FILLER_69_255 ();
 sg13g2_fill_1 FILLER_69_265 ();
 sg13g2_decap_4 FILLER_69_270 ();
 sg13g2_fill_1 FILLER_69_274 ();
 sg13g2_fill_1 FILLER_69_284 ();
 sg13g2_decap_8 FILLER_69_337 ();
 sg13g2_decap_8 FILLER_69_344 ();
 sg13g2_decap_8 FILLER_69_351 ();
 sg13g2_decap_8 FILLER_69_358 ();
 sg13g2_decap_8 FILLER_69_365 ();
 sg13g2_decap_8 FILLER_69_372 ();
 sg13g2_decap_8 FILLER_69_379 ();
 sg13g2_decap_8 FILLER_69_386 ();
 sg13g2_decap_8 FILLER_69_393 ();
 sg13g2_decap_8 FILLER_69_400 ();
 sg13g2_fill_2 FILLER_69_407 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_fill_2 FILLER_70_35 ();
 sg13g2_fill_1 FILLER_70_37 ();
 sg13g2_fill_2 FILLER_70_103 ();
 sg13g2_fill_2 FILLER_70_175 ();
 sg13g2_fill_1 FILLER_70_189 ();
 sg13g2_fill_1 FILLER_70_203 ();
 sg13g2_fill_1 FILLER_70_223 ();
 sg13g2_fill_1 FILLER_70_259 ();
 sg13g2_decap_8 FILLER_70_269 ();
 sg13g2_fill_1 FILLER_70_276 ();
 sg13g2_decap_4 FILLER_70_285 ();
 sg13g2_fill_2 FILLER_70_289 ();
 sg13g2_fill_1 FILLER_70_304 ();
 sg13g2_fill_2 FILLER_70_323 ();
 sg13g2_decap_8 FILLER_70_339 ();
 sg13g2_decap_8 FILLER_70_346 ();
 sg13g2_decap_8 FILLER_70_353 ();
 sg13g2_decap_8 FILLER_70_360 ();
 sg13g2_decap_8 FILLER_70_367 ();
 sg13g2_decap_8 FILLER_70_374 ();
 sg13g2_decap_8 FILLER_70_381 ();
 sg13g2_decap_8 FILLER_70_388 ();
 sg13g2_decap_8 FILLER_70_395 ();
 sg13g2_decap_8 FILLER_70_402 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_fill_2 FILLER_71_42 ();
 sg13g2_fill_1 FILLER_71_44 ();
 sg13g2_decap_8 FILLER_71_71 ();
 sg13g2_decap_4 FILLER_71_78 ();
 sg13g2_decap_8 FILLER_71_86 ();
 sg13g2_fill_1 FILLER_71_93 ();
 sg13g2_fill_2 FILLER_71_98 ();
 sg13g2_decap_4 FILLER_71_114 ();
 sg13g2_fill_1 FILLER_71_123 ();
 sg13g2_fill_2 FILLER_71_159 ();
 sg13g2_fill_1 FILLER_71_218 ();
 sg13g2_fill_1 FILLER_71_229 ();
 sg13g2_fill_2 FILLER_71_243 ();
 sg13g2_fill_1 FILLER_71_249 ();
 sg13g2_fill_1 FILLER_71_289 ();
 sg13g2_fill_2 FILLER_71_303 ();
 sg13g2_decap_8 FILLER_71_333 ();
 sg13g2_decap_8 FILLER_71_340 ();
 sg13g2_decap_8 FILLER_71_347 ();
 sg13g2_decap_8 FILLER_71_354 ();
 sg13g2_decap_8 FILLER_71_361 ();
 sg13g2_decap_8 FILLER_71_368 ();
 sg13g2_decap_8 FILLER_71_375 ();
 sg13g2_decap_8 FILLER_71_382 ();
 sg13g2_decap_8 FILLER_71_389 ();
 sg13g2_decap_8 FILLER_71_396 ();
 sg13g2_decap_4 FILLER_71_403 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_4 FILLER_72_56 ();
 sg13g2_fill_2 FILLER_72_72 ();
 sg13g2_fill_2 FILLER_72_100 ();
 sg13g2_fill_2 FILLER_72_107 ();
 sg13g2_decap_8 FILLER_72_114 ();
 sg13g2_decap_8 FILLER_72_121 ();
 sg13g2_fill_2 FILLER_72_132 ();
 sg13g2_fill_2 FILLER_72_142 ();
 sg13g2_fill_2 FILLER_72_167 ();
 sg13g2_decap_4 FILLER_72_201 ();
 sg13g2_fill_2 FILLER_72_222 ();
 sg13g2_fill_1 FILLER_72_250 ();
 sg13g2_fill_2 FILLER_72_286 ();
 sg13g2_fill_1 FILLER_72_288 ();
 sg13g2_decap_8 FILLER_72_328 ();
 sg13g2_decap_8 FILLER_72_335 ();
 sg13g2_decap_8 FILLER_72_342 ();
 sg13g2_decap_8 FILLER_72_349 ();
 sg13g2_decap_8 FILLER_72_356 ();
 sg13g2_decap_8 FILLER_72_363 ();
 sg13g2_decap_8 FILLER_72_370 ();
 sg13g2_decap_8 FILLER_72_377 ();
 sg13g2_decap_8 FILLER_72_384 ();
 sg13g2_decap_8 FILLER_72_391 ();
 sg13g2_decap_8 FILLER_72_398 ();
 sg13g2_decap_4 FILLER_72_405 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_fill_2 FILLER_73_49 ();
 sg13g2_fill_1 FILLER_73_51 ();
 sg13g2_fill_2 FILLER_73_149 ();
 sg13g2_fill_1 FILLER_73_151 ();
 sg13g2_decap_8 FILLER_73_196 ();
 sg13g2_fill_2 FILLER_73_203 ();
 sg13g2_fill_1 FILLER_73_205 ();
 sg13g2_fill_1 FILLER_73_211 ();
 sg13g2_decap_8 FILLER_73_320 ();
 sg13g2_decap_8 FILLER_73_327 ();
 sg13g2_decap_8 FILLER_73_334 ();
 sg13g2_decap_8 FILLER_73_341 ();
 sg13g2_decap_8 FILLER_73_348 ();
 sg13g2_decap_8 FILLER_73_355 ();
 sg13g2_decap_8 FILLER_73_362 ();
 sg13g2_decap_8 FILLER_73_369 ();
 sg13g2_decap_8 FILLER_73_376 ();
 sg13g2_decap_8 FILLER_73_383 ();
 sg13g2_decap_8 FILLER_73_390 ();
 sg13g2_decap_8 FILLER_73_397 ();
 sg13g2_decap_4 FILLER_73_404 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_4 FILLER_74_35 ();
 sg13g2_fill_1 FILLER_74_39 ();
 sg13g2_fill_1 FILLER_74_66 ();
 sg13g2_fill_2 FILLER_74_106 ();
 sg13g2_fill_1 FILLER_74_108 ();
 sg13g2_fill_2 FILLER_74_140 ();
 sg13g2_decap_4 FILLER_74_191 ();
 sg13g2_fill_2 FILLER_74_235 ();
 sg13g2_fill_1 FILLER_74_237 ();
 sg13g2_fill_1 FILLER_74_269 ();
 sg13g2_decap_8 FILLER_74_279 ();
 sg13g2_fill_1 FILLER_74_286 ();
 sg13g2_fill_2 FILLER_74_294 ();
 sg13g2_decap_8 FILLER_74_319 ();
 sg13g2_decap_8 FILLER_74_326 ();
 sg13g2_decap_8 FILLER_74_333 ();
 sg13g2_decap_8 FILLER_74_340 ();
 sg13g2_decap_8 FILLER_74_347 ();
 sg13g2_decap_8 FILLER_74_354 ();
 sg13g2_decap_8 FILLER_74_361 ();
 sg13g2_decap_8 FILLER_74_368 ();
 sg13g2_decap_8 FILLER_74_375 ();
 sg13g2_decap_8 FILLER_74_382 ();
 sg13g2_decap_8 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_74_396 ();
 sg13g2_decap_4 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_4 FILLER_75_35 ();
 sg13g2_fill_1 FILLER_75_39 ();
 sg13g2_fill_1 FILLER_75_66 ();
 sg13g2_fill_2 FILLER_75_93 ();
 sg13g2_fill_2 FILLER_75_120 ();
 sg13g2_fill_1 FILLER_75_122 ();
 sg13g2_decap_8 FILLER_75_162 ();
 sg13g2_fill_1 FILLER_75_177 ();
 sg13g2_fill_1 FILLER_75_186 ();
 sg13g2_fill_1 FILLER_75_238 ();
 sg13g2_fill_1 FILLER_75_261 ();
 sg13g2_fill_2 FILLER_75_275 ();
 sg13g2_fill_1 FILLER_75_294 ();
 sg13g2_decap_8 FILLER_75_313 ();
 sg13g2_decap_8 FILLER_75_320 ();
 sg13g2_decap_8 FILLER_75_327 ();
 sg13g2_decap_8 FILLER_75_334 ();
 sg13g2_decap_8 FILLER_75_341 ();
 sg13g2_decap_8 FILLER_75_348 ();
 sg13g2_decap_8 FILLER_75_355 ();
 sg13g2_decap_8 FILLER_75_362 ();
 sg13g2_decap_8 FILLER_75_369 ();
 sg13g2_decap_8 FILLER_75_376 ();
 sg13g2_decap_8 FILLER_75_383 ();
 sg13g2_decap_8 FILLER_75_390 ();
 sg13g2_decap_8 FILLER_75_397 ();
 sg13g2_decap_4 FILLER_75_404 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_4 FILLER_76_42 ();
 sg13g2_fill_1 FILLER_76_58 ();
 sg13g2_fill_1 FILLER_76_82 ();
 sg13g2_decap_4 FILLER_76_96 ();
 sg13g2_fill_1 FILLER_76_100 ();
 sg13g2_fill_2 FILLER_76_123 ();
 sg13g2_fill_1 FILLER_76_125 ();
 sg13g2_fill_2 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_153 ();
 sg13g2_fill_2 FILLER_76_160 ();
 sg13g2_fill_1 FILLER_76_162 ();
 sg13g2_decap_8 FILLER_76_188 ();
 sg13g2_fill_2 FILLER_76_195 ();
 sg13g2_fill_1 FILLER_76_197 ();
 sg13g2_fill_2 FILLER_76_206 ();
 sg13g2_decap_8 FILLER_76_221 ();
 sg13g2_decap_8 FILLER_76_246 ();
 sg13g2_fill_1 FILLER_76_253 ();
 sg13g2_decap_4 FILLER_76_270 ();
 sg13g2_decap_8 FILLER_76_317 ();
 sg13g2_decap_8 FILLER_76_324 ();
 sg13g2_decap_8 FILLER_76_331 ();
 sg13g2_decap_8 FILLER_76_338 ();
 sg13g2_decap_8 FILLER_76_345 ();
 sg13g2_decap_8 FILLER_76_352 ();
 sg13g2_decap_8 FILLER_76_359 ();
 sg13g2_decap_8 FILLER_76_366 ();
 sg13g2_decap_8 FILLER_76_373 ();
 sg13g2_decap_8 FILLER_76_380 ();
 sg13g2_decap_8 FILLER_76_387 ();
 sg13g2_decap_8 FILLER_76_394 ();
 sg13g2_decap_8 FILLER_76_401 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_fill_2 FILLER_77_49 ();
 sg13g2_decap_4 FILLER_77_55 ();
 sg13g2_fill_1 FILLER_77_77 ();
 sg13g2_fill_2 FILLER_77_109 ();
 sg13g2_fill_1 FILLER_77_111 ();
 sg13g2_fill_2 FILLER_77_116 ();
 sg13g2_fill_1 FILLER_77_118 ();
 sg13g2_fill_2 FILLER_77_136 ();
 sg13g2_fill_1 FILLER_77_138 ();
 sg13g2_fill_1 FILLER_77_204 ();
 sg13g2_decap_4 FILLER_77_214 ();
 sg13g2_fill_2 FILLER_77_231 ();
 sg13g2_fill_2 FILLER_77_288 ();
 sg13g2_decap_8 FILLER_77_325 ();
 sg13g2_decap_8 FILLER_77_332 ();
 sg13g2_decap_8 FILLER_77_339 ();
 sg13g2_decap_8 FILLER_77_346 ();
 sg13g2_decap_8 FILLER_77_353 ();
 sg13g2_decap_8 FILLER_77_360 ();
 sg13g2_decap_8 FILLER_77_367 ();
 sg13g2_decap_8 FILLER_77_374 ();
 sg13g2_decap_8 FILLER_77_381 ();
 sg13g2_decap_8 FILLER_77_388 ();
 sg13g2_decap_8 FILLER_77_395 ();
 sg13g2_decap_8 FILLER_77_402 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_fill_2 FILLER_78_56 ();
 sg13g2_fill_1 FILLER_78_58 ();
 sg13g2_fill_1 FILLER_78_163 ();
 sg13g2_fill_2 FILLER_78_173 ();
 sg13g2_fill_1 FILLER_78_175 ();
 sg13g2_fill_1 FILLER_78_185 ();
 sg13g2_decap_8 FILLER_78_327 ();
 sg13g2_decap_8 FILLER_78_334 ();
 sg13g2_decap_8 FILLER_78_341 ();
 sg13g2_decap_8 FILLER_78_348 ();
 sg13g2_decap_8 FILLER_78_355 ();
 sg13g2_decap_8 FILLER_78_362 ();
 sg13g2_decap_8 FILLER_78_369 ();
 sg13g2_decap_8 FILLER_78_376 ();
 sg13g2_decap_8 FILLER_78_383 ();
 sg13g2_decap_8 FILLER_78_390 ();
 sg13g2_decap_8 FILLER_78_397 ();
 sg13g2_decap_4 FILLER_78_404 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_4 FILLER_79_49 ();
 sg13g2_fill_1 FILLER_79_87 ();
 sg13g2_fill_2 FILLER_79_243 ();
 sg13g2_fill_1 FILLER_79_245 ();
 sg13g2_fill_2 FILLER_79_280 ();
 sg13g2_decap_8 FILLER_79_321 ();
 sg13g2_decap_8 FILLER_79_328 ();
 sg13g2_decap_8 FILLER_79_335 ();
 sg13g2_decap_8 FILLER_79_342 ();
 sg13g2_decap_8 FILLER_79_349 ();
 sg13g2_decap_8 FILLER_79_356 ();
 sg13g2_decap_8 FILLER_79_363 ();
 sg13g2_decap_8 FILLER_79_370 ();
 sg13g2_decap_8 FILLER_79_377 ();
 sg13g2_decap_8 FILLER_79_384 ();
 sg13g2_decap_8 FILLER_79_391 ();
 sg13g2_decap_8 FILLER_79_398 ();
 sg13g2_decap_4 FILLER_79_405 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_fill_2 FILLER_80_42 ();
 sg13g2_fill_1 FILLER_80_44 ();
 sg13g2_fill_2 FILLER_80_96 ();
 sg13g2_fill_1 FILLER_80_98 ();
 sg13g2_fill_2 FILLER_80_120 ();
 sg13g2_fill_1 FILLER_80_131 ();
 sg13g2_decap_8 FILLER_80_148 ();
 sg13g2_fill_2 FILLER_80_168 ();
 sg13g2_fill_1 FILLER_80_170 ();
 sg13g2_fill_2 FILLER_80_184 ();
 sg13g2_fill_1 FILLER_80_186 ();
 sg13g2_decap_4 FILLER_80_279 ();
 sg13g2_fill_1 FILLER_80_283 ();
 sg13g2_fill_2 FILLER_80_287 ();
 sg13g2_fill_1 FILLER_80_289 ();
 sg13g2_decap_8 FILLER_80_312 ();
 sg13g2_decap_8 FILLER_80_319 ();
 sg13g2_decap_8 FILLER_80_326 ();
 sg13g2_decap_8 FILLER_80_333 ();
 sg13g2_decap_8 FILLER_80_340 ();
 sg13g2_decap_8 FILLER_80_347 ();
 sg13g2_decap_8 FILLER_80_354 ();
 sg13g2_decap_8 FILLER_80_361 ();
 sg13g2_decap_8 FILLER_80_368 ();
 sg13g2_fill_1 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net314;
 assign uio_oe[1] = net315;
 assign uio_oe[2] = net316;
 assign uio_oe[3] = net317;
 assign uio_oe[4] = net318;
 assign uio_oe[5] = net319;
 assign uio_oe[6] = net320;
 assign uio_oe[7] = net321;
 assign uo_out[2] = net2;
 assign uo_out[3] = net3;
 assign uo_out[4] = net4;
 assign uo_out[5] = net5;
 assign uo_out[6] = net6;
 assign uo_out[7] = net7;
endmodule

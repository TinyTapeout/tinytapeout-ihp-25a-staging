module tt_um_gcd_stephan (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \C[0] ;
 wire \C[1] ;
 wire \C[2] ;
 wire \C[3] ;
 wire \C[4] ;
 wire \C[5] ;
 wire \C[6] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire ack_w;
 wire \gcd_module_inst.datapath_comp.RegA_int[0] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[10] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[11] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[12] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[13] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[14] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[15] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[1] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[2] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[3] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[4] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[5] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[6] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[7] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[8] ;
 wire \gcd_module_inst.datapath_comp.RegA_int[9] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[0] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[10] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[11] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[12] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[13] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[14] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[15] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[1] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[2] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[3] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[4] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[5] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[6] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[7] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[8] ;
 wire \gcd_module_inst.datapath_comp.RegB_int[9] ;
 wire \gcd_module_inst.fsm_comp.next_state[0] ;
 wire \gcd_module_inst.fsm_comp.next_state[1] ;
 wire \gcd_module_inst.fsm_comp.next_state[2] ;
 wire \gcd_module_inst.fsm_comp.state[0] ;
 wire \gcd_module_inst.fsm_comp.state[1] ;
 wire \gcd_module_inst.fsm_comp.state[2] ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire clknet_0_clk;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;

 sg13g2_inv_1 _365_ (.Y(_330_),
    .A(net111));
 sg13g2_inv_1 _366_ (.Y(_331_),
    .A(_000_));
 sg13g2_inv_2 _367_ (.Y(_034_),
    .A(net112));
 sg13g2_inv_1 _368_ (.Y(_035_),
    .A(net1));
 sg13g2_inv_1 _369_ (.Y(_036_),
    .A(net52));
 sg13g2_nand2b_2 _370_ (.Y(_037_),
    .B(net111),
    .A_N(\gcd_module_inst.fsm_comp.state[2] ));
 sg13g2_nor2b_2 _371_ (.A(net111),
    .B_N(\gcd_module_inst.fsm_comp.state[2] ),
    .Y(_038_));
 sg13g2_and2_2 _372_ (.A(\gcd_module_inst.fsm_comp.state[1] ),
    .B(_038_),
    .X(_039_));
 sg13g2_and2_2 _373_ (.A(net111),
    .B(net110),
    .X(_040_));
 sg13g2_and2_1 _374_ (.A(_331_),
    .B(_040_),
    .X(_041_));
 sg13g2_or2_1 _375_ (.X(_042_),
    .B(_041_),
    .A(_039_));
 sg13g2_or2_1 _376_ (.X(_043_),
    .B(_000_),
    .A(net111));
 sg13g2_nor2_1 _377_ (.A(\gcd_module_inst.fsm_comp.state[0] ),
    .B(net110),
    .Y(_044_));
 sg13g2_nor3_2 _378_ (.A(net65),
    .B(net110),
    .C(_000_),
    .Y(_045_));
 sg13g2_a221oi_1 _379_ (.B2(_331_),
    .C1(_045_),
    .B1(_040_),
    .A1(\gcd_module_inst.fsm_comp.state[1] ),
    .Y(_046_),
    .A2(_038_));
 sg13g2_nand2b_1 _380_ (.Y(_047_),
    .B(net111),
    .A_N(_001_));
 sg13g2_nand2_1 _381_ (.Y(_048_),
    .A(_043_),
    .B(_047_));
 sg13g2_nor2b_2 _382_ (.A(_046_),
    .B_N(_048_),
    .Y(_049_));
 sg13g2_nor2b_1 _383_ (.A(\gcd_module_inst.datapath_comp.RegB_int[0] ),
    .B_N(\gcd_module_inst.datapath_comp.RegA_int[0] ),
    .Y(_050_));
 sg13g2_nand2b_1 _384_ (.Y(_051_),
    .B(\gcd_module_inst.datapath_comp.RegA_int[0] ),
    .A_N(\gcd_module_inst.datapath_comp.RegB_int[0] ));
 sg13g2_nor2b_1 _385_ (.A(\gcd_module_inst.datapath_comp.RegA_int[0] ),
    .B_N(\gcd_module_inst.datapath_comp.RegB_int[0] ),
    .Y(_052_));
 sg13g2_o21ai_1 _386_ (.B1(_049_),
    .Y(_053_),
    .A1(_050_),
    .A2(_052_));
 sg13g2_a221oi_1 _387_ (.B2(_047_),
    .C1(_046_),
    .B1(_043_),
    .A1(\gcd_module_inst.fsm_comp.state[1] ),
    .Y(_054_),
    .A2(_038_));
 sg13g2_nand2b_2 _388_ (.Y(_055_),
    .B(_049_),
    .A_N(_039_));
 sg13g2_mux2_1 _389_ (.A0(_039_),
    .A1(_046_),
    .S(_048_),
    .X(_056_));
 sg13g2_nor2_1 _390_ (.A(_038_),
    .B(_040_),
    .Y(_057_));
 sg13g2_a22oi_1 _391_ (.Y(_058_),
    .B1(net105),
    .B2(\gcd_module_inst.datapath_comp.RegA_int[0] ),
    .A2(net97),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[0] ));
 sg13g2_o21ai_1 _392_ (.B1(_053_),
    .Y(_059_),
    .A1(net100),
    .A2(_058_));
 sg13g2_nand3_1 _393_ (.B(net106),
    .C(_059_),
    .A(net119),
    .Y(_060_));
 sg13g2_o21ai_1 _394_ (.B1(_060_),
    .Y(\C[0] ),
    .A1(_035_),
    .A2(net106));
 sg13g2_nor2_1 _395_ (.A(net2),
    .B(net106),
    .Y(_061_));
 sg13g2_nand4_1 _396_ (.B(_330_),
    .C(net110),
    .A(\gcd_module_inst.fsm_comp.state[2] ),
    .Y(_062_),
    .D(_331_));
 sg13g2_nor2b_1 _397_ (.A(\gcd_module_inst.datapath_comp.RegA_int[1] ),
    .B_N(\gcd_module_inst.datapath_comp.RegB_int[1] ),
    .Y(_063_));
 sg13g2_xnor2_1 _398_ (.Y(_064_),
    .A(\gcd_module_inst.datapath_comp.RegB_int[1] ),
    .B(\gcd_module_inst.datapath_comp.RegA_int[1] ));
 sg13g2_xnor2_1 _399_ (.Y(_065_),
    .A(_051_),
    .B(_064_));
 sg13g2_a221oi_1 _400_ (.B2(\gcd_module_inst.datapath_comp.RegA_int[1] ),
    .C1(net101),
    .B1(net105),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[1] ),
    .Y(_066_),
    .A2(net97));
 sg13g2_o21ai_1 _401_ (.B1(_066_),
    .Y(_067_),
    .A1(net103),
    .A2(_065_));
 sg13g2_nand2b_1 _402_ (.Y(_068_),
    .B(_064_),
    .A_N(_052_));
 sg13g2_xnor2_1 _403_ (.Y(_069_),
    .A(_052_),
    .B(_064_));
 sg13g2_o21ai_1 _404_ (.B1(net118),
    .Y(_070_),
    .A1(_055_),
    .A2(_069_));
 sg13g2_nand2b_1 _405_ (.Y(_071_),
    .B(_067_),
    .A_N(_070_));
 sg13g2_a21oi_1 _406_ (.A1(_037_),
    .A2(_071_),
    .Y(\C[1] ),
    .B1(_061_));
 sg13g2_nor2_1 _407_ (.A(net3),
    .B(net106),
    .Y(_072_));
 sg13g2_nand2b_1 _408_ (.Y(_073_),
    .B(\gcd_module_inst.datapath_comp.RegA_int[2] ),
    .A_N(\gcd_module_inst.datapath_comp.RegB_int[2] ));
 sg13g2_nand2b_1 _409_ (.Y(_074_),
    .B(\gcd_module_inst.datapath_comp.RegB_int[2] ),
    .A_N(\gcd_module_inst.datapath_comp.RegA_int[2] ));
 sg13g2_xor2_1 _410_ (.B(\gcd_module_inst.datapath_comp.RegA_int[2] ),
    .A(\gcd_module_inst.datapath_comp.RegB_int[2] ),
    .X(_075_));
 sg13g2_a21o_2 _411_ (.A2(_064_),
    .A1(_051_),
    .B1(_063_),
    .X(_076_));
 sg13g2_nand2b_1 _412_ (.Y(_077_),
    .B(_076_),
    .A_N(_075_));
 sg13g2_xor2_1 _413_ (.B(_076_),
    .A(_075_),
    .X(_078_));
 sg13g2_a221oi_1 _414_ (.B2(\gcd_module_inst.datapath_comp.RegA_int[2] ),
    .C1(net100),
    .B1(net105),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[2] ),
    .Y(_079_),
    .A2(net97));
 sg13g2_o21ai_1 _415_ (.B1(_079_),
    .Y(_080_),
    .A1(net103),
    .A2(_078_));
 sg13g2_and2_1 _416_ (.A(_068_),
    .B(_076_),
    .X(_081_));
 sg13g2_xnor2_1 _417_ (.Y(_082_),
    .A(_075_),
    .B(_081_));
 sg13g2_a21oi_1 _418_ (.A1(net100),
    .A2(_082_),
    .Y(_083_),
    .B1(_034_));
 sg13g2_nand2_1 _419_ (.Y(_084_),
    .A(_080_),
    .B(_083_));
 sg13g2_a21oi_1 _420_ (.A1(net106),
    .A2(_084_),
    .Y(\C[2] ),
    .B1(_072_));
 sg13g2_nor2_1 _421_ (.A(net4),
    .B(net106),
    .Y(_085_));
 sg13g2_nand2b_1 _422_ (.Y(_086_),
    .B(\gcd_module_inst.datapath_comp.RegB_int[3] ),
    .A_N(\gcd_module_inst.datapath_comp.RegA_int[3] ));
 sg13g2_xor2_1 _423_ (.B(\gcd_module_inst.datapath_comp.RegA_int[3] ),
    .A(\gcd_module_inst.datapath_comp.RegB_int[3] ),
    .X(_087_));
 sg13g2_o21ai_1 _424_ (.B1(_073_),
    .Y(_088_),
    .A1(_075_),
    .A2(_081_));
 sg13g2_a21oi_1 _425_ (.A1(_087_),
    .A2(_088_),
    .Y(_089_),
    .B1(_055_));
 sg13g2_o21ai_1 _426_ (.B1(_089_),
    .Y(_090_),
    .A1(_087_),
    .A2(_088_));
 sg13g2_nand3_1 _427_ (.B(_077_),
    .C(_087_),
    .A(_074_),
    .Y(_091_));
 sg13g2_nor2_1 _428_ (.A(_075_),
    .B(_087_),
    .Y(_092_));
 sg13g2_or2_1 _429_ (.X(_093_),
    .B(_087_),
    .A(_075_));
 sg13g2_a21o_1 _430_ (.A2(_077_),
    .A1(_074_),
    .B1(_087_),
    .X(_094_));
 sg13g2_nand4_1 _431_ (.B(_049_),
    .C(_091_),
    .A(_039_),
    .Y(_095_),
    .D(_094_));
 sg13g2_a221oi_1 _432_ (.B2(\gcd_module_inst.datapath_comp.RegA_int[3] ),
    .C1(net101),
    .B1(net105),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[3] ),
    .Y(_096_),
    .A2(net97));
 sg13g2_a21oi_1 _433_ (.A1(_095_),
    .A2(_096_),
    .Y(_097_),
    .B1(_034_));
 sg13g2_nand2_1 _434_ (.Y(_098_),
    .A(_090_),
    .B(_097_));
 sg13g2_a21oi_1 _435_ (.A1(net107),
    .A2(_098_),
    .Y(\C[3] ),
    .B1(_085_));
 sg13g2_nor2_1 _436_ (.A(net5),
    .B(net106),
    .Y(_099_));
 sg13g2_nand2b_1 _437_ (.Y(_100_),
    .B(\gcd_module_inst.datapath_comp.RegB_int[4] ),
    .A_N(\gcd_module_inst.datapath_comp.RegA_int[4] ));
 sg13g2_nor2b_2 _438_ (.A(\gcd_module_inst.datapath_comp.RegB_int[4] ),
    .B_N(\gcd_module_inst.datapath_comp.RegA_int[4] ),
    .Y(_101_));
 sg13g2_xor2_1 _439_ (.B(\gcd_module_inst.datapath_comp.RegA_int[4] ),
    .A(\gcd_module_inst.datapath_comp.RegB_int[4] ),
    .X(_102_));
 sg13g2_o21ai_1 _440_ (.B1(_086_),
    .Y(_103_),
    .A1(_074_),
    .A2(_087_));
 sg13g2_a21oi_2 _441_ (.B1(_103_),
    .Y(_104_),
    .A2(_092_),
    .A1(_076_));
 sg13g2_a21o_1 _442_ (.A2(_092_),
    .A1(_076_),
    .B1(_103_),
    .X(_105_));
 sg13g2_nor2_1 _443_ (.A(_081_),
    .B(_093_),
    .Y(_106_));
 sg13g2_a21o_1 _444_ (.A2(_076_),
    .A1(_068_),
    .B1(_093_),
    .X(_107_));
 sg13g2_a21oi_1 _445_ (.A1(_105_),
    .A2(_107_),
    .Y(_108_),
    .B1(_102_));
 sg13g2_and3_1 _446_ (.X(_109_),
    .A(_102_),
    .B(_105_),
    .C(_107_));
 sg13g2_o21ai_1 _447_ (.B1(net99),
    .Y(_110_),
    .A1(_108_),
    .A2(_109_));
 sg13g2_nor2_1 _448_ (.A(_102_),
    .B(_104_),
    .Y(_111_));
 sg13g2_a21o_1 _449_ (.A2(_104_),
    .A1(_102_),
    .B1(net102),
    .X(_112_));
 sg13g2_a221oi_1 _450_ (.B2(\gcd_module_inst.datapath_comp.RegA_int[4] ),
    .C1(net99),
    .B1(net104),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[4] ),
    .Y(_113_),
    .A2(net96));
 sg13g2_o21ai_1 _451_ (.B1(_113_),
    .Y(_114_),
    .A1(_111_),
    .A2(_112_));
 sg13g2_nand3_1 _452_ (.B(_110_),
    .C(_114_),
    .A(net119),
    .Y(_115_));
 sg13g2_a21oi_1 _453_ (.A1(net107),
    .A2(_115_),
    .Y(\C[4] ),
    .B1(_099_));
 sg13g2_nand2b_1 _454_ (.Y(_116_),
    .B(\gcd_module_inst.datapath_comp.RegB_int[5] ),
    .A_N(\gcd_module_inst.datapath_comp.RegA_int[5] ));
 sg13g2_nor2b_1 _455_ (.A(\gcd_module_inst.datapath_comp.RegB_int[5] ),
    .B_N(\gcd_module_inst.datapath_comp.RegA_int[5] ),
    .Y(_117_));
 sg13g2_xor2_1 _456_ (.B(\gcd_module_inst.datapath_comp.RegA_int[5] ),
    .A(\gcd_module_inst.datapath_comp.RegB_int[5] ),
    .X(_118_));
 sg13g2_o21ai_1 _457_ (.B1(_100_),
    .Y(_119_),
    .A1(_101_),
    .A2(_104_));
 sg13g2_xor2_1 _458_ (.B(_119_),
    .A(_118_),
    .X(_120_));
 sg13g2_a221oi_1 _459_ (.B2(\gcd_module_inst.datapath_comp.RegA_int[5] ),
    .C1(net99),
    .B1(net104),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[5] ),
    .Y(_121_),
    .A2(net96));
 sg13g2_o21ai_1 _460_ (.B1(_121_),
    .Y(_122_),
    .A1(net102),
    .A2(_120_));
 sg13g2_o21ai_1 _461_ (.B1(_118_),
    .Y(_123_),
    .A1(_101_),
    .A2(_108_));
 sg13g2_or3_1 _462_ (.A(_101_),
    .B(_108_),
    .C(_118_),
    .X(_124_));
 sg13g2_nand3_1 _463_ (.B(_123_),
    .C(_124_),
    .A(net99),
    .Y(_125_));
 sg13g2_nand3_1 _464_ (.B(_122_),
    .C(_125_),
    .A(net119),
    .Y(_126_));
 sg13g2_nor2_1 _465_ (.A(net6),
    .B(net107),
    .Y(_127_));
 sg13g2_a21oi_1 _466_ (.A1(net107),
    .A2(_126_),
    .Y(\C[5] ),
    .B1(_127_));
 sg13g2_nor2_1 _467_ (.A(net7),
    .B(net107),
    .Y(_128_));
 sg13g2_nor2b_1 _468_ (.A(\gcd_module_inst.datapath_comp.RegA_int[6] ),
    .B_N(\gcd_module_inst.datapath_comp.RegB_int[6] ),
    .Y(_129_));
 sg13g2_nand2b_1 _469_ (.Y(_130_),
    .B(\gcd_module_inst.datapath_comp.RegA_int[6] ),
    .A_N(\gcd_module_inst.datapath_comp.RegB_int[6] ));
 sg13g2_xor2_1 _470_ (.B(\gcd_module_inst.datapath_comp.RegA_int[6] ),
    .A(\gcd_module_inst.datapath_comp.RegB_int[6] ),
    .X(_131_));
 sg13g2_nor2_1 _471_ (.A(_102_),
    .B(_118_),
    .Y(_132_));
 sg13g2_o21ai_1 _472_ (.B1(_132_),
    .Y(_133_),
    .A1(_104_),
    .A2(_106_));
 sg13g2_o21ai_1 _473_ (.B1(_116_),
    .Y(_134_),
    .A1(_101_),
    .A2(_117_));
 sg13g2_nand3_1 _474_ (.B(_133_),
    .C(_134_),
    .A(_131_),
    .Y(_135_));
 sg13g2_a21o_1 _475_ (.A2(_134_),
    .A1(_133_),
    .B1(_131_),
    .X(_136_));
 sg13g2_a21oi_1 _476_ (.A1(_135_),
    .A2(_136_),
    .Y(_137_),
    .B1(_055_));
 sg13g2_o21ai_1 _477_ (.B1(_116_),
    .Y(_138_),
    .A1(_100_),
    .A2(_118_));
 sg13g2_a21oi_1 _478_ (.A1(_105_),
    .A2(_132_),
    .Y(_139_),
    .B1(_138_));
 sg13g2_nor2_1 _479_ (.A(_131_),
    .B(_139_),
    .Y(_140_));
 sg13g2_a21o_1 _480_ (.A2(_139_),
    .A1(_131_),
    .B1(net102),
    .X(_141_));
 sg13g2_a221oi_1 _481_ (.B2(\gcd_module_inst.datapath_comp.RegA_int[6] ),
    .C1(net99),
    .B1(net104),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[6] ),
    .Y(_142_),
    .A2(net96));
 sg13g2_o21ai_1 _482_ (.B1(_142_),
    .Y(_143_),
    .A1(_140_),
    .A2(_141_));
 sg13g2_nand3b_1 _483_ (.B(_143_),
    .C(net114),
    .Y(_144_),
    .A_N(_137_));
 sg13g2_a21oi_1 _484_ (.A1(net107),
    .A2(_144_),
    .Y(\C[6] ),
    .B1(_128_));
 sg13g2_nor2_1 _485_ (.A(_330_),
    .B(net110),
    .Y(_145_));
 sg13g2_and2_1 _486_ (.A(\gcd_module_inst.fsm_comp.state[2] ),
    .B(_145_),
    .X(_146_));
 sg13g2_o21ai_1 _487_ (.B1(_000_),
    .Y(_147_),
    .A1(net111),
    .A2(net110));
 sg13g2_nor2_1 _488_ (.A(_040_),
    .B(_147_),
    .Y(_148_));
 sg13g2_nor2_1 _489_ (.A(net110),
    .B(_038_),
    .Y(_149_));
 sg13g2_a21oi_1 _490_ (.A1(net110),
    .A2(net109),
    .Y(_150_),
    .B1(_149_));
 sg13g2_nor4_2 _491_ (.A(_042_),
    .B(_146_),
    .C(_148_),
    .Y(_151_),
    .D(_150_));
 sg13g2_nor2b_1 _492_ (.A(\gcd_module_inst.datapath_comp.RegA_int[15] ),
    .B_N(\gcd_module_inst.datapath_comp.RegB_int[15] ),
    .Y(_152_));
 sg13g2_nor2b_1 _493_ (.A(\gcd_module_inst.datapath_comp.RegB_int[15] ),
    .B_N(\gcd_module_inst.datapath_comp.RegA_int[15] ),
    .Y(_153_));
 sg13g2_nand2b_1 _494_ (.Y(_154_),
    .B(\gcd_module_inst.datapath_comp.RegB_int[14] ),
    .A_N(\gcd_module_inst.datapath_comp.RegA_int[14] ));
 sg13g2_nor2b_1 _495_ (.A(\gcd_module_inst.datapath_comp.RegB_int[14] ),
    .B_N(\gcd_module_inst.datapath_comp.RegA_int[14] ),
    .Y(_155_));
 sg13g2_xor2_1 _496_ (.B(\gcd_module_inst.datapath_comp.RegA_int[14] ),
    .A(\gcd_module_inst.datapath_comp.RegB_int[14] ),
    .X(_156_));
 sg13g2_inv_1 _497_ (.Y(_157_),
    .A(_156_));
 sg13g2_nor2b_1 _498_ (.A(\gcd_module_inst.datapath_comp.RegB_int[13] ),
    .B_N(\gcd_module_inst.datapath_comp.RegA_int[13] ),
    .Y(_158_));
 sg13g2_nand2b_1 _499_ (.Y(_159_),
    .B(\gcd_module_inst.datapath_comp.RegB_int[13] ),
    .A_N(\gcd_module_inst.datapath_comp.RegA_int[13] ));
 sg13g2_nor2b_1 _500_ (.A(_158_),
    .B_N(_159_),
    .Y(_160_));
 sg13g2_nand2b_1 _501_ (.Y(_161_),
    .B(_159_),
    .A_N(_158_));
 sg13g2_nor2b_2 _502_ (.A(\gcd_module_inst.datapath_comp.RegB_int[12] ),
    .B_N(\gcd_module_inst.datapath_comp.RegA_int[12] ),
    .Y(_162_));
 sg13g2_nand2b_1 _503_ (.Y(_163_),
    .B(\gcd_module_inst.datapath_comp.RegB_int[12] ),
    .A_N(\gcd_module_inst.datapath_comp.RegA_int[12] ));
 sg13g2_nor2b_1 _504_ (.A(_162_),
    .B_N(_163_),
    .Y(_164_));
 sg13g2_inv_1 _505_ (.Y(_165_),
    .A(_164_));
 sg13g2_nor2_1 _506_ (.A(_161_),
    .B(_165_),
    .Y(_166_));
 sg13g2_nand2b_1 _507_ (.Y(_167_),
    .B(\gcd_module_inst.datapath_comp.RegB_int[11] ),
    .A_N(\gcd_module_inst.datapath_comp.RegA_int[11] ));
 sg13g2_nor2b_1 _508_ (.A(\gcd_module_inst.datapath_comp.RegB_int[11] ),
    .B_N(\gcd_module_inst.datapath_comp.RegA_int[11] ),
    .Y(_168_));
 sg13g2_xnor2_1 _509_ (.Y(_169_),
    .A(\gcd_module_inst.datapath_comp.RegB_int[11] ),
    .B(\gcd_module_inst.datapath_comp.RegA_int[11] ));
 sg13g2_xor2_1 _510_ (.B(\gcd_module_inst.datapath_comp.RegA_int[11] ),
    .A(\gcd_module_inst.datapath_comp.RegB_int[11] ),
    .X(_170_));
 sg13g2_nand2b_1 _511_ (.Y(_171_),
    .B(\gcd_module_inst.datapath_comp.RegB_int[10] ),
    .A_N(\gcd_module_inst.datapath_comp.RegA_int[10] ));
 sg13g2_nor2b_2 _512_ (.A(\gcd_module_inst.datapath_comp.RegB_int[10] ),
    .B_N(\gcd_module_inst.datapath_comp.RegA_int[10] ),
    .Y(_172_));
 sg13g2_xor2_1 _513_ (.B(\gcd_module_inst.datapath_comp.RegA_int[10] ),
    .A(\gcd_module_inst.datapath_comp.RegB_int[10] ),
    .X(_173_));
 sg13g2_inv_1 _514_ (.Y(_174_),
    .A(_173_));
 sg13g2_nor2_1 _515_ (.A(_170_),
    .B(_173_),
    .Y(_175_));
 sg13g2_nor2b_1 _516_ (.A(\gcd_module_inst.datapath_comp.RegA_int[8] ),
    .B_N(\gcd_module_inst.datapath_comp.RegB_int[8] ),
    .Y(_176_));
 sg13g2_nand2b_1 _517_ (.Y(_177_),
    .B(\gcd_module_inst.datapath_comp.RegB_int[9] ),
    .A_N(\gcd_module_inst.datapath_comp.RegA_int[9] ));
 sg13g2_nand2b_2 _518_ (.Y(_178_),
    .B(\gcd_module_inst.datapath_comp.RegA_int[8] ),
    .A_N(\gcd_module_inst.datapath_comp.RegB_int[8] ));
 sg13g2_nand2b_1 _519_ (.Y(_179_),
    .B(\gcd_module_inst.datapath_comp.RegA_int[9] ),
    .A_N(\gcd_module_inst.datapath_comp.RegB_int[9] ));
 sg13g2_and2_1 _520_ (.A(_178_),
    .B(_179_),
    .X(_180_));
 sg13g2_nand2b_2 _521_ (.Y(_181_),
    .B(_178_),
    .A_N(_176_));
 sg13g2_nand2_1 _522_ (.Y(_182_),
    .A(_177_),
    .B(_179_));
 sg13g2_nor2_1 _523_ (.A(_181_),
    .B(_182_),
    .Y(_183_));
 sg13g2_and2_1 _524_ (.A(_175_),
    .B(_183_),
    .X(_184_));
 sg13g2_nand2_1 _525_ (.Y(_185_),
    .A(_175_),
    .B(_183_));
 sg13g2_nor2b_1 _526_ (.A(\gcd_module_inst.datapath_comp.RegA_int[7] ),
    .B_N(\gcd_module_inst.datapath_comp.RegB_int[7] ),
    .Y(_186_));
 sg13g2_nand2b_1 _527_ (.Y(_187_),
    .B(\gcd_module_inst.datapath_comp.RegA_int[7] ),
    .A_N(\gcd_module_inst.datapath_comp.RegB_int[7] ));
 sg13g2_xnor2_1 _528_ (.Y(_188_),
    .A(\gcd_module_inst.datapath_comp.RegB_int[7] ),
    .B(\gcd_module_inst.datapath_comp.RegA_int[7] ));
 sg13g2_nor2b_1 _529_ (.A(_131_),
    .B_N(_188_),
    .Y(_189_));
 sg13g2_nand2_1 _530_ (.Y(_190_),
    .A(_132_),
    .B(_189_));
 sg13g2_a221oi_1 _531_ (.B2(_138_),
    .C1(_186_),
    .B1(_189_),
    .A1(_129_),
    .Y(_191_),
    .A2(_187_));
 sg13g2_o21ai_1 _532_ (.B1(_191_),
    .Y(_192_),
    .A1(_104_),
    .A2(_190_));
 sg13g2_o21ai_1 _533_ (.B1(_167_),
    .Y(_193_),
    .A1(_168_),
    .A2(_171_));
 sg13g2_nand2_1 _534_ (.Y(_194_),
    .A(_176_),
    .B(_179_));
 sg13g2_nand2_1 _535_ (.Y(_195_),
    .A(_177_),
    .B(_194_));
 sg13g2_a221oi_1 _536_ (.B2(_175_),
    .C1(_193_),
    .B1(_195_),
    .A1(_184_),
    .Y(_196_),
    .A2(net93));
 sg13g2_nor2b_1 _537_ (.A(_196_),
    .B_N(_166_),
    .Y(_197_));
 sg13g2_a21oi_1 _538_ (.A1(_159_),
    .A2(_163_),
    .Y(_198_),
    .B1(_158_));
 sg13g2_nor2_1 _539_ (.A(_197_),
    .B(_198_),
    .Y(_199_));
 sg13g2_o21ai_1 _540_ (.B1(_157_),
    .Y(_200_),
    .A1(_197_),
    .A2(_198_));
 sg13g2_nor2b_1 _541_ (.A(_152_),
    .B_N(_154_),
    .Y(_201_));
 sg13g2_a21oi_1 _542_ (.A1(_200_),
    .A2(_201_),
    .Y(_202_),
    .B1(_153_));
 sg13g2_a21o_2 _543_ (.A2(_107_),
    .A1(_105_),
    .B1(_190_),
    .X(_203_));
 sg13g2_a21oi_2 _544_ (.B1(_185_),
    .Y(_204_),
    .A2(_203_),
    .A1(net93));
 sg13g2_a21o_1 _545_ (.A2(_203_),
    .A1(net93),
    .B1(_185_),
    .X(_205_));
 sg13g2_or2_1 _546_ (.X(_206_),
    .B(_153_),
    .A(_152_));
 sg13g2_nor2_1 _547_ (.A(_156_),
    .B(_206_),
    .Y(_207_));
 sg13g2_nand3_1 _548_ (.B(_204_),
    .C(_207_),
    .A(_166_),
    .Y(_208_));
 sg13g2_a21o_1 _549_ (.A2(_208_),
    .A1(_202_),
    .B1(_055_),
    .X(_209_));
 sg13g2_nand2_1 _550_ (.Y(_210_),
    .A(_039_),
    .B(_202_));
 sg13g2_nand4_1 _551_ (.B(_049_),
    .C(_209_),
    .A(net113),
    .Y(_211_),
    .D(_210_));
 sg13g2_and2_1 _552_ (.A(net16),
    .B(_146_),
    .X(_212_));
 sg13g2_o21ai_1 _553_ (.B1(net16),
    .Y(_213_),
    .A1(_040_),
    .A2(_044_));
 sg13g2_o21ai_1 _554_ (.B1(_213_),
    .Y(_214_),
    .A1(net16),
    .A2(_040_));
 sg13g2_inv_1 _555_ (.Y(_215_),
    .A(_214_));
 sg13g2_a221oi_1 _556_ (.B2(net68),
    .C1(_212_),
    .B1(_215_),
    .A1(_045_),
    .Y(_216_),
    .A2(_211_));
 sg13g2_nand2_1 _557_ (.Y(_217_),
    .A(net16),
    .B(_151_));
 sg13g2_o21ai_1 _558_ (.B1(_217_),
    .Y(\gcd_module_inst.fsm_comp.next_state[0] ),
    .A1(_151_),
    .A2(net69));
 sg13g2_a21oi_1 _559_ (.A1(_154_),
    .A2(_200_),
    .Y(_218_),
    .B1(_206_));
 sg13g2_nand3_1 _560_ (.B(_200_),
    .C(_206_),
    .A(_154_),
    .Y(_219_));
 sg13g2_nor2_1 _561_ (.A(net102),
    .B(_218_),
    .Y(_220_));
 sg13g2_a21oi_1 _562_ (.A1(\gcd_module_inst.datapath_comp.RegA_int[15] ),
    .A2(net104),
    .Y(_221_),
    .B1(net98));
 sg13g2_a22oi_1 _563_ (.Y(_222_),
    .B1(_219_),
    .B2(_220_),
    .A2(net96),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[15] ));
 sg13g2_a21oi_1 _564_ (.A1(\gcd_module_inst.datapath_comp.RegB_int[9] ),
    .A2(_036_),
    .Y(_223_),
    .B1(_180_));
 sg13g2_a21o_1 _565_ (.A2(_172_),
    .A1(_167_),
    .B1(_168_),
    .X(_224_));
 sg13g2_a21o_1 _566_ (.A2(_223_),
    .A1(_175_),
    .B1(_224_),
    .X(_225_));
 sg13g2_inv_1 _567_ (.Y(_226_),
    .A(_225_));
 sg13g2_o21ai_1 _568_ (.B1(_166_),
    .Y(_227_),
    .A1(_204_),
    .A2(_225_));
 sg13g2_a21oi_1 _569_ (.A1(_159_),
    .A2(_162_),
    .Y(_228_),
    .B1(_158_));
 sg13g2_a21oi_1 _570_ (.A1(_227_),
    .A2(_228_),
    .Y(_229_),
    .B1(_156_));
 sg13g2_o21ai_1 _571_ (.B1(_206_),
    .Y(_230_),
    .A1(_155_),
    .A2(_229_));
 sg13g2_nor3_1 _572_ (.A(_155_),
    .B(_206_),
    .C(_229_),
    .Y(_231_));
 sg13g2_nor2_1 _573_ (.A(_055_),
    .B(_231_),
    .Y(_232_));
 sg13g2_a221oi_1 _574_ (.B2(_232_),
    .C1(_034_),
    .B1(_230_),
    .A1(_221_),
    .Y(_233_),
    .A2(_222_));
 sg13g2_xnor2_1 _575_ (.Y(_234_),
    .A(_156_),
    .B(_199_));
 sg13g2_a221oi_1 _576_ (.B2(\gcd_module_inst.datapath_comp.RegA_int[14] ),
    .C1(net98),
    .B1(net104),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[14] ),
    .Y(_235_),
    .A2(net96));
 sg13g2_o21ai_1 _577_ (.B1(_235_),
    .Y(_236_),
    .A1(net102),
    .A2(_234_));
 sg13g2_and3_1 _578_ (.X(_237_),
    .A(_156_),
    .B(_227_),
    .C(_228_));
 sg13g2_o21ai_1 _579_ (.B1(net98),
    .Y(_238_),
    .A1(_229_),
    .A2(_237_));
 sg13g2_nand3_1 _580_ (.B(_236_),
    .C(_238_),
    .A(net113),
    .Y(_239_));
 sg13g2_a21o_1 _581_ (.A2(_203_),
    .A1(net93),
    .B1(_181_),
    .X(_240_));
 sg13g2_a221oi_1 _582_ (.B2(_203_),
    .C1(_181_),
    .B1(net93),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[9] ),
    .Y(_241_),
    .A2(_036_));
 sg13g2_a221oi_1 _583_ (.B2(_240_),
    .C1(_173_),
    .B1(_180_),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[9] ),
    .Y(_242_),
    .A2(_036_));
 sg13g2_o21ai_1 _584_ (.B1(_170_),
    .Y(_243_),
    .A1(_172_),
    .A2(_242_));
 sg13g2_nor3_1 _585_ (.A(_170_),
    .B(_172_),
    .C(_242_),
    .Y(_244_));
 sg13g2_nor2_1 _586_ (.A(_055_),
    .B(_244_),
    .Y(_245_));
 sg13g2_a21oi_1 _587_ (.A1(_183_),
    .A2(net93),
    .Y(_246_),
    .B1(_195_));
 sg13g2_o21ai_1 _588_ (.B1(_171_),
    .Y(_247_),
    .A1(_172_),
    .A2(_246_));
 sg13g2_a21oi_1 _589_ (.A1(_169_),
    .A2(_247_),
    .Y(_248_),
    .B1(net103));
 sg13g2_o21ai_1 _590_ (.B1(_248_),
    .Y(_249_),
    .A1(_169_),
    .A2(_247_));
 sg13g2_a221oi_1 _591_ (.B2(\gcd_module_inst.datapath_comp.RegA_int[11] ),
    .C1(net100),
    .B1(net105),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[11] ),
    .Y(_250_),
    .A2(net97));
 sg13g2_a221oi_1 _592_ (.B2(_250_),
    .C1(_034_),
    .B1(_249_),
    .A1(_243_),
    .Y(_251_),
    .A2(_245_));
 sg13g2_o21ai_1 _593_ (.B1(_163_),
    .Y(_252_),
    .A1(_162_),
    .A2(_196_));
 sg13g2_nor2_1 _594_ (.A(_160_),
    .B(_252_),
    .Y(_253_));
 sg13g2_a21o_1 _595_ (.A2(_252_),
    .A1(_160_),
    .B1(net102),
    .X(_254_));
 sg13g2_a221oi_1 _596_ (.B2(\gcd_module_inst.datapath_comp.RegA_int[13] ),
    .C1(net98),
    .B1(net104),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[13] ),
    .Y(_255_),
    .A2(net96));
 sg13g2_o21ai_1 _597_ (.B1(_255_),
    .Y(_256_),
    .A1(_253_),
    .A2(_254_));
 sg13g2_a21oi_1 _598_ (.A1(_205_),
    .A2(_226_),
    .Y(_257_),
    .B1(_165_));
 sg13g2_or3_1 _599_ (.A(_161_),
    .B(_162_),
    .C(_257_),
    .X(_258_));
 sg13g2_o21ai_1 _600_ (.B1(_161_),
    .Y(_259_),
    .A1(_162_),
    .A2(_257_));
 sg13g2_nand3_1 _601_ (.B(_258_),
    .C(_259_),
    .A(net98),
    .Y(_260_));
 sg13g2_nand3_1 _602_ (.B(_256_),
    .C(_260_),
    .A(net113),
    .Y(_261_));
 sg13g2_nor2b_1 _603_ (.A(_251_),
    .B_N(_261_),
    .Y(_262_));
 sg13g2_nor3_1 _604_ (.A(_174_),
    .B(_223_),
    .C(_241_),
    .Y(_263_));
 sg13g2_o21ai_1 _605_ (.B1(net100),
    .Y(_264_),
    .A1(_242_),
    .A2(_263_));
 sg13g2_xnor2_1 _606_ (.Y(_265_),
    .A(_173_),
    .B(_246_));
 sg13g2_a221oi_1 _607_ (.B2(\gcd_module_inst.datapath_comp.RegA_int[10] ),
    .C1(net100),
    .B1(net105),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[10] ),
    .Y(_266_),
    .A2(net97));
 sg13g2_o21ai_1 _608_ (.B1(_266_),
    .Y(_267_),
    .A1(net103),
    .A2(_265_));
 sg13g2_nand3_1 _609_ (.B(_264_),
    .C(_267_),
    .A(net116),
    .Y(_268_));
 sg13g2_nor2_1 _610_ (.A(_034_),
    .B(_059_),
    .Y(_269_));
 sg13g2_and3_1 _611_ (.X(_270_),
    .A(_071_),
    .B(_115_),
    .C(_269_));
 sg13g2_and4_1 _612_ (.A(_084_),
    .B(_098_),
    .C(_126_),
    .D(_270_),
    .X(_271_));
 sg13g2_nand3_1 _613_ (.B(_192_),
    .C(_203_),
    .A(_181_),
    .Y(_272_));
 sg13g2_a21oi_1 _614_ (.A1(_240_),
    .A2(_272_),
    .Y(_273_),
    .B1(_055_));
 sg13g2_xor2_1 _615_ (.B(net93),
    .A(_181_),
    .X(_274_));
 sg13g2_a221oi_1 _616_ (.B2(\gcd_module_inst.datapath_comp.RegA_int[8] ),
    .C1(net101),
    .B1(net105),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[8] ),
    .Y(_275_),
    .A2(net97));
 sg13g2_o21ai_1 _617_ (.B1(_275_),
    .Y(_276_),
    .A1(net103),
    .A2(_274_));
 sg13g2_nand3b_1 _618_ (.B(_276_),
    .C(net118),
    .Y(_277_),
    .A_N(_273_));
 sg13g2_nand3_1 _619_ (.B(_271_),
    .C(_277_),
    .A(_144_),
    .Y(_278_));
 sg13g2_a22oi_1 _620_ (.Y(_279_),
    .B1(_240_),
    .B2(_178_),
    .A2(_179_),
    .A1(_177_));
 sg13g2_nand3_1 _621_ (.B(_180_),
    .C(_240_),
    .A(_177_),
    .Y(_280_));
 sg13g2_nand3b_1 _622_ (.B(_280_),
    .C(net100),
    .Y(_281_),
    .A_N(_279_));
 sg13g2_a21oi_1 _623_ (.A1(_178_),
    .A2(net93),
    .Y(_282_),
    .B1(_176_));
 sg13g2_xnor2_1 _624_ (.Y(_283_),
    .A(_182_),
    .B(_282_));
 sg13g2_a221oi_1 _625_ (.B2(\gcd_module_inst.datapath_comp.RegA_int[9] ),
    .C1(net100),
    .B1(net105),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[9] ),
    .Y(_284_),
    .A2(net97));
 sg13g2_o21ai_1 _626_ (.B1(_284_),
    .Y(_285_),
    .A1(net103),
    .A2(_283_));
 sg13g2_nand3_1 _627_ (.B(_281_),
    .C(_285_),
    .A(net116),
    .Y(_286_));
 sg13g2_nor3_1 _628_ (.A(_164_),
    .B(_204_),
    .C(_225_),
    .Y(_287_));
 sg13g2_o21ai_1 _629_ (.B1(net98),
    .Y(_288_),
    .A1(_257_),
    .A2(_287_));
 sg13g2_xnor2_1 _630_ (.Y(_289_),
    .A(_165_),
    .B(_196_));
 sg13g2_a221oi_1 _631_ (.B2(\gcd_module_inst.datapath_comp.RegA_int[12] ),
    .C1(net98),
    .B1(net104),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[12] ),
    .Y(_290_),
    .A2(net96));
 sg13g2_o21ai_1 _632_ (.B1(_290_),
    .Y(_291_),
    .A1(net102),
    .A2(_289_));
 sg13g2_nand3_1 _633_ (.B(_288_),
    .C(_291_),
    .A(net116),
    .Y(_292_));
 sg13g2_nand3_1 _634_ (.B(_136_),
    .C(_188_),
    .A(_130_),
    .Y(_293_));
 sg13g2_a21oi_1 _635_ (.A1(_130_),
    .A2(_136_),
    .Y(_294_),
    .B1(_188_));
 sg13g2_nor2_1 _636_ (.A(_055_),
    .B(_294_),
    .Y(_295_));
 sg13g2_o21ai_1 _637_ (.B1(_188_),
    .Y(_296_),
    .A1(_129_),
    .A2(_140_));
 sg13g2_nor3_1 _638_ (.A(_129_),
    .B(_140_),
    .C(_188_),
    .Y(_297_));
 sg13g2_nor2_1 _639_ (.A(net102),
    .B(_297_),
    .Y(_298_));
 sg13g2_a21oi_1 _640_ (.A1(\gcd_module_inst.datapath_comp.RegA_int[7] ),
    .A2(net104),
    .Y(_299_),
    .B1(net98));
 sg13g2_a22oi_1 _641_ (.Y(_300_),
    .B1(_296_),
    .B2(_298_),
    .A2(net96),
    .A1(\gcd_module_inst.datapath_comp.RegB_int[7] ));
 sg13g2_a221oi_1 _642_ (.B2(_300_),
    .C1(_034_),
    .B1(_299_),
    .A1(_293_),
    .Y(_301_),
    .A2(_295_));
 sg13g2_nand3_1 _643_ (.B(_286_),
    .C(_292_),
    .A(_268_),
    .Y(_302_));
 sg13g2_nor3_1 _644_ (.A(_278_),
    .B(_301_),
    .C(_302_),
    .Y(_303_));
 sg13g2_nand4_1 _645_ (.B(_239_),
    .C(_262_),
    .A(_211_),
    .Y(_304_),
    .D(_303_));
 sg13g2_o21ai_1 _646_ (.B1(net66),
    .Y(_305_),
    .A1(_233_),
    .A2(_304_));
 sg13g2_a21o_1 _647_ (.A2(net16),
    .A1(net111),
    .B1(_147_),
    .X(_306_));
 sg13g2_a21oi_1 _648_ (.A1(_305_),
    .A2(_306_),
    .Y(\gcd_module_inst.fsm_comp.next_state[1] ),
    .B1(_151_));
 sg13g2_nand3_1 _649_ (.B(net16),
    .C(_040_),
    .A(net68),
    .Y(_307_));
 sg13g2_nor2b_1 _650_ (.A(_212_),
    .B_N(_307_),
    .Y(_308_));
 sg13g2_a21oi_1 _651_ (.A1(_046_),
    .A2(_308_),
    .Y(\gcd_module_inst.fsm_comp.next_state[2] ),
    .B1(_151_));
 sg13g2_nand2_1 _652_ (.Y(_309_),
    .A(\gcd_module_inst.fsm_comp.state[2] ),
    .B(_001_));
 sg13g2_a21oi_1 _653_ (.A1(net109),
    .A2(_309_),
    .Y(ack_w),
    .B1(_150_));
 sg13g2_nor2_1 _654_ (.A(\gcd_module_inst.fsm_comp.state[2] ),
    .B(_044_),
    .Y(_310_));
 sg13g2_nor2_1 _655_ (.A(_038_),
    .B(_310_),
    .Y(_311_));
 sg13g2_nor3_1 _656_ (.A(_045_),
    .B(_148_),
    .C(_311_),
    .Y(_312_));
 sg13g2_mux2_1 _657_ (.A0(net39),
    .A1(\C[0] ),
    .S(net92),
    .X(_002_));
 sg13g2_mux2_1 _658_ (.A0(net48),
    .A1(\C[1] ),
    .S(net92),
    .X(_003_));
 sg13g2_mux2_1 _659_ (.A0(net50),
    .A1(\C[2] ),
    .S(net92),
    .X(_004_));
 sg13g2_mux2_1 _660_ (.A0(net41),
    .A1(\C[3] ),
    .S(net92),
    .X(_005_));
 sg13g2_mux2_1 _661_ (.A0(net61),
    .A1(\C[4] ),
    .S(net91),
    .X(_006_));
 sg13g2_mux2_1 _662_ (.A0(net47),
    .A1(\C[5] ),
    .S(net91),
    .X(_007_));
 sg13g2_mux2_1 _663_ (.A0(net43),
    .A1(\C[6] ),
    .S(net91),
    .X(_008_));
 sg13g2_mux2_1 _664_ (.A0(net8),
    .A1(_301_),
    .S(net108),
    .X(_313_));
 sg13g2_mux2_1 _665_ (.A0(net42),
    .A1(_313_),
    .S(net91),
    .X(_009_));
 sg13g2_nor2_1 _666_ (.A(net9),
    .B(net106),
    .Y(_314_));
 sg13g2_a21oi_1 _667_ (.A1(net108),
    .A2(_277_),
    .Y(_315_),
    .B1(_314_));
 sg13g2_mux2_1 _668_ (.A0(net33),
    .A1(_315_),
    .S(net92),
    .X(_010_));
 sg13g2_nor2_1 _669_ (.A(net10),
    .B(net107),
    .Y(_316_));
 sg13g2_a21oi_1 _670_ (.A1(net108),
    .A2(_286_),
    .Y(_317_),
    .B1(_316_));
 sg13g2_mux2_1 _671_ (.A0(net56),
    .A1(_317_),
    .S(net92),
    .X(_011_));
 sg13g2_nor2_1 _672_ (.A(net11),
    .B(net107),
    .Y(_318_));
 sg13g2_a21oi_1 _673_ (.A1(net108),
    .A2(_268_),
    .Y(_319_),
    .B1(_318_));
 sg13g2_mux2_1 _674_ (.A0(net51),
    .A1(_319_),
    .S(net92),
    .X(_012_));
 sg13g2_mux2_1 _675_ (.A0(net12),
    .A1(_251_),
    .S(net108),
    .X(_320_));
 sg13g2_mux2_1 _676_ (.A0(net64),
    .A1(_320_),
    .S(net92),
    .X(_013_));
 sg13g2_nor2_1 _677_ (.A(net13),
    .B(net109),
    .Y(_321_));
 sg13g2_a21oi_1 _678_ (.A1(net108),
    .A2(_292_),
    .Y(_322_),
    .B1(_321_));
 sg13g2_mux2_1 _679_ (.A0(net37),
    .A1(_322_),
    .S(net91),
    .X(_014_));
 sg13g2_nor2_1 _680_ (.A(net14),
    .B(net109),
    .Y(_323_));
 sg13g2_a21oi_1 _681_ (.A1(net109),
    .A2(_261_),
    .Y(_324_),
    .B1(_323_));
 sg13g2_mux2_1 _682_ (.A0(net35),
    .A1(_324_),
    .S(net91),
    .X(_015_));
 sg13g2_nor2_1 _683_ (.A(net15),
    .B(net109),
    .Y(_325_));
 sg13g2_a21oi_1 _684_ (.A1(net109),
    .A2(_239_),
    .Y(_326_),
    .B1(_325_));
 sg13g2_mux2_1 _685_ (.A0(net45),
    .A1(_326_),
    .S(net91),
    .X(_016_));
 sg13g2_and2_1 _686_ (.A(net109),
    .B(_233_),
    .X(_327_));
 sg13g2_mux2_1 _687_ (.A0(net34),
    .A1(_327_),
    .S(net91),
    .X(_017_));
 sg13g2_a21oi_2 _688_ (.B1(_041_),
    .Y(_328_),
    .A2(_145_),
    .A1(_000_));
 sg13g2_mux2_1 _689_ (.A0(\C[0] ),
    .A1(net49),
    .S(_328_),
    .X(_018_));
 sg13g2_mux2_1 _690_ (.A0(\C[1] ),
    .A1(net60),
    .S(net95),
    .X(_019_));
 sg13g2_mux2_1 _691_ (.A0(\C[2] ),
    .A1(net54),
    .S(_328_),
    .X(_020_));
 sg13g2_mux2_1 _692_ (.A0(\C[3] ),
    .A1(net46),
    .S(net95),
    .X(_021_));
 sg13g2_mux2_1 _693_ (.A0(\C[4] ),
    .A1(net55),
    .S(net94),
    .X(_022_));
 sg13g2_mux2_1 _694_ (.A0(\C[5] ),
    .A1(net57),
    .S(net94),
    .X(_023_));
 sg13g2_mux2_1 _695_ (.A0(\C[6] ),
    .A1(net62),
    .S(net94),
    .X(_024_));
 sg13g2_mux2_1 _696_ (.A0(_313_),
    .A1(net59),
    .S(net94),
    .X(_025_));
 sg13g2_mux2_1 _697_ (.A0(_315_),
    .A1(net36),
    .S(net95),
    .X(_026_));
 sg13g2_nor2_1 _698_ (.A(_317_),
    .B(net95),
    .Y(_329_));
 sg13g2_a21oi_1 _699_ (.A1(_036_),
    .A2(net95),
    .Y(_027_),
    .B1(_329_));
 sg13g2_mux2_1 _700_ (.A0(_319_),
    .A1(net58),
    .S(net95),
    .X(_028_));
 sg13g2_mux2_1 _701_ (.A0(_320_),
    .A1(net63),
    .S(net95),
    .X(_029_));
 sg13g2_mux2_1 _702_ (.A0(_322_),
    .A1(net44),
    .S(net94),
    .X(_030_));
 sg13g2_mux2_1 _703_ (.A0(_324_),
    .A1(net40),
    .S(net94),
    .X(_031_));
 sg13g2_mux2_1 _704_ (.A0(_326_),
    .A1(net53),
    .S(net94),
    .X(_032_));
 sg13g2_mux2_1 _705_ (.A0(_327_),
    .A1(net38),
    .S(net94),
    .X(_033_));
 sg13g2_dfrbp_1 _706_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net118),
    .D(_002_),
    .Q_N(_362_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[0] ));
 sg13g2_dfrbp_1 _707_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net118),
    .D(_003_),
    .Q_N(_361_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[1] ));
 sg13g2_dfrbp_1 _708_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net119),
    .D(_004_),
    .Q_N(_360_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[2] ));
 sg13g2_dfrbp_1 _709_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net119),
    .D(_005_),
    .Q_N(_359_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[3] ));
 sg13g2_dfrbp_1 _710_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net115),
    .D(_006_),
    .Q_N(_358_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[4] ));
 sg13g2_dfrbp_1 _711_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net114),
    .D(_007_),
    .Q_N(_357_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[5] ));
 sg13g2_dfrbp_1 _712_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net114),
    .D(_008_),
    .Q_N(_356_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[6] ));
 sg13g2_dfrbp_1 _713_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net112),
    .D(_009_),
    .Q_N(_355_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[7] ));
 sg13g2_dfrbp_1 _714_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net118),
    .D(_010_),
    .Q_N(_354_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[8] ));
 sg13g2_dfrbp_1 _715_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net117),
    .D(_011_),
    .Q_N(_353_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[9] ));
 sg13g2_dfrbp_1 _716_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net117),
    .D(_012_),
    .Q_N(_352_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[10] ));
 sg13g2_dfrbp_1 _717_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net116),
    .D(_013_),
    .Q_N(_351_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[11] ));
 sg13g2_dfrbp_1 _718_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net116),
    .D(_014_),
    .Q_N(_350_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[12] ));
 sg13g2_dfrbp_1 _719_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net113),
    .D(_015_),
    .Q_N(_349_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[13] ));
 sg13g2_dfrbp_1 _720_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net112),
    .D(_016_),
    .Q_N(_348_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[14] ));
 sg13g2_dfrbp_1 _721_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net112),
    .D(_017_),
    .Q_N(_347_),
    .Q(\gcd_module_inst.datapath_comp.RegB_int[15] ));
 sg13g2_dfrbp_1 _722_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net118),
    .D(_018_),
    .Q_N(_346_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[0] ));
 sg13g2_dfrbp_1 _723_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net118),
    .D(_019_),
    .Q_N(_345_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[1] ));
 sg13g2_dfrbp_1 _724_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net119),
    .D(_020_),
    .Q_N(_344_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[2] ));
 sg13g2_dfrbp_1 _725_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net119),
    .D(_021_),
    .Q_N(_343_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[3] ));
 sg13g2_dfrbp_1 _726_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net114),
    .D(_022_),
    .Q_N(_342_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[4] ));
 sg13g2_dfrbp_1 _727_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net114),
    .D(_023_),
    .Q_N(_341_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[5] ));
 sg13g2_dfrbp_1 _728_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net114),
    .D(_024_),
    .Q_N(_340_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[6] ));
 sg13g2_dfrbp_1 _729_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net116),
    .D(_025_),
    .Q_N(_339_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[7] ));
 sg13g2_dfrbp_1 _730_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net118),
    .D(_026_),
    .Q_N(_338_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[8] ));
 sg13g2_dfrbp_1 _731_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net117),
    .D(_027_),
    .Q_N(_337_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[9] ));
 sg13g2_dfrbp_1 _732_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net117),
    .D(_028_),
    .Q_N(_336_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[10] ));
 sg13g2_dfrbp_1 _733_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net116),
    .D(_029_),
    .Q_N(_335_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[11] ));
 sg13g2_dfrbp_1 _734_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net116),
    .D(_030_),
    .Q_N(_334_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[12] ));
 sg13g2_dfrbp_1 _735_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net112),
    .D(_031_),
    .Q_N(_333_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[13] ));
 sg13g2_dfrbp_1 _736_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net112),
    .D(_032_),
    .Q_N(_332_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[14] ));
 sg13g2_dfrbp_1 _737_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net112),
    .D(_033_),
    .Q_N(_363_),
    .Q(\gcd_module_inst.datapath_comp.RegA_int[15] ));
 sg13g2_dfrbp_1 _738_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net112),
    .D(\gcd_module_inst.fsm_comp.next_state[0] ),
    .Q_N(_364_),
    .Q(\gcd_module_inst.fsm_comp.state[0] ));
 sg13g2_dfrbp_1 _739_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net114),
    .D(net67),
    .Q_N(_001_),
    .Q(\gcd_module_inst.fsm_comp.state[1] ));
 sg13g2_dfrbp_1 _740_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net114),
    .D(\gcd_module_inst.fsm_comp.next_state[2] ),
    .Q_N(_000_),
    .Q(\gcd_module_inst.fsm_comp.state[2] ));
 sg13g2_tielo tt_um_gcd_stephan_18 (.L_LO(net18));
 sg13g2_tielo tt_um_gcd_stephan_19 (.L_LO(net19));
 sg13g2_tielo tt_um_gcd_stephan_20 (.L_LO(net20));
 sg13g2_tielo tt_um_gcd_stephan_21 (.L_LO(net21));
 sg13g2_tielo tt_um_gcd_stephan_22 (.L_LO(net22));
 sg13g2_tielo tt_um_gcd_stephan_23 (.L_LO(net23));
 sg13g2_tielo tt_um_gcd_stephan_24 (.L_LO(net24));
 sg13g2_tielo tt_um_gcd_stephan_25 (.L_LO(net25));
 sg13g2_tielo tt_um_gcd_stephan_26 (.L_LO(net26));
 sg13g2_tielo tt_um_gcd_stephan_27 (.L_LO(net27));
 sg13g2_tielo tt_um_gcd_stephan_28 (.L_LO(net28));
 sg13g2_tielo tt_um_gcd_stephan_29 (.L_LO(net29));
 sg13g2_tielo tt_um_gcd_stephan_30 (.L_LO(net30));
 sg13g2_tielo tt_um_gcd_stephan_31 (.L_LO(net31));
 sg13g2_tielo tt_um_gcd_stephan_32 (.L_LO(net32));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _757_ (.A(\C[0] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _758_ (.A(\C[1] ),
    .X(uo_out[1]));
 sg13g2_buf_1 _759_ (.A(\C[2] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _760_ (.A(\C[3] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _761_ (.A(\C[4] ),
    .X(uo_out[4]));
 sg13g2_buf_1 _762_ (.A(\C[5] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _763_ (.A(\C[6] ),
    .X(uo_out[6]));
 sg13g2_buf_1 _764_ (.A(ack_w),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout91 (.X(net91),
    .A(_312_));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(_312_));
 sg13g2_buf_2 fanout93 (.A(_192_),
    .X(net93));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(net95));
 sg13g2_buf_4 fanout95 (.X(net95),
    .A(_328_));
 sg13g2_buf_2 fanout96 (.A(_056_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_056_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(net101),
    .X(net98));
 sg13g2_buf_1 fanout99 (.A(net101),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(net101),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_054_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_062_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_062_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_057_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_057_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(net108),
    .X(net106));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(net108));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(_037_));
 sg13g2_buf_2 fanout109 (.A(_037_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(\gcd_module_inst.fsm_comp.state[1] ),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(\gcd_module_inst.fsm_comp.state[0] ),
    .X(net111));
 sg13g2_buf_4 fanout112 (.X(net112),
    .A(net115));
 sg13g2_buf_2 fanout113 (.A(net115),
    .X(net113));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(net115));
 sg13g2_buf_2 fanout115 (.A(net120),
    .X(net115));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(net120));
 sg13g2_buf_2 fanout117 (.A(net120),
    .X(net117));
 sg13g2_buf_4 fanout118 (.X(net118),
    .A(net119));
 sg13g2_buf_4 fanout119 (.X(net119),
    .A(net120));
 sg13g2_buf_2 fanout120 (.A(rst_n),
    .X(net120));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_2 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_tielo tt_um_gcd_stephan_17 (.L_LO(net17));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\gcd_module_inst.datapath_comp.RegB_int[8] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold2 (.A(\gcd_module_inst.datapath_comp.RegB_int[15] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold3 (.A(\gcd_module_inst.datapath_comp.RegB_int[13] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold4 (.A(\gcd_module_inst.datapath_comp.RegA_int[8] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold5 (.A(\gcd_module_inst.datapath_comp.RegB_int[12] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold6 (.A(\gcd_module_inst.datapath_comp.RegA_int[15] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold7 (.A(\gcd_module_inst.datapath_comp.RegB_int[0] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold8 (.A(\gcd_module_inst.datapath_comp.RegA_int[13] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold9 (.A(\gcd_module_inst.datapath_comp.RegB_int[3] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold10 (.A(\gcd_module_inst.datapath_comp.RegB_int[7] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold11 (.A(\gcd_module_inst.datapath_comp.RegB_int[6] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold12 (.A(\gcd_module_inst.datapath_comp.RegA_int[12] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold13 (.A(\gcd_module_inst.datapath_comp.RegB_int[14] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold14 (.A(\gcd_module_inst.datapath_comp.RegA_int[3] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold15 (.A(\gcd_module_inst.datapath_comp.RegB_int[5] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold16 (.A(\gcd_module_inst.datapath_comp.RegB_int[1] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold17 (.A(\gcd_module_inst.datapath_comp.RegA_int[0] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold18 (.A(\gcd_module_inst.datapath_comp.RegB_int[2] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold19 (.A(\gcd_module_inst.datapath_comp.RegB_int[10] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold20 (.A(\gcd_module_inst.datapath_comp.RegA_int[9] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold21 (.A(\gcd_module_inst.datapath_comp.RegA_int[14] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold22 (.A(\gcd_module_inst.datapath_comp.RegA_int[2] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold23 (.A(\gcd_module_inst.datapath_comp.RegA_int[4] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold24 (.A(\gcd_module_inst.datapath_comp.RegB_int[9] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold25 (.A(\gcd_module_inst.datapath_comp.RegA_int[5] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold26 (.A(\gcd_module_inst.datapath_comp.RegA_int[10] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold27 (.A(\gcd_module_inst.datapath_comp.RegA_int[7] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold28 (.A(\gcd_module_inst.datapath_comp.RegA_int[1] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold29 (.A(\gcd_module_inst.datapath_comp.RegB_int[4] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold30 (.A(\gcd_module_inst.datapath_comp.RegA_int[6] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold31 (.A(\gcd_module_inst.datapath_comp.RegA_int[11] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold32 (.A(\gcd_module_inst.datapath_comp.RegB_int[11] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold33 (.A(\gcd_module_inst.fsm_comp.state[0] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold34 (.A(_045_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold35 (.A(\gcd_module_inst.fsm_comp.next_state[1] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold36 (.A(_000_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold37 (.A(_216_),
    .X(net69));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_fill_2 FILLER_19_231 ();
 sg13g2_fill_1 FILLER_19_233 ();
 sg13g2_decap_8 FILLER_19_260 ();
 sg13g2_decap_8 FILLER_19_267 ();
 sg13g2_decap_8 FILLER_19_274 ();
 sg13g2_fill_2 FILLER_19_281 ();
 sg13g2_fill_1 FILLER_19_283 ();
 sg13g2_decap_8 FILLER_19_310 ();
 sg13g2_decap_8 FILLER_19_317 ();
 sg13g2_decap_8 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_331 ();
 sg13g2_decap_8 FILLER_19_338 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_fill_2 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_233 ();
 sg13g2_decap_4 FILLER_20_260 ();
 sg13g2_fill_2 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_302 ();
 sg13g2_decap_8 FILLER_20_309 ();
 sg13g2_decap_4 FILLER_20_316 ();
 sg13g2_decap_8 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_353 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_fill_2 FILLER_21_182 ();
 sg13g2_fill_1 FILLER_21_184 ();
 sg13g2_decap_4 FILLER_21_221 ();
 sg13g2_decap_4 FILLER_21_239 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_decap_8 FILLER_21_262 ();
 sg13g2_decap_4 FILLER_21_269 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_fill_2 FILLER_21_315 ();
 sg13g2_fill_1 FILLER_21_317 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_168 ();
 sg13g2_fill_1 FILLER_22_224 ();
 sg13g2_fill_2 FILLER_22_235 ();
 sg13g2_decap_8 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_255 ();
 sg13g2_decap_4 FILLER_22_275 ();
 sg13g2_decap_4 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_295 ();
 sg13g2_decap_4 FILLER_22_302 ();
 sg13g2_fill_1 FILLER_22_306 ();
 sg13g2_fill_1 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_fill_2 FILLER_22_378 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_fill_2 FILLER_23_189 ();
 sg13g2_fill_1 FILLER_23_196 ();
 sg13g2_fill_2 FILLER_23_206 ();
 sg13g2_fill_1 FILLER_23_208 ();
 sg13g2_fill_2 FILLER_23_245 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_fill_1 FILLER_23_311 ();
 sg13g2_decap_4 FILLER_23_322 ();
 sg13g2_fill_2 FILLER_23_326 ();
 sg13g2_fill_2 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_368 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_4 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_fill_1 FILLER_24_203 ();
 sg13g2_decap_4 FILLER_24_214 ();
 sg13g2_fill_2 FILLER_24_218 ();
 sg13g2_decap_8 FILLER_24_232 ();
 sg13g2_fill_2 FILLER_24_239 ();
 sg13g2_fill_2 FILLER_24_283 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_310 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_fill_2 FILLER_24_325 ();
 sg13g2_fill_1 FILLER_24_327 ();
 sg13g2_fill_2 FILLER_24_358 ();
 sg13g2_fill_2 FILLER_24_368 ();
 sg13g2_fill_1 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_fill_2 FILLER_24_388 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_4 FILLER_25_154 ();
 sg13g2_fill_1 FILLER_25_158 ();
 sg13g2_decap_4 FILLER_25_185 ();
 sg13g2_decap_4 FILLER_25_208 ();
 sg13g2_fill_1 FILLER_25_262 ();
 sg13g2_fill_1 FILLER_25_278 ();
 sg13g2_decap_4 FILLER_25_304 ();
 sg13g2_fill_1 FILLER_25_336 ();
 sg13g2_fill_1 FILLER_25_352 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_168 ();
 sg13g2_decap_4 FILLER_26_173 ();
 sg13g2_decap_4 FILLER_26_181 ();
 sg13g2_decap_4 FILLER_26_199 ();
 sg13g2_fill_2 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_fill_2 FILLER_26_238 ();
 sg13g2_decap_4 FILLER_26_245 ();
 sg13g2_fill_2 FILLER_26_257 ();
 sg13g2_decap_4 FILLER_26_262 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_fill_2 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_299 ();
 sg13g2_decap_4 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_decap_8 FILLER_26_323 ();
 sg13g2_fill_2 FILLER_26_330 ();
 sg13g2_fill_2 FILLER_26_363 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_fill_2 FILLER_26_383 ();
 sg13g2_fill_1 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_fill_1 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_174 ();
 sg13g2_fill_1 FILLER_27_198 ();
 sg13g2_decap_4 FILLER_27_215 ();
 sg13g2_fill_1 FILLER_27_219 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_2 FILLER_27_271 ();
 sg13g2_decap_4 FILLER_27_283 ();
 sg13g2_fill_2 FILLER_27_301 ();
 sg13g2_decap_4 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_315 ();
 sg13g2_fill_2 FILLER_27_333 ();
 sg13g2_fill_2 FILLER_27_357 ();
 sg13g2_decap_4 FILLER_27_367 ();
 sg13g2_fill_1 FILLER_27_371 ();
 sg13g2_fill_1 FILLER_27_380 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_4 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_137 ();
 sg13g2_fill_1 FILLER_28_161 ();
 sg13g2_fill_2 FILLER_28_180 ();
 sg13g2_decap_4 FILLER_28_218 ();
 sg13g2_fill_2 FILLER_28_227 ();
 sg13g2_decap_4 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_251 ();
 sg13g2_fill_2 FILLER_28_317 ();
 sg13g2_fill_1 FILLER_28_319 ();
 sg13g2_decap_4 FILLER_28_351 ();
 sg13g2_fill_1 FILLER_28_360 ();
 sg13g2_fill_2 FILLER_28_369 ();
 sg13g2_decap_4 FILLER_28_379 ();
 sg13g2_fill_1 FILLER_28_383 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_4 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_fill_2 FILLER_29_161 ();
 sg13g2_fill_1 FILLER_29_168 ();
 sg13g2_fill_1 FILLER_29_203 ();
 sg13g2_fill_2 FILLER_29_209 ();
 sg13g2_fill_1 FILLER_29_211 ();
 sg13g2_decap_8 FILLER_29_216 ();
 sg13g2_decap_4 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_237 ();
 sg13g2_decap_4 FILLER_29_244 ();
 sg13g2_fill_1 FILLER_29_248 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_276 ();
 sg13g2_decap_8 FILLER_29_283 ();
 sg13g2_decap_8 FILLER_29_290 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_299 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_fill_2 FILLER_29_322 ();
 sg13g2_decap_4 FILLER_29_339 ();
 sg13g2_fill_2 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_fill_1 FILLER_29_370 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_135 ();
 sg13g2_fill_1 FILLER_30_161 ();
 sg13g2_fill_1 FILLER_30_189 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_decap_4 FILLER_30_290 ();
 sg13g2_fill_2 FILLER_30_294 ();
 sg13g2_fill_2 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_303 ();
 sg13g2_decap_8 FILLER_30_309 ();
 sg13g2_decap_4 FILLER_30_316 ();
 sg13g2_fill_1 FILLER_30_325 ();
 sg13g2_decap_4 FILLER_30_331 ();
 sg13g2_fill_2 FILLER_30_335 ();
 sg13g2_fill_2 FILLER_30_342 ();
 sg13g2_fill_2 FILLER_30_351 ();
 sg13g2_fill_1 FILLER_30_353 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_fill_1 FILLER_31_147 ();
 sg13g2_fill_1 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_212 ();
 sg13g2_decap_4 FILLER_31_219 ();
 sg13g2_fill_1 FILLER_31_223 ();
 sg13g2_decap_8 FILLER_31_229 ();
 sg13g2_fill_1 FILLER_31_236 ();
 sg13g2_fill_2 FILLER_31_247 ();
 sg13g2_fill_1 FILLER_31_249 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_fill_1 FILLER_31_266 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_fill_2 FILLER_31_281 ();
 sg13g2_fill_1 FILLER_31_283 ();
 sg13g2_decap_4 FILLER_31_327 ();
 sg13g2_fill_2 FILLER_31_331 ();
 sg13g2_decap_4 FILLER_31_338 ();
 sg13g2_decap_8 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_31_354 ();
 sg13g2_decap_4 FILLER_31_361 ();
 sg13g2_fill_2 FILLER_31_381 ();
 sg13g2_fill_2 FILLER_31_388 ();
 sg13g2_fill_1 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_4 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_fill_2 FILLER_32_221 ();
 sg13g2_fill_1 FILLER_32_223 ();
 sg13g2_fill_1 FILLER_32_233 ();
 sg13g2_fill_2 FILLER_32_254 ();
 sg13g2_fill_2 FILLER_32_268 ();
 sg13g2_fill_1 FILLER_32_285 ();
 sg13g2_fill_1 FILLER_32_301 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_fill_1 FILLER_32_321 ();
 sg13g2_decap_4 FILLER_32_327 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_fill_1 FILLER_32_369 ();
 sg13g2_fill_2 FILLER_32_383 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_182 ();
 sg13g2_fill_1 FILLER_33_184 ();
 sg13g2_fill_1 FILLER_33_230 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_262 ();
 sg13g2_decap_4 FILLER_33_269 ();
 sg13g2_fill_1 FILLER_33_273 ();
 sg13g2_fill_2 FILLER_33_278 ();
 sg13g2_fill_1 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_293 ();
 sg13g2_fill_2 FILLER_33_341 ();
 sg13g2_fill_2 FILLER_33_351 ();
 sg13g2_fill_1 FILLER_33_353 ();
 sg13g2_decap_8 FILLER_33_359 ();
 sg13g2_fill_2 FILLER_33_366 ();
 sg13g2_decap_4 FILLER_33_382 ();
 sg13g2_fill_2 FILLER_33_386 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_4 FILLER_34_168 ();
 sg13g2_fill_1 FILLER_34_172 ();
 sg13g2_fill_2 FILLER_34_199 ();
 sg13g2_fill_1 FILLER_34_201 ();
 sg13g2_fill_1 FILLER_34_252 ();
 sg13g2_decap_4 FILLER_34_268 ();
 sg13g2_fill_2 FILLER_34_272 ();
 sg13g2_decap_8 FILLER_34_291 ();
 sg13g2_decap_8 FILLER_34_298 ();
 sg13g2_fill_2 FILLER_34_313 ();
 sg13g2_decap_4 FILLER_34_319 ();
 sg13g2_fill_1 FILLER_34_323 ();
 sg13g2_fill_1 FILLER_34_361 ();
 sg13g2_fill_1 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_4 FILLER_35_168 ();
 sg13g2_decap_4 FILLER_35_198 ();
 sg13g2_fill_1 FILLER_35_202 ();
 sg13g2_fill_2 FILLER_35_233 ();
 sg13g2_fill_1 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_383 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_4 FILLER_36_189 ();
 sg13g2_fill_2 FILLER_36_193 ();
 sg13g2_decap_4 FILLER_36_214 ();
 sg13g2_fill_1 FILLER_36_218 ();
 sg13g2_decap_4 FILLER_36_233 ();
 sg13g2_decap_4 FILLER_36_245 ();
 sg13g2_fill_2 FILLER_36_249 ();
 sg13g2_fill_2 FILLER_36_266 ();
 sg13g2_fill_1 FILLER_36_268 ();
 sg13g2_fill_2 FILLER_36_290 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_fill_2 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_fill_1 FILLER_37_224 ();
 sg13g2_fill_2 FILLER_37_265 ();
 sg13g2_fill_1 FILLER_37_267 ();
 sg13g2_fill_2 FILLER_37_277 ();
 sg13g2_fill_1 FILLER_37_279 ();
 sg13g2_fill_2 FILLER_37_300 ();
 sg13g2_fill_1 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_313 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_4 FILLER_38_236 ();
 sg13g2_fill_2 FILLER_38_240 ();
 sg13g2_fill_2 FILLER_38_282 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_1 FILLER_38_348 ();
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net25;
 assign uio_out[1] = net26;
 assign uio_out[2] = net27;
 assign uio_out[3] = net28;
 assign uio_out[4] = net29;
 assign uio_out[5] = net30;
 assign uio_out[6] = net31;
 assign uio_out[7] = net32;
endmodule

module tt_um_MichaelBell_tinyQV (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire clk_regs;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire \addr[0] ;
 wire \addr[10] ;
 wire \addr[11] ;
 wire \addr[12] ;
 wire \addr[13] ;
 wire \addr[14] ;
 wire \addr[15] ;
 wire \addr[16] ;
 wire \addr[17] ;
 wire \addr[18] ;
 wire \addr[19] ;
 wire \addr[1] ;
 wire \addr[20] ;
 wire \addr[21] ;
 wire \addr[22] ;
 wire \addr[23] ;
 wire \addr[24] ;
 wire \addr[25] ;
 wire \addr[26] ;
 wire \addr[27] ;
 wire \addr[2] ;
 wire \addr[3] ;
 wire \addr[4] ;
 wire \addr[5] ;
 wire \addr[6] ;
 wire \addr[7] ;
 wire \addr[8] ;
 wire \addr[9] ;
 wire \controller1_data[0] ;
 wire \controller1_data[10] ;
 wire \controller1_data[11] ;
 wire \controller1_data[1] ;
 wire \controller1_data[2] ;
 wire \controller1_data[3] ;
 wire \controller1_data[4] ;
 wire \controller1_data[5] ;
 wire \controller1_data[6] ;
 wire \controller1_data[7] ;
 wire \controller1_data[8] ;
 wire \controller1_data[9] ;
 wire \controller2_data[0] ;
 wire \controller2_data[10] ;
 wire \controller2_data[11] ;
 wire \controller2_data[1] ;
 wire \controller2_data[2] ;
 wire \controller2_data[3] ;
 wire \controller2_data[4] ;
 wire \controller2_data[5] ;
 wire \controller2_data[6] ;
 wire \controller2_data[7] ;
 wire \controller2_data[8] ;
 wire \controller2_data[9] ;
 wire \data_to_write[0] ;
 wire \data_to_write[10] ;
 wire \data_to_write[11] ;
 wire \data_to_write[12] ;
 wire \data_to_write[13] ;
 wire \data_to_write[14] ;
 wire \data_to_write[15] ;
 wire \data_to_write[16] ;
 wire \data_to_write[17] ;
 wire \data_to_write[18] ;
 wire \data_to_write[19] ;
 wire \data_to_write[1] ;
 wire \data_to_write[20] ;
 wire \data_to_write[21] ;
 wire \data_to_write[22] ;
 wire \data_to_write[23] ;
 wire \data_to_write[24] ;
 wire \data_to_write[25] ;
 wire \data_to_write[26] ;
 wire \data_to_write[27] ;
 wire \data_to_write[28] ;
 wire \data_to_write[29] ;
 wire \data_to_write[2] ;
 wire \data_to_write[30] ;
 wire \data_to_write[31] ;
 wire \data_to_write[3] ;
 wire \data_to_write[4] ;
 wire \data_to_write[5] ;
 wire \data_to_write[6] ;
 wire \data_to_write[7] ;
 wire \data_to_write[8] ;
 wire \data_to_write[9] ;
 wire debug_data_continue;
 wire debug_instr_valid;
 wire \debug_rd[0] ;
 wire \debug_rd[1] ;
 wire \debug_rd[2] ;
 wire \debug_rd[3] ;
 wire \debug_rd_r[0] ;
 wire \debug_rd_r[1] ;
 wire \debug_rd_r[2] ;
 wire \debug_rd_r[3] ;
 wire debug_register_data;
 wire debug_uart_txd;
 wire game_clk;
 wire \gpio_out[0] ;
 wire \gpio_out[1] ;
 wire \gpio_out[2] ;
 wire \gpio_out[3] ;
 wire \gpio_out[4] ;
 wire \gpio_out[5] ;
 wire \gpio_out[6] ;
 wire \gpio_out[7] ;
 wire \gpio_out_sel[0] ;
 wire \gpio_out_sel[1] ;
 wire \gpio_out_sel[2] ;
 wire \gpio_out_sel[3] ;
 wire \gpio_out_sel[4] ;
 wire \gpio_out_sel[5] ;
 wire \gpio_out_sel[6] ;
 wire \gpio_out_sel[7] ;
 wire \gpio_out_sel[8] ;
 wire \gpio_out_sel[9] ;
 wire \i_debug_uart_tx.cycle_counter[0] ;
 wire \i_debug_uart_tx.cycle_counter[1] ;
 wire \i_debug_uart_tx.cycle_counter[2] ;
 wire \i_debug_uart_tx.cycle_counter[3] ;
 wire \i_debug_uart_tx.cycle_counter[4] ;
 wire \i_debug_uart_tx.data_to_send[0] ;
 wire \i_debug_uart_tx.data_to_send[1] ;
 wire \i_debug_uart_tx.data_to_send[2] ;
 wire \i_debug_uart_tx.data_to_send[3] ;
 wire \i_debug_uart_tx.data_to_send[4] ;
 wire \i_debug_uart_tx.data_to_send[5] ;
 wire \i_debug_uart_tx.data_to_send[6] ;
 wire \i_debug_uart_tx.data_to_send[7] ;
 wire \i_debug_uart_tx.fsm_state[0] ;
 wire \i_debug_uart_tx.fsm_state[1] ;
 wire \i_debug_uart_tx.fsm_state[2] ;
 wire \i_debug_uart_tx.fsm_state[3] ;
 wire \i_debug_uart_tx.resetn ;
 wire \i_game.data_latch_wen ;
 wire net656;
 wire \i_game.game_latch_sync[0] ;
 wire \i_game.game_latch_sync[1] ;
 wire \i_game.l_data.data_in[0] ;
 wire \i_game.l_data.data_in[10] ;
 wire \i_game.l_data.data_in[11] ;
 wire \i_game.l_data.data_in[12] ;
 wire \i_game.l_data.data_in[13] ;
 wire \i_game.l_data.data_in[14] ;
 wire \i_game.l_data.data_in[15] ;
 wire \i_game.l_data.data_in[16] ;
 wire \i_game.l_data.data_in[17] ;
 wire \i_game.l_data.data_in[18] ;
 wire \i_game.l_data.data_in[19] ;
 wire \i_game.l_data.data_in[1] ;
 wire \i_game.l_data.data_in[20] ;
 wire \i_game.l_data.data_in[21] ;
 wire \i_game.l_data.data_in[22] ;
 wire \i_game.l_data.data_in[23] ;
 wire \i_game.l_data.data_in[2] ;
 wire \i_game.l_data.data_in[3] ;
 wire \i_game.l_data.data_in[4] ;
 wire \i_game.l_data.data_in[5] ;
 wire \i_game.l_data.data_in[6] ;
 wire \i_game.l_data.data_in[7] ;
 wire \i_game.l_data.data_in[8] ;
 wire \i_game.l_data.data_in[9] ;
 wire \i_latch_mem.cycle[0] ;
 wire \i_latch_mem.cycle[1] ;
 wire \i_latch_mem.data_out[0] ;
 wire \i_latch_mem.data_out[10] ;
 wire \i_latch_mem.data_out[11] ;
 wire \i_latch_mem.data_out[12] ;
 wire \i_latch_mem.data_out[13] ;
 wire \i_latch_mem.data_out[14] ;
 wire \i_latch_mem.data_out[15] ;
 wire \i_latch_mem.data_out[16] ;
 wire \i_latch_mem.data_out[17] ;
 wire \i_latch_mem.data_out[18] ;
 wire \i_latch_mem.data_out[19] ;
 wire \i_latch_mem.data_out[1] ;
 wire \i_latch_mem.data_out[20] ;
 wire \i_latch_mem.data_out[21] ;
 wire \i_latch_mem.data_out[22] ;
 wire \i_latch_mem.data_out[23] ;
 wire \i_latch_mem.data_out[24] ;
 wire \i_latch_mem.data_out[25] ;
 wire \i_latch_mem.data_out[26] ;
 wire \i_latch_mem.data_out[27] ;
 wire \i_latch_mem.data_out[28] ;
 wire \i_latch_mem.data_out[29] ;
 wire \i_latch_mem.data_out[2] ;
 wire \i_latch_mem.data_out[30] ;
 wire \i_latch_mem.data_out[31] ;
 wire \i_latch_mem.data_out[3] ;
 wire \i_latch_mem.data_out[4] ;
 wire \i_latch_mem.data_out[5] ;
 wire \i_latch_mem.data_out[6] ;
 wire \i_latch_mem.data_out[7] ;
 wire \i_latch_mem.data_out[8] ;
 wire \i_latch_mem.data_out[9] ;
 wire \i_latch_mem.data_ready ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[7] ;
 wire \i_pwm.l_pwm_level.data_out[0] ;
 wire \i_pwm.l_pwm_level.data_out[1] ;
 wire \i_pwm.l_pwm_level.data_out[2] ;
 wire \i_pwm.l_pwm_level.data_out[3] ;
 wire \i_pwm.l_pwm_level.data_out[4] ;
 wire \i_pwm.l_pwm_level.data_out[5] ;
 wire \i_pwm.l_pwm_level.data_out[6] ;
 wire \i_pwm.l_pwm_level.data_out[7] ;
 wire \i_pwm.pwm ;
 wire \i_pwm.pwm_count[0] ;
 wire \i_pwm.pwm_count[1] ;
 wire \i_pwm.pwm_count[2] ;
 wire \i_pwm.pwm_count[3] ;
 wire \i_pwm.pwm_count[4] ;
 wire \i_pwm.pwm_count[5] ;
 wire \i_pwm.pwm_count[6] ;
 wire \i_pwm.pwm_count[7] ;
 wire \i_spi.bits_remaining[0] ;
 wire \i_spi.bits_remaining[1] ;
 wire \i_spi.bits_remaining[2] ;
 wire \i_spi.bits_remaining[3] ;
 wire \i_spi.busy ;
 wire \i_spi.clock_count[0] ;
 wire \i_spi.clock_count[1] ;
 wire \i_spi.clock_count[2] ;
 wire \i_spi.clock_count[3] ;
 wire \i_spi.clock_divider[0] ;
 wire \i_spi.clock_divider[1] ;
 wire \i_spi.clock_divider[2] ;
 wire \i_spi.clock_divider[3] ;
 wire \i_spi.data[0] ;
 wire \i_spi.data[1] ;
 wire \i_spi.data[2] ;
 wire \i_spi.data[3] ;
 wire \i_spi.data[4] ;
 wire \i_spi.data[5] ;
 wire \i_spi.data[6] ;
 wire \i_spi.data[7] ;
 wire \i_spi.end_txn_reg ;
 wire \i_spi.read_latency ;
 wire \i_spi.spi_clk_out ;
 wire \i_spi.spi_dc ;
 wire \i_spi.spi_select ;
 wire \i_time.l_mtimecmp.data_out[0] ;
 wire \i_time.l_mtimecmp.data_out[10] ;
 wire \i_time.l_mtimecmp.data_out[11] ;
 wire \i_time.l_mtimecmp.data_out[12] ;
 wire \i_time.l_mtimecmp.data_out[13] ;
 wire \i_time.l_mtimecmp.data_out[14] ;
 wire \i_time.l_mtimecmp.data_out[15] ;
 wire \i_time.l_mtimecmp.data_out[16] ;
 wire \i_time.l_mtimecmp.data_out[17] ;
 wire \i_time.l_mtimecmp.data_out[18] ;
 wire \i_time.l_mtimecmp.data_out[19] ;
 wire \i_time.l_mtimecmp.data_out[1] ;
 wire \i_time.l_mtimecmp.data_out[20] ;
 wire \i_time.l_mtimecmp.data_out[21] ;
 wire \i_time.l_mtimecmp.data_out[22] ;
 wire \i_time.l_mtimecmp.data_out[23] ;
 wire \i_time.l_mtimecmp.data_out[24] ;
 wire \i_time.l_mtimecmp.data_out[25] ;
 wire \i_time.l_mtimecmp.data_out[26] ;
 wire \i_time.l_mtimecmp.data_out[27] ;
 wire \i_time.l_mtimecmp.data_out[28] ;
 wire \i_time.l_mtimecmp.data_out[29] ;
 wire \i_time.l_mtimecmp.data_out[2] ;
 wire \i_time.l_mtimecmp.data_out[30] ;
 wire \i_time.l_mtimecmp.data_out[31] ;
 wire \i_time.l_mtimecmp.data_out[3] ;
 wire \i_time.l_mtimecmp.data_out[4] ;
 wire \i_time.l_mtimecmp.data_out[5] ;
 wire \i_time.l_mtimecmp.data_out[6] ;
 wire \i_time.l_mtimecmp.data_out[7] ;
 wire \i_time.l_mtimecmp.data_out[8] ;
 wire \i_time.l_mtimecmp.data_out[9] ;
 wire \i_time.mtime[0] ;
 wire \i_time.mtime[10] ;
 wire \i_time.mtime[11] ;
 wire \i_time.mtime[12] ;
 wire \i_time.mtime[13] ;
 wire \i_time.mtime[14] ;
 wire \i_time.mtime[15] ;
 wire \i_time.mtime[16] ;
 wire \i_time.mtime[17] ;
 wire \i_time.mtime[18] ;
 wire \i_time.mtime[19] ;
 wire \i_time.mtime[1] ;
 wire \i_time.mtime[20] ;
 wire \i_time.mtime[21] ;
 wire \i_time.mtime[22] ;
 wire \i_time.mtime[23] ;
 wire \i_time.mtime[24] ;
 wire \i_time.mtime[25] ;
 wire \i_time.mtime[26] ;
 wire \i_time.mtime[27] ;
 wire \i_time.mtime[28] ;
 wire \i_time.mtime[29] ;
 wire \i_time.mtime[2] ;
 wire \i_time.mtime[30] ;
 wire \i_time.mtime[31] ;
 wire \i_time.mtime[3] ;
 wire \i_time.mtime[4] ;
 wire \i_time.mtime[5] ;
 wire \i_time.mtime[6] ;
 wire \i_time.mtime[7] ;
 wire \i_time.mtime[8] ;
 wire \i_time.mtime[9] ;
 wire \i_time.time_pulse ;
 wire \i_time.timer_interrupt ;
 wire \i_tinyqv.cpu.additional_mem_ops[0] ;
 wire \i_tinyqv.cpu.additional_mem_ops[1] ;
 wire \i_tinyqv.cpu.additional_mem_ops[2] ;
 wire \i_tinyqv.cpu.alu_op[0] ;
 wire \i_tinyqv.cpu.alu_op[1] ;
 wire \i_tinyqv.cpu.alu_op[2] ;
 wire \i_tinyqv.cpu.alu_op[3] ;
 wire \i_tinyqv.cpu.counter[2] ;
 wire \i_tinyqv.cpu.counter[3] ;
 wire \i_tinyqv.cpu.counter[4] ;
 wire \i_tinyqv.cpu.data_read_n[0] ;
 wire \i_tinyqv.cpu.data_read_n[1] ;
 wire \i_tinyqv.cpu.data_ready_latch ;
 wire \i_tinyqv.cpu.data_ready_sync ;
 wire \i_tinyqv.cpu.data_write_n[0] ;
 wire \i_tinyqv.cpu.data_write_n[1] ;
 wire \i_tinyqv.cpu.i_core.cmp ;
 wire \i_tinyqv.cpu.i_core.cmp_out ;
 wire \i_tinyqv.cpu.i_core.cy ;
 wire \i_tinyqv.cpu.i_core.cy_out ;
 wire \i_tinyqv.cpu.i_core.cycle[0] ;
 wire \i_tinyqv.cpu.i_core.cycle[1] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[0] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[1] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[2] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[3] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[4] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[5] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[6] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.cy ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.rstn ;
 wire \i_tinyqv.cpu.i_core.i_instrret.add ;
 wire \i_tinyqv.cpu.i_core.i_instrret.cy ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[0] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[1] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[2] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[3] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[0] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[10] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[11] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[12] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[13] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[14] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[15] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[16] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[17] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[18] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[19] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[1] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[20] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[21] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[22] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[23] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[24] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[25] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[26] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[27] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[28] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[29] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[2] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[30] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[31] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[4] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[5] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[6] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[7] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[8] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[9] ;
 wire \i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ;
 wire \i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[2] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[4] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[0] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[10] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[11] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[1] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[2] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[3] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[4] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[5] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[6] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[7] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[8] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[9] ;
 wire \i_tinyqv.cpu.i_core.interrupt_req[0] ;
 wire \i_tinyqv.cpu.i_core.interrupt_req[1] ;
 wire \i_tinyqv.cpu.i_core.is_double_fault_r ;
 wire \i_tinyqv.cpu.i_core.is_interrupt ;
 wire \i_tinyqv.cpu.i_core.last_interrupt_req[0] ;
 wire \i_tinyqv.cpu.i_core.last_interrupt_req[1] ;
 wire \i_tinyqv.cpu.i_core.load_done ;
 wire \i_tinyqv.cpu.i_core.load_top_bit ;
 wire \i_tinyqv.cpu.i_core.mcause[0] ;
 wire \i_tinyqv.cpu.i_core.mcause[1] ;
 wire \i_tinyqv.cpu.i_core.mcause[2] ;
 wire \i_tinyqv.cpu.i_core.mcause[3] ;
 wire \i_tinyqv.cpu.i_core.mcause[4] ;
 wire \i_tinyqv.cpu.i_core.mcause[5] ;
 wire \i_tinyqv.cpu.i_core.mem_op[0] ;
 wire \i_tinyqv.cpu.i_core.mem_op[1] ;
 wire \i_tinyqv.cpu.i_core.mem_op[2] ;
 wire \i_tinyqv.cpu.i_core.mepc[0] ;
 wire \i_tinyqv.cpu.i_core.mepc[10] ;
 wire \i_tinyqv.cpu.i_core.mepc[11] ;
 wire \i_tinyqv.cpu.i_core.mepc[12] ;
 wire \i_tinyqv.cpu.i_core.mepc[13] ;
 wire \i_tinyqv.cpu.i_core.mepc[14] ;
 wire \i_tinyqv.cpu.i_core.mepc[15] ;
 wire \i_tinyqv.cpu.i_core.mepc[16] ;
 wire \i_tinyqv.cpu.i_core.mepc[17] ;
 wire \i_tinyqv.cpu.i_core.mepc[18] ;
 wire \i_tinyqv.cpu.i_core.mepc[19] ;
 wire \i_tinyqv.cpu.i_core.mepc[1] ;
 wire \i_tinyqv.cpu.i_core.mepc[20] ;
 wire \i_tinyqv.cpu.i_core.mepc[21] ;
 wire \i_tinyqv.cpu.i_core.mepc[22] ;
 wire \i_tinyqv.cpu.i_core.mepc[23] ;
 wire \i_tinyqv.cpu.i_core.mepc[2] ;
 wire \i_tinyqv.cpu.i_core.mepc[3] ;
 wire \i_tinyqv.cpu.i_core.mepc[4] ;
 wire \i_tinyqv.cpu.i_core.mepc[5] ;
 wire \i_tinyqv.cpu.i_core.mepc[6] ;
 wire \i_tinyqv.cpu.i_core.mepc[7] ;
 wire \i_tinyqv.cpu.i_core.mepc[8] ;
 wire \i_tinyqv.cpu.i_core.mepc[9] ;
 wire \i_tinyqv.cpu.i_core.mie[0] ;
 wire \i_tinyqv.cpu.i_core.mie[1] ;
 wire \i_tinyqv.cpu.i_core.mie[2] ;
 wire \i_tinyqv.cpu.i_core.mie[3] ;
 wire \i_tinyqv.cpu.i_core.mie[4] ;
 wire \i_tinyqv.cpu.i_core.mip[0] ;
 wire \i_tinyqv.cpu.i_core.mip[1] ;
 wire \i_tinyqv.cpu.i_core.mstatus_mie ;
 wire \i_tinyqv.cpu.i_core.mstatus_mpie ;
 wire \i_tinyqv.cpu.i_core.mstatus_mte ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[0] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[10] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[11] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[12] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[13] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[14] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[15] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[1] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[2] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[3] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[4] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[5] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[6] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[7] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[8] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[9] ;
 wire \i_tinyqv.cpu.i_core.time_hi[0] ;
 wire \i_tinyqv.cpu.i_core.time_hi[1] ;
 wire \i_tinyqv.cpu.i_core.time_hi[2] ;
 wire \i_tinyqv.cpu.imm[12] ;
 wire \i_tinyqv.cpu.imm[13] ;
 wire \i_tinyqv.cpu.imm[14] ;
 wire \i_tinyqv.cpu.imm[15] ;
 wire \i_tinyqv.cpu.imm[16] ;
 wire \i_tinyqv.cpu.imm[17] ;
 wire \i_tinyqv.cpu.imm[18] ;
 wire \i_tinyqv.cpu.imm[19] ;
 wire \i_tinyqv.cpu.imm[20] ;
 wire \i_tinyqv.cpu.imm[21] ;
 wire \i_tinyqv.cpu.imm[22] ;
 wire \i_tinyqv.cpu.imm[23] ;
 wire \i_tinyqv.cpu.imm[24] ;
 wire \i_tinyqv.cpu.imm[25] ;
 wire \i_tinyqv.cpu.imm[26] ;
 wire \i_tinyqv.cpu.imm[27] ;
 wire \i_tinyqv.cpu.imm[28] ;
 wire \i_tinyqv.cpu.imm[29] ;
 wire \i_tinyqv.cpu.imm[30] ;
 wire \i_tinyqv.cpu.imm[31] ;
 wire \i_tinyqv.cpu.instr_data[0][0] ;
 wire \i_tinyqv.cpu.instr_data[0][10] ;
 wire \i_tinyqv.cpu.instr_data[0][11] ;
 wire \i_tinyqv.cpu.instr_data[0][12] ;
 wire \i_tinyqv.cpu.instr_data[0][13] ;
 wire \i_tinyqv.cpu.instr_data[0][14] ;
 wire \i_tinyqv.cpu.instr_data[0][15] ;
 wire \i_tinyqv.cpu.instr_data[0][1] ;
 wire \i_tinyqv.cpu.instr_data[0][2] ;
 wire \i_tinyqv.cpu.instr_data[0][3] ;
 wire \i_tinyqv.cpu.instr_data[0][4] ;
 wire \i_tinyqv.cpu.instr_data[0][5] ;
 wire \i_tinyqv.cpu.instr_data[0][6] ;
 wire \i_tinyqv.cpu.instr_data[0][7] ;
 wire \i_tinyqv.cpu.instr_data[0][8] ;
 wire \i_tinyqv.cpu.instr_data[0][9] ;
 wire \i_tinyqv.cpu.instr_data[1][0] ;
 wire \i_tinyqv.cpu.instr_data[1][10] ;
 wire \i_tinyqv.cpu.instr_data[1][11] ;
 wire \i_tinyqv.cpu.instr_data[1][12] ;
 wire \i_tinyqv.cpu.instr_data[1][13] ;
 wire \i_tinyqv.cpu.instr_data[1][14] ;
 wire \i_tinyqv.cpu.instr_data[1][15] ;
 wire \i_tinyqv.cpu.instr_data[1][1] ;
 wire \i_tinyqv.cpu.instr_data[1][2] ;
 wire \i_tinyqv.cpu.instr_data[1][3] ;
 wire \i_tinyqv.cpu.instr_data[1][4] ;
 wire \i_tinyqv.cpu.instr_data[1][5] ;
 wire \i_tinyqv.cpu.instr_data[1][6] ;
 wire \i_tinyqv.cpu.instr_data[1][7] ;
 wire \i_tinyqv.cpu.instr_data[1][8] ;
 wire \i_tinyqv.cpu.instr_data[1][9] ;
 wire \i_tinyqv.cpu.instr_data[2][0] ;
 wire \i_tinyqv.cpu.instr_data[2][10] ;
 wire \i_tinyqv.cpu.instr_data[2][11] ;
 wire \i_tinyqv.cpu.instr_data[2][12] ;
 wire \i_tinyqv.cpu.instr_data[2][13] ;
 wire \i_tinyqv.cpu.instr_data[2][14] ;
 wire \i_tinyqv.cpu.instr_data[2][15] ;
 wire \i_tinyqv.cpu.instr_data[2][1] ;
 wire \i_tinyqv.cpu.instr_data[2][2] ;
 wire \i_tinyqv.cpu.instr_data[2][3] ;
 wire \i_tinyqv.cpu.instr_data[2][4] ;
 wire \i_tinyqv.cpu.instr_data[2][5] ;
 wire \i_tinyqv.cpu.instr_data[2][6] ;
 wire \i_tinyqv.cpu.instr_data[2][7] ;
 wire \i_tinyqv.cpu.instr_data[2][8] ;
 wire \i_tinyqv.cpu.instr_data[2][9] ;
 wire \i_tinyqv.cpu.instr_data[3][0] ;
 wire \i_tinyqv.cpu.instr_data[3][10] ;
 wire \i_tinyqv.cpu.instr_data[3][11] ;
 wire \i_tinyqv.cpu.instr_data[3][12] ;
 wire \i_tinyqv.cpu.instr_data[3][13] ;
 wire \i_tinyqv.cpu.instr_data[3][14] ;
 wire \i_tinyqv.cpu.instr_data[3][15] ;
 wire \i_tinyqv.cpu.instr_data[3][1] ;
 wire \i_tinyqv.cpu.instr_data[3][2] ;
 wire \i_tinyqv.cpu.instr_data[3][3] ;
 wire \i_tinyqv.cpu.instr_data[3][4] ;
 wire \i_tinyqv.cpu.instr_data[3][5] ;
 wire \i_tinyqv.cpu.instr_data[3][6] ;
 wire \i_tinyqv.cpu.instr_data[3][7] ;
 wire \i_tinyqv.cpu.instr_data[3][8] ;
 wire \i_tinyqv.cpu.instr_data[3][9] ;
 wire \i_tinyqv.cpu.instr_data_in[0] ;
 wire \i_tinyqv.cpu.instr_data_in[10] ;
 wire \i_tinyqv.cpu.instr_data_in[11] ;
 wire \i_tinyqv.cpu.instr_data_in[12] ;
 wire \i_tinyqv.cpu.instr_data_in[13] ;
 wire \i_tinyqv.cpu.instr_data_in[14] ;
 wire \i_tinyqv.cpu.instr_data_in[15] ;
 wire \i_tinyqv.cpu.instr_data_in[1] ;
 wire \i_tinyqv.cpu.instr_data_in[2] ;
 wire \i_tinyqv.cpu.instr_data_in[3] ;
 wire \i_tinyqv.cpu.instr_data_in[4] ;
 wire \i_tinyqv.cpu.instr_data_in[5] ;
 wire \i_tinyqv.cpu.instr_data_in[6] ;
 wire \i_tinyqv.cpu.instr_data_in[7] ;
 wire \i_tinyqv.cpu.instr_data_in[8] ;
 wire \i_tinyqv.cpu.instr_data_in[9] ;
 wire \i_tinyqv.cpu.instr_data_start[10] ;
 wire \i_tinyqv.cpu.instr_data_start[11] ;
 wire \i_tinyqv.cpu.instr_data_start[12] ;
 wire \i_tinyqv.cpu.instr_data_start[13] ;
 wire \i_tinyqv.cpu.instr_data_start[14] ;
 wire \i_tinyqv.cpu.instr_data_start[15] ;
 wire \i_tinyqv.cpu.instr_data_start[16] ;
 wire \i_tinyqv.cpu.instr_data_start[17] ;
 wire \i_tinyqv.cpu.instr_data_start[18] ;
 wire \i_tinyqv.cpu.instr_data_start[19] ;
 wire \i_tinyqv.cpu.instr_data_start[20] ;
 wire \i_tinyqv.cpu.instr_data_start[21] ;
 wire \i_tinyqv.cpu.instr_data_start[22] ;
 wire \i_tinyqv.cpu.instr_data_start[23] ;
 wire \i_tinyqv.cpu.instr_data_start[3] ;
 wire \i_tinyqv.cpu.instr_data_start[4] ;
 wire \i_tinyqv.cpu.instr_data_start[5] ;
 wire \i_tinyqv.cpu.instr_data_start[6] ;
 wire \i_tinyqv.cpu.instr_data_start[7] ;
 wire \i_tinyqv.cpu.instr_data_start[8] ;
 wire \i_tinyqv.cpu.instr_data_start[9] ;
 wire \i_tinyqv.cpu.instr_fetch_running ;
 wire \i_tinyqv.cpu.instr_fetch_started ;
 wire \i_tinyqv.cpu.instr_fetch_stopped ;
 wire \i_tinyqv.cpu.instr_len[1] ;
 wire \i_tinyqv.cpu.instr_len[2] ;
 wire \i_tinyqv.cpu.instr_write_offset[1] ;
 wire \i_tinyqv.cpu.instr_write_offset[2] ;
 wire \i_tinyqv.cpu.instr_write_offset[3] ;
 wire \i_tinyqv.cpu.is_alu_imm ;
 wire \i_tinyqv.cpu.is_alu_reg ;
 wire \i_tinyqv.cpu.is_auipc ;
 wire \i_tinyqv.cpu.is_branch ;
 wire \i_tinyqv.cpu.is_jal ;
 wire \i_tinyqv.cpu.is_jalr ;
 wire \i_tinyqv.cpu.is_load ;
 wire \i_tinyqv.cpu.is_lui ;
 wire \i_tinyqv.cpu.is_store ;
 wire \i_tinyqv.cpu.is_system ;
 wire \i_tinyqv.cpu.load_started ;
 wire \i_tinyqv.cpu.mem_op_increment_reg ;
 wire \i_tinyqv.cpu.no_write_in_progress ;
 wire \i_tinyqv.cpu.pc[1] ;
 wire \i_tinyqv.cpu.pc[2] ;
 wire \i_tinyqv.cpu.was_early_branch ;
 wire \i_tinyqv.mem.data_from_read[16] ;
 wire \i_tinyqv.mem.data_from_read[17] ;
 wire \i_tinyqv.mem.data_from_read[18] ;
 wire \i_tinyqv.mem.data_from_read[19] ;
 wire \i_tinyqv.mem.data_from_read[20] ;
 wire \i_tinyqv.mem.data_from_read[21] ;
 wire \i_tinyqv.mem.data_from_read[22] ;
 wire \i_tinyqv.mem.data_from_read[23] ;
 wire \i_tinyqv.mem.data_stall ;
 wire \i_tinyqv.mem.instr_active ;
 wire \i_tinyqv.mem.q_ctrl.addr[0] ;
 wire \i_tinyqv.mem.q_ctrl.addr[10] ;
 wire \i_tinyqv.mem.q_ctrl.addr[11] ;
 wire \i_tinyqv.mem.q_ctrl.addr[12] ;
 wire \i_tinyqv.mem.q_ctrl.addr[13] ;
 wire \i_tinyqv.mem.q_ctrl.addr[14] ;
 wire \i_tinyqv.mem.q_ctrl.addr[15] ;
 wire \i_tinyqv.mem.q_ctrl.addr[16] ;
 wire \i_tinyqv.mem.q_ctrl.addr[17] ;
 wire \i_tinyqv.mem.q_ctrl.addr[18] ;
 wire \i_tinyqv.mem.q_ctrl.addr[19] ;
 wire \i_tinyqv.mem.q_ctrl.addr[1] ;
 wire \i_tinyqv.mem.q_ctrl.addr[20] ;
 wire \i_tinyqv.mem.q_ctrl.addr[21] ;
 wire \i_tinyqv.mem.q_ctrl.addr[22] ;
 wire \i_tinyqv.mem.q_ctrl.addr[23] ;
 wire \i_tinyqv.mem.q_ctrl.addr[2] ;
 wire \i_tinyqv.mem.q_ctrl.addr[3] ;
 wire \i_tinyqv.mem.q_ctrl.addr[4] ;
 wire \i_tinyqv.mem.q_ctrl.addr[5] ;
 wire \i_tinyqv.mem.q_ctrl.addr[6] ;
 wire \i_tinyqv.mem.q_ctrl.addr[7] ;
 wire \i_tinyqv.mem.q_ctrl.addr[8] ;
 wire \i_tinyqv.mem.q_ctrl.addr[9] ;
 wire \i_tinyqv.mem.q_ctrl.data_ready ;
 wire \i_tinyqv.mem.q_ctrl.data_req ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[0] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[1] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[2] ;
 wire \i_tinyqv.mem.q_ctrl.is_writing ;
 wire \i_tinyqv.mem.q_ctrl.last_ram_a_sel ;
 wire \i_tinyqv.mem.q_ctrl.last_ram_b_sel ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[0] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[1] ;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_neg ;
 wire net654;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_pos ;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_use_neg ;
 wire \i_tinyqv.mem.q_ctrl.spi_data_oe[0] ;
 wire net655;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ;
 wire net653;
 wire \i_tinyqv.mem.q_ctrl.spi_ram_b_select ;
 wire \i_tinyqv.mem.q_ctrl.stop_txn_reg ;
 wire \i_tinyqv.mem.qspi_data_buf[10] ;
 wire \i_tinyqv.mem.qspi_data_buf[11] ;
 wire \i_tinyqv.mem.qspi_data_buf[12] ;
 wire \i_tinyqv.mem.qspi_data_buf[13] ;
 wire \i_tinyqv.mem.qspi_data_buf[14] ;
 wire \i_tinyqv.mem.qspi_data_buf[15] ;
 wire \i_tinyqv.mem.qspi_data_buf[24] ;
 wire \i_tinyqv.mem.qspi_data_buf[25] ;
 wire \i_tinyqv.mem.qspi_data_buf[26] ;
 wire \i_tinyqv.mem.qspi_data_buf[27] ;
 wire \i_tinyqv.mem.qspi_data_buf[28] ;
 wire \i_tinyqv.mem.qspi_data_buf[29] ;
 wire \i_tinyqv.mem.qspi_data_buf[30] ;
 wire \i_tinyqv.mem.qspi_data_buf[31] ;
 wire \i_tinyqv.mem.qspi_data_buf[8] ;
 wire \i_tinyqv.mem.qspi_data_buf[9] ;
 wire \i_tinyqv.mem.qspi_data_byte_idx[0] ;
 wire \i_tinyqv.mem.qspi_data_byte_idx[1] ;
 wire \i_tinyqv.mem.qspi_write_done ;
 wire \i_uart_rx.bit_sample ;
 wire \i_uart_rx.cycle_counter[0] ;
 wire \i_uart_rx.cycle_counter[10] ;
 wire \i_uart_rx.cycle_counter[1] ;
 wire \i_uart_rx.cycle_counter[2] ;
 wire \i_uart_rx.cycle_counter[3] ;
 wire \i_uart_rx.cycle_counter[4] ;
 wire \i_uart_rx.cycle_counter[5] ;
 wire \i_uart_rx.cycle_counter[6] ;
 wire \i_uart_rx.cycle_counter[7] ;
 wire \i_uart_rx.cycle_counter[8] ;
 wire \i_uart_rx.cycle_counter[9] ;
 wire \i_uart_rx.fsm_state[0] ;
 wire \i_uart_rx.fsm_state[1] ;
 wire \i_uart_rx.fsm_state[2] ;
 wire \i_uart_rx.fsm_state[3] ;
 wire \i_uart_rx.recieved_data[0] ;
 wire \i_uart_rx.recieved_data[1] ;
 wire \i_uart_rx.recieved_data[2] ;
 wire \i_uart_rx.recieved_data[3] ;
 wire \i_uart_rx.recieved_data[4] ;
 wire \i_uart_rx.recieved_data[5] ;
 wire \i_uart_rx.recieved_data[6] ;
 wire \i_uart_rx.recieved_data[7] ;
 wire \i_uart_rx.rxd_reg[0] ;
 wire \i_uart_rx.rxd_reg[1] ;
 wire \i_uart_rx.uart_rts ;
 wire \i_uart_tx.cycle_counter[0] ;
 wire \i_uart_tx.cycle_counter[10] ;
 wire \i_uart_tx.cycle_counter[1] ;
 wire \i_uart_tx.cycle_counter[2] ;
 wire \i_uart_tx.cycle_counter[3] ;
 wire \i_uart_tx.cycle_counter[4] ;
 wire \i_uart_tx.cycle_counter[5] ;
 wire \i_uart_tx.cycle_counter[6] ;
 wire \i_uart_tx.cycle_counter[7] ;
 wire \i_uart_tx.cycle_counter[8] ;
 wire \i_uart_tx.cycle_counter[9] ;
 wire \i_uart_tx.data_to_send[0] ;
 wire \i_uart_tx.data_to_send[1] ;
 wire \i_uart_tx.data_to_send[2] ;
 wire \i_uart_tx.data_to_send[3] ;
 wire \i_uart_tx.data_to_send[4] ;
 wire \i_uart_tx.data_to_send[5] ;
 wire \i_uart_tx.data_to_send[6] ;
 wire \i_uart_tx.data_to_send[7] ;
 wire \i_uart_tx.fsm_state[0] ;
 wire \i_uart_tx.fsm_state[1] ;
 wire \i_uart_tx.fsm_state[2] ;
 wire \i_uart_tx.fsm_state[3] ;
 wire \i_uart_tx.txd_reg ;
 wire \mhz_clk_sync[0] ;
 wire \mhz_clk_sync[1] ;
 wire \mhz_clk_sync[2] ;
 wire net652;
 wire net651;
 wire net650;
 wire net649;
 wire net648;
 wire net647;
 wire net646;
 wire net645;
 wire net644;
 wire net643;
 wire net642;
 wire net641;
 wire net640;
 wire net639;
 wire net638;
 wire net637;
 wire net636;
 wire net635;
 wire net634;
 wire net633;
 wire net632;
 wire net631;
 wire net630;
 wire net629;
 wire net628;
 wire net627;
 wire net626;
 wire net625;
 wire net624;
 wire net623;
 wire net622;
 wire net621;
 wire net620;
 wire net619;
 wire net618;
 wire net617;
 wire net616;
 wire net615;
 wire net614;
 wire net613;
 wire net612;
 wire net611;
 wire net610;
 wire net609;
 wire net608;
 wire net607;
 wire net606;
 wire net605;
 wire net604;
 wire net603;
 wire net602;
 wire net601;
 wire net600;
 wire net599;
 wire net598;
 wire net597;
 wire net596;
 wire net595;
 wire net594;
 wire net593;
 wire net592;
 wire net591;
 wire net590;
 wire net589;
 wire net588;
 wire net587;
 wire net586;
 wire net585;
 wire net584;
 wire net583;
 wire net582;
 wire net581;
 wire net580;
 wire net579;
 wire net578;
 wire net577;
 wire net576;
 wire net575;
 wire net574;
 wire net573;
 wire net572;
 wire net571;
 wire net570;
 wire net569;
 wire net568;
 wire net567;
 wire net566;
 wire net565;
 wire net564;
 wire net563;
 wire net562;
 wire net561;
 wire net560;
 wire net559;
 wire net558;
 wire net557;
 wire net556;
 wire net555;
 wire net554;
 wire net553;
 wire net552;
 wire net551;
 wire net550;
 wire net549;
 wire net548;
 wire net547;
 wire net546;
 wire net545;
 wire net544;
 wire net543;
 wire net542;
 wire net541;
 wire net540;
 wire net539;
 wire net538;
 wire net537;
 wire net536;
 wire net535;
 wire net534;
 wire net533;
 wire net532;
 wire net531;
 wire net530;
 wire net529;
 wire net528;
 wire net527;
 wire net526;
 wire net525;
 wire net524;
 wire net523;
 wire net522;
 wire net521;
 wire net520;
 wire net519;
 wire net518;
 wire net517;
 wire net516;
 wire net515;
 wire net514;
 wire net513;
 wire net512;
 wire net511;
 wire net510;
 wire net509;
 wire net508;
 wire net507;
 wire net506;
 wire net505;
 wire net504;
 wire net503;
 wire net502;
 wire net501;
 wire net500;
 wire net499;
 wire net498;
 wire net497;
 wire net496;
 wire net495;
 wire net494;
 wire net493;
 wire net492;
 wire net491;
 wire net490;
 wire net489;
 wire net488;
 wire net487;
 wire net486;
 wire net485;
 wire net484;
 wire net483;
 wire net482;
 wire net481;
 wire net480;
 wire net479;
 wire net478;
 wire net477;
 wire net476;
 wire net475;
 wire net474;
 wire net473;
 wire net472;
 wire net471;
 wire net470;
 wire net469;
 wire net468;
 wire net467;
 wire net466;
 wire net465;
 wire net464;
 wire net463;
 wire net462;
 wire net461;
 wire net460;
 wire net459;
 wire net458;
 wire net457;
 wire net456;
 wire net455;
 wire net454;
 wire net453;
 wire net452;
 wire net451;
 wire net450;
 wire net449;
 wire net448;
 wire net447;
 wire net446;
 wire net445;
 wire net444;
 wire net443;
 wire net442;
 wire net441;
 wire net440;
 wire net439;
 wire net438;
 wire net437;
 wire net436;
 wire net435;
 wire net434;
 wire net433;
 wire net432;
 wire net431;
 wire net430;
 wire net429;
 wire net428;
 wire net427;
 wire net426;
 wire net425;
 wire net424;
 wire net423;
 wire net422;
 wire net421;
 wire net420;
 wire net419;
 wire net418;
 wire net417;
 wire net416;
 wire net415;
 wire net414;
 wire net413;
 wire net412;
 wire net411;
 wire net410;
 wire net409;
 wire net408;
 wire net407;
 wire net406;
 wire net405;
 wire net404;
 wire net403;
 wire net402;
 wire net401;
 wire net400;
 wire net399;
 wire net398;
 wire net397;
 wire net396;
 wire net395;
 wire net394;
 wire net393;
 wire net392;
 wire net391;
 wire net390;
 wire net389;
 wire net388;
 wire net387;
 wire net386;
 wire net385;
 wire net384;
 wire net383;
 wire net382;
 wire net381;
 wire net380;
 wire net379;
 wire net378;
 wire net377;
 wire net376;
 wire net375;
 wire net374;
 wire net373;
 wire net372;
 wire net371;
 wire net370;
 wire net369;
 wire net368;
 wire net367;
 wire net366;
 wire net365;
 wire net364;
 wire net363;
 wire net362;
 wire net361;
 wire net360;
 wire net359;
 wire net358;
 wire net357;
 wire net356;
 wire net355;
 wire net354;
 wire net353;
 wire net352;
 wire net351;
 wire net350;
 wire net349;
 wire net348;
 wire net347;
 wire net346;
 wire net345;
 wire net344;
 wire net343;
 wire net342;
 wire net341;
 wire net340;
 wire net339;
 wire net338;
 wire net337;
 wire net336;
 wire net335;
 wire net334;
 wire net333;
 wire net332;
 wire net331;
 wire net330;
 wire net329;
 wire net328;
 wire net327;
 wire net326;
 wire net325;
 wire net324;
 wire net323;
 wire net322;
 wire net321;
 wire net320;
 wire net319;
 wire net318;
 wire net317;
 wire net316;
 wire net315;
 wire net314;
 wire net313;
 wire net312;
 wire net311;
 wire net310;
 wire net309;
 wire net308;
 wire net307;
 wire net306;
 wire net305;
 wire net304;
 wire net303;
 wire net302;
 wire net301;
 wire net300;
 wire net299;
 wire net298;
 wire net297;
 wire net296;
 wire net295;
 wire net294;
 wire net293;
 wire net292;
 wire net291;
 wire net290;
 wire net289;
 wire net288;
 wire net287;
 wire net286;
 wire net285;
 wire net284;
 wire net283;
 wire net282;
 wire net281;
 wire net280;
 wire net279;
 wire net278;
 wire net277;
 wire net276;
 wire net275;
 wire net274;
 wire net273;
 wire net272;
 wire net271;
 wire net270;
 wire net269;
 wire net268;
 wire net267;
 wire net266;
 wire net265;
 wire net264;
 wire net263;
 wire net262;
 wire net261;
 wire net260;
 wire net259;
 wire net258;
 wire net257;
 wire net256;
 wire net255;
 wire net254;
 wire net253;
 wire net252;
 wire net251;
 wire net250;
 wire net249;
 wire net248;
 wire net247;
 wire net246;
 wire net245;
 wire net244;
 wire net243;
 wire net242;
 wire net241;
 wire net240;
 wire net239;
 wire net238;
 wire net237;
 wire net236;
 wire net235;
 wire net234;
 wire net233;
 wire net232;
 wire net231;
 wire net230;
 wire net229;
 wire net228;
 wire net227;
 wire net226;
 wire net225;
 wire net224;
 wire net223;
 wire net222;
 wire net221;
 wire net220;
 wire net219;
 wire net218;
 wire net217;
 wire net216;
 wire net215;
 wire net214;
 wire net213;
 wire net212;
 wire net211;
 wire net210;
 wire net209;
 wire net208;
 wire net207;
 wire net206;
 wire net205;
 wire net204;
 wire net203;
 wire net202;
 wire net201;
 wire net200;
 wire net199;
 wire net198;
 wire net197;
 wire net196;
 wire net195;
 wire net194;
 wire net193;
 wire net192;
 wire net191;
 wire net190;
 wire net189;
 wire net188;
 wire net187;
 wire net186;
 wire net185;
 wire net184;
 wire net183;
 wire net182;
 wire net181;
 wire net180;
 wire net179;
 wire net178;
 wire net177;
 wire net176;
 wire net175;
 wire net174;
 wire net173;
 wire net172;
 wire net171;
 wire net170;
 wire net169;
 wire net168;
 wire net167;
 wire net166;
 wire net165;
 wire net164;
 wire net163;
 wire net162;
 wire net161;
 wire net160;
 wire net159;
 wire net158;
 wire net157;
 wire net156;
 wire net155;
 wire net154;
 wire net153;
 wire net152;
 wire net151;
 wire net150;
 wire net149;
 wire net148;
 wire net147;
 wire net146;
 wire net145;
 wire net144;
 wire net143;
 wire net142;
 wire net141;
 wire net140;
 wire net139;
 wire net138;
 wire net137;
 wire net136;
 wire net135;
 wire net134;
 wire net133;
 wire net132;
 wire net131;
 wire net130;
 wire net129;
 wire net128;
 wire net127;
 wire net126;
 wire net125;
 wire net124;
 wire net123;
 wire net122;
 wire net121;
 wire net120;
 wire net119;
 wire net118;
 wire net117;
 wire net116;
 wire net115;
 wire net114;
 wire net113;
 wire net112;
 wire net111;
 wire net110;
 wire net109;
 wire net108;
 wire net107;
 wire net106;
 wire net105;
 wire net104;
 wire net103;
 wire net102;
 wire net101;
 wire net100;
 wire net99;
 wire net98;
 wire net97;
 wire net96;
 wire net95;
 wire net94;
 wire net93;
 wire net92;
 wire net91;
 wire net90;
 wire net89;
 wire net88;
 wire net87;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net72;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire net67;
 wire net66;
 wire net65;
 wire net64;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire net51;
 wire net50;
 wire net49;
 wire net48;
 wire net47;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_leaf_36_clk_regs;
 wire clknet_leaf_37_clk_regs;
 wire clknet_leaf_38_clk_regs;
 wire clknet_leaf_39_clk_regs;
 wire clknet_leaf_40_clk_regs;
 wire clknet_leaf_41_clk_regs;
 wire clknet_leaf_42_clk_regs;
 wire clknet_leaf_43_clk_regs;
 wire clknet_leaf_44_clk_regs;
 wire clknet_leaf_45_clk_regs;
 wire clknet_leaf_46_clk_regs;
 wire clknet_leaf_47_clk_regs;
 wire clknet_leaf_48_clk_regs;
 wire clknet_leaf_49_clk_regs;
 wire clknet_leaf_50_clk_regs;
 wire clknet_leaf_51_clk_regs;
 wire clknet_leaf_52_clk_regs;
 wire clknet_leaf_53_clk_regs;
 wire clknet_leaf_54_clk_regs;
 wire clknet_leaf_55_clk_regs;
 wire clknet_leaf_56_clk_regs;
 wire clknet_leaf_58_clk_regs;
 wire clknet_leaf_59_clk_regs;
 wire clknet_leaf_60_clk_regs;
 wire clknet_leaf_61_clk_regs;
 wire clknet_leaf_62_clk_regs;
 wire clknet_leaf_63_clk_regs;
 wire clknet_leaf_64_clk_regs;
 wire clknet_leaf_65_clk_regs;
 wire clknet_leaf_66_clk_regs;
 wire clknet_leaf_67_clk_regs;
 wire clknet_leaf_68_clk_regs;
 wire clknet_leaf_69_clk_regs;
 wire clknet_leaf_70_clk_regs;
 wire clknet_leaf_71_clk_regs;
 wire clknet_leaf_72_clk_regs;
 wire clknet_leaf_73_clk_regs;
 wire clknet_leaf_74_clk_regs;
 wire clknet_leaf_75_clk_regs;
 wire clknet_leaf_76_clk_regs;
 wire clknet_leaf_77_clk_regs;
 wire clknet_leaf_78_clk_regs;
 wire clknet_leaf_79_clk_regs;
 wire clknet_leaf_80_clk_regs;
 wire clknet_leaf_81_clk_regs;
 wire clknet_leaf_82_clk_regs;
 wire clknet_leaf_83_clk_regs;
 wire clknet_leaf_84_clk_regs;
 wire clknet_leaf_85_clk_regs;
 wire clknet_leaf_86_clk_regs;
 wire clknet_leaf_87_clk_regs;
 wire clknet_leaf_88_clk_regs;
 wire clknet_leaf_89_clk_regs;
 wire clknet_leaf_90_clk_regs;
 wire clknet_leaf_91_clk_regs;
 wire clknet_leaf_92_clk_regs;
 wire clknet_leaf_93_clk_regs;
 wire clknet_leaf_94_clk_regs;
 wire clknet_leaf_95_clk_regs;
 wire clknet_leaf_96_clk_regs;
 wire clknet_leaf_97_clk_regs;
 wire clknet_leaf_98_clk_regs;
 wire clknet_leaf_99_clk_regs;
 wire clknet_leaf_100_clk_regs;
 wire clknet_leaf_101_clk_regs;
 wire clknet_leaf_102_clk_regs;
 wire clknet_leaf_103_clk_regs;
 wire clknet_leaf_104_clk_regs;
 wire clknet_leaf_105_clk_regs;
 wire clknet_leaf_106_clk_regs;
 wire clknet_leaf_107_clk_regs;
 wire clknet_leaf_108_clk_regs;
 wire clknet_leaf_109_clk_regs;
 wire clknet_leaf_110_clk_regs;
 wire clknet_leaf_111_clk_regs;
 wire clknet_leaf_112_clk_regs;
 wire clknet_leaf_113_clk_regs;
 wire clknet_leaf_114_clk_regs;
 wire clknet_leaf_115_clk_regs;
 wire clknet_leaf_116_clk_regs;
 wire clknet_leaf_117_clk_regs;
 wire clknet_leaf_118_clk_regs;
 wire clknet_leaf_119_clk_regs;
 wire clknet_leaf_120_clk_regs;
 wire clknet_leaf_121_clk_regs;
 wire clknet_leaf_122_clk_regs;
 wire clknet_leaf_123_clk_regs;
 wire clknet_leaf_124_clk_regs;
 wire clknet_leaf_125_clk_regs;
 wire clknet_leaf_126_clk_regs;
 wire clknet_leaf_127_clk_regs;
 wire clknet_leaf_128_clk_regs;
 wire clknet_leaf_129_clk_regs;
 wire clknet_leaf_130_clk_regs;
 wire clknet_leaf_131_clk_regs;
 wire clknet_leaf_132_clk_regs;
 wire clknet_leaf_133_clk_regs;
 wire clknet_leaf_134_clk_regs;
 wire clknet_leaf_135_clk_regs;
 wire clknet_leaf_136_clk_regs;
 wire clknet_leaf_137_clk_regs;
 wire clknet_leaf_138_clk_regs;
 wire clknet_leaf_139_clk_regs;
 wire clknet_leaf_140_clk_regs;
 wire clknet_leaf_141_clk_regs;
 wire clknet_leaf_142_clk_regs;
 wire clknet_leaf_143_clk_regs;
 wire clknet_leaf_144_clk_regs;
 wire clknet_leaf_145_clk_regs;
 wire clknet_leaf_146_clk_regs;
 wire clknet_leaf_147_clk_regs;
 wire clknet_leaf_148_clk_regs;
 wire clknet_leaf_149_clk_regs;
 wire clknet_leaf_150_clk_regs;
 wire clknet_leaf_151_clk_regs;
 wire clknet_leaf_152_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;

 sg13g2_inv_2 _08710_ (.Y(_01487_),
    .A(net568));
 sg13g2_inv_1 _08711_ (.Y(_01488_),
    .A(net3444));
 sg13g2_inv_1 _08712_ (.Y(_01489_),
    .A(net3590));
 sg13g2_inv_1 _08713_ (.Y(_01490_),
    .A(net3678));
 sg13g2_inv_1 _08714_ (.Y(_01491_),
    .A(\i_tinyqv.cpu.is_branch ));
 sg13g2_inv_1 _08715_ (.Y(_01492_),
    .A(net3932));
 sg13g2_inv_1 _08716_ (.Y(_01493_),
    .A(\i_tinyqv.cpu.is_load ));
 sg13g2_inv_1 _08717_ (.Y(_01494_),
    .A(net3178));
 sg13g2_inv_1 _08718_ (.Y(_01495_),
    .A(\i_tinyqv.cpu.data_write_n[1] ));
 sg13g2_inv_1 _08719_ (.Y(_01496_),
    .A(net3771));
 sg13g2_inv_1 _08720_ (.Y(_01497_),
    .A(net3920));
 sg13g2_inv_1 _08721_ (.Y(_01498_),
    .A(net3909));
 sg13g2_inv_1 _08722_ (.Y(_01499_),
    .A(net3842));
 sg13g2_inv_1 _08723_ (.Y(_01500_),
    .A(net3873));
 sg13g2_inv_1 _08724_ (.Y(_01501_),
    .A(net3882));
 sg13g2_inv_1 _08725_ (.Y(_01502_),
    .A(net3835));
 sg13g2_inv_1 _08726_ (.Y(_01503_),
    .A(net3800));
 sg13g2_inv_1 _08727_ (.Y(_01504_),
    .A(\data_to_write[7] ));
 sg13g2_inv_1 _08728_ (.Y(_01505_),
    .A(net597));
 sg13g2_inv_1 _08729_ (.Y(_01506_),
    .A(net598));
 sg13g2_inv_1 _08730_ (.Y(_01507_),
    .A(net599));
 sg13g2_inv_4 _08731_ (.A(\data_to_write[3] ),
    .Y(_01508_));
 sg13g2_inv_2 _08732_ (.Y(_01509_),
    .A(net600));
 sg13g2_inv_2 _08733_ (.Y(_01510_),
    .A(net601));
 sg13g2_inv_4 _08734_ (.A(\data_to_write[0] ),
    .Y(_01511_));
 sg13g2_inv_1 _08735_ (.Y(_01512_),
    .A(net607));
 sg13g2_inv_2 _08736_ (.Y(_01513_),
    .A(\i_tinyqv.cpu.instr_data_start[18] ));
 sg13g2_inv_1 _08737_ (.Y(_01514_),
    .A(net3927));
 sg13g2_inv_1 _08738_ (.Y(_01515_),
    .A(net3938));
 sg13g2_inv_1 _08739_ (.Y(_01516_),
    .A(net4121));
 sg13g2_inv_1 _08740_ (.Y(_01517_),
    .A(net4110));
 sg13g2_inv_2 _08741_ (.Y(_01518_),
    .A(net4058));
 sg13g2_inv_1 _08742_ (.Y(_01519_),
    .A(\i_tinyqv.cpu.instr_data_start[5] ));
 sg13g2_inv_1 _08743_ (.Y(_01520_),
    .A(net615));
 sg13g2_inv_2 _08744_ (.Y(_01521_),
    .A(net4054));
 sg13g2_inv_1 _08745_ (.Y(_01522_),
    .A(net618));
 sg13g2_inv_2 _08746_ (.Y(_01523_),
    .A(net3799));
 sg13g2_inv_1 _08747_ (.Y(_01524_),
    .A(\i_tinyqv.mem.instr_active ));
 sg13g2_inv_1 _08748_ (.Y(_01525_),
    .A(net635));
 sg13g2_inv_1 _08749_ (.Y(_01526_),
    .A(net3763));
 sg13g2_inv_1 _08750_ (.Y(_01527_),
    .A(net538));
 sg13g2_inv_1 _08751_ (.Y(_00340_),
    .A(net2745));
 sg13g2_inv_1 _08752_ (.Y(_00339_),
    .A(net2678));
 sg13g2_inv_1 _08753_ (.Y(_00338_),
    .A(net2771));
 sg13g2_inv_1 _08754_ (.Y(_00337_),
    .A(net2780));
 sg13g2_inv_1 _08755_ (.Y(_00336_),
    .A(net2803));
 sg13g2_inv_1 _08756_ (.Y(_00335_),
    .A(net2775));
 sg13g2_inv_1 _08757_ (.Y(_00334_),
    .A(net2717));
 sg13g2_inv_1 _08758_ (.Y(_00333_),
    .A(net2527));
 sg13g2_inv_1 _08759_ (.Y(_00332_),
    .A(net2628));
 sg13g2_inv_1 _08760_ (.Y(_00331_),
    .A(net2720));
 sg13g2_inv_1 _08761_ (.Y(_00330_),
    .A(net2789));
 sg13g2_inv_1 _08762_ (.Y(_00329_),
    .A(net2801));
 sg13g2_inv_1 _08763_ (.Y(_00328_),
    .A(net2749));
 sg13g2_inv_1 _08764_ (.Y(_00327_),
    .A(net2772));
 sg13g2_inv_1 _08765_ (.Y(_00326_),
    .A(net2705));
 sg13g2_inv_1 _08766_ (.Y(_00325_),
    .A(net2735));
 sg13g2_inv_1 _08767_ (.Y(_00324_),
    .A(net2804));
 sg13g2_inv_1 _08768_ (.Y(_00323_),
    .A(net2790));
 sg13g2_inv_1 _08769_ (.Y(_00322_),
    .A(net2642));
 sg13g2_inv_1 _08770_ (.Y(_00321_),
    .A(net2787));
 sg13g2_inv_1 _08771_ (.Y(_00320_),
    .A(net2619));
 sg13g2_inv_1 _08772_ (.Y(_00319_),
    .A(net2755));
 sg13g2_inv_1 _08773_ (.Y(_00318_),
    .A(net2548));
 sg13g2_inv_1 _08774_ (.Y(_00317_),
    .A(net8));
 sg13g2_inv_1 _08775_ (.Y(_01528_),
    .A(net3928));
 sg13g2_inv_1 _08776_ (.Y(_01529_),
    .A(net3959));
 sg13g2_inv_1 _08777_ (.Y(_01530_),
    .A(\i_time.mtime[26] ));
 sg13g2_inv_1 _08778_ (.Y(_01531_),
    .A(\i_time.mtime[25] ));
 sg13g2_inv_1 _08779_ (.Y(_01532_),
    .A(net4029));
 sg13g2_inv_1 _08780_ (.Y(_01533_),
    .A(net4067));
 sg13g2_inv_1 _08781_ (.Y(_01534_),
    .A(\i_time.mtime[20] ));
 sg13g2_inv_1 _08782_ (.Y(_01535_),
    .A(net4049));
 sg13g2_inv_1 _08783_ (.Y(_01536_),
    .A(\i_time.mtime[16] ));
 sg13g2_inv_1 _08784_ (.Y(_01537_),
    .A(net4012));
 sg13g2_inv_1 _08785_ (.Y(_01538_),
    .A(\i_time.mtime[13] ));
 sg13g2_inv_1 _08786_ (.Y(_01539_),
    .A(net3943));
 sg13g2_inv_1 _08787_ (.Y(_01540_),
    .A(\i_time.mtime[10] ));
 sg13g2_inv_1 _08788_ (.Y(_01541_),
    .A(net4107));
 sg13g2_inv_1 _08789_ (.Y(_01542_),
    .A(net4114));
 sg13g2_inv_1 _08790_ (.Y(_01543_),
    .A(net4115));
 sg13g2_inv_1 _08791_ (.Y(_01544_),
    .A(\i_time.mtime[4] ));
 sg13g2_inv_1 _08792_ (.Y(_01545_),
    .A(\i_time.mtime[3] ));
 sg13g2_inv_1 _08793_ (.Y(_01546_),
    .A(net4119));
 sg13g2_inv_1 _08794_ (.Y(_01547_),
    .A(\i_time.mtime[1] ));
 sg13g2_inv_1 _08795_ (.Y(_01548_),
    .A(\i_time.mtime[0] ));
 sg13g2_inv_1 _08796_ (.Y(_01549_),
    .A(net3188));
 sg13g2_inv_1 _08797_ (.Y(_01550_),
    .A(net3265));
 sg13g2_inv_1 _08798_ (.Y(_01551_),
    .A(net3246));
 sg13g2_inv_1 _08799_ (.Y(_01552_),
    .A(net3327));
 sg13g2_inv_1 _08800_ (.Y(_01553_),
    .A(net3186));
 sg13g2_inv_1 _08801_ (.Y(_01554_),
    .A(\i_spi.spi_clk_out ));
 sg13g2_inv_1 _08802_ (.Y(_01555_),
    .A(\i_spi.bits_remaining[3] ));
 sg13g2_inv_1 _08803_ (.Y(_01556_),
    .A(net3723));
 sg13g2_inv_1 _08804_ (.Y(_01557_),
    .A(net3365));
 sg13g2_inv_1 _08805_ (.Y(_01558_),
    .A(\i_debug_uart_tx.data_to_send[6] ));
 sg13g2_inv_1 _08806_ (.Y(_01559_),
    .A(net3402));
 sg13g2_inv_1 _08807_ (.Y(_01560_),
    .A(net3432));
 sg13g2_inv_1 _08808_ (.Y(_01561_),
    .A(\i_debug_uart_tx.data_to_send[3] ));
 sg13g2_inv_1 _08809_ (.Y(_01562_),
    .A(net3446));
 sg13g2_inv_1 _08810_ (.Y(_01563_),
    .A(\i_debug_uart_tx.data_to_send[1] ));
 sg13g2_inv_1 _08811_ (.Y(_01564_),
    .A(net3642));
 sg13g2_inv_1 _08812_ (.Y(_01565_),
    .A(net3317));
 sg13g2_inv_1 _08813_ (.Y(_01566_),
    .A(\i_uart_tx.fsm_state[3] ));
 sg13g2_inv_1 _08814_ (.Y(_01567_),
    .A(net3983));
 sg13g2_inv_1 _08815_ (.Y(_01568_),
    .A(net4135));
 sg13g2_inv_1 _08816_ (.Y(_01569_),
    .A(\i_uart_tx.data_to_send[7] ));
 sg13g2_inv_1 _08817_ (.Y(_01570_),
    .A(net3452));
 sg13g2_inv_1 _08818_ (.Y(_01571_),
    .A(\i_uart_tx.data_to_send[5] ));
 sg13g2_inv_1 _08819_ (.Y(_01572_),
    .A(net3428));
 sg13g2_inv_1 _08820_ (.Y(_01573_),
    .A(net3472));
 sg13g2_inv_1 _08821_ (.Y(_01574_),
    .A(net3494));
 sg13g2_inv_1 _08822_ (.Y(_01575_),
    .A(\i_uart_tx.data_to_send[1] ));
 sg13g2_inv_1 _08823_ (.Y(_01576_),
    .A(net3525));
 sg13g2_inv_2 _08824_ (.Y(_01577_),
    .A(net656));
 sg13g2_inv_1 _08825_ (.Y(_01578_),
    .A(net3423));
 sg13g2_inv_1 _08826_ (.Y(_01579_),
    .A(net2831));
 sg13g2_inv_1 _08827_ (.Y(_01580_),
    .A(net584));
 sg13g2_inv_2 _08828_ (.Y(_01581_),
    .A(net588));
 sg13g2_inv_4 _08829_ (.A(net596),
    .Y(_01582_));
 sg13g2_inv_1 _08830_ (.Y(_01583_),
    .A(net4117));
 sg13g2_inv_1 _08831_ (.Y(_01584_),
    .A(net4103));
 sg13g2_inv_1 _08832_ (.Y(_01585_),
    .A(net3970));
 sg13g2_inv_1 _08833_ (.Y(_01586_),
    .A(net4002));
 sg13g2_inv_1 _08834_ (.Y(_01587_),
    .A(net3314));
 sg13g2_inv_1 _08835_ (.Y(_01588_),
    .A(net4010));
 sg13g2_inv_1 _08836_ (.Y(_01589_),
    .A(net4086));
 sg13g2_inv_1 _08837_ (.Y(_01590_),
    .A(net3963));
 sg13g2_inv_1 _08838_ (.Y(_01591_),
    .A(net3588));
 sg13g2_inv_1 _08839_ (.Y(_01592_),
    .A(net3939));
 sg13g2_inv_1 _08840_ (.Y(_01593_),
    .A(net3185));
 sg13g2_inv_1 _08841_ (.Y(_01594_),
    .A(net3192));
 sg13g2_inv_2 _08842_ (.Y(_01595_),
    .A(net581));
 sg13g2_inv_1 _08843_ (.Y(_01596_),
    .A(_00122_));
 sg13g2_inv_1 _08844_ (.Y(_01597_),
    .A(\i_tinyqv.cpu.instr_write_offset[2] ));
 sg13g2_inv_1 _08845_ (.Y(_01598_),
    .A(\i_tinyqv.cpu.instr_write_offset[1] ));
 sg13g2_inv_1 _08846_ (.Y(_01599_),
    .A(\i_pwm.pwm_count[0] ));
 sg13g2_inv_1 _08847_ (.Y(_01600_),
    .A(net3386));
 sg13g2_inv_1 _08848_ (.Y(_01601_),
    .A(net3199));
 sg13g2_inv_1 _08849_ (.Y(_01602_),
    .A(net3377));
 sg13g2_inv_1 _08850_ (.Y(_01603_),
    .A(_00184_));
 sg13g2_inv_2 _08851_ (.Y(_01604_),
    .A(_00133_));
 sg13g2_inv_1 _08852_ (.Y(_01605_),
    .A(\i_uart_rx.cycle_counter[0] ));
 sg13g2_inv_1 _08853_ (.Y(_01606_),
    .A(\i_uart_rx.cycle_counter[2] ));
 sg13g2_inv_1 _08854_ (.Y(_01607_),
    .A(\i_uart_rx.cycle_counter[9] ));
 sg13g2_inv_1 _08855_ (.Y(_01608_),
    .A(\i_uart_rx.cycle_counter[8] ));
 sg13g2_inv_1 _08856_ (.Y(_01609_),
    .A(_00196_));
 sg13g2_inv_1 _08857_ (.Y(_01610_),
    .A(net3349));
 sg13g2_inv_1 _08858_ (.Y(_01611_),
    .A(\i_tinyqv.cpu.instr_fetch_started ));
 sg13g2_inv_1 _08859_ (.Y(_01612_),
    .A(\addr[9] ));
 sg13g2_inv_1 _08860_ (.Y(_01613_),
    .A(net3626));
 sg13g2_inv_1 _08861_ (.Y(_01614_),
    .A(net3548));
 sg13g2_inv_1 _08862_ (.Y(_01615_),
    .A(net3664));
 sg13g2_inv_4 _08863_ (.A(\addr[4] ),
    .Y(_01616_));
 sg13g2_inv_1 _08864_ (.Y(_01617_),
    .A(net4060));
 sg13g2_inv_1 _08865_ (.Y(_01618_),
    .A(\i_pwm.pwm_count[1] ));
 sg13g2_inv_1 _08866_ (.Y(_01619_),
    .A(\i_pwm.pwm_count[3] ));
 sg13g2_inv_1 _08867_ (.Y(_01620_),
    .A(\i_pwm.pwm_count[6] ));
 sg13g2_inv_1 _08868_ (.Y(_01621_),
    .A(net4099));
 sg13g2_inv_1 _08869_ (.Y(_01622_),
    .A(\i_latch_mem.data_ready ));
 sg13g2_inv_1 _08870_ (.Y(_01623_),
    .A(net3656));
 sg13g2_inv_1 _08871_ (.Y(_01624_),
    .A(net3592));
 sg13g2_inv_1 _08872_ (.Y(_01625_),
    .A(net3725));
 sg13g2_inv_1 _08873_ (.Y(_01626_),
    .A(net3701));
 sg13g2_inv_1 _08874_ (.Y(_01627_),
    .A(net3721));
 sg13g2_inv_1 _08875_ (.Y(_01628_),
    .A(net3630));
 sg13g2_inv_1 _08876_ (.Y(_01629_),
    .A(net3636));
 sg13g2_inv_1 _08877_ (.Y(_01630_),
    .A(net3757));
 sg13g2_inv_1 _08878_ (.Y(_01631_),
    .A(net3571));
 sg13g2_inv_1 _08879_ (.Y(_01632_),
    .A(net3647));
 sg13g2_inv_1 _08880_ (.Y(_01633_),
    .A(net3660));
 sg13g2_inv_1 _08881_ (.Y(_01634_),
    .A(net3695));
 sg13g2_inv_1 _08882_ (.Y(_01635_),
    .A(net3544));
 sg13g2_inv_1 _08883_ (.Y(_01636_),
    .A(net3814));
 sg13g2_inv_1 _08884_ (.Y(_01637_),
    .A(net3728));
 sg13g2_inv_1 _08885_ (.Y(_01638_),
    .A(net3834));
 sg13g2_inv_1 _08886_ (.Y(_01639_),
    .A(\i_time.l_mtimecmp.data_out[11] ));
 sg13g2_inv_1 _08887_ (.Y(_01640_),
    .A(\i_time.l_mtimecmp.data_out[9] ));
 sg13g2_inv_1 _08888_ (.Y(_01641_),
    .A(net3662));
 sg13g2_inv_1 _08889_ (.Y(_01642_),
    .A(net3674));
 sg13g2_inv_1 _08890_ (.Y(_01643_),
    .A(net3483));
 sg13g2_inv_1 _08891_ (.Y(_01644_),
    .A(net3568));
 sg13g2_inv_1 _08892_ (.Y(_01645_),
    .A(net3618));
 sg13g2_inv_1 _08893_ (.Y(_01646_),
    .A(net3473));
 sg13g2_inv_1 _08894_ (.Y(_01647_),
    .A(net3989));
 sg13g2_inv_1 _08895_ (.Y(_01648_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[4] ));
 sg13g2_inv_1 _08896_ (.Y(_01649_),
    .A(_00206_));
 sg13g2_inv_1 _08897_ (.Y(_01650_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[5] ));
 sg13g2_inv_1 _08898_ (.Y(_01651_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[6] ));
 sg13g2_inv_1 _08899_ (.Y(_01652_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[7] ));
 sg13g2_inv_1 _08900_ (.Y(_01653_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[9] ));
 sg13g2_inv_1 _08901_ (.Y(_01654_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[11] ));
 sg13g2_inv_1 _08902_ (.Y(_01655_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[12] ));
 sg13g2_inv_1 _08903_ (.Y(_01656_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[13] ));
 sg13g2_inv_1 _08904_ (.Y(_01657_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[14] ));
 sg13g2_inv_1 _08905_ (.Y(_01658_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[14] ));
 sg13g2_inv_1 _08906_ (.Y(_01659_),
    .A(\i_tinyqv.cpu.i_core.mepc[0] ));
 sg13g2_inv_1 _08907_ (.Y(_01660_),
    .A(net3914));
 sg13g2_inv_1 _08908_ (.Y(_01661_),
    .A(\i_tinyqv.cpu.instr_data_in[8] ));
 sg13g2_inv_4 _08909_ (.A(net3788),
    .Y(_01662_));
 sg13g2_inv_1 _08910_ (.Y(_01663_),
    .A(\i_latch_mem.data_out[12] ));
 sg13g2_inv_1 _08911_ (.Y(_01664_),
    .A(\i_tinyqv.mem.data_from_read[16] ));
 sg13g2_inv_1 _08912_ (.Y(_01665_),
    .A(\i_tinyqv.mem.data_from_read[20] ));
 sg13g2_inv_1 _08913_ (.Y(_01666_),
    .A(\i_latch_mem.data_out[24] ));
 sg13g2_inv_1 _08914_ (.Y(_01667_),
    .A(net621));
 sg13g2_inv_1 _08915_ (.Y(_01668_),
    .A(net4087));
 sg13g2_inv_2 _08916_ (.Y(_01669_),
    .A(net3689));
 sg13g2_inv_1 _08917_ (.Y(_01670_),
    .A(\i_tinyqv.cpu.instr_data_in[9] ));
 sg13g2_inv_4 _08918_ (.A(net3786),
    .Y(_01671_));
 sg13g2_inv_1 _08919_ (.Y(_01672_),
    .A(net4040));
 sg13g2_inv_1 _08920_ (.Y(_01673_),
    .A(net7));
 sg13g2_inv_1 _08921_ (.Y(_01674_),
    .A(\i_tinyqv.mem.data_from_read[17] ));
 sg13g2_inv_2 _08922_ (.Y(_01675_),
    .A(net4079));
 sg13g2_inv_1 _08923_ (.Y(_01676_),
    .A(\i_latch_mem.data_out[10] ));
 sg13g2_inv_1 _08924_ (.Y(_01677_),
    .A(\i_latch_mem.data_out[18] ));
 sg13g2_inv_1 _08925_ (.Y(_01678_),
    .A(\i_tinyqv.mem.data_from_read[18] ));
 sg13g2_inv_1 _08926_ (.Y(_01679_),
    .A(\i_latch_mem.data_out[22] ));
 sg13g2_inv_1 _08927_ (.Y(_01680_),
    .A(\i_tinyqv.mem.data_from_read[22] ));
 sg13g2_inv_1 _08928_ (.Y(_01681_),
    .A(\i_latch_mem.data_out[26] ));
 sg13g2_inv_1 _08929_ (.Y(_01682_),
    .A(net3884));
 sg13g2_inv_1 _08930_ (.Y(_01683_),
    .A(\i_tinyqv.cpu.i_core.mepc[3] ));
 sg13g2_inv_2 _08931_ (.Y(_01684_),
    .A(net3940));
 sg13g2_inv_2 _08932_ (.Y(_01685_),
    .A(net5));
 sg13g2_inv_1 _08933_ (.Y(_01686_),
    .A(\i_latch_mem.data_out[3] ));
 sg13g2_inv_2 _08934_ (.Y(_01687_),
    .A(net4100));
 sg13g2_inv_1 _08935_ (.Y(_01688_),
    .A(\gpio_out_sel[7] ));
 sg13g2_inv_1 _08936_ (.Y(_01689_),
    .A(\gpio_out[7] ));
 sg13g2_inv_1 _08937_ (.Y(_01690_),
    .A(\i_latch_mem.data_out[7] ));
 sg13g2_inv_1 _08938_ (.Y(_01691_),
    .A(\i_tinyqv.mem.qspi_data_buf[11] ));
 sg13g2_inv_1 _08939_ (.Y(_01692_),
    .A(\i_latch_mem.data_out[11] ));
 sg13g2_inv_1 _08940_ (.Y(_01693_),
    .A(\i_latch_mem.data_out[15] ));
 sg13g2_inv_1 _08941_ (.Y(_01694_),
    .A(\i_latch_mem.data_out[27] ));
 sg13g2_inv_1 _08942_ (.Y(_01695_),
    .A(net3301));
 sg13g2_inv_1 _08943_ (.Y(_01696_),
    .A(net3682));
 sg13g2_inv_1 _08944_ (.Y(_01697_),
    .A(net3279));
 sg13g2_inv_1 _08945_ (.Y(_01698_),
    .A(net3451));
 sg13g2_inv_1 _08946_ (.Y(_01699_),
    .A(net3457));
 sg13g2_inv_1 _08947_ (.Y(_01700_),
    .A(\i_tinyqv.mem.q_ctrl.addr[7] ));
 sg13g2_inv_1 _08948_ (.Y(_01701_),
    .A(net3354));
 sg13g2_inv_1 _08949_ (.Y(_01702_),
    .A(net3468));
 sg13g2_inv_1 _08950_ (.Y(_01703_),
    .A(\i_tinyqv.mem.q_ctrl.addr[18] ));
 sg13g2_inv_1 _08951_ (.Y(_01704_),
    .A(\i_tinyqv.mem.q_ctrl.addr[19] ));
 sg13g2_inv_1 _08952_ (.Y(_01705_),
    .A(net3893));
 sg13g2_inv_1 _08953_ (.Y(_01706_),
    .A(\i_spi.end_txn_reg ));
 sg13g2_inv_1 _08954_ (.Y(_01707_),
    .A(net2822));
 sg13g2_inv_1 _14256__2 (.Y(net2109),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _08956_ (.Y(_01708_),
    .A(net2823));
 sg13g2_nand2_2 _08957_ (.Y(_01709_),
    .A(\i_tinyqv.cpu.data_write_n[1] ),
    .B(\i_tinyqv.cpu.data_write_n[0] ));
 sg13g2_and2_2 _08958_ (.A(net636),
    .B(_01709_),
    .X(_01710_));
 sg13g2_nand2_1 _08959_ (.Y(_01711_),
    .A(net636),
    .B(_01709_));
 sg13g2_nand2_1 _08960_ (.Y(_01712_),
    .A(\addr[0] ),
    .B(net639));
 sg13g2_xnor2_1 _08961_ (.Y(_01713_),
    .A(\addr[0] ),
    .B(net639));
 sg13g2_xnor2_1 _08962_ (.Y(_01714_),
    .A(net2380),
    .B(net640));
 sg13g2_or2_2 _08963_ (.X(_01715_),
    .B(net2385),
    .A(_01713_));
 sg13g2_nor2_1 _08964_ (.A(_01712_),
    .B(_01714_),
    .Y(_01716_));
 sg13g2_a21oi_1 _08965_ (.A1(net640),
    .A2(net2380),
    .Y(_01717_),
    .B1(_01716_));
 sg13g2_nor2b_1 _08966_ (.A(_01717_),
    .B_N(net632),
    .Y(_01718_));
 sg13g2_xnor2_1 _08967_ (.Y(_01719_),
    .A(net632),
    .B(_01717_));
 sg13g2_xnor2_1 _08968_ (.Y(_01720_),
    .A(_00198_),
    .B(_01718_));
 sg13g2_or2_2 _08969_ (.X(_01721_),
    .B(_01720_),
    .A(_01719_));
 sg13g2_nand2_1 _08970_ (.Y(_01722_),
    .A(\addr[3] ),
    .B(_01718_));
 sg13g2_xnor2_1 _08971_ (.Y(_01723_),
    .A(_01616_),
    .B(_01722_));
 sg13g2_xnor2_1 _08972_ (.Y(_01724_),
    .A(\addr[4] ),
    .B(_01722_));
 sg13g2_nor3_2 _08973_ (.A(_01715_),
    .B(_01721_),
    .C(net319),
    .Y(_01725_));
 sg13g2_and2_1 _08974_ (.A(net424),
    .B(net260),
    .X(_01726_));
 sg13g2_nor2b_1 _08975_ (.A(net639),
    .B_N(net640),
    .Y(_01727_));
 sg13g2_nor2b_2 _08976_ (.A(net640),
    .B_N(net639),
    .Y(_01728_));
 sg13g2_nand2b_2 _08977_ (.Y(_01729_),
    .B(net2386),
    .A_N(\i_latch_mem.cycle[1] ));
 sg13g2_a22oi_1 _08978_ (.Y(_01730_),
    .B1(_01728_),
    .B2(\data_to_write[15] ),
    .A2(net500),
    .A1(\data_to_write[23] ));
 sg13g2_and2_1 _08979_ (.A(net640),
    .B(net639),
    .X(_01731_));
 sg13g2_nand2_1 _08980_ (.Y(_01732_),
    .A(net640),
    .B(net639));
 sg13g2_nor2_1 _08981_ (.A(net640),
    .B(net639),
    .Y(_01733_));
 sg13g2_a22oi_1 _08982_ (.Y(_01734_),
    .B1(net490),
    .B2(\data_to_write[7] ),
    .A2(net495),
    .A1(\data_to_write[31] ));
 sg13g2_and2_1 _08983_ (.A(_01730_),
    .B(_01734_),
    .X(_01735_));
 sg13g2_nor2_1 _08984_ (.A(net3135),
    .B(net166),
    .Y(_01736_));
 sg13g2_a21oi_1 _08985_ (.A1(net166),
    .A2(net391),
    .Y(_01057_),
    .B1(_01736_));
 sg13g2_a22oi_1 _08986_ (.Y(_01737_),
    .B1(_01728_),
    .B2(\data_to_write[14] ),
    .A2(net500),
    .A1(\data_to_write[22] ));
 sg13g2_a22oi_1 _08987_ (.Y(_01738_),
    .B1(net490),
    .B2(net597),
    .A2(net495),
    .A1(\data_to_write[30] ));
 sg13g2_and2_1 _08988_ (.A(_01737_),
    .B(_01738_),
    .X(_01739_));
 sg13g2_nor2_1 _08989_ (.A(net3166),
    .B(net166),
    .Y(_01740_));
 sg13g2_a21oi_1 _08990_ (.A1(net166),
    .A2(net385),
    .Y(_01056_),
    .B1(_01740_));
 sg13g2_a22oi_1 _08991_ (.Y(_01741_),
    .B1(net490),
    .B2(net598),
    .A2(_01728_),
    .A1(\data_to_write[13] ));
 sg13g2_a22oi_1 _08992_ (.Y(_01742_),
    .B1(net495),
    .B2(\data_to_write[29] ),
    .A2(net500),
    .A1(\data_to_write[21] ));
 sg13g2_and2_1 _08993_ (.A(_01741_),
    .B(_01742_),
    .X(_01743_));
 sg13g2_nor2_1 _08994_ (.A(net3015),
    .B(net165),
    .Y(_01744_));
 sg13g2_a21oi_1 _08995_ (.A1(net165),
    .A2(net381),
    .Y(_01055_),
    .B1(_01744_));
 sg13g2_a22oi_1 _08996_ (.Y(_01745_),
    .B1(net490),
    .B2(net599),
    .A2(_01728_),
    .A1(\data_to_write[12] ));
 sg13g2_a22oi_1 _08997_ (.Y(_01746_),
    .B1(net495),
    .B2(\data_to_write[28] ),
    .A2(net500),
    .A1(\data_to_write[20] ));
 sg13g2_and2_1 _08998_ (.A(_01745_),
    .B(_01746_),
    .X(_01747_));
 sg13g2_nor2_1 _08999_ (.A(net3112),
    .B(net166),
    .Y(_01748_));
 sg13g2_a21oi_1 _09000_ (.A1(net166),
    .A2(net374),
    .Y(_01054_),
    .B1(_01748_));
 sg13g2_a22oi_1 _09001_ (.Y(_01749_),
    .B1(net490),
    .B2(\data_to_write[3] ),
    .A2(_01728_),
    .A1(\data_to_write[11] ));
 sg13g2_a22oi_1 _09002_ (.Y(_01750_),
    .B1(net495),
    .B2(\data_to_write[27] ),
    .A2(net500),
    .A1(\data_to_write[19] ));
 sg13g2_and2_2 _09003_ (.A(_01749_),
    .B(_01750_),
    .X(_01751_));
 sg13g2_nor2_1 _09004_ (.A(net3064),
    .B(net165),
    .Y(_01752_));
 sg13g2_a21oi_1 _09005_ (.A1(net165),
    .A2(net371),
    .Y(_01053_),
    .B1(_01752_));
 sg13g2_a22oi_1 _09006_ (.Y(_01753_),
    .B1(net490),
    .B2(net600),
    .A2(_01728_),
    .A1(\data_to_write[10] ));
 sg13g2_a22oi_1 _09007_ (.Y(_01754_),
    .B1(_01731_),
    .B2(\data_to_write[26] ),
    .A2(net500),
    .A1(\data_to_write[18] ));
 sg13g2_and2_2 _09008_ (.A(_01753_),
    .B(_01754_),
    .X(_01755_));
 sg13g2_nor2_1 _09009_ (.A(net3047),
    .B(net165),
    .Y(_01756_));
 sg13g2_a21oi_1 _09010_ (.A1(net165),
    .A2(net365),
    .Y(_01052_),
    .B1(_01756_));
 sg13g2_a22oi_1 _09011_ (.Y(_01757_),
    .B1(_01733_),
    .B2(net601),
    .A2(_01728_),
    .A1(\data_to_write[9] ));
 sg13g2_a22oi_1 _09012_ (.Y(_01758_),
    .B1(_01731_),
    .B2(\data_to_write[25] ),
    .A2(_01727_),
    .A1(\data_to_write[17] ));
 sg13g2_and2_1 _09013_ (.A(_01757_),
    .B(_01758_),
    .X(_01759_));
 sg13g2_nor2_1 _09014_ (.A(net2986),
    .B(net165),
    .Y(_01760_));
 sg13g2_a21oi_1 _09015_ (.A1(net165),
    .A2(net360),
    .Y(_01051_),
    .B1(_01760_));
 sg13g2_a22oi_1 _09016_ (.Y(_01761_),
    .B1(net490),
    .B2(\data_to_write[0] ),
    .A2(_01728_),
    .A1(\data_to_write[8] ));
 sg13g2_a22oi_1 _09017_ (.Y(_01762_),
    .B1(_01731_),
    .B2(\data_to_write[24] ),
    .A2(net500),
    .A1(\data_to_write[16] ));
 sg13g2_and2_2 _09018_ (.A(_01761_),
    .B(_01762_),
    .X(_01763_));
 sg13g2_nor2_1 _09019_ (.A(net3117),
    .B(net166),
    .Y(_01764_));
 sg13g2_a21oi_1 _09020_ (.A1(net166),
    .A2(net356),
    .Y(_01050_),
    .B1(_01764_));
 sg13g2_nand2b_2 _09021_ (.Y(_01765_),
    .B(_01719_),
    .A_N(_00198_));
 sg13g2_nand2b_2 _09022_ (.Y(_01766_),
    .B(net2384),
    .A_N(_01713_));
 sg13g2_nor3_2 _09023_ (.A(net320),
    .B(_01765_),
    .C(_01766_),
    .Y(_01767_));
 sg13g2_nand2_1 _09024_ (.Y(_01768_),
    .A(net426),
    .B(net259));
 sg13g2_nand2_1 _09025_ (.Y(_01769_),
    .A(net2991),
    .B(net200));
 sg13g2_o21ai_1 _09026_ (.B1(_01769_),
    .Y(_01049_),
    .A1(net395),
    .A2(net200));
 sg13g2_nand2_1 _09027_ (.Y(_01770_),
    .A(net2918),
    .B(net201));
 sg13g2_o21ai_1 _09028_ (.B1(_01770_),
    .Y(_01048_),
    .A1(net388),
    .A2(_01768_));
 sg13g2_nand2_1 _09029_ (.Y(_01771_),
    .A(net2916),
    .B(net201));
 sg13g2_o21ai_1 _09030_ (.B1(_01771_),
    .Y(_01047_),
    .A1(net383),
    .A2(net201));
 sg13g2_nand2_1 _09031_ (.Y(_01772_),
    .A(net2984),
    .B(net201));
 sg13g2_o21ai_1 _09032_ (.B1(_01772_),
    .Y(_01046_),
    .A1(net377),
    .A2(net201));
 sg13g2_nand2_1 _09033_ (.Y(_01773_),
    .A(net2946),
    .B(net200));
 sg13g2_o21ai_1 _09034_ (.B1(_01773_),
    .Y(_01045_),
    .A1(net373),
    .A2(net200));
 sg13g2_nand2_1 _09035_ (.Y(_01774_),
    .A(net3110),
    .B(net200));
 sg13g2_o21ai_1 _09036_ (.B1(_01774_),
    .Y(_01044_),
    .A1(net369),
    .A2(net200));
 sg13g2_nand2_1 _09037_ (.Y(_01775_),
    .A(net2985),
    .B(net200));
 sg13g2_o21ai_1 _09038_ (.B1(_01775_),
    .Y(_01043_),
    .A1(net363),
    .A2(net200));
 sg13g2_nand2_1 _09039_ (.Y(_01776_),
    .A(net2875),
    .B(net201));
 sg13g2_o21ai_1 _09040_ (.B1(_01776_),
    .Y(_01042_),
    .A1(net358),
    .A2(net201));
 sg13g2_nor3_2 _09041_ (.A(_01715_),
    .B(net320),
    .C(_01765_),
    .Y(_01777_));
 sg13g2_nand2_1 _09042_ (.Y(_01778_),
    .A(net425),
    .B(net258));
 sg13g2_nand2_1 _09043_ (.Y(_01779_),
    .A(net3006),
    .B(net199));
 sg13g2_o21ai_1 _09044_ (.B1(_01779_),
    .Y(_01041_),
    .A1(net394),
    .A2(net198));
 sg13g2_nand2_1 _09045_ (.Y(_01780_),
    .A(net2980),
    .B(net199));
 sg13g2_o21ai_1 _09046_ (.B1(_01780_),
    .Y(_01040_),
    .A1(net388),
    .A2(net198));
 sg13g2_nand2_1 _09047_ (.Y(_01781_),
    .A(net2973),
    .B(net199));
 sg13g2_o21ai_1 _09048_ (.B1(_01781_),
    .Y(_01039_),
    .A1(net383),
    .A2(net199));
 sg13g2_nand2_1 _09049_ (.Y(_01782_),
    .A(net2994),
    .B(net198));
 sg13g2_o21ai_1 _09050_ (.B1(_01782_),
    .Y(_01038_),
    .A1(net377),
    .A2(net198));
 sg13g2_nand2_1 _09051_ (.Y(_01783_),
    .A(net2968),
    .B(net199));
 sg13g2_o21ai_1 _09052_ (.B1(_01783_),
    .Y(_01037_),
    .A1(net373),
    .A2(net199));
 sg13g2_nand2_1 _09053_ (.Y(_01784_),
    .A(net2907),
    .B(net198));
 sg13g2_o21ai_1 _09054_ (.B1(_01784_),
    .Y(_01036_),
    .A1(net368),
    .A2(net198));
 sg13g2_nand2_1 _09055_ (.Y(_01785_),
    .A(net2870),
    .B(net198));
 sg13g2_o21ai_1 _09056_ (.B1(_01785_),
    .Y(_01035_),
    .A1(net363),
    .A2(net198));
 sg13g2_nand2_1 _09057_ (.Y(_01786_),
    .A(net2849),
    .B(_01778_));
 sg13g2_o21ai_1 _09058_ (.B1(_01786_),
    .Y(_01034_),
    .A1(net358),
    .A2(net199));
 sg13g2_nor3_2 _09059_ (.A(_01715_),
    .B(_01721_),
    .C(net317),
    .Y(_01787_));
 sg13g2_and2_1 _09060_ (.A(net422),
    .B(_01787_),
    .X(_01788_));
 sg13g2_nor2_1 _09061_ (.A(net3245),
    .B(net163),
    .Y(_01789_));
 sg13g2_a21oi_1 _09062_ (.A1(net391),
    .A2(net163),
    .Y(_01033_),
    .B1(_01789_));
 sg13g2_nor2_1 _09063_ (.A(net3000),
    .B(net164),
    .Y(_01790_));
 sg13g2_a21oi_1 _09064_ (.A1(net386),
    .A2(_01788_),
    .Y(_01032_),
    .B1(_01790_));
 sg13g2_nor2_1 _09065_ (.A(net3040),
    .B(net163),
    .Y(_01791_));
 sg13g2_a21oi_1 _09066_ (.A1(net382),
    .A2(net163),
    .Y(_01031_),
    .B1(_01791_));
 sg13g2_nor2_1 _09067_ (.A(net3174),
    .B(net163),
    .Y(_01792_));
 sg13g2_a21oi_1 _09068_ (.A1(net374),
    .A2(net163),
    .Y(_01030_),
    .B1(_01792_));
 sg13g2_nor2_1 _09069_ (.A(net3184),
    .B(net164),
    .Y(_01793_));
 sg13g2_a21oi_1 _09070_ (.A1(net371),
    .A2(net164),
    .Y(_01029_),
    .B1(_01793_));
 sg13g2_nor2_1 _09071_ (.A(net3133),
    .B(net164),
    .Y(_01794_));
 sg13g2_a21oi_1 _09072_ (.A1(net365),
    .A2(net164),
    .Y(_01028_),
    .B1(_01794_));
 sg13g2_nor2_1 _09073_ (.A(net3171),
    .B(net163),
    .Y(_01795_));
 sg13g2_a21oi_1 _09074_ (.A1(net361),
    .A2(net163),
    .Y(_01027_),
    .B1(_01795_));
 sg13g2_nor2_1 _09075_ (.A(net3005),
    .B(net164),
    .Y(_01796_));
 sg13g2_a21oi_1 _09076_ (.A1(net354),
    .A2(net164),
    .Y(_01026_),
    .B1(_01796_));
 sg13g2_xnor2_1 _09077_ (.Y(_01797_),
    .A(_01712_),
    .B(net2384));
 sg13g2_nand2_2 _09078_ (.Y(_01798_),
    .A(_01713_),
    .B(_01797_));
 sg13g2_nand2_2 _09079_ (.Y(_01799_),
    .A(_00198_),
    .B(_01719_));
 sg13g2_nor3_1 _09080_ (.A(net318),
    .B(_01798_),
    .C(_01799_),
    .Y(_01800_));
 sg13g2_and2_1 _09081_ (.A(net425),
    .B(_01800_),
    .X(_01801_));
 sg13g2_nor2_1 _09082_ (.A(net3013),
    .B(net161),
    .Y(_01802_));
 sg13g2_a21oi_1 _09083_ (.A1(net394),
    .A2(net161),
    .Y(_01025_),
    .B1(_01802_));
 sg13g2_nor2_1 _09084_ (.A(net3203),
    .B(net161),
    .Y(_01803_));
 sg13g2_a21oi_1 _09085_ (.A1(net388),
    .A2(net161),
    .Y(_01024_),
    .B1(_01803_));
 sg13g2_nor2_1 _09086_ (.A(net3172),
    .B(net162),
    .Y(_01804_));
 sg13g2_a21oi_1 _09087_ (.A1(net381),
    .A2(net162),
    .Y(_01023_),
    .B1(_01804_));
 sg13g2_nor2_1 _09088_ (.A(net3086),
    .B(net161),
    .Y(_01805_));
 sg13g2_a21oi_1 _09089_ (.A1(net377),
    .A2(net161),
    .Y(_01022_),
    .B1(_01805_));
 sg13g2_nor2_1 _09090_ (.A(net3037),
    .B(net162),
    .Y(_01806_));
 sg13g2_a21oi_1 _09091_ (.A1(net372),
    .A2(net162),
    .Y(_01021_),
    .B1(_01806_));
 sg13g2_nor2_1 _09092_ (.A(net3225),
    .B(net162),
    .Y(_01807_));
 sg13g2_a21oi_1 _09093_ (.A1(net368),
    .A2(net161),
    .Y(_01020_),
    .B1(_01807_));
 sg13g2_nor2_1 _09094_ (.A(net3216),
    .B(_01801_),
    .Y(_01808_));
 sg13g2_a21oi_1 _09095_ (.A1(net363),
    .A2(net161),
    .Y(_01019_),
    .B1(_01808_));
 sg13g2_nor2_1 _09096_ (.A(net3096),
    .B(net162),
    .Y(_01809_));
 sg13g2_a21oi_1 _09097_ (.A1(net354),
    .A2(net162),
    .Y(_01018_),
    .B1(_01809_));
 sg13g2_nor3_1 _09098_ (.A(net318),
    .B(_01766_),
    .C(_01799_),
    .Y(_01810_));
 sg13g2_and2_1 _09099_ (.A(net424),
    .B(_01810_),
    .X(_01811_));
 sg13g2_nor2_1 _09100_ (.A(net2981),
    .B(net158),
    .Y(_01812_));
 sg13g2_a21oi_1 _09101_ (.A1(net393),
    .A2(net158),
    .Y(_01017_),
    .B1(_01812_));
 sg13g2_nor2_1 _09102_ (.A(net3094),
    .B(net158),
    .Y(_01813_));
 sg13g2_a21oi_1 _09103_ (.A1(net387),
    .A2(net158),
    .Y(_01016_),
    .B1(_01813_));
 sg13g2_nor2_1 _09104_ (.A(net3291),
    .B(net160),
    .Y(_01814_));
 sg13g2_a21oi_1 _09105_ (.A1(net380),
    .A2(net160),
    .Y(_01015_),
    .B1(_01814_));
 sg13g2_nor2_1 _09106_ (.A(net3004),
    .B(net160),
    .Y(_01815_));
 sg13g2_a21oi_1 _09107_ (.A1(net376),
    .A2(net160),
    .Y(_01014_),
    .B1(_01815_));
 sg13g2_nor2_1 _09108_ (.A(net3163),
    .B(net159),
    .Y(_01816_));
 sg13g2_a21oi_1 _09109_ (.A1(net370),
    .A2(net160),
    .Y(_01013_),
    .B1(_01816_));
 sg13g2_nor2_1 _09110_ (.A(net3045),
    .B(net158),
    .Y(_01817_));
 sg13g2_a21oi_1 _09111_ (.A1(net366),
    .A2(net159),
    .Y(_01012_),
    .B1(_01817_));
 sg13g2_nor2_1 _09112_ (.A(net3169),
    .B(net158),
    .Y(_01818_));
 sg13g2_a21oi_1 _09113_ (.A1(net359),
    .A2(net158),
    .Y(_01011_),
    .B1(_01818_));
 sg13g2_nor2_1 _09114_ (.A(net2993),
    .B(net158),
    .Y(_01819_));
 sg13g2_a21oi_1 _09115_ (.A1(net355),
    .A2(net159),
    .Y(_01010_),
    .B1(_01819_));
 sg13g2_nand2b_2 _09116_ (.Y(_01820_),
    .B(_01713_),
    .A_N(_01797_));
 sg13g2_nor3_1 _09117_ (.A(net318),
    .B(_01799_),
    .C(_01820_),
    .Y(_01821_));
 sg13g2_and2_1 _09118_ (.A(net424),
    .B(_01821_),
    .X(_01822_));
 sg13g2_nor2_1 _09119_ (.A(net3016),
    .B(net155),
    .Y(_01823_));
 sg13g2_a21oi_1 _09120_ (.A1(net393),
    .A2(net155),
    .Y(_01009_),
    .B1(_01823_));
 sg13g2_nor2_1 _09121_ (.A(net3028),
    .B(net155),
    .Y(_01824_));
 sg13g2_a21oi_1 _09122_ (.A1(net387),
    .A2(net155),
    .Y(_01008_),
    .B1(_01824_));
 sg13g2_nor2_1 _09123_ (.A(net3111),
    .B(net157),
    .Y(_01825_));
 sg13g2_a21oi_1 _09124_ (.A1(net381),
    .A2(net157),
    .Y(_01007_),
    .B1(_01825_));
 sg13g2_nor2_1 _09125_ (.A(net3003),
    .B(net155),
    .Y(_01826_));
 sg13g2_a21oi_1 _09126_ (.A1(net376),
    .A2(net155),
    .Y(_01006_),
    .B1(_01826_));
 sg13g2_nor2_1 _09127_ (.A(net3127),
    .B(net156),
    .Y(_01827_));
 sg13g2_a21oi_1 _09128_ (.A1(net371),
    .A2(net155),
    .Y(_01005_),
    .B1(_01827_));
 sg13g2_nor2_1 _09129_ (.A(net3167),
    .B(net156),
    .Y(_01828_));
 sg13g2_a21oi_1 _09130_ (.A1(net366),
    .A2(net156),
    .Y(_01004_),
    .B1(_01828_));
 sg13g2_nor2_1 _09131_ (.A(net3208),
    .B(net155),
    .Y(_01829_));
 sg13g2_a21oi_1 _09132_ (.A1(net359),
    .A2(net156),
    .Y(_01003_),
    .B1(_01829_));
 sg13g2_nor2_1 _09133_ (.A(net3087),
    .B(net157),
    .Y(_01830_));
 sg13g2_a21oi_1 _09134_ (.A1(net354),
    .A2(net157),
    .Y(_01002_),
    .B1(_01830_));
 sg13g2_nor3_2 _09135_ (.A(_01715_),
    .B(net318),
    .C(_01799_),
    .Y(_01831_));
 sg13g2_and2_1 _09136_ (.A(net424),
    .B(net253),
    .X(_01832_));
 sg13g2_nor2_1 _09137_ (.A(net3030),
    .B(net153),
    .Y(_01833_));
 sg13g2_a21oi_1 _09138_ (.A1(net393),
    .A2(net153),
    .Y(_01001_),
    .B1(_01833_));
 sg13g2_nor2_1 _09139_ (.A(net3252),
    .B(net154),
    .Y(_01834_));
 sg13g2_a21oi_1 _09140_ (.A1(net387),
    .A2(net154),
    .Y(_01000_),
    .B1(_01834_));
 sg13g2_nor2_1 _09141_ (.A(net3165),
    .B(net154),
    .Y(_01835_));
 sg13g2_a21oi_1 _09142_ (.A1(net380),
    .A2(net154),
    .Y(_00999_),
    .B1(_01835_));
 sg13g2_nor2_1 _09143_ (.A(net3153),
    .B(net153),
    .Y(_01836_));
 sg13g2_a21oi_1 _09144_ (.A1(net376),
    .A2(net153),
    .Y(_00998_),
    .B1(_01836_));
 sg13g2_nor2_1 _09145_ (.A(net3170),
    .B(net154),
    .Y(_01837_));
 sg13g2_a21oi_1 _09146_ (.A1(net370),
    .A2(net154),
    .Y(_00997_),
    .B1(_01837_));
 sg13g2_nor2_1 _09147_ (.A(net3168),
    .B(net153),
    .Y(_01838_));
 sg13g2_a21oi_1 _09148_ (.A1(net365),
    .A2(net153),
    .Y(_00996_),
    .B1(_01838_));
 sg13g2_nor2_1 _09149_ (.A(net3076),
    .B(net153),
    .Y(_01839_));
 sg13g2_a21oi_1 _09150_ (.A1(net359),
    .A2(net153),
    .Y(_00995_),
    .B1(_01839_));
 sg13g2_nor2_1 _09151_ (.A(net3244),
    .B(net154),
    .Y(_01840_));
 sg13g2_a21oi_1 _09152_ (.A1(net354),
    .A2(net154),
    .Y(_00994_),
    .B1(_01840_));
 sg13g2_nand2b_2 _09153_ (.Y(_01841_),
    .B(_01720_),
    .A_N(_01719_));
 sg13g2_nor3_2 _09154_ (.A(net317),
    .B(_01798_),
    .C(_01841_),
    .Y(_01842_));
 sg13g2_nand2_1 _09155_ (.Y(_01843_),
    .A(net422),
    .B(_01842_));
 sg13g2_nand2_1 _09156_ (.Y(_01844_),
    .A(net2926),
    .B(net151));
 sg13g2_o21ai_1 _09157_ (.B1(_01844_),
    .Y(_00993_),
    .A1(net391),
    .A2(net151));
 sg13g2_nand2_1 _09158_ (.Y(_01845_),
    .A(net2886),
    .B(net151));
 sg13g2_o21ai_1 _09159_ (.B1(_01845_),
    .Y(_00992_),
    .A1(net385),
    .A2(net151));
 sg13g2_nand2_1 _09160_ (.Y(_01846_),
    .A(net2851),
    .B(net151));
 sg13g2_o21ai_1 _09161_ (.B1(_01846_),
    .Y(_00991_),
    .A1(net382),
    .A2(_01843_));
 sg13g2_nand2_1 _09162_ (.Y(_01847_),
    .A(net2868),
    .B(net151));
 sg13g2_o21ai_1 _09163_ (.B1(_01847_),
    .Y(_00990_),
    .A1(net374),
    .A2(net151));
 sg13g2_nand2_1 _09164_ (.Y(_01848_),
    .A(net2905),
    .B(net152));
 sg13g2_o21ai_1 _09165_ (.B1(_01848_),
    .Y(_00989_),
    .A1(net371),
    .A2(net152));
 sg13g2_nand2_1 _09166_ (.Y(_01849_),
    .A(net2930),
    .B(net152));
 sg13g2_o21ai_1 _09167_ (.B1(_01849_),
    .Y(_00988_),
    .A1(net366),
    .A2(net152));
 sg13g2_nand2_1 _09168_ (.Y(_01850_),
    .A(net2942),
    .B(net152));
 sg13g2_o21ai_1 _09169_ (.B1(_01850_),
    .Y(_00987_),
    .A1(net360),
    .A2(net151));
 sg13g2_nand2_1 _09170_ (.Y(_01851_),
    .A(net2937),
    .B(net152));
 sg13g2_o21ai_1 _09171_ (.B1(_01851_),
    .Y(_00986_),
    .A1(net354),
    .A2(net152));
 sg13g2_or2_1 _09172_ (.X(_01852_),
    .B(_01798_),
    .A(_01721_));
 sg13g2_nor2_2 _09173_ (.A(net317),
    .B(_01852_),
    .Y(_01853_));
 sg13g2_nor3_1 _09174_ (.A(_01711_),
    .B(_01724_),
    .C(_01852_),
    .Y(_01854_));
 sg13g2_nor2_1 _09175_ (.A(net2949),
    .B(net249),
    .Y(_01855_));
 sg13g2_a21oi_1 _09176_ (.A1(net396),
    .A2(net249),
    .Y(_00985_),
    .B1(_01855_));
 sg13g2_nor2_1 _09177_ (.A(net3009),
    .B(net249),
    .Y(_01856_));
 sg13g2_a21oi_1 _09178_ (.A1(net389),
    .A2(_01854_),
    .Y(_00984_),
    .B1(_01856_));
 sg13g2_nor2_1 _09179_ (.A(net2957),
    .B(net248),
    .Y(_01857_));
 sg13g2_a21oi_1 _09180_ (.A1(net384),
    .A2(net248),
    .Y(_00983_),
    .B1(_01857_));
 sg13g2_nor2_1 _09181_ (.A(net2962),
    .B(net249),
    .Y(_01858_));
 sg13g2_a21oi_1 _09182_ (.A1(net378),
    .A2(net249),
    .Y(_00982_),
    .B1(_01858_));
 sg13g2_nor2_1 _09183_ (.A(net3041),
    .B(net248),
    .Y(_01859_));
 sg13g2_a21oi_1 _09184_ (.A1(_01751_),
    .A2(net248),
    .Y(_00981_),
    .B1(_01859_));
 sg13g2_nor2_1 _09185_ (.A(net2979),
    .B(net248),
    .Y(_01860_));
 sg13g2_a21oi_1 _09186_ (.A1(net368),
    .A2(net248),
    .Y(_00980_),
    .B1(_01860_));
 sg13g2_nor2_1 _09187_ (.A(net3029),
    .B(net249),
    .Y(_01861_));
 sg13g2_a21oi_1 _09188_ (.A1(net364),
    .A2(net249),
    .Y(_00979_),
    .B1(_01861_));
 sg13g2_nor2_1 _09189_ (.A(net2928),
    .B(net248),
    .Y(_01862_));
 sg13g2_a21oi_1 _09190_ (.A1(net358),
    .A2(net248),
    .Y(_00978_),
    .B1(_01862_));
 sg13g2_nor3_1 _09191_ (.A(net317),
    .B(_01820_),
    .C(_01841_),
    .Y(_01863_));
 sg13g2_nand2_1 _09192_ (.Y(_01864_),
    .A(net423),
    .B(_01863_));
 sg13g2_nand2_1 _09193_ (.Y(_01865_),
    .A(net2869),
    .B(net149));
 sg13g2_o21ai_1 _09194_ (.B1(_01865_),
    .Y(_00977_),
    .A1(net393),
    .A2(net149));
 sg13g2_nand2_1 _09195_ (.Y(_01866_),
    .A(net2895),
    .B(net149));
 sg13g2_o21ai_1 _09196_ (.B1(_01866_),
    .Y(_00976_),
    .A1(net387),
    .A2(net149));
 sg13g2_nand2_1 _09197_ (.Y(_01867_),
    .A(net2892),
    .B(net149));
 sg13g2_o21ai_1 _09198_ (.B1(_01867_),
    .Y(_00975_),
    .A1(net381),
    .A2(net149));
 sg13g2_nand2_1 _09199_ (.Y(_01868_),
    .A(net2959),
    .B(net150));
 sg13g2_o21ai_1 _09200_ (.B1(_01868_),
    .Y(_00974_),
    .A1(net375),
    .A2(net150));
 sg13g2_nand2_1 _09201_ (.Y(_01869_),
    .A(net2860),
    .B(net149));
 sg13g2_o21ai_1 _09202_ (.B1(_01869_),
    .Y(_00973_),
    .A1(net370),
    .A2(net149));
 sg13g2_nand2_1 _09203_ (.Y(_01870_),
    .A(net3027),
    .B(net150));
 sg13g2_o21ai_1 _09204_ (.B1(_01870_),
    .Y(_00972_),
    .A1(net367),
    .A2(net150));
 sg13g2_nand2_1 _09205_ (.Y(_01871_),
    .A(net2879),
    .B(net150));
 sg13g2_o21ai_1 _09206_ (.B1(_01871_),
    .Y(_00971_),
    .A1(net361),
    .A2(_01864_));
 sg13g2_nand2_1 _09207_ (.Y(_01872_),
    .A(net2861),
    .B(net150));
 sg13g2_o21ai_1 _09208_ (.B1(_01872_),
    .Y(_00970_),
    .A1(net354),
    .A2(net150));
 sg13g2_nor3_1 _09209_ (.A(_01715_),
    .B(net317),
    .C(_01841_),
    .Y(_01873_));
 sg13g2_nand2_1 _09210_ (.Y(_01874_),
    .A(net423),
    .B(net246));
 sg13g2_nand2_1 _09211_ (.Y(_01875_),
    .A(net2953),
    .B(net147));
 sg13g2_o21ai_1 _09212_ (.B1(_01875_),
    .Y(_00969_),
    .A1(net391),
    .A2(net147));
 sg13g2_nand2_1 _09213_ (.Y(_01876_),
    .A(net2922),
    .B(net148));
 sg13g2_o21ai_1 _09214_ (.B1(_01876_),
    .Y(_00968_),
    .A1(net386),
    .A2(net148));
 sg13g2_nand2_1 _09215_ (.Y(_01877_),
    .A(net2909),
    .B(net148));
 sg13g2_o21ai_1 _09216_ (.B1(_01877_),
    .Y(_00967_),
    .A1(net382),
    .A2(net148));
 sg13g2_nand2_1 _09217_ (.Y(_01878_),
    .A(net2978),
    .B(net147));
 sg13g2_o21ai_1 _09218_ (.B1(_01878_),
    .Y(_00966_),
    .A1(net374),
    .A2(net147));
 sg13g2_nand2_1 _09219_ (.Y(_01879_),
    .A(net2931),
    .B(net148));
 sg13g2_o21ai_1 _09220_ (.B1(_01879_),
    .Y(_00965_),
    .A1(net372),
    .A2(net148));
 sg13g2_nand2_1 _09221_ (.Y(_01880_),
    .A(net2943),
    .B(net148));
 sg13g2_o21ai_1 _09222_ (.B1(_01880_),
    .Y(_00964_),
    .A1(net367),
    .A2(net148));
 sg13g2_nand2_1 _09223_ (.Y(_01881_),
    .A(net2924),
    .B(net147));
 sg13g2_o21ai_1 _09224_ (.B1(_01881_),
    .Y(_00963_),
    .A1(net361),
    .A2(net147));
 sg13g2_nand2_1 _09225_ (.Y(_01882_),
    .A(net2890),
    .B(net147));
 sg13g2_o21ai_1 _09226_ (.B1(_01882_),
    .Y(_00962_),
    .A1(net357),
    .A2(net147));
 sg13g2_nor3_2 _09227_ (.A(net318),
    .B(_01765_),
    .C(_01798_),
    .Y(_01883_));
 sg13g2_nand2_1 _09228_ (.Y(_01884_),
    .A(net424),
    .B(net245));
 sg13g2_nand2_1 _09229_ (.Y(_01885_),
    .A(net2972),
    .B(net146));
 sg13g2_o21ai_1 _09230_ (.B1(_01885_),
    .Y(_00961_),
    .A1(net394),
    .A2(net146));
 sg13g2_nand2_1 _09231_ (.Y(_01886_),
    .A(net2867),
    .B(net145));
 sg13g2_o21ai_1 _09232_ (.B1(_01886_),
    .Y(_00960_),
    .A1(net387),
    .A2(net145));
 sg13g2_nand2_1 _09233_ (.Y(_01887_),
    .A(net2948),
    .B(net145));
 sg13g2_o21ai_1 _09234_ (.B1(_01887_),
    .Y(_00959_),
    .A1(net380),
    .A2(net145));
 sg13g2_nand2_1 _09235_ (.Y(_01888_),
    .A(net2992),
    .B(net146));
 sg13g2_o21ai_1 _09236_ (.B1(_01888_),
    .Y(_00958_),
    .A1(net377),
    .A2(net146));
 sg13g2_nand2_1 _09237_ (.Y(_01889_),
    .A(net2945),
    .B(net145));
 sg13g2_o21ai_1 _09238_ (.B1(_01889_),
    .Y(_00957_),
    .A1(net370),
    .A2(net145));
 sg13g2_nand2_1 _09239_ (.Y(_01890_),
    .A(net2902),
    .B(net146));
 sg13g2_o21ai_1 _09240_ (.B1(_01890_),
    .Y(_00956_),
    .A1(net368),
    .A2(net146));
 sg13g2_nand2_1 _09241_ (.Y(_01891_),
    .A(net2947),
    .B(net146));
 sg13g2_o21ai_1 _09242_ (.B1(_01891_),
    .Y(_00955_),
    .A1(net359),
    .A2(net146));
 sg13g2_nand2_1 _09243_ (.Y(_01892_),
    .A(net2855),
    .B(net145));
 sg13g2_o21ai_1 _09244_ (.B1(_01892_),
    .Y(_00954_),
    .A1(net355),
    .A2(net145));
 sg13g2_nor3_2 _09245_ (.A(net318),
    .B(_01765_),
    .C(_01766_),
    .Y(_01893_));
 sg13g2_nand2_2 _09246_ (.Y(_01894_),
    .A(net425),
    .B(net244));
 sg13g2_nand2_1 _09247_ (.Y(_01895_),
    .A(net2966),
    .B(net144));
 sg13g2_o21ai_1 _09248_ (.B1(_01895_),
    .Y(_00953_),
    .A1(net394),
    .A2(net144));
 sg13g2_nand2_1 _09249_ (.Y(_01896_),
    .A(net2903),
    .B(net144));
 sg13g2_o21ai_1 _09250_ (.B1(_01896_),
    .Y(_00952_),
    .A1(net388),
    .A2(net144));
 sg13g2_nand2_1 _09251_ (.Y(_01897_),
    .A(net2983),
    .B(net143));
 sg13g2_o21ai_1 _09252_ (.B1(_01897_),
    .Y(_00951_),
    .A1(net380),
    .A2(net143));
 sg13g2_nand2_1 _09253_ (.Y(_01898_),
    .A(net2858),
    .B(net144));
 sg13g2_o21ai_1 _09254_ (.B1(_01898_),
    .Y(_00950_),
    .A1(net378),
    .A2(net144));
 sg13g2_nand2_1 _09255_ (.Y(_01899_),
    .A(net2896),
    .B(net143));
 sg13g2_o21ai_1 _09256_ (.B1(_01899_),
    .Y(_00949_),
    .A1(net370),
    .A2(net143));
 sg13g2_nand2_1 _09257_ (.Y(_01900_),
    .A(net2852),
    .B(net143));
 sg13g2_o21ai_1 _09258_ (.B1(_01900_),
    .Y(_00948_),
    .A1(net365),
    .A2(net143));
 sg13g2_nand2_1 _09259_ (.Y(_01901_),
    .A(net2863),
    .B(net144));
 sg13g2_o21ai_1 _09260_ (.B1(_01901_),
    .Y(_00947_),
    .A1(net363),
    .A2(net144));
 sg13g2_nand2_1 _09261_ (.Y(_01902_),
    .A(net2933),
    .B(net143));
 sg13g2_o21ai_1 _09262_ (.B1(_01902_),
    .Y(_00946_),
    .A1(net355),
    .A2(net143));
 sg13g2_nor3_2 _09263_ (.A(net318),
    .B(_01765_),
    .C(_01820_),
    .Y(_01903_));
 sg13g2_nand2_2 _09264_ (.Y(_01904_),
    .A(net425),
    .B(net243));
 sg13g2_nand2_1 _09265_ (.Y(_01905_),
    .A(net2848),
    .B(net197));
 sg13g2_o21ai_1 _09266_ (.B1(_01905_),
    .Y(_00945_),
    .A1(net394),
    .A2(net197));
 sg13g2_nand2_1 _09267_ (.Y(_01906_),
    .A(net2872),
    .B(net196));
 sg13g2_o21ai_1 _09268_ (.B1(_01906_),
    .Y(_00944_),
    .A1(net387),
    .A2(net196));
 sg13g2_nand2_1 _09269_ (.Y(_01907_),
    .A(net2915),
    .B(net196));
 sg13g2_o21ai_1 _09270_ (.B1(_01907_),
    .Y(_00943_),
    .A1(net380),
    .A2(net196));
 sg13g2_nand2_1 _09271_ (.Y(_01908_),
    .A(net2865),
    .B(net197));
 sg13g2_o21ai_1 _09272_ (.B1(_01908_),
    .Y(_00942_),
    .A1(net377),
    .A2(net197));
 sg13g2_nand2_1 _09273_ (.Y(_01909_),
    .A(net2956),
    .B(net197));
 sg13g2_o21ai_1 _09274_ (.B1(_01909_),
    .Y(_00941_),
    .A1(net371),
    .A2(net197));
 sg13g2_nand2_1 _09275_ (.Y(_01910_),
    .A(net2908),
    .B(net196));
 sg13g2_o21ai_1 _09276_ (.B1(_01910_),
    .Y(_00940_),
    .A1(net365),
    .A2(net196));
 sg13g2_nand2_1 _09277_ (.Y(_01911_),
    .A(net2850),
    .B(net197));
 sg13g2_o21ai_1 _09278_ (.B1(_01911_),
    .Y(_00939_),
    .A1(net363),
    .A2(net197));
 sg13g2_nand2_1 _09279_ (.Y(_01912_),
    .A(net2912),
    .B(net196));
 sg13g2_o21ai_1 _09280_ (.B1(_01912_),
    .Y(_00938_),
    .A1(net355),
    .A2(net196));
 sg13g2_nor3_2 _09281_ (.A(_01715_),
    .B(net318),
    .C(_01765_),
    .Y(_01913_));
 sg13g2_nand2_1 _09282_ (.Y(_01914_),
    .A(net425),
    .B(net242));
 sg13g2_nand2_1 _09283_ (.Y(_01915_),
    .A(net2847),
    .B(net194));
 sg13g2_o21ai_1 _09284_ (.B1(_01915_),
    .Y(_00937_),
    .A1(net394),
    .A2(net194));
 sg13g2_nand2_1 _09285_ (.Y(_01916_),
    .A(net2938),
    .B(net193));
 sg13g2_o21ai_1 _09286_ (.B1(_01916_),
    .Y(_00936_),
    .A1(net387),
    .A2(net193));
 sg13g2_nand2_1 _09287_ (.Y(_01917_),
    .A(net2934),
    .B(net195));
 sg13g2_o21ai_1 _09288_ (.B1(_01917_),
    .Y(_00935_),
    .A1(net383),
    .A2(net195));
 sg13g2_nand2_1 _09289_ (.Y(_01918_),
    .A(net2876),
    .B(net194));
 sg13g2_o21ai_1 _09290_ (.B1(_01918_),
    .Y(_00934_),
    .A1(net376),
    .A2(net193));
 sg13g2_nand2_1 _09291_ (.Y(_01919_),
    .A(net2929),
    .B(net193));
 sg13g2_o21ai_1 _09292_ (.B1(_01919_),
    .Y(_00933_),
    .A1(net371),
    .A2(net193));
 sg13g2_nand2_1 _09293_ (.Y(_01920_),
    .A(net2971),
    .B(net193));
 sg13g2_o21ai_1 _09294_ (.B1(_01920_),
    .Y(_00932_),
    .A1(net368),
    .A2(net194));
 sg13g2_nand2_1 _09295_ (.Y(_01921_),
    .A(net2914),
    .B(net193));
 sg13g2_o21ai_1 _09296_ (.B1(_01921_),
    .Y(_00931_),
    .A1(net359),
    .A2(net193));
 sg13g2_nand2_1 _09297_ (.Y(_01922_),
    .A(net2877),
    .B(net195));
 sg13g2_o21ai_1 _09298_ (.B1(_01922_),
    .Y(_00930_),
    .A1(net358),
    .A2(net195));
 sg13g2_nor2_2 _09299_ (.A(net319),
    .B(_01852_),
    .Y(_01923_));
 sg13g2_nor3_1 _09300_ (.A(_01711_),
    .B(_01723_),
    .C(_01852_),
    .Y(_01924_));
 sg13g2_nor2_1 _09301_ (.A(net3400),
    .B(net241),
    .Y(_01925_));
 sg13g2_a21oi_1 _09302_ (.A1(net396),
    .A2(net241),
    .Y(_00929_),
    .B1(_01925_));
 sg13g2_nor2_1 _09303_ (.A(net3046),
    .B(net241),
    .Y(_01926_));
 sg13g2_a21oi_1 _09304_ (.A1(net389),
    .A2(net241),
    .Y(_00928_),
    .B1(_01926_));
 sg13g2_nor2_1 _09305_ (.A(net3214),
    .B(net241),
    .Y(_01927_));
 sg13g2_a21oi_1 _09306_ (.A1(net384),
    .A2(net241),
    .Y(_00927_),
    .B1(_01927_));
 sg13g2_nor2_1 _09307_ (.A(net3196),
    .B(net240),
    .Y(_01928_));
 sg13g2_a21oi_1 _09308_ (.A1(net377),
    .A2(net240),
    .Y(_00926_),
    .B1(_01928_));
 sg13g2_nor2_1 _09309_ (.A(net3173),
    .B(net241),
    .Y(_01929_));
 sg13g2_a21oi_1 _09310_ (.A1(_01751_),
    .A2(net241),
    .Y(_00925_),
    .B1(_01929_));
 sg13g2_nor2_1 _09311_ (.A(net3152),
    .B(net240),
    .Y(_01930_));
 sg13g2_a21oi_1 _09312_ (.A1(net368),
    .A2(net240),
    .Y(_00924_),
    .B1(_01930_));
 sg13g2_nor2_1 _09313_ (.A(net3113),
    .B(net240),
    .Y(_01931_));
 sg13g2_a21oi_1 _09314_ (.A1(net364),
    .A2(net240),
    .Y(_00923_),
    .B1(_01931_));
 sg13g2_nor2_1 _09315_ (.A(net3223),
    .B(net240),
    .Y(_01932_));
 sg13g2_a21oi_1 _09316_ (.A1(_01763_),
    .A2(net240),
    .Y(_00922_),
    .B1(_01932_));
 sg13g2_nor3_2 _09317_ (.A(_01721_),
    .B(net319),
    .C(_01766_),
    .Y(_01933_));
 sg13g2_and2_1 _09318_ (.A(net424),
    .B(net239),
    .X(_01934_));
 sg13g2_nor2_1 _09319_ (.A(net3100),
    .B(net141),
    .Y(_01935_));
 sg13g2_a21oi_1 _09320_ (.A1(net391),
    .A2(net141),
    .Y(_00921_),
    .B1(_01935_));
 sg13g2_nor2_1 _09321_ (.A(net3149),
    .B(net141),
    .Y(_01936_));
 sg13g2_a21oi_1 _09322_ (.A1(net385),
    .A2(net141),
    .Y(_00920_),
    .B1(_01936_));
 sg13g2_nor2_1 _09323_ (.A(net3193),
    .B(net142),
    .Y(_01937_));
 sg13g2_a21oi_1 _09324_ (.A1(net380),
    .A2(net142),
    .Y(_00919_),
    .B1(_01937_));
 sg13g2_nor2_1 _09325_ (.A(net3052),
    .B(net142),
    .Y(_01938_));
 sg13g2_a21oi_1 _09326_ (.A1(net376),
    .A2(net142),
    .Y(_00918_),
    .B1(_01938_));
 sg13g2_nor2_1 _09327_ (.A(net3187),
    .B(_01934_),
    .Y(_01939_));
 sg13g2_a21oi_1 _09328_ (.A1(net370),
    .A2(net142),
    .Y(_00917_),
    .B1(_01939_));
 sg13g2_nor2_1 _09329_ (.A(net3242),
    .B(net142),
    .Y(_01940_));
 sg13g2_a21oi_1 _09330_ (.A1(net366),
    .A2(net142),
    .Y(_00916_),
    .B1(_01940_));
 sg13g2_nor2_1 _09331_ (.A(net3116),
    .B(net141),
    .Y(_01941_));
 sg13g2_a21oi_1 _09332_ (.A1(net360),
    .A2(net141),
    .Y(_00915_),
    .B1(_01941_));
 sg13g2_nor2_1 _09333_ (.A(net3051),
    .B(net141),
    .Y(_01942_));
 sg13g2_a21oi_1 _09334_ (.A1(net356),
    .A2(net141),
    .Y(_00914_),
    .B1(_01942_));
 sg13g2_nor3_2 _09335_ (.A(_01721_),
    .B(net319),
    .C(_01820_),
    .Y(_01943_));
 sg13g2_and2_1 _09336_ (.A(net422),
    .B(net238),
    .X(_01944_));
 sg13g2_nor2_1 _09337_ (.A(net3053),
    .B(net140),
    .Y(_01945_));
 sg13g2_a21oi_1 _09338_ (.A1(net392),
    .A2(net140),
    .Y(_00913_),
    .B1(_01945_));
 sg13g2_nor2_1 _09339_ (.A(net3115),
    .B(net139),
    .Y(_01946_));
 sg13g2_a21oi_1 _09340_ (.A1(net385),
    .A2(net139),
    .Y(_00912_),
    .B1(_01946_));
 sg13g2_nor2_1 _09341_ (.A(net3022),
    .B(net139),
    .Y(_01947_));
 sg13g2_a21oi_1 _09342_ (.A1(net382),
    .A2(net139),
    .Y(_00911_),
    .B1(_01947_));
 sg13g2_nor2_1 _09343_ (.A(net3305),
    .B(net140),
    .Y(_01948_));
 sg13g2_a21oi_1 _09344_ (.A1(net375),
    .A2(net140),
    .Y(_00910_),
    .B1(_01948_));
 sg13g2_nor2_1 _09345_ (.A(net3209),
    .B(net140),
    .Y(_01949_));
 sg13g2_a21oi_1 _09346_ (.A1(net373),
    .A2(net140),
    .Y(_00909_),
    .B1(_01949_));
 sg13g2_nor2_1 _09347_ (.A(net3233),
    .B(net139),
    .Y(_01950_));
 sg13g2_a21oi_1 _09348_ (.A1(net367),
    .A2(net139),
    .Y(_00908_),
    .B1(_01950_));
 sg13g2_nor2_1 _09349_ (.A(net3137),
    .B(net140),
    .Y(_01951_));
 sg13g2_a21oi_1 _09350_ (.A1(net360),
    .A2(net140),
    .Y(_00907_),
    .B1(_01951_));
 sg13g2_nor2_1 _09351_ (.A(net3048),
    .B(net139),
    .Y(_01952_));
 sg13g2_a21oi_1 _09352_ (.A1(net356),
    .A2(net139),
    .Y(_00906_),
    .B1(_01952_));
 sg13g2_nor3_2 _09353_ (.A(_01721_),
    .B(net317),
    .C(_01766_),
    .Y(_01953_));
 sg13g2_and2_1 _09354_ (.A(net423),
    .B(net237),
    .X(_01954_));
 sg13g2_nor2_1 _09355_ (.A(net3105),
    .B(net191),
    .Y(_01955_));
 sg13g2_a21oi_1 _09356_ (.A1(net392),
    .A2(net191),
    .Y(_00905_),
    .B1(_01955_));
 sg13g2_nor2_1 _09357_ (.A(net3260),
    .B(net192),
    .Y(_01956_));
 sg13g2_a21oi_1 _09358_ (.A1(net386),
    .A2(net192),
    .Y(_00904_),
    .B1(_01956_));
 sg13g2_nor2_1 _09359_ (.A(net3456),
    .B(net191),
    .Y(_01957_));
 sg13g2_a21oi_1 _09360_ (.A1(net384),
    .A2(net191),
    .Y(_00903_),
    .B1(_01957_));
 sg13g2_nor2_1 _09361_ (.A(net3104),
    .B(net192),
    .Y(_01958_));
 sg13g2_a21oi_1 _09362_ (.A1(net375),
    .A2(_01954_),
    .Y(_00902_),
    .B1(_01958_));
 sg13g2_nor2_1 _09363_ (.A(net3042),
    .B(net192),
    .Y(_01959_));
 sg13g2_a21oi_1 _09364_ (.A1(net372),
    .A2(net192),
    .Y(_00901_),
    .B1(_01959_));
 sg13g2_nor2_1 _09365_ (.A(net3316),
    .B(net191),
    .Y(_01960_));
 sg13g2_a21oi_1 _09366_ (.A1(net367),
    .A2(net191),
    .Y(_00900_),
    .B1(_01960_));
 sg13g2_nor2_1 _09367_ (.A(net3131),
    .B(net191),
    .Y(_01961_));
 sg13g2_a21oi_1 _09368_ (.A1(net360),
    .A2(net191),
    .Y(_00899_),
    .B1(_01961_));
 sg13g2_nor2_1 _09369_ (.A(net3132),
    .B(net192),
    .Y(_01962_));
 sg13g2_a21oi_1 _09370_ (.A1(net357),
    .A2(net192),
    .Y(_00898_),
    .B1(_01962_));
 sg13g2_nor3_2 _09371_ (.A(net320),
    .B(_01798_),
    .C(_01799_),
    .Y(_01963_));
 sg13g2_and2_1 _09372_ (.A(net424),
    .B(net236),
    .X(_01964_));
 sg13g2_nor2_1 _09373_ (.A(net3597),
    .B(net137),
    .Y(_01965_));
 sg13g2_a21oi_1 _09374_ (.A1(net393),
    .A2(net137),
    .Y(_00897_),
    .B1(_01965_));
 sg13g2_nor2_1 _09375_ (.A(net3160),
    .B(net138),
    .Y(_01966_));
 sg13g2_a21oi_1 _09376_ (.A1(net387),
    .A2(net138),
    .Y(_00896_),
    .B1(_01966_));
 sg13g2_nor2_1 _09377_ (.A(net3287),
    .B(net138),
    .Y(_01967_));
 sg13g2_a21oi_1 _09378_ (.A1(net380),
    .A2(net138),
    .Y(_00895_),
    .B1(_01967_));
 sg13g2_nor2_1 _09379_ (.A(net3467),
    .B(net138),
    .Y(_01968_));
 sg13g2_a21oi_1 _09380_ (.A1(net376),
    .A2(net138),
    .Y(_00894_),
    .B1(_01968_));
 sg13g2_nor2_1 _09381_ (.A(net3065),
    .B(net137),
    .Y(_01969_));
 sg13g2_a21oi_1 _09382_ (.A1(net370),
    .A2(net137),
    .Y(_00893_),
    .B1(_01969_));
 sg13g2_nor2_1 _09383_ (.A(net3282),
    .B(net137),
    .Y(_01970_));
 sg13g2_a21oi_1 _09384_ (.A1(net365),
    .A2(net137),
    .Y(_00892_),
    .B1(_01970_));
 sg13g2_nor2_1 _09385_ (.A(net3114),
    .B(net137),
    .Y(_01971_));
 sg13g2_a21oi_1 _09386_ (.A1(net359),
    .A2(net137),
    .Y(_00891_),
    .B1(_01971_));
 sg13g2_nor2_1 _09387_ (.A(net3226),
    .B(net138),
    .Y(_01972_));
 sg13g2_a21oi_1 _09388_ (.A1(net354),
    .A2(_01964_),
    .Y(_00890_),
    .B1(_01972_));
 sg13g2_nor3_2 _09389_ (.A(net320),
    .B(_01766_),
    .C(_01799_),
    .Y(_01973_));
 sg13g2_and2_2 _09390_ (.A(net425),
    .B(net235),
    .X(_01974_));
 sg13g2_nor2_1 _09391_ (.A(net3012),
    .B(net189),
    .Y(_01975_));
 sg13g2_a21oi_1 _09392_ (.A1(net393),
    .A2(net189),
    .Y(_00889_),
    .B1(_01975_));
 sg13g2_nor2_1 _09393_ (.A(net3101),
    .B(net190),
    .Y(_01976_));
 sg13g2_a21oi_1 _09394_ (.A1(net388),
    .A2(net190),
    .Y(_00888_),
    .B1(_01976_));
 sg13g2_nor2_1 _09395_ (.A(net3088),
    .B(net190),
    .Y(_01977_));
 sg13g2_a21oi_1 _09396_ (.A1(net383),
    .A2(net190),
    .Y(_00887_),
    .B1(_01977_));
 sg13g2_nor2_1 _09397_ (.A(net3083),
    .B(net189),
    .Y(_01978_));
 sg13g2_a21oi_1 _09398_ (.A1(net376),
    .A2(net189),
    .Y(_00886_),
    .B1(_01978_));
 sg13g2_nor2_1 _09399_ (.A(net3091),
    .B(net190),
    .Y(_01979_));
 sg13g2_a21oi_1 _09400_ (.A1(net373),
    .A2(net190),
    .Y(_00885_),
    .B1(_01979_));
 sg13g2_nor2_1 _09401_ (.A(net3202),
    .B(net189),
    .Y(_01980_));
 sg13g2_a21oi_1 _09402_ (.A1(net365),
    .A2(net189),
    .Y(_00884_),
    .B1(_01980_));
 sg13g2_nor2_1 _09403_ (.A(net3552),
    .B(net189),
    .Y(_01981_));
 sg13g2_a21oi_1 _09404_ (.A1(net359),
    .A2(net189),
    .Y(_00883_),
    .B1(_01981_));
 sg13g2_nor2_1 _09405_ (.A(net3345),
    .B(net190),
    .Y(_01982_));
 sg13g2_a21oi_1 _09406_ (.A1(net358),
    .A2(net190),
    .Y(_00882_),
    .B1(_01982_));
 sg13g2_nor3_2 _09407_ (.A(net320),
    .B(_01799_),
    .C(_01820_),
    .Y(_01983_));
 sg13g2_and2_1 _09408_ (.A(net425),
    .B(net234),
    .X(_01984_));
 sg13g2_nor2_1 _09409_ (.A(net3324),
    .B(net136),
    .Y(_01985_));
 sg13g2_a21oi_1 _09410_ (.A1(net395),
    .A2(net136),
    .Y(_00881_),
    .B1(_01985_));
 sg13g2_nor2_1 _09411_ (.A(net3205),
    .B(net135),
    .Y(_01986_));
 sg13g2_a21oi_1 _09412_ (.A1(net388),
    .A2(net135),
    .Y(_00880_),
    .B1(_01986_));
 sg13g2_nor2_1 _09413_ (.A(net3072),
    .B(net136),
    .Y(_01987_));
 sg13g2_a21oi_1 _09414_ (.A1(net383),
    .A2(net136),
    .Y(_00879_),
    .B1(_01987_));
 sg13g2_nor2_1 _09415_ (.A(net3277),
    .B(net136),
    .Y(_01988_));
 sg13g2_a21oi_1 _09416_ (.A1(net378),
    .A2(net136),
    .Y(_00878_),
    .B1(_01988_));
 sg13g2_nor2_1 _09417_ (.A(net3311),
    .B(net135),
    .Y(_01989_));
 sg13g2_a21oi_1 _09418_ (.A1(net373),
    .A2(net135),
    .Y(_00877_),
    .B1(_01989_));
 sg13g2_nor2_1 _09419_ (.A(net3237),
    .B(net135),
    .Y(_01990_));
 sg13g2_a21oi_1 _09420_ (.A1(net369),
    .A2(net135),
    .Y(_00876_),
    .B1(_01990_));
 sg13g2_nor2_1 _09421_ (.A(net3141),
    .B(net135),
    .Y(_01991_));
 sg13g2_a21oi_1 _09422_ (.A1(net363),
    .A2(net135),
    .Y(_00875_),
    .B1(_01991_));
 sg13g2_nor2_1 _09423_ (.A(net3134),
    .B(net136),
    .Y(_01992_));
 sg13g2_a21oi_1 _09424_ (.A1(net358),
    .A2(net136),
    .Y(_00874_),
    .B1(_01992_));
 sg13g2_nor3_2 _09425_ (.A(_01715_),
    .B(net320),
    .C(_01799_),
    .Y(_01993_));
 sg13g2_and2_1 _09426_ (.A(net426),
    .B(net233),
    .X(_01994_));
 sg13g2_nor2_1 _09427_ (.A(net3328),
    .B(net134),
    .Y(_01995_));
 sg13g2_a21oi_1 _09428_ (.A1(net395),
    .A2(_01994_),
    .Y(_00873_),
    .B1(_01995_));
 sg13g2_nor2_1 _09429_ (.A(net3422),
    .B(net133),
    .Y(_01996_));
 sg13g2_a21oi_1 _09430_ (.A1(net389),
    .A2(net133),
    .Y(_00872_),
    .B1(_01996_));
 sg13g2_nor2_1 _09431_ (.A(net3191),
    .B(net133),
    .Y(_01997_));
 sg13g2_a21oi_1 _09432_ (.A1(net383),
    .A2(net133),
    .Y(_00871_),
    .B1(_01997_));
 sg13g2_nor2_1 _09433_ (.A(net3362),
    .B(net134),
    .Y(_01998_));
 sg13g2_a21oi_1 _09434_ (.A1(net378),
    .A2(net134),
    .Y(_00870_),
    .B1(_01998_));
 sg13g2_nor2_1 _09435_ (.A(net3262),
    .B(net133),
    .Y(_01999_));
 sg13g2_a21oi_1 _09436_ (.A1(_01751_),
    .A2(net133),
    .Y(_00869_),
    .B1(_01999_));
 sg13g2_nor2_1 _09437_ (.A(net3414),
    .B(net133),
    .Y(_02000_));
 sg13g2_a21oi_1 _09438_ (.A1(net369),
    .A2(net133),
    .Y(_00868_),
    .B1(_02000_));
 sg13g2_nor2_1 _09439_ (.A(net3296),
    .B(net134),
    .Y(_02001_));
 sg13g2_a21oi_1 _09440_ (.A1(net363),
    .A2(net134),
    .Y(_00867_),
    .B1(_02001_));
 sg13g2_nor2_1 _09441_ (.A(net3315),
    .B(net134),
    .Y(_02002_));
 sg13g2_a21oi_1 _09442_ (.A1(net358),
    .A2(net134),
    .Y(_00866_),
    .B1(_02002_));
 sg13g2_nor3_2 _09443_ (.A(net319),
    .B(_01798_),
    .C(_01841_),
    .Y(_02003_));
 sg13g2_nand2_1 _09444_ (.Y(_02004_),
    .A(net422),
    .B(net232));
 sg13g2_nand2_1 _09445_ (.Y(_02005_),
    .A(net2990),
    .B(net132));
 sg13g2_o21ai_1 _09446_ (.B1(_02005_),
    .Y(_00865_),
    .A1(net391),
    .A2(_02004_));
 sg13g2_nand2_1 _09447_ (.Y(_02006_),
    .A(net2955),
    .B(net132));
 sg13g2_o21ai_1 _09448_ (.B1(_02006_),
    .Y(_00864_),
    .A1(net385),
    .A2(net132));
 sg13g2_nand2_1 _09449_ (.Y(_02007_),
    .A(net2871),
    .B(net131));
 sg13g2_o21ai_1 _09450_ (.B1(_02007_),
    .Y(_00863_),
    .A1(net380),
    .A2(net131));
 sg13g2_nand2_1 _09451_ (.Y(_02008_),
    .A(net2995),
    .B(net131));
 sg13g2_o21ai_1 _09452_ (.B1(_02008_),
    .Y(_00862_),
    .A1(net376),
    .A2(net131));
 sg13g2_nand2_1 _09453_ (.Y(_02009_),
    .A(net2960),
    .B(net132));
 sg13g2_o21ai_1 _09454_ (.B1(_02009_),
    .Y(_00861_),
    .A1(net370),
    .A2(net132));
 sg13g2_nand2_1 _09455_ (.Y(_02010_),
    .A(net2976),
    .B(net131));
 sg13g2_o21ai_1 _09456_ (.B1(_02010_),
    .Y(_00860_),
    .A1(net365),
    .A2(net131));
 sg13g2_nand2_1 _09457_ (.Y(_02011_),
    .A(net3201),
    .B(net131));
 sg13g2_o21ai_1 _09458_ (.B1(_02011_),
    .Y(_00859_),
    .A1(net359),
    .A2(net131));
 sg13g2_nand2_1 _09459_ (.Y(_02012_),
    .A(net2864),
    .B(net132));
 sg13g2_o21ai_1 _09460_ (.B1(_02012_),
    .Y(_00858_),
    .A1(net356),
    .A2(net132));
 sg13g2_nor3_2 _09461_ (.A(net319),
    .B(_01766_),
    .C(_01841_),
    .Y(_02013_));
 sg13g2_nand2_1 _09462_ (.Y(_02014_),
    .A(net422),
    .B(net231));
 sg13g2_nand2_1 _09463_ (.Y(_02015_),
    .A(net2965),
    .B(net129));
 sg13g2_o21ai_1 _09464_ (.B1(_02015_),
    .Y(_00857_),
    .A1(net391),
    .A2(net130));
 sg13g2_nand2_1 _09465_ (.Y(_02016_),
    .A(net3274),
    .B(net129));
 sg13g2_o21ai_1 _09466_ (.B1(_02016_),
    .Y(_00856_),
    .A1(net385),
    .A2(net129));
 sg13g2_nand2_1 _09467_ (.Y(_02017_),
    .A(net2954),
    .B(net129));
 sg13g2_o21ai_1 _09468_ (.B1(_02017_),
    .Y(_00855_),
    .A1(net382),
    .A2(net129));
 sg13g2_nand2_1 _09469_ (.Y(_02018_),
    .A(net3227),
    .B(net130));
 sg13g2_o21ai_1 _09470_ (.B1(_02018_),
    .Y(_00854_),
    .A1(net374),
    .A2(net130));
 sg13g2_nand2_1 _09471_ (.Y(_02019_),
    .A(net2883),
    .B(net129));
 sg13g2_o21ai_1 _09472_ (.B1(_02019_),
    .Y(_00853_),
    .A1(net372),
    .A2(_02014_));
 sg13g2_nand2_1 _09473_ (.Y(_02020_),
    .A(net2891),
    .B(net130));
 sg13g2_o21ai_1 _09474_ (.B1(_02020_),
    .Y(_00852_),
    .A1(net367),
    .A2(net130));
 sg13g2_nand2_1 _09475_ (.Y(_02021_),
    .A(net2923),
    .B(net130));
 sg13g2_o21ai_1 _09476_ (.B1(_02021_),
    .Y(_00851_),
    .A1(net360),
    .A2(net130));
 sg13g2_nand2_1 _09477_ (.Y(_02022_),
    .A(net2894),
    .B(net129));
 sg13g2_o21ai_1 _09478_ (.B1(_02022_),
    .Y(_00850_),
    .A1(net356),
    .A2(net129));
 sg13g2_nor3_2 _09479_ (.A(net319),
    .B(_01820_),
    .C(_01841_),
    .Y(_02023_));
 sg13g2_nand2_1 _09480_ (.Y(_02024_),
    .A(net422),
    .B(_02023_));
 sg13g2_nand2_1 _09481_ (.Y(_02025_),
    .A(net2932),
    .B(net128));
 sg13g2_o21ai_1 _09482_ (.B1(_02025_),
    .Y(_00849_),
    .A1(net392),
    .A2(net128));
 sg13g2_nand2_1 _09483_ (.Y(_02026_),
    .A(net2987),
    .B(net127));
 sg13g2_o21ai_1 _09484_ (.B1(_02026_),
    .Y(_00848_),
    .A1(net385),
    .A2(net127));
 sg13g2_nand2_1 _09485_ (.Y(_02027_),
    .A(net2969),
    .B(net128));
 sg13g2_o21ai_1 _09486_ (.B1(_02027_),
    .Y(_00847_),
    .A1(net382),
    .A2(net128));
 sg13g2_nand2_1 _09487_ (.Y(_02028_),
    .A(net2940),
    .B(net128));
 sg13g2_o21ai_1 _09488_ (.B1(_02028_),
    .Y(_00846_),
    .A1(net374),
    .A2(_02024_));
 sg13g2_nand2_1 _09489_ (.Y(_02029_),
    .A(net2904),
    .B(net128));
 sg13g2_o21ai_1 _09490_ (.B1(_02029_),
    .Y(_00845_),
    .A1(net372),
    .A2(net128));
 sg13g2_nand2_1 _09491_ (.Y(_02030_),
    .A(net2964),
    .B(net127));
 sg13g2_o21ai_1 _09492_ (.B1(_02030_),
    .Y(_00844_),
    .A1(net367),
    .A2(net127));
 sg13g2_nand2_1 _09493_ (.Y(_02031_),
    .A(net3130),
    .B(net127));
 sg13g2_o21ai_1 _09494_ (.B1(_02031_),
    .Y(_00843_),
    .A1(net360),
    .A2(net127));
 sg13g2_nand2_1 _09495_ (.Y(_02032_),
    .A(net2874),
    .B(net127));
 sg13g2_o21ai_1 _09496_ (.B1(_02032_),
    .Y(_00842_),
    .A1(net356),
    .A2(net127));
 sg13g2_nor3_2 _09497_ (.A(_01715_),
    .B(net319),
    .C(_01841_),
    .Y(_02033_));
 sg13g2_nand2_1 _09498_ (.Y(_02034_),
    .A(net422),
    .B(net229));
 sg13g2_nand2_1 _09499_ (.Y(_02035_),
    .A(net2967),
    .B(_02034_));
 sg13g2_o21ai_1 _09500_ (.B1(_02035_),
    .Y(_00841_),
    .A1(net392),
    .A2(net126));
 sg13g2_nand2_1 _09501_ (.Y(_02036_),
    .A(net2927),
    .B(net125));
 sg13g2_o21ai_1 _09502_ (.B1(_02036_),
    .Y(_00840_),
    .A1(net385),
    .A2(net125));
 sg13g2_nand2_1 _09503_ (.Y(_02037_),
    .A(net3215),
    .B(net126));
 sg13g2_o21ai_1 _09504_ (.B1(_02037_),
    .Y(_00839_),
    .A1(net382),
    .A2(net126));
 sg13g2_nand2_1 _09505_ (.Y(_02038_),
    .A(net2982),
    .B(net125));
 sg13g2_o21ai_1 _09506_ (.B1(_02038_),
    .Y(_00838_),
    .A1(net374),
    .A2(net125));
 sg13g2_nand2_1 _09507_ (.Y(_02039_),
    .A(net3081),
    .B(net125));
 sg13g2_o21ai_1 _09508_ (.B1(_02039_),
    .Y(_00837_),
    .A1(net372),
    .A2(net125));
 sg13g2_nand2_1 _09509_ (.Y(_02040_),
    .A(net2919),
    .B(net125));
 sg13g2_o21ai_1 _09510_ (.B1(_02040_),
    .Y(_00836_),
    .A1(net367),
    .A2(net125));
 sg13g2_nand2_1 _09511_ (.Y(_02041_),
    .A(net3272),
    .B(net126));
 sg13g2_o21ai_1 _09512_ (.B1(_02041_),
    .Y(_00835_),
    .A1(net360),
    .A2(net126));
 sg13g2_nand2_1 _09513_ (.Y(_02042_),
    .A(net3007),
    .B(net126));
 sg13g2_o21ai_1 _09514_ (.B1(_02042_),
    .Y(_00834_),
    .A1(net356),
    .A2(net126));
 sg13g2_nor3_2 _09515_ (.A(net320),
    .B(_01765_),
    .C(_01798_),
    .Y(_02043_));
 sg13g2_nand2_1 _09516_ (.Y(_02044_),
    .A(net425),
    .B(net228));
 sg13g2_nand2_1 _09517_ (.Y(_02045_),
    .A(net2970),
    .B(net188));
 sg13g2_o21ai_1 _09518_ (.B1(_02045_),
    .Y(_00833_),
    .A1(net394),
    .A2(net188));
 sg13g2_nand2_1 _09519_ (.Y(_02046_),
    .A(net2939),
    .B(net188));
 sg13g2_o21ai_1 _09520_ (.B1(_02046_),
    .Y(_00832_),
    .A1(net388),
    .A2(net188));
 sg13g2_nand2_1 _09521_ (.Y(_02047_),
    .A(net2963),
    .B(net188));
 sg13g2_o21ai_1 _09522_ (.B1(_02047_),
    .Y(_00831_),
    .A1(net383),
    .A2(net188));
 sg13g2_nand2_1 _09523_ (.Y(_02048_),
    .A(net2917),
    .B(net188));
 sg13g2_o21ai_1 _09524_ (.B1(_02048_),
    .Y(_00830_),
    .A1(net377),
    .A2(net188));
 sg13g2_nand2_1 _09525_ (.Y(_02049_),
    .A(net2936),
    .B(net187));
 sg13g2_o21ai_1 _09526_ (.B1(_02049_),
    .Y(_00829_),
    .A1(net371),
    .A2(net187));
 sg13g2_nand2_1 _09527_ (.Y(_02050_),
    .A(net2941),
    .B(net187));
 sg13g2_o21ai_1 _09528_ (.B1(_02050_),
    .Y(_00828_),
    .A1(net368),
    .A2(net187));
 sg13g2_nand2_1 _09529_ (.Y(_02051_),
    .A(net2885),
    .B(net187));
 sg13g2_o21ai_1 _09530_ (.B1(_02051_),
    .Y(_00827_),
    .A1(net362),
    .A2(net187));
 sg13g2_nand2_1 _09531_ (.Y(_02052_),
    .A(net2901),
    .B(net187));
 sg13g2_o21ai_1 _09532_ (.B1(_02052_),
    .Y(_00826_),
    .A1(net354),
    .A2(net187));
 sg13g2_nor3_2 _09533_ (.A(_01721_),
    .B(net317),
    .C(_01820_),
    .Y(_02053_));
 sg13g2_and2_1 _09534_ (.A(net422),
    .B(net227),
    .X(_02054_));
 sg13g2_nor2_1 _09535_ (.A(net3082),
    .B(net123),
    .Y(_02055_));
 sg13g2_a21oi_1 _09536_ (.A1(net391),
    .A2(net123),
    .Y(_00825_),
    .B1(_02055_));
 sg13g2_nor2_1 _09537_ (.A(net3294),
    .B(net123),
    .Y(_02056_));
 sg13g2_a21oi_1 _09538_ (.A1(net386),
    .A2(net123),
    .Y(_00824_),
    .B1(_02056_));
 sg13g2_nor2_1 _09539_ (.A(net3164),
    .B(net123),
    .Y(_02057_));
 sg13g2_a21oi_1 _09540_ (.A1(net382),
    .A2(net123),
    .Y(_00823_),
    .B1(_02057_));
 sg13g2_nor2_1 _09541_ (.A(net3234),
    .B(net124),
    .Y(_02058_));
 sg13g2_a21oi_1 _09542_ (.A1(net374),
    .A2(net124),
    .Y(_00822_),
    .B1(_02058_));
 sg13g2_nor2_1 _09543_ (.A(net3120),
    .B(net124),
    .Y(_02059_));
 sg13g2_a21oi_1 _09544_ (.A1(net373),
    .A2(net124),
    .Y(_00821_),
    .B1(_02059_));
 sg13g2_nor2_1 _09545_ (.A(net3204),
    .B(net124),
    .Y(_02060_));
 sg13g2_a21oi_1 _09546_ (.A1(_01755_),
    .A2(net124),
    .Y(_00820_),
    .B1(_02060_));
 sg13g2_nor2_1 _09547_ (.A(net3236),
    .B(net124),
    .Y(_02061_));
 sg13g2_a21oi_1 _09548_ (.A1(net361),
    .A2(net124),
    .Y(_00819_),
    .B1(_02061_));
 sg13g2_nor2_1 _09549_ (.A(net3175),
    .B(net123),
    .Y(_02062_));
 sg13g2_a21oi_1 _09550_ (.A1(net356),
    .A2(net123),
    .Y(_00818_),
    .B1(_02062_));
 sg13g2_nor3_2 _09551_ (.A(net320),
    .B(_01765_),
    .C(_01820_),
    .Y(_02063_));
 sg13g2_nand2_1 _09552_ (.Y(_02064_),
    .A(net426),
    .B(net226));
 sg13g2_nand2_1 _09553_ (.Y(_02065_),
    .A(net2893),
    .B(net186));
 sg13g2_o21ai_1 _09554_ (.B1(_02065_),
    .Y(_00817_),
    .A1(net394),
    .A2(net186));
 sg13g2_nand2_1 _09555_ (.Y(_02066_),
    .A(net2884),
    .B(net185));
 sg13g2_o21ai_1 _09556_ (.B1(_02066_),
    .Y(_00816_),
    .A1(net388),
    .A2(net185));
 sg13g2_nand2_1 _09557_ (.Y(_02067_),
    .A(net2952),
    .B(net185));
 sg13g2_o21ai_1 _09558_ (.B1(_02067_),
    .Y(_00815_),
    .A1(net383),
    .A2(net185));
 sg13g2_nand2_1 _09559_ (.Y(_02068_),
    .A(net2944),
    .B(net186));
 sg13g2_o21ai_1 _09560_ (.B1(_02068_),
    .Y(_00814_),
    .A1(net377),
    .A2(net186));
 sg13g2_nand2_1 _09561_ (.Y(_02069_),
    .A(net2889),
    .B(net185));
 sg13g2_o21ai_1 _09562_ (.B1(_02069_),
    .Y(_00813_),
    .A1(net373),
    .A2(net186));
 sg13g2_nand2_1 _09563_ (.Y(_02070_),
    .A(net2878),
    .B(net186));
 sg13g2_o21ai_1 _09564_ (.B1(_02070_),
    .Y(_00812_),
    .A1(net368),
    .A2(net186));
 sg13g2_nand2_1 _09565_ (.Y(_02071_),
    .A(net2862),
    .B(net185));
 sg13g2_o21ai_1 _09566_ (.B1(_02071_),
    .Y(_00811_),
    .A1(net363),
    .A2(net185));
 sg13g2_nand2_1 _09567_ (.Y(_02072_),
    .A(net2866),
    .B(_02064_));
 sg13g2_o21ai_1 _09568_ (.B1(_02072_),
    .Y(_00810_),
    .A1(net358),
    .A2(net185));
 sg13g2_nand2b_1 _09569_ (.Y(_00808_),
    .B(net526),
    .A_N(\i_game.game_latch_sync[1] ));
 sg13g2_nor2_1 _09570_ (.A(net637),
    .B(\addr[25] ),
    .Y(_02073_));
 sg13g2_and2_1 _09571_ (.A(_00191_),
    .B(_02073_),
    .X(_02074_));
 sg13g2_nand2_2 _09572_ (.Y(_02075_),
    .A(_00191_),
    .B(_02073_));
 sg13g2_and2_2 _09573_ (.A(_01709_),
    .B(net417),
    .X(_02076_));
 sg13g2_nand2_2 _09574_ (.Y(_02077_),
    .A(_01709_),
    .B(_02075_));
 sg13g2_nor2b_2 _09575_ (.A(\addr[4] ),
    .B_N(\addr[5] ),
    .Y(_02078_));
 sg13g2_nor4_1 _09576_ (.A(_00191_),
    .B(net2380),
    .C(\addr[8] ),
    .D(\addr[7] ),
    .Y(_02079_));
 sg13g2_nor4_1 _09577_ (.A(net637),
    .B(\addr[25] ),
    .C(\addr[24] ),
    .D(net2387),
    .Y(_02080_));
 sg13g2_nor3_1 _09578_ (.A(\addr[22] ),
    .B(\addr[21] ),
    .C(\addr[23] ),
    .Y(_02081_));
 sg13g2_nor4_1 _09579_ (.A(\addr[18] ),
    .B(\addr[17] ),
    .C(\addr[20] ),
    .D(\addr[19] ),
    .Y(_02082_));
 sg13g2_nand2_2 _09580_ (.Y(_02083_),
    .A(_02081_),
    .B(_02082_));
 sg13g2_nor4_2 _09581_ (.A(\addr[14] ),
    .B(\addr[13] ),
    .C(\addr[16] ),
    .Y(_02084_),
    .D(\addr[15] ));
 sg13g2_nor4_2 _09582_ (.A(\addr[10] ),
    .B(\addr[9] ),
    .C(\addr[12] ),
    .Y(_02085_),
    .D(\addr[11] ));
 sg13g2_nand4_1 _09583_ (.B(_02079_),
    .C(_02084_),
    .A(_02080_),
    .Y(_02086_),
    .D(_02085_));
 sg13g2_nor2_1 _09584_ (.A(_02083_),
    .B(net2381),
    .Y(_02087_));
 sg13g2_and2_1 _09585_ (.A(_00198_),
    .B(_02087_),
    .X(_02088_));
 sg13g2_nand2_1 _09586_ (.Y(_02089_),
    .A(_00198_),
    .B(_02087_));
 sg13g2_nor2b_1 _09587_ (.A(\addr[6] ),
    .B_N(net633),
    .Y(_02090_));
 sg13g2_nand2_1 _09588_ (.Y(_02091_),
    .A(net633),
    .B(_02088_));
 sg13g2_nor2_2 _09589_ (.A(\addr[6] ),
    .B(_02091_),
    .Y(_02092_));
 sg13g2_inv_1 _09590_ (.Y(_02093_),
    .A(_02092_));
 sg13g2_and2_1 _09591_ (.A(_02078_),
    .B(_02092_),
    .X(_02094_));
 sg13g2_nor3_1 _09592_ (.A(\addr[6] ),
    .B(_02083_),
    .C(net2381),
    .Y(_02095_));
 sg13g2_nand2_1 _09593_ (.Y(_02096_),
    .A(net632),
    .B(_02095_));
 sg13g2_a21oi_2 _09594_ (.B1(net516),
    .Y(_02097_),
    .A2(_02094_),
    .A1(_02076_));
 sg13g2_nand2_1 _09595_ (.Y(_02098_),
    .A(net3146),
    .B(net184));
 sg13g2_o21ai_1 _09596_ (.B1(_02098_),
    .Y(_00773_),
    .A1(_01508_),
    .A2(net184));
 sg13g2_nand2_1 _09597_ (.Y(_02099_),
    .A(net3075),
    .B(net184));
 sg13g2_o21ai_1 _09598_ (.B1(_02099_),
    .Y(_00772_),
    .A1(_01509_),
    .A2(net184));
 sg13g2_nand2_1 _09599_ (.Y(_02100_),
    .A(net3095),
    .B(net184));
 sg13g2_o21ai_1 _09600_ (.B1(_02100_),
    .Y(_00771_),
    .A1(_01510_),
    .A2(net184));
 sg13g2_nand2_1 _09601_ (.Y(_02101_),
    .A(net3008),
    .B(net184));
 sg13g2_o21ai_1 _09602_ (.B1(_02101_),
    .Y(_00770_),
    .A1(_01511_),
    .A2(net184));
 sg13g2_mux2_1 _09603_ (.A0(\data_to_write[8] ),
    .A1(net3401),
    .S(_02097_),
    .X(_00769_));
 sg13g2_nor3_1 _09604_ (.A(net317),
    .B(_01766_),
    .C(_01841_),
    .Y(_02102_));
 sg13g2_nand2_1 _09605_ (.Y(_02103_),
    .A(net423),
    .B(_02102_));
 sg13g2_nand2_1 _09606_ (.Y(_02104_),
    .A(net2925),
    .B(net121));
 sg13g2_o21ai_1 _09607_ (.B1(_02104_),
    .Y(_00752_),
    .A1(net392),
    .A2(net121));
 sg13g2_nand2_1 _09608_ (.Y(_02105_),
    .A(net3014),
    .B(net122));
 sg13g2_o21ai_1 _09609_ (.B1(_02105_),
    .Y(_00751_),
    .A1(net386),
    .A2(net121));
 sg13g2_nand2_1 _09610_ (.Y(_02106_),
    .A(net2977),
    .B(net122));
 sg13g2_o21ai_1 _09611_ (.B1(_02106_),
    .Y(_00750_),
    .A1(net381),
    .A2(net122));
 sg13g2_nand2_1 _09612_ (.Y(_02107_),
    .A(net2961),
    .B(net121));
 sg13g2_o21ai_1 _09613_ (.B1(_02107_),
    .Y(_00749_),
    .A1(net375),
    .A2(_02103_));
 sg13g2_nand2_1 _09614_ (.Y(_02108_),
    .A(net2859),
    .B(net122));
 sg13g2_o21ai_1 _09615_ (.B1(_02108_),
    .Y(_00748_),
    .A1(net372),
    .A2(net122));
 sg13g2_nand2_1 _09616_ (.Y(_02109_),
    .A(net2873),
    .B(net122));
 sg13g2_o21ai_1 _09617_ (.B1(_02109_),
    .Y(_00747_),
    .A1(net366),
    .A2(net122));
 sg13g2_nand2_1 _09618_ (.Y(_02110_),
    .A(net2906),
    .B(net121));
 sg13g2_o21ai_1 _09619_ (.B1(_02110_),
    .Y(_00746_),
    .A1(net361),
    .A2(net121));
 sg13g2_nand2_1 _09620_ (.Y(_02111_),
    .A(net2882),
    .B(net121));
 sg13g2_o21ai_1 _09621_ (.B1(_02111_),
    .Y(_00745_),
    .A1(net357),
    .A2(net121));
 sg13g2_nor2b_1 _09622_ (.A(_00198_),
    .B_N(_02095_),
    .Y(_02112_));
 sg13g2_nor2b_2 _09623_ (.A(net632),
    .B_N(_02112_),
    .Y(_02113_));
 sg13g2_and2_1 _09624_ (.A(_02076_),
    .B(_02078_),
    .X(_02114_));
 sg13g2_a21oi_2 _09625_ (.B1(net516),
    .Y(_02115_),
    .A2(_02114_),
    .A1(_02113_));
 sg13g2_nor2_1 _09626_ (.A(\data_to_write[7] ),
    .B(net223),
    .Y(_02116_));
 sg13g2_a21oi_1 _09627_ (.A1(_01549_),
    .A2(net223),
    .Y(_00736_),
    .B1(_02116_));
 sg13g2_nor2_1 _09628_ (.A(net597),
    .B(net223),
    .Y(_02117_));
 sg13g2_a21oi_1 _09629_ (.A1(_01550_),
    .A2(net223),
    .Y(_00735_),
    .B1(_02117_));
 sg13g2_nor2_1 _09630_ (.A(net598),
    .B(net223),
    .Y(_02118_));
 sg13g2_a21oi_1 _09631_ (.A1(_01551_),
    .A2(net223),
    .Y(_00734_),
    .B1(_02118_));
 sg13g2_nor2_1 _09632_ (.A(net599),
    .B(net224),
    .Y(_02119_));
 sg13g2_a21oi_1 _09633_ (.A1(_01552_),
    .A2(net224),
    .Y(_00733_),
    .B1(_02119_));
 sg13g2_nor2_1 _09634_ (.A(\data_to_write[3] ),
    .B(net223),
    .Y(_02120_));
 sg13g2_a21oi_1 _09635_ (.A1(_01553_),
    .A2(net223),
    .Y(_00732_),
    .B1(_02120_));
 sg13g2_nand2_1 _09636_ (.Y(_02121_),
    .A(net3021),
    .B(net224));
 sg13g2_o21ai_1 _09637_ (.B1(_02121_),
    .Y(_00731_),
    .A1(_01509_),
    .A2(net224));
 sg13g2_nand2_1 _09638_ (.Y(_02122_),
    .A(net3084),
    .B(net224));
 sg13g2_o21ai_1 _09639_ (.B1(_02122_),
    .Y(_00730_),
    .A1(_01510_),
    .A2(_02115_));
 sg13g2_nand2_1 _09640_ (.Y(_02123_),
    .A(net2958),
    .B(net224));
 sg13g2_o21ai_1 _09641_ (.B1(_02123_),
    .Y(_00729_),
    .A1(_01511_),
    .A2(net224));
 sg13g2_and2_2 _09642_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .X(_02124_));
 sg13g2_nor2_2 _09643_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .Y(_02125_));
 sg13g2_and2_1 _09644_ (.A(_02124_),
    .B(_02125_),
    .X(_02126_));
 sg13g2_nand2_1 _09645_ (.Y(_02127_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .B(_02126_));
 sg13g2_nor2b_1 _09646_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .Y(_02128_));
 sg13g2_and2_1 _09647_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .X(_02129_));
 sg13g2_and2_1 _09648_ (.A(net566),
    .B(net565),
    .X(_02130_));
 sg13g2_nand3_1 _09649_ (.B(net566),
    .C(net565),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .Y(_02131_));
 sg13g2_nor2b_1 _09650_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .Y(_02132_));
 sg13g2_and2_1 _09651_ (.A(net566),
    .B(net564),
    .X(_02133_));
 sg13g2_nand3_1 _09652_ (.B(net566),
    .C(net564),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .Y(_02134_));
 sg13g2_nor2b_1 _09653_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .Y(_02135_));
 sg13g2_nand3_1 _09654_ (.B(net566),
    .C(net561),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .Y(_02136_));
 sg13g2_nor2_2 _09655_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .Y(_02137_));
 sg13g2_nand3_1 _09656_ (.B(net561),
    .C(net560),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .Y(_02138_));
 sg13g2_nand3_1 _09657_ (.B(net563),
    .C(net560),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .Y(_02139_));
 sg13g2_nor2b_1 _09658_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .Y(_02140_));
 sg13g2_and2_1 _09659_ (.A(net561),
    .B(net559),
    .X(_02141_));
 sg13g2_nand3_1 _09660_ (.B(net562),
    .C(net558),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .Y(_02142_));
 sg13g2_and2_1 _09661_ (.A(net565),
    .B(net558),
    .X(_02143_));
 sg13g2_nand3_1 _09662_ (.B(net565),
    .C(net558),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .Y(_02144_));
 sg13g2_nand3_1 _09663_ (.B(_02125_),
    .C(net558),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .Y(_02145_));
 sg13g2_nand3_1 _09664_ (.B(net564),
    .C(net558),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .Y(_02146_));
 sg13g2_and2_1 _09665_ (.A(_02124_),
    .B(net564),
    .X(_02147_));
 sg13g2_nand4_1 _09666_ (.B(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .C(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .Y(_02148_),
    .D(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ));
 sg13g2_nor2_1 _09667_ (.A(_00127_),
    .B(_02148_),
    .Y(_02149_));
 sg13g2_and2_1 _09668_ (.A(_02124_),
    .B(net562),
    .X(_02150_));
 sg13g2_nand4_1 _09669_ (.B(_02136_),
    .C(_02142_),
    .A(_02134_),
    .Y(_02151_),
    .D(_02144_));
 sg13g2_nand3_1 _09670_ (.B(_02145_),
    .C(_02146_),
    .A(_02131_),
    .Y(_02152_));
 sg13g2_nor2_2 _09671_ (.A(_02151_),
    .B(_02152_),
    .Y(_02153_));
 sg13g2_a221oi_1 _09672_ (.B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .C1(_02149_),
    .B1(_02150_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .Y(_02154_),
    .A2(_02147_));
 sg13g2_and4_1 _09673_ (.A(_02127_),
    .B(_02138_),
    .C(_02139_),
    .D(_02154_),
    .X(_02155_));
 sg13g2_nand2_2 _09674_ (.Y(_02156_),
    .A(_02153_),
    .B(_02155_));
 sg13g2_nand2_2 _09675_ (.Y(_02157_),
    .A(net569),
    .B(\i_tinyqv.cpu.is_auipc ));
 sg13g2_o21ai_1 _09676_ (.B1(net569),
    .Y(_02158_),
    .A1(\i_tinyqv.cpu.is_jal ),
    .A2(\i_tinyqv.cpu.is_auipc ));
 sg13g2_inv_2 _09677_ (.Y(_02159_),
    .A(_02158_));
 sg13g2_nand2_2 _09678_ (.Y(_02160_),
    .A(\i_tinyqv.cpu.alu_op[1] ),
    .B(net574));
 sg13g2_nor2_2 _09679_ (.A(_00121_),
    .B(_02160_),
    .Y(_02161_));
 sg13g2_or2_2 _09680_ (.X(_02162_),
    .B(_02160_),
    .A(_00121_));
 sg13g2_nor2b_1 _09681_ (.A(net589),
    .B_N(net595),
    .Y(_02163_));
 sg13g2_nand2_2 _09682_ (.Y(_02164_),
    .A(_01581_),
    .B(net590));
 sg13g2_nor2b_1 _09683_ (.A(net595),
    .B_N(\i_tinyqv.cpu.counter[3] ),
    .Y(_02165_));
 sg13g2_nand2b_2 _09684_ (.Y(_02166_),
    .B(net588),
    .A_N(net595));
 sg13g2_a22oi_1 _09685_ (.Y(_02167_),
    .B1(net466),
    .B2(\i_tinyqv.cpu.instr_data_start[9] ),
    .A2(net469),
    .A1(\i_tinyqv.cpu.instr_data_start[5] ));
 sg13g2_nor2_1 _09686_ (.A(net588),
    .B(net595),
    .Y(_02168_));
 sg13g2_nand2_2 _09687_ (.Y(_02169_),
    .A(_01581_),
    .B(net472));
 sg13g2_and2_1 _09688_ (.A(net589),
    .B(net591),
    .X(_02170_));
 sg13g2_nand2_2 _09689_ (.Y(_02171_),
    .A(net589),
    .B(net595));
 sg13g2_a22oi_1 _09690_ (.Y(_02172_),
    .B1(net458),
    .B2(net614),
    .A2(net462),
    .A1(\i_tinyqv.cpu.pc[1] ));
 sg13g2_nand2_1 _09691_ (.Y(_02173_),
    .A(_02167_),
    .B(_02172_));
 sg13g2_nor2_2 _09692_ (.A(net474),
    .B(net589),
    .Y(_02174_));
 sg13g2_mux2_1 _09693_ (.A0(net611),
    .A1(net609),
    .S(net594),
    .X(_02175_));
 sg13g2_a22oi_1 _09694_ (.Y(_02176_),
    .B1(_02174_),
    .B2(_02175_),
    .A2(_02173_),
    .A1(net474));
 sg13g2_a21oi_1 _09695_ (.A1(_02159_),
    .A2(_02176_),
    .Y(_02177_),
    .B1(_02161_));
 sg13g2_o21ai_1 _09696_ (.B1(_02177_),
    .Y(_02178_),
    .A1(_02156_),
    .A2(_02159_));
 sg13g2_nor2_1 _09697_ (.A(\i_tinyqv.cpu.alu_op[3] ),
    .B(_00125_),
    .Y(_02179_));
 sg13g2_a21oi_2 _09698_ (.B1(_02179_),
    .Y(_02180_),
    .A2(_02160_),
    .A1(\i_tinyqv.cpu.alu_op[3] ));
 sg13g2_a21o_1 _09699_ (.A2(_02160_),
    .A1(\i_tinyqv.cpu.alu_op[3] ),
    .B1(_02179_),
    .X(_02181_));
 sg13g2_nor2_1 _09700_ (.A(_01487_),
    .B(_01491_),
    .Y(_02182_));
 sg13g2_nand2_1 _09701_ (.Y(_02183_),
    .A(net570),
    .B(\i_tinyqv.cpu.is_branch ));
 sg13g2_o21ai_1 _09702_ (.B1(net569),
    .Y(_02184_),
    .A1(\i_tinyqv.cpu.is_branch ),
    .A2(\i_tinyqv.cpu.is_alu_reg ));
 sg13g2_and2_1 _09703_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .X(_02185_));
 sg13g2_nor2b_1 _09704_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .Y(_02186_));
 sg13g2_and2_1 _09705_ (.A(net556),
    .B(net555),
    .X(_02187_));
 sg13g2_nor2b_2 _09706_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .Y(_02188_));
 sg13g2_nor2b_1 _09707_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .Y(_02189_));
 sg13g2_and2_1 _09708_ (.A(_02188_),
    .B(net552),
    .X(_02190_));
 sg13g2_a22oi_1 _09709_ (.Y(_02191_),
    .B1(_02190_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .A2(_02187_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ));
 sg13g2_nor2_1 _09710_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .Y(_02192_));
 sg13g2_nor2b_1 _09711_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .Y(_02193_));
 sg13g2_nand3_1 _09712_ (.B(net551),
    .C(net550),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .Y(_02194_));
 sg13g2_nand3_1 _09713_ (.B(net553),
    .C(net551),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .Y(_02195_));
 sg13g2_and2_1 _09714_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .X(_02196_));
 sg13g2_and2_1 _09715_ (.A(net550),
    .B(net548),
    .X(_02197_));
 sg13g2_and2_1 _09716_ (.A(net552),
    .B(net548),
    .X(_02198_));
 sg13g2_a22oi_1 _09717_ (.Y(_02199_),
    .B1(_02198_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .A2(_02197_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ));
 sg13g2_nand4_1 _09718_ (.B(_02194_),
    .C(_02195_),
    .A(_02191_),
    .Y(_02200_),
    .D(_02199_));
 sg13g2_nor2_2 _09719_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .Y(_02201_));
 sg13g2_and2_1 _09720_ (.A(net548),
    .B(_02201_),
    .X(_02202_));
 sg13g2_and2_1 _09721_ (.A(_02188_),
    .B(net549),
    .X(_02203_));
 sg13g2_and2_1 _09722_ (.A(net556),
    .B(net548),
    .X(_02204_));
 sg13g2_nand4_1 _09723_ (.B(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .C(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .Y(_02205_),
    .D(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ));
 sg13g2_nor2_1 _09724_ (.A(_00127_),
    .B(_02205_),
    .Y(_02206_));
 sg13g2_a221oi_1 _09725_ (.B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .C1(_02206_),
    .B1(_02203_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .Y(_02207_),
    .A2(_02202_));
 sg13g2_and2_1 _09726_ (.A(net556),
    .B(_02188_),
    .X(_02208_));
 sg13g2_and2_1 _09727_ (.A(_02188_),
    .B(_02201_),
    .X(_02209_));
 sg13g2_a22oi_1 _09728_ (.Y(_02210_),
    .B1(_02209_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .A2(_02208_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ));
 sg13g2_nand3_1 _09729_ (.B(net554),
    .C(net552),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .Y(_02211_));
 sg13g2_nand3_1 _09730_ (.B(net554),
    .C(net549),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .Y(_02212_));
 sg13g2_nand4_1 _09731_ (.B(_02210_),
    .C(_02211_),
    .A(_02207_),
    .Y(_02213_),
    .D(_02212_));
 sg13g2_or2_2 _09732_ (.X(_02214_),
    .B(_02213_),
    .A(_02200_));
 sg13g2_a21oi_1 _09733_ (.A1(\i_tinyqv.cpu.imm[25] ),
    .A2(net465),
    .Y(_02215_),
    .B1(net475));
 sg13g2_and2_1 _09734_ (.A(\i_tinyqv.cpu.imm[17] ),
    .B(net462),
    .X(_02216_));
 sg13g2_a221oi_1 _09735_ (.B2(\i_tinyqv.cpu.imm[29] ),
    .C1(_02216_),
    .B1(net457),
    .A1(\i_tinyqv.cpu.imm[21] ),
    .Y(_02217_),
    .A2(net468));
 sg13g2_nor2_1 _09736_ (.A(_01590_),
    .B(_02171_),
    .Y(_02218_));
 sg13g2_a221oi_1 _09737_ (.B2(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .C1(_02218_),
    .B1(net465),
    .A1(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .Y(_02219_),
    .A2(net468));
 sg13g2_a21oi_1 _09738_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .A2(net461),
    .Y(_02220_),
    .B1(net585));
 sg13g2_a22oi_1 _09739_ (.Y(_02221_),
    .B1(_02219_),
    .B2(_02220_),
    .A2(_02217_),
    .A1(_02215_));
 sg13g2_mux2_1 _09740_ (.A0(_02214_),
    .A1(_02221_),
    .S(_02184_),
    .X(_02222_));
 sg13g2_inv_1 _09741_ (.Y(_02223_),
    .A(_02222_));
 sg13g2_xnor2_1 _09742_ (.Y(_02224_),
    .A(_02180_),
    .B(_02222_));
 sg13g2_nor2b_1 _09743_ (.A(_02178_),
    .B_N(_02224_),
    .Y(_02225_));
 sg13g2_nand3_1 _09744_ (.B(net563),
    .C(net560),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .Y(_02226_));
 sg13g2_nand3_1 _09745_ (.B(net561),
    .C(net560),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .Y(_02227_));
 sg13g2_nand3_1 _09746_ (.B(_02125_),
    .C(net559),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .Y(_02228_));
 sg13g2_nand3_1 _09747_ (.B(net565),
    .C(net559),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .Y(_02229_));
 sg13g2_nand3_1 _09748_ (.B(_02124_),
    .C(_02125_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .Y(_02230_));
 sg13g2_and2_1 _09749_ (.A(net586),
    .B(net589),
    .X(_02231_));
 sg13g2_nand2_1 _09750_ (.Y(_02232_),
    .A(net586),
    .B(net589));
 sg13g2_and2_1 _09751_ (.A(_02129_),
    .B(net560),
    .X(_02233_));
 sg13g2_nand4_1 _09752_ (.B(net565),
    .C(net560),
    .A(net473),
    .Y(_02234_),
    .D(net456));
 sg13g2_nand3_1 _09753_ (.B(_02124_),
    .C(net563),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .Y(_02235_));
 sg13g2_nand3_1 _09754_ (.B(net567),
    .C(net563),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .Y(_02236_));
 sg13g2_nand3_1 _09755_ (.B(net567),
    .C(net565),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .Y(_02237_));
 sg13g2_nand3_1 _09756_ (.B(net561),
    .C(net559),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .Y(_02238_));
 sg13g2_nand3_1 _09757_ (.B(_02124_),
    .C(net562),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .Y(_02239_));
 sg13g2_nand3_1 _09758_ (.B(net563),
    .C(net559),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .Y(_02240_));
 sg13g2_nand3_1 _09759_ (.B(net567),
    .C(net561),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .Y(_02241_));
 sg13g2_nand4_1 _09760_ (.B(_02237_),
    .C(_02238_),
    .A(_02235_),
    .Y(_02242_),
    .D(_02240_));
 sg13g2_nand4_1 _09761_ (.B(_02227_),
    .C(_02228_),
    .A(_02226_),
    .Y(_02243_),
    .D(_02234_));
 sg13g2_nor2_1 _09762_ (.A(_02242_),
    .B(_02243_),
    .Y(_02244_));
 sg13g2_o21ai_1 _09763_ (.B1(_02230_),
    .Y(_02245_),
    .A1(_01591_),
    .A2(_02148_));
 sg13g2_nand4_1 _09764_ (.B(_02236_),
    .C(_02239_),
    .A(_02229_),
    .Y(_02246_),
    .D(_02241_));
 sg13g2_nor2_2 _09765_ (.A(_02245_),
    .B(_02246_),
    .Y(_02247_));
 sg13g2_nand2_2 _09766_ (.Y(_02248_),
    .A(_02244_),
    .B(_02247_));
 sg13g2_nor2_2 _09767_ (.A(net583),
    .B(net588),
    .Y(_02249_));
 sg13g2_nor2_2 _09768_ (.A(net583),
    .B(_02164_),
    .Y(_02250_));
 sg13g2_a22oi_1 _09769_ (.Y(_02251_),
    .B1(net458),
    .B2(\i_tinyqv.cpu.instr_data_start[12] ),
    .A2(net469),
    .A1(\i_tinyqv.cpu.instr_data_start[4] ));
 sg13g2_nor2_1 _09770_ (.A(net585),
    .B(_02251_),
    .Y(_02252_));
 sg13g2_mux2_1 _09771_ (.A0(net612),
    .A1(net610),
    .S(net594),
    .X(_02253_));
 sg13g2_nor2_2 _09772_ (.A(net583),
    .B(net464),
    .Y(_02254_));
 sg13g2_a221oi_1 _09773_ (.B2(\i_tinyqv.cpu.instr_data_start[8] ),
    .C1(_02252_),
    .B1(_02254_),
    .A1(_02174_),
    .Y(_02255_),
    .A2(_02253_));
 sg13g2_a21oi_1 _09774_ (.A1(_02159_),
    .A2(_02255_),
    .Y(_02256_),
    .B1(_02161_));
 sg13g2_o21ai_1 _09775_ (.B1(_02256_),
    .Y(_02257_),
    .A1(_02159_),
    .A2(_02248_));
 sg13g2_inv_1 _09776_ (.Y(_02258_),
    .A(_02257_));
 sg13g2_nand3_1 _09777_ (.B(net548),
    .C(_02201_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .Y(_02259_));
 sg13g2_a22oi_1 _09778_ (.Y(_02260_),
    .B1(_02203_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .A2(_02198_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ));
 sg13g2_nand3_1 _09779_ (.B(net556),
    .C(net554),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .Y(_02261_));
 sg13g2_nand3_1 _09780_ (.B(net555),
    .C(net550),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .Y(_02262_));
 sg13g2_a22oi_1 _09781_ (.Y(_02263_),
    .B1(_02204_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .A2(_02190_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ));
 sg13g2_nand3_1 _09782_ (.B(net553),
    .C(net551),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .Y(_02264_));
 sg13g2_nand3_1 _09783_ (.B(net555),
    .C(net553),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .Y(_02265_));
 sg13g2_nand4_1 _09784_ (.B(net556),
    .C(net551),
    .A(net473),
    .Y(_02266_),
    .D(net456));
 sg13g2_nand2_1 _09785_ (.Y(_02267_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .B(_02197_));
 sg13g2_nand3_1 _09786_ (.B(net551),
    .C(net549),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .Y(_02268_));
 sg13g2_and4_2 _09787_ (.A(_02259_),
    .B(_02260_),
    .C(_02263_),
    .D(_02264_),
    .X(_02269_));
 sg13g2_a22oi_1 _09788_ (.Y(_02270_),
    .B1(_02209_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .A2(_02208_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ));
 sg13g2_and4_1 _09789_ (.A(_02261_),
    .B(_02262_),
    .C(_02266_),
    .D(_02268_),
    .X(_02271_));
 sg13g2_and4_2 _09790_ (.A(_02265_),
    .B(_02267_),
    .C(_02270_),
    .D(_02271_),
    .X(_02272_));
 sg13g2_nand2_1 _09791_ (.Y(_02273_),
    .A(_02269_),
    .B(_02272_));
 sg13g2_and2_1 _09792_ (.A(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .B(net468),
    .X(_02274_));
 sg13g2_a221oi_1 _09793_ (.B2(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .C1(_02274_),
    .B1(net461),
    .A1(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .Y(_02275_),
    .A2(net465));
 sg13g2_a21oi_1 _09794_ (.A1(\i_tinyqv.cpu.imm[12] ),
    .A2(net457),
    .Y(_02276_),
    .B1(net585));
 sg13g2_a22oi_1 _09795_ (.Y(_02277_),
    .B1(net462),
    .B2(\i_tinyqv.cpu.imm[16] ),
    .A2(net465),
    .A1(\i_tinyqv.cpu.imm[24] ));
 sg13g2_a221oi_1 _09796_ (.B2(\i_tinyqv.cpu.imm[28] ),
    .C1(net475),
    .B1(net459),
    .A1(\i_tinyqv.cpu.imm[20] ),
    .Y(_02278_),
    .A2(net470));
 sg13g2_a22oi_1 _09797_ (.Y(_02279_),
    .B1(_02277_),
    .B2(_02278_),
    .A2(_02276_),
    .A1(_02275_));
 sg13g2_inv_2 _09798_ (.Y(_02280_),
    .A(_02279_));
 sg13g2_nand2_1 _09799_ (.Y(_02281_),
    .A(_02184_),
    .B(_02279_));
 sg13g2_a21o_1 _09800_ (.A2(_02272_),
    .A1(_02269_),
    .B1(_02184_),
    .X(_02282_));
 sg13g2_nand2_1 _09801_ (.Y(_02283_),
    .A(_02281_),
    .B(_02282_));
 sg13g2_and3_1 _09802_ (.X(_02284_),
    .A(_02180_),
    .B(_02281_),
    .C(_02282_));
 sg13g2_a21oi_1 _09803_ (.A1(_02281_),
    .A2(_02282_),
    .Y(_02285_),
    .B1(_02180_));
 sg13g2_nor3_1 _09804_ (.A(_02257_),
    .B(_02284_),
    .C(_02285_),
    .Y(_02286_));
 sg13g2_o21ai_1 _09805_ (.B1(_02257_),
    .Y(_02287_),
    .A1(_02284_),
    .A2(_02285_));
 sg13g2_nor2b_1 _09806_ (.A(_02286_),
    .B_N(_02287_),
    .Y(_02288_));
 sg13g2_nor2_1 _09807_ (.A(net586),
    .B(_02169_),
    .Y(_02289_));
 sg13g2_nand2_2 _09808_ (.Y(_02290_),
    .A(net474),
    .B(net462));
 sg13g2_nor2_1 _09809_ (.A(_02181_),
    .B(net335),
    .Y(_02291_));
 sg13g2_a21oi_1 _09810_ (.A1(_00128_),
    .A2(net335),
    .Y(_02292_),
    .B1(_02291_));
 sg13g2_a21o_1 _09811_ (.A2(_02292_),
    .A1(_02287_),
    .B1(_02286_),
    .X(_02293_));
 sg13g2_xnor2_1 _09812_ (.Y(_02294_),
    .A(_02178_),
    .B(_02224_));
 sg13g2_a21oi_2 _09813_ (.B1(_02225_),
    .Y(_02295_),
    .A2(_02294_),
    .A1(_02293_));
 sg13g2_nand3_1 _09814_ (.B(net563),
    .C(net560),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .Y(_02296_));
 sg13g2_nand3_1 _09815_ (.B(net567),
    .C(net561),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .Y(_02297_));
 sg13g2_nor2_1 _09816_ (.A(_00123_),
    .B(_02148_),
    .Y(_02298_));
 sg13g2_nand3_1 _09817_ (.B(net563),
    .C(net559),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .Y(_02299_));
 sg13g2_nand3_1 _09818_ (.B(net561),
    .C(net560),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .Y(_02300_));
 sg13g2_and2_1 _09819_ (.A(_02299_),
    .B(_02300_),
    .X(_02301_));
 sg13g2_nand4_1 _09820_ (.B(_02125_),
    .C(net567),
    .A(net473),
    .Y(_02302_),
    .D(net456));
 sg13g2_a22oi_1 _09821_ (.Y(_02303_),
    .B1(_02147_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .A2(_02130_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ));
 sg13g2_nand3_1 _09822_ (.B(_02125_),
    .C(net558),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .Y(_02304_));
 sg13g2_and2_1 _09823_ (.A(_02296_),
    .B(_02304_),
    .X(_02305_));
 sg13g2_a22oi_1 _09824_ (.Y(_02306_),
    .B1(_02143_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .A2(_02126_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ));
 sg13g2_a22oi_1 _09825_ (.Y(_02307_),
    .B1(_02150_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .A2(_02133_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ));
 sg13g2_and4_2 _09826_ (.A(_02303_),
    .B(_02305_),
    .C(_02306_),
    .D(_02307_),
    .X(_02308_));
 sg13g2_a21oi_1 _09827_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .A2(_02141_),
    .Y(_02309_),
    .B1(_02298_));
 sg13g2_and4_2 _09828_ (.A(_02297_),
    .B(_02301_),
    .C(_02302_),
    .D(_02309_),
    .X(_02310_));
 sg13g2_nand2_2 _09829_ (.Y(_02311_),
    .A(_02308_),
    .B(_02310_));
 sg13g2_a22oi_1 _09830_ (.Y(_02312_),
    .B1(net466),
    .B2(\i_tinyqv.cpu.instr_data_start[11] ),
    .A2(net469),
    .A1(\i_tinyqv.cpu.instr_data_start[7] ));
 sg13g2_a22oi_1 _09831_ (.Y(_02313_),
    .B1(net458),
    .B2(\i_tinyqv.cpu.instr_data_start[15] ),
    .A2(net461),
    .A1(\i_tinyqv.cpu.instr_data_start[3] ));
 sg13g2_nand2_1 _09832_ (.Y(_02314_),
    .A(_02312_),
    .B(_02313_));
 sg13g2_mux2_1 _09833_ (.A0(\i_tinyqv.cpu.instr_data_start[19] ),
    .A1(\i_tinyqv.cpu.instr_data_start[23] ),
    .S(net593),
    .X(_02315_));
 sg13g2_a22oi_1 _09834_ (.Y(_02316_),
    .B1(_02315_),
    .B2(_02174_),
    .A2(_02314_),
    .A1(net475));
 sg13g2_a21oi_1 _09835_ (.A1(_02159_),
    .A2(_02316_),
    .Y(_02317_),
    .B1(_02161_));
 sg13g2_o21ai_1 _09836_ (.B1(_02317_),
    .Y(_02318_),
    .A1(_02159_),
    .A2(_02311_));
 sg13g2_nand4_1 _09837_ (.B(net554),
    .C(_02201_),
    .A(net473),
    .Y(_02319_),
    .D(net456));
 sg13g2_nand3_1 _09838_ (.B(net548),
    .C(_02201_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .Y(_02320_));
 sg13g2_nand3_1 _09839_ (.B(net552),
    .C(net548),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .Y(_02321_));
 sg13g2_nand3_1 _09840_ (.B(net550),
    .C(_02196_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .Y(_02322_));
 sg13g2_or2_1 _09841_ (.X(_02323_),
    .B(_02205_),
    .A(_00123_));
 sg13g2_nand3_1 _09842_ (.B(net552),
    .C(_02192_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .Y(_02324_));
 sg13g2_nand3_1 _09843_ (.B(net554),
    .C(net549),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .Y(_02325_));
 sg13g2_nand3_1 _09844_ (.B(net556),
    .C(net555),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .Y(_02326_));
 sg13g2_nand3_1 _09845_ (.B(net556),
    .C(_02188_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .Y(_02327_));
 sg13g2_nand3_1 _09846_ (.B(_02188_),
    .C(net549),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .Y(_02328_));
 sg13g2_nand4_1 _09847_ (.B(_02326_),
    .C(_02327_),
    .A(_02325_),
    .Y(_02329_),
    .D(_02328_));
 sg13g2_nand3_1 _09848_ (.B(net551),
    .C(net549),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .Y(_02330_));
 sg13g2_nand3_1 _09849_ (.B(_02188_),
    .C(_02201_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .Y(_02331_));
 sg13g2_nand3_1 _09850_ (.B(net555),
    .C(net553),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .Y(_02332_));
 sg13g2_nand3_1 _09851_ (.B(_02188_),
    .C(net552),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .Y(_02333_));
 sg13g2_nand3_1 _09852_ (.B(_02323_),
    .C(_02333_),
    .A(_02319_),
    .Y(_02334_));
 sg13g2_nand4_1 _09853_ (.B(_02322_),
    .C(_02330_),
    .A(_02321_),
    .Y(_02335_),
    .D(_02332_));
 sg13g2_nand3_1 _09854_ (.B(_02324_),
    .C(_02331_),
    .A(_02320_),
    .Y(_02336_));
 sg13g2_nor4_2 _09855_ (.A(_02329_),
    .B(_02334_),
    .C(_02335_),
    .Y(_02337_),
    .D(_02336_));
 sg13g2_a21oi_1 _09856_ (.A1(\i_tinyqv.cpu.imm[31] ),
    .A2(net457),
    .Y(_02338_),
    .B1(net474));
 sg13g2_and2_1 _09857_ (.A(\i_tinyqv.cpu.imm[19] ),
    .B(net462),
    .X(_02339_));
 sg13g2_a221oi_1 _09858_ (.B2(\i_tinyqv.cpu.imm[27] ),
    .C1(_02339_),
    .B1(net466),
    .A1(\i_tinyqv.cpu.imm[23] ),
    .Y(_02340_),
    .A2(net470));
 sg13g2_a22oi_1 _09859_ (.Y(_02341_),
    .B1(net457),
    .B2(\i_tinyqv.cpu.imm[15] ),
    .A2(net468),
    .A1(\i_tinyqv.cpu.i_core.imm_lo[7] ));
 sg13g2_a221oi_1 _09860_ (.B2(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .C1(net585),
    .B1(net461),
    .A1(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .Y(_02342_),
    .A2(net465));
 sg13g2_a22oi_1 _09861_ (.Y(_02343_),
    .B1(_02341_),
    .B2(_02342_),
    .A2(_02340_),
    .A1(_02338_));
 sg13g2_nor2_1 _09862_ (.A(_02184_),
    .B(_02337_),
    .Y(_02344_));
 sg13g2_a21oi_2 _09863_ (.B1(_02344_),
    .Y(_02345_),
    .A2(_02343_),
    .A1(_02184_));
 sg13g2_xnor2_1 _09864_ (.Y(_02346_),
    .A(_02181_),
    .B(_02345_));
 sg13g2_nor2b_1 _09865_ (.A(_02318_),
    .B_N(_02346_),
    .Y(_02347_));
 sg13g2_nand2b_1 _09866_ (.Y(_02348_),
    .B(_02318_),
    .A_N(_02346_));
 sg13g2_xor2_1 _09867_ (.B(_02346_),
    .A(_02318_),
    .X(_02349_));
 sg13g2_inv_1 _09868_ (.Y(_02350_),
    .A(_02349_));
 sg13g2_nand3_1 _09869_ (.B(_02124_),
    .C(_02125_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .Y(_02351_));
 sg13g2_nand3_1 _09870_ (.B(net563),
    .C(_02137_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .Y(_02352_));
 sg13g2_nand3_1 _09871_ (.B(_02125_),
    .C(net558),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .Y(_02353_));
 sg13g2_nand3_1 _09872_ (.B(net566),
    .C(net565),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .Y(_02354_));
 sg13g2_nand3_1 _09873_ (.B(net564),
    .C(net558),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .Y(_02355_));
 sg13g2_nand3_1 _09874_ (.B(net566),
    .C(net564),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .Y(_02356_));
 sg13g2_or2_1 _09875_ (.X(_02357_),
    .B(_02148_),
    .A(_00126_));
 sg13g2_nand2_1 _09876_ (.Y(_02358_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .B(_02141_));
 sg13g2_nand3_1 _09877_ (.B(net562),
    .C(_02137_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .Y(_02359_));
 sg13g2_nand3_1 _09878_ (.B(net566),
    .C(net562),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .Y(_02360_));
 sg13g2_nand4_1 _09879_ (.B(_02357_),
    .C(_02358_),
    .A(_02355_),
    .Y(_02361_),
    .D(_02359_));
 sg13g2_a221oi_1 _09880_ (.B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .C1(_02361_),
    .B1(_02150_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .Y(_02362_),
    .A2(_02143_));
 sg13g2_nand4_1 _09881_ (.B(_02354_),
    .C(_02356_),
    .A(_02351_),
    .Y(_02363_),
    .D(_02360_));
 sg13g2_a221oi_1 _09882_ (.B2(_02254_),
    .C1(_02363_),
    .B1(_02233_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .Y(_02364_),
    .A2(_02147_));
 sg13g2_nand4_1 _09883_ (.B(_02353_),
    .C(_02362_),
    .A(_02352_),
    .Y(_02365_),
    .D(_02364_));
 sg13g2_a22oi_1 _09884_ (.Y(_02366_),
    .B1(net465),
    .B2(\i_tinyqv.cpu.instr_data_start[10] ),
    .A2(net469),
    .A1(\i_tinyqv.cpu.instr_data_start[6] ));
 sg13g2_a22oi_1 _09885_ (.Y(_02367_),
    .B1(net458),
    .B2(net613),
    .A2(net461),
    .A1(\i_tinyqv.cpu.pc[2] ));
 sg13g2_nand2_1 _09886_ (.Y(_02368_),
    .A(_02366_),
    .B(_02367_));
 sg13g2_nand2_1 _09887_ (.Y(_02369_),
    .A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(net593));
 sg13g2_o21ai_1 _09888_ (.B1(_02369_),
    .Y(_02370_),
    .A1(_01513_),
    .A2(net593));
 sg13g2_a22oi_1 _09889_ (.Y(_02371_),
    .B1(_02370_),
    .B2(_02174_),
    .A2(_02368_),
    .A1(net474));
 sg13g2_a21oi_1 _09890_ (.A1(_02159_),
    .A2(_02371_),
    .Y(_02372_),
    .B1(_02161_));
 sg13g2_o21ai_1 _09891_ (.B1(_02372_),
    .Y(_02373_),
    .A1(_02159_),
    .A2(_02365_));
 sg13g2_nand3_1 _09892_ (.B(net548),
    .C(_02201_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .Y(_02374_));
 sg13g2_nand3_1 _09893_ (.B(net556),
    .C(net554),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .Y(_02375_));
 sg13g2_nand3_1 _09894_ (.B(net551),
    .C(_02254_),
    .A(net557),
    .Y(_02376_));
 sg13g2_nand3_1 _09895_ (.B(net554),
    .C(net549),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .Y(_02377_));
 sg13g2_nand3_1 _09896_ (.B(net554),
    .C(net552),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .Y(_02378_));
 sg13g2_nand3_1 _09897_ (.B(net552),
    .C(_02192_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .Y(_02379_));
 sg13g2_nand3_1 _09898_ (.B(net551),
    .C(net549),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .Y(_02380_));
 sg13g2_or2_1 _09899_ (.X(_02381_),
    .B(_02205_),
    .A(_00126_));
 sg13g2_a22oi_1 _09900_ (.Y(_02382_),
    .B1(_02198_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .A2(_02197_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ));
 sg13g2_a22oi_1 _09901_ (.Y(_02383_),
    .B1(_02203_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .A2(_02190_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ));
 sg13g2_and4_1 _09902_ (.A(_02374_),
    .B(_02377_),
    .C(_02378_),
    .D(_02381_),
    .X(_02384_));
 sg13g2_nand4_1 _09903_ (.B(_02379_),
    .C(_02383_),
    .A(_02375_),
    .Y(_02385_),
    .D(_02384_));
 sg13g2_a22oi_1 _09904_ (.Y(_02386_),
    .B1(_02209_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .A2(_02208_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ));
 sg13g2_nand4_1 _09905_ (.B(_02380_),
    .C(_02382_),
    .A(_02376_),
    .Y(_02387_),
    .D(_02386_));
 sg13g2_or2_2 _09906_ (.X(_02388_),
    .B(_02387_),
    .A(_02385_));
 sg13g2_a21oi_1 _09907_ (.A1(\i_tinyqv.cpu.imm[14] ),
    .A2(net457),
    .Y(_02389_),
    .B1(net585));
 sg13g2_nand2_1 _09908_ (.Y(_02390_),
    .A(net582),
    .B(net461));
 sg13g2_a22oi_1 _09909_ (.Y(_02391_),
    .B1(net465),
    .B2(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .A2(net468),
    .A1(\i_tinyqv.cpu.i_core.imm_lo[6] ));
 sg13g2_nand3_1 _09910_ (.B(_02390_),
    .C(_02391_),
    .A(_02389_),
    .Y(_02392_));
 sg13g2_a22oi_1 _09911_ (.Y(_02393_),
    .B1(net459),
    .B2(\i_tinyqv.cpu.imm[30] ),
    .A2(net462),
    .A1(\i_tinyqv.cpu.imm[18] ));
 sg13g2_a221oi_1 _09912_ (.B2(\i_tinyqv.cpu.imm[26] ),
    .C1(net475),
    .B1(net466),
    .A1(\i_tinyqv.cpu.imm[22] ),
    .Y(_02394_),
    .A2(net470));
 sg13g2_nand2_2 _09913_ (.Y(_02395_),
    .A(_02393_),
    .B(_02394_));
 sg13g2_nand2_2 _09914_ (.Y(_02396_),
    .A(_02392_),
    .B(_02395_));
 sg13g2_nand2_1 _09915_ (.Y(_02397_),
    .A(_02184_),
    .B(_02396_));
 sg13g2_o21ai_1 _09916_ (.B1(_02397_),
    .Y(_02398_),
    .A1(_02184_),
    .A2(_02388_));
 sg13g2_xnor2_1 _09917_ (.Y(_02399_),
    .A(_02181_),
    .B(_02398_));
 sg13g2_nor2b_1 _09918_ (.A(_02373_),
    .B_N(_02399_),
    .Y(_02400_));
 sg13g2_xor2_1 _09919_ (.B(_02399_),
    .A(_02373_),
    .X(_02401_));
 sg13g2_or2_1 _09920_ (.X(_02402_),
    .B(_02401_),
    .A(_02349_));
 sg13g2_o21ai_1 _09921_ (.B1(_02348_),
    .Y(_02403_),
    .A1(_02347_),
    .A2(_02400_));
 sg13g2_o21ai_1 _09922_ (.B1(_02403_),
    .Y(\i_tinyqv.cpu.i_core.cy_out ),
    .A1(_02295_),
    .A2(_02402_));
 sg13g2_nand2b_1 _09923_ (.Y(_02404_),
    .B(\i_time.l_mtimecmp.data_out[29] ),
    .A_N(\i_time.mtime[29] ));
 sg13g2_nand2b_1 _09924_ (.Y(_02405_),
    .B(\i_time.mtime[27] ),
    .A_N(\i_time.l_mtimecmp.data_out[27] ));
 sg13g2_o21ai_1 _09925_ (.B1(_02405_),
    .Y(_02406_),
    .A1(_01530_),
    .A2(\i_time.l_mtimecmp.data_out[26] ));
 sg13g2_nand2_1 _09926_ (.Y(_02407_),
    .A(_01529_),
    .B(\i_time.l_mtimecmp.data_out[27] ));
 sg13g2_nand2b_1 _09927_ (.Y(_02408_),
    .B(_02407_),
    .A_N(_02406_));
 sg13g2_a221oi_1 _09928_ (.B2(_01531_),
    .C1(_02408_),
    .B1(\i_time.l_mtimecmp.data_out[25] ),
    .A1(_01530_),
    .Y(_02409_),
    .A2(\i_time.l_mtimecmp.data_out[26] ));
 sg13g2_a22oi_1 _09929_ (.Y(_02410_),
    .B1(_01627_),
    .B2(\i_time.mtime[24] ),
    .A2(_01626_),
    .A1(\i_time.mtime[25] ));
 sg13g2_nand2_1 _09930_ (.Y(_02411_),
    .A(_01537_),
    .B(\i_time.l_mtimecmp.data_out[15] ));
 sg13g2_a22oi_1 _09931_ (.Y(_02412_),
    .B1(_01636_),
    .B2(\i_time.mtime[14] ),
    .A2(_01635_),
    .A1(\i_time.mtime[15] ));
 sg13g2_nand2_1 _09932_ (.Y(_02413_),
    .A(\i_time.mtime[12] ),
    .B(_01638_));
 sg13g2_a22oi_1 _09933_ (.Y(_02414_),
    .B1(_01638_),
    .B2(\i_time.mtime[12] ),
    .A2(_01637_),
    .A1(\i_time.mtime[13] ));
 sg13g2_o21ai_1 _09934_ (.B1(_02413_),
    .Y(_02415_),
    .A1(_01538_),
    .A2(\i_time.l_mtimecmp.data_out[13] ));
 sg13g2_nand2_1 _09935_ (.Y(_02416_),
    .A(_01538_),
    .B(\i_time.l_mtimecmp.data_out[13] ));
 sg13g2_o21ai_1 _09936_ (.B1(_02416_),
    .Y(_02417_),
    .A1(\i_time.mtime[14] ),
    .A2(_01636_));
 sg13g2_o21ai_1 _09937_ (.B1(_02412_),
    .Y(_02418_),
    .A1(_02414_),
    .A2(_02417_));
 sg13g2_nand2b_1 _09938_ (.Y(_02419_),
    .B(\i_time.l_mtimecmp.data_out[8] ),
    .A_N(\i_time.mtime[8] ));
 sg13g2_a22oi_1 _09939_ (.Y(_02420_),
    .B1(\i_time.l_mtimecmp.data_out[0] ),
    .B2(_01548_),
    .A2(\i_time.l_mtimecmp.data_out[1] ),
    .A1(_01547_));
 sg13g2_a221oi_1 _09940_ (.B2(\i_time.mtime[1] ),
    .C1(_02420_),
    .B1(_01646_),
    .A1(\i_time.mtime[2] ),
    .Y(_02421_),
    .A2(_01645_));
 sg13g2_a21o_1 _09941_ (.A2(\i_time.l_mtimecmp.data_out[2] ),
    .A1(_01546_),
    .B1(_02421_),
    .X(_02422_));
 sg13g2_o21ai_1 _09942_ (.B1(_02422_),
    .Y(_02423_),
    .A1(_01545_),
    .A2(\i_time.l_mtimecmp.data_out[3] ));
 sg13g2_a22oi_1 _09943_ (.Y(_02424_),
    .B1(\i_time.l_mtimecmp.data_out[3] ),
    .B2(_01545_),
    .A2(\i_time.l_mtimecmp.data_out[4] ),
    .A1(_01544_));
 sg13g2_nor2_1 _09944_ (.A(_01543_),
    .B(\i_time.l_mtimecmp.data_out[5] ),
    .Y(_02425_));
 sg13g2_a221oi_1 _09945_ (.B2(_02424_),
    .C1(_02425_),
    .B1(_02423_),
    .A1(\i_time.mtime[4] ),
    .Y(_02426_),
    .A2(_01644_));
 sg13g2_a221oi_1 _09946_ (.B2(_01543_),
    .C1(_02426_),
    .B1(\i_time.l_mtimecmp.data_out[5] ),
    .A1(_01542_),
    .Y(_02427_),
    .A2(\i_time.l_mtimecmp.data_out[6] ));
 sg13g2_a221oi_1 _09947_ (.B2(\i_time.mtime[6] ),
    .C1(_02427_),
    .B1(_01643_),
    .A1(\i_time.mtime[7] ),
    .Y(_02428_),
    .A2(_01642_));
 sg13g2_o21ai_1 _09948_ (.B1(_02419_),
    .Y(_02429_),
    .A1(\i_time.mtime[7] ),
    .A2(_01642_));
 sg13g2_a22oi_1 _09949_ (.Y(_02430_),
    .B1(_01641_),
    .B2(\i_time.mtime[8] ),
    .A2(_01640_),
    .A1(\i_time.mtime[9] ));
 sg13g2_o21ai_1 _09950_ (.B1(_02430_),
    .Y(_02431_),
    .A1(_02428_),
    .A2(_02429_));
 sg13g2_nand2b_1 _09951_ (.Y(_02432_),
    .B(\i_time.l_mtimecmp.data_out[11] ),
    .A_N(\i_time.mtime[11] ));
 sg13g2_a22oi_1 _09952_ (.Y(_02433_),
    .B1(\i_time.l_mtimecmp.data_out[9] ),
    .B2(_01541_),
    .A2(\i_time.l_mtimecmp.data_out[10] ),
    .A1(_01540_));
 sg13g2_nand3_1 _09953_ (.B(_02432_),
    .C(_02433_),
    .A(_02431_),
    .Y(_02434_));
 sg13g2_nand2b_1 _09954_ (.Y(_02435_),
    .B(\i_time.mtime[10] ),
    .A_N(\i_time.l_mtimecmp.data_out[10] ));
 sg13g2_nand2_1 _09955_ (.Y(_02436_),
    .A(\i_time.mtime[11] ),
    .B(_01639_));
 sg13g2_nand3_1 _09956_ (.B(_02435_),
    .C(_02436_),
    .A(_02434_),
    .Y(_02437_));
 sg13g2_nand2_1 _09957_ (.Y(_02438_),
    .A(_01539_),
    .B(\i_time.l_mtimecmp.data_out[12] ));
 sg13g2_nand3_1 _09958_ (.B(_02412_),
    .C(_02438_),
    .A(_02411_),
    .Y(_02439_));
 sg13g2_nor2_1 _09959_ (.A(_02432_),
    .B(_02435_),
    .Y(_02440_));
 sg13g2_nor4_1 _09960_ (.A(_02415_),
    .B(_02417_),
    .C(_02439_),
    .D(_02440_),
    .Y(_02441_));
 sg13g2_a22oi_1 _09961_ (.Y(_02442_),
    .B1(_02437_),
    .B2(_02441_),
    .A2(_02418_),
    .A1(_02411_));
 sg13g2_a22oi_1 _09962_ (.Y(_02443_),
    .B1(_01630_),
    .B2(\i_time.mtime[21] ),
    .A2(_01629_),
    .A1(\i_time.mtime[22] ));
 sg13g2_a22oi_1 _09963_ (.Y(_02444_),
    .B1(\i_time.l_mtimecmp.data_out[20] ),
    .B2(_01534_),
    .A2(\i_time.l_mtimecmp.data_out[21] ),
    .A1(_01533_));
 sg13g2_a22oi_1 _09964_ (.Y(_02445_),
    .B1(_01634_),
    .B2(\i_time.mtime[16] ),
    .A2(_01633_),
    .A1(\i_time.mtime[17] ));
 sg13g2_nand2b_1 _09965_ (.Y(_02446_),
    .B(\i_time.mtime[19] ),
    .A_N(\i_time.l_mtimecmp.data_out[19] ));
 sg13g2_o21ai_1 _09966_ (.B1(_02446_),
    .Y(_02447_),
    .A1(\i_time.mtime[18] ),
    .A2(_01632_));
 sg13g2_nand2b_1 _09967_ (.Y(_02448_),
    .B(\i_time.l_mtimecmp.data_out[22] ),
    .A_N(\i_time.mtime[22] ));
 sg13g2_o21ai_1 _09968_ (.B1(_02448_),
    .Y(_02449_),
    .A1(\i_time.mtime[23] ),
    .A2(_01628_));
 sg13g2_nor2b_1 _09969_ (.A(\i_time.mtime[19] ),
    .B_N(\i_time.l_mtimecmp.data_out[19] ),
    .Y(_02450_));
 sg13g2_nor2_1 _09970_ (.A(_01535_),
    .B(\i_time.l_mtimecmp.data_out[18] ),
    .Y(_02451_));
 sg13g2_nor3_1 _09971_ (.A(_02449_),
    .B(_02450_),
    .C(_02451_),
    .Y(_02452_));
 sg13g2_nor2_1 _09972_ (.A(\i_time.mtime[17] ),
    .B(_01633_),
    .Y(_02453_));
 sg13g2_nand2_1 _09973_ (.Y(_02454_),
    .A(\i_time.mtime[20] ),
    .B(_01631_));
 sg13g2_nor2b_1 _09974_ (.A(_02453_),
    .B_N(_02454_),
    .Y(_02455_));
 sg13g2_nor2b_1 _09975_ (.A(\i_time.l_mtimecmp.data_out[23] ),
    .B_N(\i_time.mtime[23] ),
    .Y(_02456_));
 sg13g2_a21oi_1 _09976_ (.A1(_01536_),
    .A2(\i_time.l_mtimecmp.data_out[16] ),
    .Y(_02457_),
    .B1(_02456_));
 sg13g2_nand2_1 _09977_ (.Y(_02458_),
    .A(_02444_),
    .B(_02452_));
 sg13g2_nand4_1 _09978_ (.B(_02445_),
    .C(_02455_),
    .A(_02443_),
    .Y(_02459_),
    .D(_02457_));
 sg13g2_nor4_1 _09979_ (.A(_02442_),
    .B(_02447_),
    .C(_02458_),
    .D(_02459_),
    .Y(_02460_));
 sg13g2_nor3_1 _09980_ (.A(_02445_),
    .B(_02447_),
    .C(_02453_),
    .Y(_02461_));
 sg13g2_nor2_1 _09981_ (.A(_02451_),
    .B(_02461_),
    .Y(_02462_));
 sg13g2_or2_1 _09982_ (.X(_02463_),
    .B(_02462_),
    .A(_02450_));
 sg13g2_nand3_1 _09983_ (.B(_02454_),
    .C(_02463_),
    .A(_02446_),
    .Y(_02464_));
 sg13g2_nand2_1 _09984_ (.Y(_02465_),
    .A(_02444_),
    .B(_02464_));
 sg13g2_a21oi_1 _09985_ (.A1(_02443_),
    .A2(_02465_),
    .Y(_02466_),
    .B1(_02449_));
 sg13g2_nor3_1 _09986_ (.A(_02456_),
    .B(_02460_),
    .C(_02466_),
    .Y(_02467_));
 sg13g2_nor2_1 _09987_ (.A(\i_time.mtime[24] ),
    .B(_01627_),
    .Y(_02468_));
 sg13g2_o21ai_1 _09988_ (.B1(_02410_),
    .Y(_02469_),
    .A1(_02467_),
    .A2(_02468_));
 sg13g2_a22oi_1 _09989_ (.Y(_02470_),
    .B1(_02409_),
    .B2(_02469_),
    .A2(_02407_),
    .A1(_02406_));
 sg13g2_nor2_1 _09990_ (.A(\i_time.mtime[28] ),
    .B(_01625_),
    .Y(_02471_));
 sg13g2_a22oi_1 _09991_ (.Y(_02472_),
    .B1(_01625_),
    .B2(\i_time.mtime[28] ),
    .A2(_01624_),
    .A1(\i_time.mtime[29] ));
 sg13g2_o21ai_1 _09992_ (.B1(_02472_),
    .Y(_02473_),
    .A1(_02470_),
    .A2(_02471_));
 sg13g2_xor2_1 _09993_ (.B(\i_time.l_mtimecmp.data_out[31] ),
    .A(\i_time.mtime[31] ),
    .X(_02474_));
 sg13g2_a21o_1 _09994_ (.A2(_02473_),
    .A1(_02404_),
    .B1(_02474_),
    .X(_02475_));
 sg13g2_o21ai_1 _09995_ (.B1(_02475_),
    .Y(_02476_),
    .A1(\i_time.mtime[30] ),
    .A2(_01623_));
 sg13g2_a21oi_1 _09996_ (.A1(net3928),
    .A2(_01623_),
    .Y(_02477_),
    .B1(_02474_));
 sg13g2_a21oi_1 _09997_ (.A1(_02404_),
    .A2(_02473_),
    .Y(_02478_),
    .B1(_02477_));
 sg13g2_mux2_2 _09998_ (.A0(_02477_),
    .A1(_02478_),
    .S(_02476_),
    .X(_00063_));
 sg13g2_nand2b_2 _09999_ (.Y(_02479_),
    .B(net568),
    .A_N(_00119_));
 sg13g2_nand3b_1 _10000_ (.B(_01493_),
    .C(net571),
    .Y(_02480_),
    .A_N(\i_tinyqv.cpu.is_store ));
 sg13g2_and2_1 _10001_ (.A(_02479_),
    .B(_02480_),
    .X(_02481_));
 sg13g2_nor2_2 _10002_ (.A(_00120_),
    .B(_02171_),
    .Y(_02482_));
 sg13g2_nand2b_1 _10003_ (.Y(_02483_),
    .B(net457),
    .A_N(_00120_));
 sg13g2_nor3_1 _10004_ (.A(_01595_),
    .B(_02161_),
    .C(\i_tinyqv.cpu.i_core.cy_out ),
    .Y(_02484_));
 sg13g2_nand2b_1 _10005_ (.Y(_02485_),
    .B(_02162_),
    .A_N(_00125_));
 sg13g2_nand2b_1 _10006_ (.Y(_02486_),
    .B(_02348_),
    .A_N(_02485_));
 sg13g2_a21o_1 _10007_ (.A2(\i_tinyqv.cpu.i_core.cy_out ),
    .A1(_02350_),
    .B1(_02486_),
    .X(_02487_));
 sg13g2_o21ai_1 _10008_ (.B1(_02485_),
    .Y(_02488_),
    .A1(\i_tinyqv.cpu.i_core.cmp ),
    .A2(net315));
 sg13g2_nor2_1 _10009_ (.A(_02318_),
    .B(_02345_),
    .Y(_02489_));
 sg13g2_xnor2_1 _10010_ (.Y(_02490_),
    .A(_02318_),
    .B(_02345_));
 sg13g2_nand2_1 _10011_ (.Y(_02491_),
    .A(_02373_),
    .B(_02398_));
 sg13g2_xnor2_1 _10012_ (.Y(_02492_),
    .A(_02373_),
    .B(_02398_));
 sg13g2_nor2_1 _10013_ (.A(_02258_),
    .B(_02283_),
    .Y(_02493_));
 sg13g2_nand2_1 _10014_ (.Y(_02494_),
    .A(_02258_),
    .B(_02283_));
 sg13g2_nor2b_1 _10015_ (.A(_02493_),
    .B_N(_02494_),
    .Y(_02495_));
 sg13g2_nand2_1 _10016_ (.Y(_02496_),
    .A(_02178_),
    .B(_02223_));
 sg13g2_xor2_1 _10017_ (.B(_02222_),
    .A(_02178_),
    .X(_02497_));
 sg13g2_inv_1 _10018_ (.Y(_02498_),
    .A(_02497_));
 sg13g2_nor2_1 _10019_ (.A(_02488_),
    .B(_02495_),
    .Y(_02499_));
 sg13g2_nand4_1 _10020_ (.B(_02492_),
    .C(_02497_),
    .A(_02490_),
    .Y(_02500_),
    .D(_02499_));
 sg13g2_a22oi_1 _10021_ (.Y(_02501_),
    .B1(_02487_),
    .B2(_02500_),
    .A2(_02162_),
    .A1(net581));
 sg13g2_or2_2 _10022_ (.X(\i_tinyqv.cpu.i_core.cmp_out ),
    .B(_02501_),
    .A(_02484_));
 sg13g2_nor3_1 _10023_ (.A(_01595_),
    .B(_02484_),
    .C(_02501_),
    .Y(_02502_));
 sg13g2_o21ai_1 _10024_ (.B1(_02161_),
    .Y(_02503_),
    .A1(net581),
    .A2(_02500_));
 sg13g2_or2_1 _10025_ (.X(_02504_),
    .B(_02503_),
    .A(_01596_));
 sg13g2_nor2_2 _10026_ (.A(\i_tinyqv.cpu.alu_op[1] ),
    .B(net581),
    .Y(_02505_));
 sg13g2_nor2_2 _10027_ (.A(_01584_),
    .B(net574),
    .Y(_02506_));
 sg13g2_nand2_2 _10028_ (.Y(_02507_),
    .A(_01584_),
    .B(net581));
 sg13g2_nand2b_1 _10029_ (.Y(_02508_),
    .B(_02507_),
    .A_N(_02506_));
 sg13g2_nand2_2 _10030_ (.Y(_02509_),
    .A(net569),
    .B(\i_tinyqv.cpu.is_alu_imm ));
 sg13g2_o21ai_1 _10031_ (.B1(net569),
    .Y(_02510_),
    .A1(\i_tinyqv.cpu.is_alu_reg ),
    .A2(\i_tinyqv.cpu.is_alu_imm ));
 sg13g2_inv_1 _10032_ (.Y(_02511_),
    .A(_02510_));
 sg13g2_a21oi_1 _10033_ (.A1(_00122_),
    .A2(_02508_),
    .Y(_02512_),
    .B1(_02510_));
 sg13g2_o21ai_1 _10034_ (.B1(_02512_),
    .Y(_02513_),
    .A1(_00122_),
    .A2(_02508_));
 sg13g2_nor2_2 _10035_ (.A(_01493_),
    .B(_02479_),
    .Y(_02514_));
 sg13g2_nand3_1 _10036_ (.B(_02510_),
    .C(_02514_),
    .A(\i_tinyqv.cpu.i_core.load_done ),
    .Y(_02515_));
 sg13g2_nand3_1 _10037_ (.B(_02513_),
    .C(_02515_),
    .A(_02162_),
    .Y(_02516_));
 sg13g2_o21ai_1 _10038_ (.B1(_02516_),
    .Y(_02517_),
    .A1(_02502_),
    .A2(_02504_));
 sg13g2_o21ai_1 _10039_ (.B1(net570),
    .Y(_02518_),
    .A1(\i_tinyqv.cpu.is_jal ),
    .A2(\i_tinyqv.cpu.is_jalr ));
 sg13g2_nand2_2 _10040_ (.Y(_02519_),
    .A(net569),
    .B(\i_tinyqv.cpu.is_lui ));
 sg13g2_nand3_1 _10041_ (.B(_02518_),
    .C(_02519_),
    .A(_02157_),
    .Y(_02520_));
 sg13g2_and2_2 _10042_ (.A(\i_tinyqv.cpu.is_store ),
    .B(\i_tinyqv.cpu.no_write_in_progress ),
    .X(_02521_));
 sg13g2_nand2_2 _10043_ (.Y(_02522_),
    .A(\i_tinyqv.cpu.is_store ),
    .B(net3790));
 sg13g2_nand2_1 _10044_ (.Y(_02523_),
    .A(net570),
    .B(_02521_));
 sg13g2_and2_1 _10045_ (.A(net569),
    .B(\i_tinyqv.cpu.is_system ),
    .X(_02524_));
 sg13g2_nand2_2 _10046_ (.Y(_02525_),
    .A(net569),
    .B(\i_tinyqv.cpu.is_system ));
 sg13g2_nand4_1 _10047_ (.B(_00129_),
    .C(_02523_),
    .A(_01491_),
    .Y(_02526_),
    .D(_02525_));
 sg13g2_nor3_2 _10048_ (.A(_02481_),
    .B(_02520_),
    .C(_02526_),
    .Y(_02527_));
 sg13g2_a21oi_2 _10049_ (.B1(net314),
    .Y(_02528_),
    .A2(_02527_),
    .A1(_02517_));
 sg13g2_a221oi_1 _10050_ (.B2(_02527_),
    .C1(net313),
    .B1(_02517_),
    .A1(_02479_),
    .Y(_02529_),
    .A2(_02480_));
 sg13g2_a221oi_1 _10051_ (.B2(_02527_),
    .C1(net314),
    .B1(_02517_),
    .A1(net4133),
    .Y(_00065_),
    .A2(_02481_));
 sg13g2_and2_2 _10052_ (.A(\i_tinyqv.cpu.data_read_n[0] ),
    .B(\i_tinyqv.cpu.data_write_n[0] ),
    .X(_02530_));
 sg13g2_nand2_2 _10053_ (.Y(_02531_),
    .A(net3846),
    .B(\i_tinyqv.cpu.data_write_n[0] ));
 sg13g2_nand2_2 _10054_ (.Y(_02532_),
    .A(\i_tinyqv.cpu.data_read_n[1] ),
    .B(\i_tinyqv.cpu.data_write_n[1] ));
 sg13g2_and2_1 _10055_ (.A(net420),
    .B(_02532_),
    .X(_02533_));
 sg13g2_nand2_2 _10056_ (.Y(_02534_),
    .A(net420),
    .B(_02532_));
 sg13g2_nor2_2 _10057_ (.A(_02530_),
    .B(_02534_),
    .Y(_02535_));
 sg13g2_nand2_1 _10058_ (.Y(_02536_),
    .A(_02531_),
    .B(_02533_));
 sg13g2_nand2_1 _10059_ (.Y(_02537_),
    .A(net619),
    .B(_02533_));
 sg13g2_a21oi_1 _10060_ (.A1(_01609_),
    .A2(_02531_),
    .Y(_02538_),
    .B1(_02534_));
 sg13g2_o21ai_1 _10061_ (.B1(_02537_),
    .Y(_02539_),
    .A1(net619),
    .A2(_02538_));
 sg13g2_a21oi_2 _10062_ (.B1(_02539_),
    .Y(_02540_),
    .A2(_02536_),
    .A1(_00196_));
 sg13g2_and2_1 _10063_ (.A(net3854),
    .B(_02540_),
    .X(_00118_));
 sg13g2_and2_2 _10064_ (.A(_01596_),
    .B(_02365_),
    .X(_02541_));
 sg13g2_and2_1 _10065_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .B(net306),
    .X(_02542_));
 sg13g2_a21oi_2 _10066_ (.B1(_00122_),
    .Y(_02543_),
    .A2(_02155_),
    .A1(_02153_));
 sg13g2_and2_1 _10067_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .B(net311),
    .X(_02544_));
 sg13g2_a21oi_2 _10068_ (.B1(_00122_),
    .Y(_02545_),
    .A2(_02247_),
    .A1(_02244_));
 sg13g2_nand2_2 _10069_ (.Y(_02546_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .B(net302));
 sg13g2_nand2_1 _10070_ (.Y(_02547_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .B(net311));
 sg13g2_nor2_1 _10071_ (.A(_02546_),
    .B(_02547_),
    .Y(_02548_));
 sg13g2_nand2_1 _10072_ (.Y(_02549_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .B(net311));
 sg13g2_nand2_1 _10073_ (.Y(_02550_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .B(net302));
 sg13g2_xnor2_1 _10074_ (.Y(_02551_),
    .A(_02544_),
    .B(_02550_));
 sg13g2_nand4_1 _10075_ (.B(_02544_),
    .C(net302),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .Y(_02552_),
    .D(_02550_));
 sg13g2_inv_1 _10076_ (.Y(_02553_),
    .A(_02552_));
 sg13g2_xor2_1 _10077_ (.B(_02551_),
    .A(_02548_),
    .X(_02554_));
 sg13g2_xor2_1 _10078_ (.B(_02554_),
    .A(_02542_),
    .X(_02555_));
 sg13g2_nand2_1 _10079_ (.Y(_02556_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[2] ),
    .B(_02555_));
 sg13g2_xnor2_1 _10080_ (.Y(_02557_),
    .A(_02546_),
    .B(_02547_));
 sg13g2_inv_1 _10081_ (.Y(_02558_),
    .A(_02557_));
 sg13g2_nand3_1 _10082_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[0] ),
    .C(net302),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .Y(_02559_));
 sg13g2_xnor2_1 _10083_ (.Y(_02560_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[1] ),
    .B(_02557_));
 sg13g2_nor2b_1 _10084_ (.A(_02559_),
    .B_N(_02560_),
    .Y(_02561_));
 sg13g2_a21oi_1 _10085_ (.A1(\i_tinyqv.cpu.i_core.multiplier.accum[1] ),
    .A2(_02558_),
    .Y(_02562_),
    .B1(_02561_));
 sg13g2_xnor2_1 _10086_ (.Y(_02563_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[2] ),
    .B(_02555_));
 sg13g2_o21ai_1 _10087_ (.B1(_02556_),
    .Y(_02564_),
    .A1(_02562_),
    .A2(_02563_));
 sg13g2_a21oi_1 _10088_ (.A1(_02542_),
    .A2(_02554_),
    .Y(_02565_),
    .B1(_02553_));
 sg13g2_nand2_1 _10089_ (.Y(_02566_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .B(net306));
 sg13g2_a21oi_2 _10090_ (.B1(_00122_),
    .Y(_02567_),
    .A2(_02310_),
    .A1(_02308_));
 sg13g2_a22oi_1 _10091_ (.Y(_02568_),
    .B1(net308),
    .B2(_01649_),
    .A2(net302),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[3] ));
 sg13g2_nand4_1 _10092_ (.B(_01649_),
    .C(net302),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .Y(_02569_),
    .D(net308));
 sg13g2_nor2b_1 _10093_ (.A(_02568_),
    .B_N(_02569_),
    .Y(_02570_));
 sg13g2_nor2b_1 _10094_ (.A(_02549_),
    .B_N(_02546_),
    .Y(_02571_));
 sg13g2_xnor2_1 _10095_ (.Y(_02572_),
    .A(_02570_),
    .B(_02571_));
 sg13g2_xnor2_1 _10096_ (.Y(_02573_),
    .A(_02566_),
    .B(_02572_));
 sg13g2_nor2_1 _10097_ (.A(_02565_),
    .B(_02573_),
    .Y(_02574_));
 sg13g2_xor2_1 _10098_ (.B(_02573_),
    .A(_02565_),
    .X(_02575_));
 sg13g2_xnor2_1 _10099_ (.Y(_02576_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[3] ),
    .B(_02575_));
 sg13g2_nor2b_2 _10100_ (.A(_02576_),
    .B_N(_02564_),
    .Y(_02577_));
 sg13g2_a21oi_1 _10101_ (.A1(\i_tinyqv.cpu.i_core.multiplier.accum[3] ),
    .A2(_02575_),
    .Y(_02578_),
    .B1(_02574_));
 sg13g2_or3_1 _10102_ (.A(_02546_),
    .B(_02549_),
    .C(_02570_),
    .X(_02579_));
 sg13g2_o21ai_1 _10103_ (.B1(_02579_),
    .Y(_02580_),
    .A1(_02566_),
    .A2(_02572_));
 sg13g2_nand2_1 _10104_ (.Y(_02581_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .B(net306));
 sg13g2_nand2_1 _10105_ (.Y(_02582_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(net311));
 sg13g2_nand2_1 _10106_ (.Y(_02583_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .B(net308));
 sg13g2_and4_1 _10107_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .C(net302),
    .D(net308),
    .X(_02584_));
 sg13g2_a22oi_1 _10108_ (.Y(_02585_),
    .B1(net308),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .A2(net303),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[4] ));
 sg13g2_or3_1 _10109_ (.A(_02582_),
    .B(_02584_),
    .C(_02585_),
    .X(_02586_));
 sg13g2_o21ai_1 _10110_ (.B1(_02582_),
    .Y(_02587_),
    .A1(_02584_),
    .A2(_02585_));
 sg13g2_a21oi_1 _10111_ (.A1(_02549_),
    .A2(_02569_),
    .Y(_02588_),
    .B1(_02568_));
 sg13g2_and3_1 _10112_ (.X(_02589_),
    .A(_02586_),
    .B(_02587_),
    .C(_02588_));
 sg13g2_a21oi_1 _10113_ (.A1(_02586_),
    .A2(_02587_),
    .Y(_02590_),
    .B1(_02588_));
 sg13g2_or3_1 _10114_ (.A(_02581_),
    .B(_02589_),
    .C(_02590_),
    .X(_02591_));
 sg13g2_o21ai_1 _10115_ (.B1(_02581_),
    .Y(_02592_),
    .A1(_02589_),
    .A2(_02590_));
 sg13g2_nand3_1 _10116_ (.B(_02591_),
    .C(_02592_),
    .A(_02580_),
    .Y(_02593_));
 sg13g2_a21o_1 _10117_ (.A2(_02592_),
    .A1(_02591_),
    .B1(_02580_),
    .X(_02594_));
 sg13g2_and3_1 _10118_ (.X(_02595_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .B(_02593_),
    .C(_02594_));
 sg13g2_nand3_1 _10119_ (.B(_02593_),
    .C(_02594_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .Y(_02596_));
 sg13g2_a21oi_1 _10120_ (.A1(_02593_),
    .A2(_02594_),
    .Y(_02597_),
    .B1(net4128));
 sg13g2_nor3_1 _10121_ (.A(_02578_),
    .B(_02595_),
    .C(_02597_),
    .Y(_02598_));
 sg13g2_o21ai_1 _10122_ (.B1(_02578_),
    .Y(_02599_),
    .A1(_02595_),
    .A2(_02597_));
 sg13g2_nor2b_1 _10123_ (.A(_02598_),
    .B_N(_02599_),
    .Y(_02600_));
 sg13g2_xor2_1 _10124_ (.B(_02600_),
    .A(_02577_),
    .X(_00019_));
 sg13g2_a21oi_1 _10125_ (.A1(_02577_),
    .A2(_02599_),
    .Y(_02601_),
    .B1(_02598_));
 sg13g2_nand2b_1 _10126_ (.Y(_02602_),
    .B(_02591_),
    .A_N(_02589_));
 sg13g2_nand2_1 _10127_ (.Y(_02603_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(net306));
 sg13g2_nand2b_1 _10128_ (.Y(_02604_),
    .B(_02586_),
    .A_N(_02584_));
 sg13g2_nand2_1 _10129_ (.Y(_02605_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .B(net311));
 sg13g2_nand2_1 _10130_ (.Y(_02606_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .B(net310));
 sg13g2_and4_1 _10131_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .C(net303),
    .D(net308),
    .X(_02607_));
 sg13g2_a22oi_1 _10132_ (.Y(_02608_),
    .B1(net308),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .A2(net303),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[5] ));
 sg13g2_nor3_1 _10133_ (.A(_02605_),
    .B(_02607_),
    .C(_02608_),
    .Y(_02609_));
 sg13g2_o21ai_1 _10134_ (.B1(_02605_),
    .Y(_02610_),
    .A1(_02607_),
    .A2(_02608_));
 sg13g2_nor2b_1 _10135_ (.A(_02609_),
    .B_N(_02610_),
    .Y(_02611_));
 sg13g2_nand2_1 _10136_ (.Y(_02612_),
    .A(_02604_),
    .B(_02611_));
 sg13g2_xnor2_1 _10137_ (.Y(_02613_),
    .A(_02604_),
    .B(_02611_));
 sg13g2_xor2_1 _10138_ (.B(_02613_),
    .A(_02603_),
    .X(_02614_));
 sg13g2_nand2_1 _10139_ (.Y(_02615_),
    .A(_02602_),
    .B(_02614_));
 sg13g2_xnor2_1 _10140_ (.Y(_02616_),
    .A(_02602_),
    .B(_02614_));
 sg13g2_xnor2_1 _10141_ (.Y(_02617_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[5] ),
    .B(_02616_));
 sg13g2_nand2_1 _10142_ (.Y(_02618_),
    .A(_02593_),
    .B(_02596_));
 sg13g2_nor2_1 _10143_ (.A(_02617_),
    .B(_02618_),
    .Y(_02619_));
 sg13g2_xor2_1 _10144_ (.B(_02618_),
    .A(_02617_),
    .X(_02620_));
 sg13g2_xnor2_1 _10145_ (.Y(_00022_),
    .A(_02601_),
    .B(_02620_));
 sg13g2_o21ai_1 _10146_ (.B1(_02615_),
    .Y(_02621_),
    .A1(_01650_),
    .A2(_02616_));
 sg13g2_o21ai_1 _10147_ (.B1(_02612_),
    .Y(_02622_),
    .A1(_02603_),
    .A2(_02613_));
 sg13g2_nand2_1 _10148_ (.Y(_02623_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .B(net306));
 sg13g2_or2_1 _10149_ (.X(_02624_),
    .B(_02609_),
    .A(_02607_));
 sg13g2_nand2_1 _10150_ (.Y(_02625_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .B(net311));
 sg13g2_nand2_1 _10151_ (.Y(_02626_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .B(net309));
 sg13g2_nand2_1 _10152_ (.Y(_02627_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(net308));
 sg13g2_nand2_1 _10153_ (.Y(_02628_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .B(net303));
 sg13g2_xor2_1 _10154_ (.B(_02628_),
    .A(_02627_),
    .X(_02629_));
 sg13g2_nand2b_1 _10155_ (.Y(_02630_),
    .B(_02629_),
    .A_N(_02625_));
 sg13g2_xnor2_1 _10156_ (.Y(_02631_),
    .A(_02625_),
    .B(_02629_));
 sg13g2_nand2_1 _10157_ (.Y(_02632_),
    .A(_02624_),
    .B(_02631_));
 sg13g2_xnor2_1 _10158_ (.Y(_02633_),
    .A(_02624_),
    .B(_02631_));
 sg13g2_xor2_1 _10159_ (.B(_02633_),
    .A(_02623_),
    .X(_02634_));
 sg13g2_nand2_1 _10160_ (.Y(_02635_),
    .A(_02622_),
    .B(_02634_));
 sg13g2_xnor2_1 _10161_ (.Y(_02636_),
    .A(_02622_),
    .B(_02634_));
 sg13g2_xnor2_1 _10162_ (.Y(_02637_),
    .A(_01651_),
    .B(_02636_));
 sg13g2_nor2b_1 _10163_ (.A(_02637_),
    .B_N(_02621_),
    .Y(_02638_));
 sg13g2_xor2_1 _10164_ (.B(_02637_),
    .A(_02621_),
    .X(_02639_));
 sg13g2_a221oi_1 _10165_ (.B2(_02618_),
    .C1(_02598_),
    .B1(_02617_),
    .A1(_02577_),
    .Y(_02640_),
    .A2(_02599_));
 sg13g2_nor3_1 _10166_ (.A(_02619_),
    .B(_02639_),
    .C(_02640_),
    .Y(_02641_));
 sg13g2_o21ai_1 _10167_ (.B1(_02639_),
    .Y(_02642_),
    .A1(_02619_),
    .A2(_02640_));
 sg13g2_nor2b_1 _10168_ (.A(_02641_),
    .B_N(_02642_),
    .Y(_00023_));
 sg13g2_or2_1 _10169_ (.X(_02643_),
    .B(_02641_),
    .A(_02638_));
 sg13g2_o21ai_1 _10170_ (.B1(_02635_),
    .Y(_02644_),
    .A1(_01651_),
    .A2(_02636_));
 sg13g2_o21ai_1 _10171_ (.B1(_02632_),
    .Y(_02645_),
    .A1(_02623_),
    .A2(_02633_));
 sg13g2_nand2_1 _10172_ (.Y(_02646_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .B(net306));
 sg13g2_o21ai_1 _10173_ (.B1(_02630_),
    .Y(_02647_),
    .A1(_02627_),
    .A2(_02628_));
 sg13g2_nand2_1 _10174_ (.Y(_02648_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .B(net311));
 sg13g2_nand2_1 _10175_ (.Y(_02649_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .B(net309));
 sg13g2_nand2_1 _10176_ (.Y(_02650_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .B(net303));
 sg13g2_xor2_1 _10177_ (.B(_02650_),
    .A(_02583_),
    .X(_02651_));
 sg13g2_nand2b_1 _10178_ (.Y(_02652_),
    .B(_02651_),
    .A_N(_02648_));
 sg13g2_xnor2_1 _10179_ (.Y(_02653_),
    .A(_02648_),
    .B(_02651_));
 sg13g2_nand2_1 _10180_ (.Y(_02654_),
    .A(_02647_),
    .B(_02653_));
 sg13g2_xnor2_1 _10181_ (.Y(_02655_),
    .A(_02647_),
    .B(_02653_));
 sg13g2_xor2_1 _10182_ (.B(_02655_),
    .A(_02646_),
    .X(_02656_));
 sg13g2_nand2_1 _10183_ (.Y(_02657_),
    .A(_02645_),
    .B(_02656_));
 sg13g2_xnor2_1 _10184_ (.Y(_02658_),
    .A(_02645_),
    .B(_02656_));
 sg13g2_xnor2_1 _10185_ (.Y(_02659_),
    .A(_01652_),
    .B(_02658_));
 sg13g2_nor2b_1 _10186_ (.A(_02659_),
    .B_N(_02644_),
    .Y(_02660_));
 sg13g2_xnor2_1 _10187_ (.Y(_02661_),
    .A(_02644_),
    .B(_02659_));
 sg13g2_xor2_1 _10188_ (.B(_02661_),
    .A(_02643_),
    .X(_00024_));
 sg13g2_a21oi_1 _10189_ (.A1(_02643_),
    .A2(_02661_),
    .Y(_02662_),
    .B1(_02660_));
 sg13g2_o21ai_1 _10190_ (.B1(_02657_),
    .Y(_02663_),
    .A1(_01652_),
    .A2(_02658_));
 sg13g2_o21ai_1 _10191_ (.B1(_02654_),
    .Y(_02664_),
    .A1(_02646_),
    .A2(_02655_));
 sg13g2_nand2_1 _10192_ (.Y(_02665_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .B(net306));
 sg13g2_o21ai_1 _10193_ (.B1(_02652_),
    .Y(_02666_),
    .A1(_02583_),
    .A2(_02650_));
 sg13g2_nand2_1 _10194_ (.Y(_02667_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .B(net311));
 sg13g2_nand2_1 _10195_ (.Y(_02668_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .B(net309));
 sg13g2_nand2_1 _10196_ (.Y(_02669_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .B(_02545_));
 sg13g2_xor2_1 _10197_ (.B(_02669_),
    .A(_02606_),
    .X(_02670_));
 sg13g2_nand2b_1 _10198_ (.Y(_02671_),
    .B(_02670_),
    .A_N(_02667_));
 sg13g2_xnor2_1 _10199_ (.Y(_02672_),
    .A(_02667_),
    .B(_02670_));
 sg13g2_nand2_1 _10200_ (.Y(_02673_),
    .A(_02666_),
    .B(_02672_));
 sg13g2_xnor2_1 _10201_ (.Y(_02674_),
    .A(_02666_),
    .B(_02672_));
 sg13g2_xor2_1 _10202_ (.B(_02674_),
    .A(_02665_),
    .X(_02675_));
 sg13g2_nand2_1 _10203_ (.Y(_02676_),
    .A(_02664_),
    .B(_02675_));
 sg13g2_xnor2_1 _10204_ (.Y(_02677_),
    .A(_02664_),
    .B(_02675_));
 sg13g2_inv_1 _10205_ (.Y(_02678_),
    .A(_02677_));
 sg13g2_nand2_1 _10206_ (.Y(_02679_),
    .A(net3925),
    .B(_02678_));
 sg13g2_xor2_1 _10207_ (.B(_02677_),
    .A(net3925),
    .X(_02680_));
 sg13g2_nor2b_1 _10208_ (.A(_02680_),
    .B_N(_02663_),
    .Y(_02681_));
 sg13g2_xor2_1 _10209_ (.B(_02680_),
    .A(_02663_),
    .X(_02682_));
 sg13g2_nor2_1 _10210_ (.A(_02662_),
    .B(_02682_),
    .Y(_02683_));
 sg13g2_xor2_1 _10211_ (.B(_02682_),
    .A(_02662_),
    .X(_00025_));
 sg13g2_nor2_1 _10212_ (.A(_02681_),
    .B(_02683_),
    .Y(_02684_));
 sg13g2_o21ai_1 _10213_ (.B1(_02673_),
    .Y(_02685_),
    .A1(_02665_),
    .A2(_02674_));
 sg13g2_nand2_1 _10214_ (.Y(_02686_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .B(net305));
 sg13g2_o21ai_1 _10215_ (.B1(_02671_),
    .Y(_02687_),
    .A1(_02606_),
    .A2(_02669_));
 sg13g2_nand2_1 _10216_ (.Y(_02688_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .B(net312));
 sg13g2_nand2_1 _10217_ (.Y(_02689_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .B(net310));
 sg13g2_nand2_1 _10218_ (.Y(_02690_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .B(net304));
 sg13g2_xor2_1 _10219_ (.B(_02690_),
    .A(_02626_),
    .X(_02691_));
 sg13g2_nand2b_1 _10220_ (.Y(_02692_),
    .B(_02691_),
    .A_N(_02688_));
 sg13g2_xnor2_1 _10221_ (.Y(_02693_),
    .A(_02688_),
    .B(_02691_));
 sg13g2_nand2_1 _10222_ (.Y(_02694_),
    .A(_02687_),
    .B(_02693_));
 sg13g2_xnor2_1 _10223_ (.Y(_02695_),
    .A(_02687_),
    .B(_02693_));
 sg13g2_xor2_1 _10224_ (.B(_02695_),
    .A(_02686_),
    .X(_02696_));
 sg13g2_nand2_1 _10225_ (.Y(_02697_),
    .A(_02685_),
    .B(_02696_));
 sg13g2_xnor2_1 _10226_ (.Y(_02698_),
    .A(_02685_),
    .B(_02696_));
 sg13g2_xnor2_1 _10227_ (.Y(_02699_),
    .A(_01653_),
    .B(_02698_));
 sg13g2_nand3_1 _10228_ (.B(_02679_),
    .C(_02699_),
    .A(_02676_),
    .Y(_02700_));
 sg13g2_inv_1 _10229_ (.Y(_02701_),
    .A(_02700_));
 sg13g2_a21o_1 _10230_ (.A2(_02679_),
    .A1(_02676_),
    .B1(_02699_),
    .X(_02702_));
 sg13g2_nand2_1 _10231_ (.Y(_02703_),
    .A(_02700_),
    .B(_02702_));
 sg13g2_xor2_1 _10232_ (.B(_02703_),
    .A(_02684_),
    .X(_00026_));
 sg13g2_o21ai_1 _10233_ (.B1(_02697_),
    .Y(_02704_),
    .A1(_01653_),
    .A2(_02698_));
 sg13g2_o21ai_1 _10234_ (.B1(_02694_),
    .Y(_02705_),
    .A1(_02686_),
    .A2(_02695_));
 sg13g2_nand2_1 _10235_ (.Y(_02706_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .B(net305));
 sg13g2_o21ai_1 _10236_ (.B1(_02692_),
    .Y(_02707_),
    .A1(_02626_),
    .A2(_02690_));
 sg13g2_nand2_1 _10237_ (.Y(_02708_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .B(net312));
 sg13g2_nand2_1 _10238_ (.Y(_02709_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .B(net310));
 sg13g2_nand2_1 _10239_ (.Y(_02710_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .B(net304));
 sg13g2_xor2_1 _10240_ (.B(_02710_),
    .A(_02649_),
    .X(_02711_));
 sg13g2_nand2b_1 _10241_ (.Y(_02712_),
    .B(_02711_),
    .A_N(_02708_));
 sg13g2_xnor2_1 _10242_ (.Y(_02713_),
    .A(_02708_),
    .B(_02711_));
 sg13g2_nand2_1 _10243_ (.Y(_02714_),
    .A(_02707_),
    .B(_02713_));
 sg13g2_xnor2_1 _10244_ (.Y(_02715_),
    .A(_02707_),
    .B(_02713_));
 sg13g2_xor2_1 _10245_ (.B(_02715_),
    .A(_02706_),
    .X(_02716_));
 sg13g2_nand2_1 _10246_ (.Y(_02717_),
    .A(_02705_),
    .B(_02716_));
 sg13g2_xnor2_1 _10247_ (.Y(_02718_),
    .A(_02705_),
    .B(_02716_));
 sg13g2_inv_1 _10248_ (.Y(_02719_),
    .A(_02718_));
 sg13g2_nand2_1 _10249_ (.Y(_02720_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[10] ),
    .B(_02719_));
 sg13g2_xor2_1 _10250_ (.B(_02718_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[10] ),
    .X(_02721_));
 sg13g2_nor2b_1 _10251_ (.A(_02721_),
    .B_N(_02704_),
    .Y(_02722_));
 sg13g2_nand2b_1 _10252_ (.Y(_02723_),
    .B(_02721_),
    .A_N(_02704_));
 sg13g2_nand2b_1 _10253_ (.Y(_02724_),
    .B(_02723_),
    .A_N(_02722_));
 sg13g2_o21ai_1 _10254_ (.B1(_02702_),
    .Y(_02725_),
    .A1(_02684_),
    .A2(_02701_));
 sg13g2_xnor2_1 _10255_ (.Y(_00027_),
    .A(_02724_),
    .B(_02725_));
 sg13g2_a21o_1 _10256_ (.A2(_02725_),
    .A1(_02723_),
    .B1(_02722_),
    .X(_02726_));
 sg13g2_o21ai_1 _10257_ (.B1(_02714_),
    .Y(_02727_),
    .A1(_02706_),
    .A2(_02715_));
 sg13g2_nand2_1 _10258_ (.Y(_02728_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .B(net305));
 sg13g2_o21ai_1 _10259_ (.B1(_02712_),
    .Y(_02729_),
    .A1(_02649_),
    .A2(_02710_));
 sg13g2_nand2_1 _10260_ (.Y(_02730_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .B(net312));
 sg13g2_nand2_1 _10261_ (.Y(_02731_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .B(net309));
 sg13g2_nand2_1 _10262_ (.Y(_02732_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .B(net304));
 sg13g2_xor2_1 _10263_ (.B(_02732_),
    .A(_02668_),
    .X(_02733_));
 sg13g2_nand2b_1 _10264_ (.Y(_02734_),
    .B(_02733_),
    .A_N(_02730_));
 sg13g2_xnor2_1 _10265_ (.Y(_02735_),
    .A(_02730_),
    .B(_02733_));
 sg13g2_nand2_1 _10266_ (.Y(_02736_),
    .A(_02729_),
    .B(_02735_));
 sg13g2_xnor2_1 _10267_ (.Y(_02737_),
    .A(_02729_),
    .B(_02735_));
 sg13g2_xor2_1 _10268_ (.B(_02737_),
    .A(_02728_),
    .X(_02738_));
 sg13g2_nand2_1 _10269_ (.Y(_02739_),
    .A(_02727_),
    .B(_02738_));
 sg13g2_xnor2_1 _10270_ (.Y(_02740_),
    .A(_02727_),
    .B(_02738_));
 sg13g2_xnor2_1 _10271_ (.Y(_02741_),
    .A(_01654_),
    .B(_02740_));
 sg13g2_nand3_1 _10272_ (.B(_02720_),
    .C(_02741_),
    .A(_02717_),
    .Y(_02742_));
 sg13g2_a21oi_1 _10273_ (.A1(_02717_),
    .A2(_02720_),
    .Y(_02743_),
    .B1(_02741_));
 sg13g2_a21o_1 _10274_ (.A2(_02720_),
    .A1(_02717_),
    .B1(_02741_),
    .X(_02744_));
 sg13g2_nand2_1 _10275_ (.Y(_02745_),
    .A(_02742_),
    .B(_02744_));
 sg13g2_xnor2_1 _10276_ (.Y(_00028_),
    .A(_02726_),
    .B(_02745_));
 sg13g2_o21ai_1 _10277_ (.B1(_02739_),
    .Y(_02746_),
    .A1(_01654_),
    .A2(_02740_));
 sg13g2_o21ai_1 _10278_ (.B1(_02736_),
    .Y(_02747_),
    .A1(_02728_),
    .A2(_02737_));
 sg13g2_nand2_1 _10279_ (.Y(_02748_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .B(net305));
 sg13g2_o21ai_1 _10280_ (.B1(_02734_),
    .Y(_02749_),
    .A1(_02668_),
    .A2(_02732_));
 sg13g2_nand2_1 _10281_ (.Y(_02750_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .B(net312));
 sg13g2_nand2_2 _10282_ (.Y(_02751_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .B(net304));
 sg13g2_xor2_1 _10283_ (.B(_02751_),
    .A(_02689_),
    .X(_02752_));
 sg13g2_nand2b_1 _10284_ (.Y(_02753_),
    .B(_02752_),
    .A_N(_02750_));
 sg13g2_xnor2_1 _10285_ (.Y(_02754_),
    .A(_02750_),
    .B(_02752_));
 sg13g2_nand2_1 _10286_ (.Y(_02755_),
    .A(_02749_),
    .B(_02754_));
 sg13g2_xnor2_1 _10287_ (.Y(_02756_),
    .A(_02749_),
    .B(_02754_));
 sg13g2_xor2_1 _10288_ (.B(_02756_),
    .A(_02748_),
    .X(_02757_));
 sg13g2_nand2_1 _10289_ (.Y(_02758_),
    .A(_02747_),
    .B(_02757_));
 sg13g2_xnor2_1 _10290_ (.Y(_02759_),
    .A(_02747_),
    .B(_02757_));
 sg13g2_xnor2_1 _10291_ (.Y(_02760_),
    .A(_01655_),
    .B(_02759_));
 sg13g2_nor2b_1 _10292_ (.A(_02760_),
    .B_N(_02746_),
    .Y(_02761_));
 sg13g2_xor2_1 _10293_ (.B(_02760_),
    .A(_02746_),
    .X(_02762_));
 sg13g2_inv_1 _10294_ (.Y(_02763_),
    .A(_02762_));
 sg13g2_a21o_1 _10295_ (.A2(_02742_),
    .A1(_02726_),
    .B1(_02743_),
    .X(_02764_));
 sg13g2_xnor2_1 _10296_ (.Y(_00029_),
    .A(_02762_),
    .B(_02764_));
 sg13g2_a21oi_1 _10297_ (.A1(_02763_),
    .A2(_02764_),
    .Y(_02765_),
    .B1(_02761_));
 sg13g2_o21ai_1 _10298_ (.B1(_02758_),
    .Y(_02766_),
    .A1(_01655_),
    .A2(_02759_));
 sg13g2_o21ai_1 _10299_ (.B1(_02755_),
    .Y(_02767_),
    .A1(_02748_),
    .A2(_02756_));
 sg13g2_nand2_1 _10300_ (.Y(_02768_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .B(net305));
 sg13g2_o21ai_1 _10301_ (.B1(_02753_),
    .Y(_02769_),
    .A1(_02689_),
    .A2(_02751_));
 sg13g2_nand2_1 _10302_ (.Y(_02770_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .B(net312));
 sg13g2_nand2_1 _10303_ (.Y(_02771_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .B(net304));
 sg13g2_xor2_1 _10304_ (.B(_02771_),
    .A(_02709_),
    .X(_02772_));
 sg13g2_nand2b_1 _10305_ (.Y(_02773_),
    .B(_02772_),
    .A_N(_02770_));
 sg13g2_xnor2_1 _10306_ (.Y(_02774_),
    .A(_02770_),
    .B(_02772_));
 sg13g2_nand2_1 _10307_ (.Y(_02775_),
    .A(_02769_),
    .B(_02774_));
 sg13g2_xnor2_1 _10308_ (.Y(_02776_),
    .A(_02769_),
    .B(_02774_));
 sg13g2_xor2_1 _10309_ (.B(_02776_),
    .A(_02768_),
    .X(_02777_));
 sg13g2_nand2_1 _10310_ (.Y(_02778_),
    .A(_02767_),
    .B(_02777_));
 sg13g2_xnor2_1 _10311_ (.Y(_02779_),
    .A(_02767_),
    .B(_02777_));
 sg13g2_xnor2_1 _10312_ (.Y(_02780_),
    .A(_01656_),
    .B(_02779_));
 sg13g2_nand2b_1 _10313_ (.Y(_02781_),
    .B(_02766_),
    .A_N(_02780_));
 sg13g2_xor2_1 _10314_ (.B(_02780_),
    .A(_02766_),
    .X(_02782_));
 sg13g2_xor2_1 _10315_ (.B(_02782_),
    .A(_02765_),
    .X(_00030_));
 sg13g2_o21ai_1 _10316_ (.B1(_02781_),
    .Y(_02783_),
    .A1(_02765_),
    .A2(_02782_));
 sg13g2_o21ai_1 _10317_ (.B1(_02778_),
    .Y(_02784_),
    .A1(_01656_),
    .A2(_02779_));
 sg13g2_o21ai_1 _10318_ (.B1(_02775_),
    .Y(_02785_),
    .A1(_02768_),
    .A2(_02776_));
 sg13g2_nand2_1 _10319_ (.Y(_02786_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .B(net305));
 sg13g2_o21ai_1 _10320_ (.B1(_02773_),
    .Y(_02787_),
    .A1(_02709_),
    .A2(_02771_));
 sg13g2_nand2_1 _10321_ (.Y(_02788_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .B(net312));
 sg13g2_nand2_1 _10322_ (.Y(_02789_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .B(net304));
 sg13g2_xor2_1 _10323_ (.B(_02789_),
    .A(_02731_),
    .X(_02790_));
 sg13g2_nand2b_1 _10324_ (.Y(_02791_),
    .B(_02790_),
    .A_N(_02788_));
 sg13g2_xnor2_1 _10325_ (.Y(_02792_),
    .A(_02788_),
    .B(_02790_));
 sg13g2_nand2_1 _10326_ (.Y(_02793_),
    .A(_02787_),
    .B(_02792_));
 sg13g2_xnor2_1 _10327_ (.Y(_02794_),
    .A(_02787_),
    .B(_02792_));
 sg13g2_xor2_1 _10328_ (.B(_02794_),
    .A(_02786_),
    .X(_02795_));
 sg13g2_nand2_1 _10329_ (.Y(_02796_),
    .A(_02785_),
    .B(_02795_));
 sg13g2_xnor2_1 _10330_ (.Y(_02797_),
    .A(_02785_),
    .B(_02795_));
 sg13g2_xnor2_1 _10331_ (.Y(_02798_),
    .A(_01658_),
    .B(_02797_));
 sg13g2_nor2b_1 _10332_ (.A(_02798_),
    .B_N(_02784_),
    .Y(_02799_));
 sg13g2_xor2_1 _10333_ (.B(_02798_),
    .A(_02784_),
    .X(_02800_));
 sg13g2_inv_1 _10334_ (.Y(_02801_),
    .A(_02800_));
 sg13g2_xnor2_1 _10335_ (.Y(_00020_),
    .A(_02783_),
    .B(_02800_));
 sg13g2_a21o_1 _10336_ (.A2(_02801_),
    .A1(_02783_),
    .B1(_02799_),
    .X(_02802_));
 sg13g2_o21ai_1 _10337_ (.B1(_02796_),
    .Y(_02803_),
    .A1(_01658_),
    .A2(_02797_));
 sg13g2_o21ai_1 _10338_ (.B1(_02793_),
    .Y(_02804_),
    .A1(_02786_),
    .A2(_02794_));
 sg13g2_nand2_1 _10339_ (.Y(_02805_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .B(_02541_));
 sg13g2_o21ai_1 _10340_ (.B1(_02791_),
    .Y(_02806_),
    .A1(_02731_),
    .A2(_02789_));
 sg13g2_nand2_1 _10341_ (.Y(_02807_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .B(net312));
 sg13g2_nand2_2 _10342_ (.Y(_02808_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[15] ),
    .B(net309));
 sg13g2_nor2_1 _10343_ (.A(_02751_),
    .B(_02808_),
    .Y(_02809_));
 sg13g2_a22oi_1 _10344_ (.Y(_02810_),
    .B1(net309),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .A2(net304),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[15] ));
 sg13g2_nor2_1 _10345_ (.A(_02809_),
    .B(_02810_),
    .Y(_02811_));
 sg13g2_nand2b_1 _10346_ (.Y(_02812_),
    .B(_02811_),
    .A_N(_02807_));
 sg13g2_xnor2_1 _10347_ (.Y(_02813_),
    .A(_02807_),
    .B(_02811_));
 sg13g2_nand2_1 _10348_ (.Y(_02814_),
    .A(_02806_),
    .B(_02813_));
 sg13g2_xnor2_1 _10349_ (.Y(_02815_),
    .A(_02806_),
    .B(_02813_));
 sg13g2_xor2_1 _10350_ (.B(_02815_),
    .A(_02805_),
    .X(_02816_));
 sg13g2_nand2_1 _10351_ (.Y(_02817_),
    .A(_02804_),
    .B(_02816_));
 sg13g2_xnor2_1 _10352_ (.Y(_02818_),
    .A(_02804_),
    .B(_02816_));
 sg13g2_inv_1 _10353_ (.Y(_02819_),
    .A(_02818_));
 sg13g2_nand2_1 _10354_ (.Y(_02820_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[15] ),
    .B(_02819_));
 sg13g2_xor2_1 _10355_ (.B(_02818_),
    .A(net4130),
    .X(_02821_));
 sg13g2_nand2b_1 _10356_ (.Y(_02822_),
    .B(_02803_),
    .A_N(_02821_));
 sg13g2_xor2_1 _10357_ (.B(_02821_),
    .A(_02803_),
    .X(_02823_));
 sg13g2_nand2b_1 _10358_ (.Y(_02824_),
    .B(_02802_),
    .A_N(_02823_));
 sg13g2_xnor2_1 _10359_ (.Y(_00021_),
    .A(_02802_),
    .B(_02823_));
 sg13g2_mux2_2 _10360_ (.A0(\i_uart_tx.txd_reg ),
    .A1(\gpio_out[0] ),
    .S(\gpio_out_sel[0] ),
    .X(uo_out[0]));
 sg13g2_mux2_1 _10361_ (.A0(\i_spi.spi_select ),
    .A1(\debug_rd_r[2] ),
    .S(debug_register_data),
    .X(_02825_));
 sg13g2_mux2_2 _10362_ (.A0(_02825_),
    .A1(\gpio_out[4] ),
    .S(\gpio_out_sel[4] ),
    .X(uo_out[4]));
 sg13g2_nand2_2 _10363_ (.Y(_02826_),
    .A(_02157_),
    .B(_02510_));
 sg13g2_nor2b_2 _10364_ (.A(\i_tinyqv.cpu.i_core.cycle[1] ),
    .B_N(\i_tinyqv.cpu.i_core.cycle[0] ),
    .Y(_02827_));
 sg13g2_nand2b_2 _10365_ (.Y(_02828_),
    .B(\i_tinyqv.cpu.i_core.cycle[0] ),
    .A_N(\i_tinyqv.cpu.i_core.cycle[1] ));
 sg13g2_nand2_2 _10366_ (.Y(_02829_),
    .A(_02161_),
    .B(_02827_));
 sg13g2_and2_2 _10367_ (.A(\i_tinyqv.cpu.alu_op[3] ),
    .B(_02506_),
    .X(_02830_));
 sg13g2_nand2_1 _10368_ (.Y(_02831_),
    .A(\i_tinyqv.cpu.alu_op[3] ),
    .B(_02506_));
 sg13g2_nand2_1 _10369_ (.Y(_02832_),
    .A(_00125_),
    .B(_01595_));
 sg13g2_nand4_1 _10370_ (.B(_01595_),
    .C(_00130_),
    .A(_00125_),
    .Y(_02833_),
    .D(_02162_));
 sg13g2_a21oi_1 _10371_ (.A1(_02288_),
    .A2(_02292_),
    .Y(_02834_),
    .B1(_02833_));
 sg13g2_o21ai_1 _10372_ (.B1(_02834_),
    .Y(_02835_),
    .A1(_02288_),
    .A2(_02292_));
 sg13g2_o21ai_1 _10373_ (.B1(_02162_),
    .Y(_02836_),
    .A1(_00130_),
    .A2(_02832_));
 sg13g2_nor2_2 _10374_ (.A(_00130_),
    .B(_02485_),
    .Y(_02837_));
 sg13g2_nand2_1 _10375_ (.Y(_02838_),
    .A(net581),
    .B(_02494_));
 sg13g2_a22oi_1 _10376_ (.Y(_02839_),
    .B1(_02837_),
    .B2(_02838_),
    .A2(_02836_),
    .A1(_02494_));
 sg13g2_o21ai_1 _10377_ (.B1(_02835_),
    .Y(_02840_),
    .A1(_02493_),
    .A2(_02839_));
 sg13g2_nor2_1 _10378_ (.A(_02507_),
    .B(_02828_),
    .Y(_02841_));
 sg13g2_nand2b_2 _10379_ (.Y(_02842_),
    .B(_02827_),
    .A_N(_02507_));
 sg13g2_a21o_1 _10380_ (.A2(net302),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[0] ),
    .X(_02843_));
 sg13g2_a21oi_1 _10381_ (.A1(_02559_),
    .A2(_02843_),
    .Y(_02844_),
    .B1(net406));
 sg13g2_o21ai_1 _10382_ (.B1(_02842_),
    .Y(_02845_),
    .A1(_02830_),
    .A2(_02840_));
 sg13g2_nand2_1 _10383_ (.Y(_02846_),
    .A(\i_tinyqv.cpu.alu_op[3] ),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[31] ));
 sg13g2_xnor2_1 _10384_ (.Y(_02847_),
    .A(net586),
    .B(net575));
 sg13g2_nor2_1 _10385_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .B(_02847_),
    .Y(_02848_));
 sg13g2_nand2_1 _10386_ (.Y(_02849_),
    .A(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .B(_02847_));
 sg13g2_xnor2_1 _10387_ (.Y(_02850_),
    .A(net589),
    .B(net575));
 sg13g2_xnor2_1 _10388_ (.Y(_02851_),
    .A(net596),
    .B(net575));
 sg13g2_nand2_2 _10389_ (.Y(_02852_),
    .A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .B(_02851_));
 sg13g2_xor2_1 _10390_ (.B(_02850_),
    .A(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .X(_02853_));
 sg13g2_nor2b_1 _10391_ (.A(_02852_),
    .B_N(_02853_),
    .Y(_02854_));
 sg13g2_a21oi_2 _10392_ (.B1(_02854_),
    .Y(_02855_),
    .A2(_02850_),
    .A1(\i_tinyqv.cpu.i_core.i_shift.b[3] ));
 sg13g2_o21ai_1 _10393_ (.B1(_02849_),
    .Y(_02856_),
    .A1(_02848_),
    .A2(_02855_));
 sg13g2_and2_1 _10394_ (.A(_02846_),
    .B(_02856_),
    .X(_02857_));
 sg13g2_nor2b_1 _10395_ (.A(net578),
    .B_N(_00229_),
    .Y(_02858_));
 sg13g2_a21oi_1 _10396_ (.A1(net578),
    .A2(_00228_),
    .Y(_02859_),
    .B1(_02858_));
 sg13g2_mux2_1 _10397_ (.A0(_00227_),
    .A1(_00226_),
    .S(net578),
    .X(_02860_));
 sg13g2_nand2_1 _10398_ (.Y(_02861_),
    .A(net629),
    .B(_02860_));
 sg13g2_o21ai_1 _10399_ (.B1(_02861_),
    .Y(_02862_),
    .A1(net629),
    .A2(_02859_));
 sg13g2_nand2_1 _10400_ (.Y(_02863_),
    .A(net624),
    .B(_02862_));
 sg13g2_xnor2_1 _10401_ (.Y(_02864_),
    .A(_01668_),
    .B(_02851_));
 sg13g2_xnor2_1 _10402_ (.Y(_02865_),
    .A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .B(_02851_));
 sg13g2_nor2b_1 _10403_ (.A(net579),
    .B_N(_00233_),
    .Y(_02866_));
 sg13g2_a21oi_1 _10404_ (.A1(net579),
    .A2(_00232_),
    .Y(_02867_),
    .B1(_02866_));
 sg13g2_mux2_1 _10405_ (.A0(_00231_),
    .A1(_00230_),
    .S(net578),
    .X(_02868_));
 sg13g2_nand2_1 _10406_ (.Y(_02869_),
    .A(net628),
    .B(_02868_));
 sg13g2_o21ai_1 _10407_ (.B1(_02869_),
    .Y(_02870_),
    .A1(net628),
    .A2(_02867_));
 sg13g2_a21oi_1 _10408_ (.A1(net502),
    .A2(_02870_),
    .Y(_02871_),
    .B1(net352));
 sg13g2_xnor2_1 _10409_ (.Y(_02872_),
    .A(_02852_),
    .B(_02853_));
 sg13g2_xor2_1 _10410_ (.B(_02853_),
    .A(_02852_),
    .X(_02873_));
 sg13g2_mux4_1 _10411_ (.S0(net577),
    .A0(_00221_),
    .A1(_00220_),
    .A2(_00219_),
    .A3(_00218_),
    .S1(net631),
    .X(_02874_));
 sg13g2_nand2_1 _10412_ (.Y(_02875_),
    .A(net622),
    .B(_02874_));
 sg13g2_mux4_1 _10413_ (.S0(net577),
    .A0(_00225_),
    .A1(_00224_),
    .A2(_00223_),
    .A3(_00222_),
    .S1(net630),
    .X(_02876_));
 sg13g2_a21oi_1 _10414_ (.A1(net502),
    .A2(_02876_),
    .Y(_02877_),
    .B1(net349));
 sg13g2_a221oi_1 _10415_ (.B2(_02877_),
    .C1(_02872_),
    .B1(_02875_),
    .A1(_02863_),
    .Y(_02878_),
    .A2(_02871_));
 sg13g2_nand2b_1 _10416_ (.Y(_02879_),
    .B(_02849_),
    .A_N(_02848_));
 sg13g2_and2_2 _10417_ (.A(_02855_),
    .B(_02879_),
    .X(_02880_));
 sg13g2_nand2_2 _10418_ (.Y(_02881_),
    .A(_02855_),
    .B(_02879_));
 sg13g2_mux2_1 _10419_ (.A0(_00209_),
    .A1(_00208_),
    .S(net580),
    .X(_02882_));
 sg13g2_mux2_1 _10420_ (.A0(_00235_),
    .A1(_00234_),
    .S(net573),
    .X(_02883_));
 sg13g2_mux2_1 _10421_ (.A0(_02882_),
    .A1(_02883_),
    .S(net625),
    .X(_02884_));
 sg13g2_nand2_1 _10422_ (.Y(_02885_),
    .A(net501),
    .B(_02884_));
 sg13g2_nor2b_1 _10423_ (.A(net573),
    .B_N(_00237_),
    .Y(_02886_));
 sg13g2_a21oi_1 _10424_ (.A1(net573),
    .A2(_00236_),
    .Y(_02887_),
    .B1(_02886_));
 sg13g2_nand2_1 _10425_ (.Y(_02888_),
    .A(net573),
    .B(_00238_));
 sg13g2_o21ai_1 _10426_ (.B1(_02888_),
    .Y(_02889_),
    .A1(net573),
    .A2(_01649_));
 sg13g2_nand2_1 _10427_ (.Y(_02890_),
    .A(net626),
    .B(_02889_));
 sg13g2_o21ai_1 _10428_ (.B1(_02890_),
    .Y(_02891_),
    .A1(net625),
    .A2(_02887_));
 sg13g2_a21oi_1 _10429_ (.A1(net624),
    .A2(_02891_),
    .Y(_02892_),
    .B1(net350));
 sg13g2_mux2_1 _10430_ (.A0(_00213_),
    .A1(_00212_),
    .S(net575),
    .X(_02893_));
 sg13g2_nor2_1 _10431_ (.A(net627),
    .B(_02893_),
    .Y(_02894_));
 sg13g2_nor2b_1 _10432_ (.A(net575),
    .B_N(_00211_),
    .Y(_02895_));
 sg13g2_a21oi_1 _10433_ (.A1(net575),
    .A2(_00210_),
    .Y(_02896_),
    .B1(_02895_));
 sg13g2_a21oi_1 _10434_ (.A1(net627),
    .A2(_02896_),
    .Y(_02897_),
    .B1(_02894_));
 sg13g2_nand2_1 _10435_ (.Y(_02898_),
    .A(net621),
    .B(_02897_));
 sg13g2_mux4_1 _10436_ (.S0(net576),
    .A0(_00217_),
    .A1(_00216_),
    .A2(_00215_),
    .A3(_00214_),
    .S1(net631),
    .X(_02899_));
 sg13g2_a21oi_1 _10437_ (.A1(net504),
    .A2(_02899_),
    .Y(_02900_),
    .B1(net351));
 sg13g2_a221oi_1 _10438_ (.B2(_02900_),
    .C1(_02873_),
    .B1(_02898_),
    .A1(_02885_),
    .Y(_02901_),
    .A2(_02892_));
 sg13g2_nor3_1 _10439_ (.A(_02878_),
    .B(_02880_),
    .C(_02901_),
    .Y(_02902_));
 sg13g2_mux4_1 _10440_ (.S0(net575),
    .A0(_00210_),
    .A1(_00211_),
    .A2(_00212_),
    .A3(_00213_),
    .S1(net627),
    .X(_02903_));
 sg13g2_mux4_1 _10441_ (.S0(net576),
    .A0(_00214_),
    .A1(_00215_),
    .A2(_00216_),
    .A3(_00217_),
    .S1(net631),
    .X(_02904_));
 sg13g2_mux4_1 _10442_ (.S0(net572),
    .A0(_00234_),
    .A1(_00235_),
    .A2(_00208_),
    .A3(_00209_),
    .S1(net626),
    .X(_02905_));
 sg13g2_mux4_1 _10443_ (.S0(net626),
    .A0(_00238_),
    .A1(_00236_),
    .A2(_00206_),
    .A3(_00237_),
    .S1(net573),
    .X(_02906_));
 sg13g2_mux4_1 _10444_ (.S0(net621),
    .A0(_02903_),
    .A1(_02904_),
    .A2(_02906_),
    .A3(_02905_),
    .S1(net350),
    .X(_02907_));
 sg13g2_mux2_1 _10445_ (.A0(_00230_),
    .A1(_00231_),
    .S(net578),
    .X(_02908_));
 sg13g2_mux2_1 _10446_ (.A0(_00232_),
    .A1(_00233_),
    .S(net579),
    .X(_02909_));
 sg13g2_mux2_1 _10447_ (.A0(_02908_),
    .A1(_02909_),
    .S(net628),
    .X(_02910_));
 sg13g2_inv_1 _10448_ (.Y(_02911_),
    .A(_02910_));
 sg13g2_mux2_1 _10449_ (.A0(_00226_),
    .A1(_00227_),
    .S(net579),
    .X(_02912_));
 sg13g2_nor2_1 _10450_ (.A(net629),
    .B(_02912_),
    .Y(_02913_));
 sg13g2_nor2b_1 _10451_ (.A(net578),
    .B_N(_00228_),
    .Y(_02914_));
 sg13g2_a21oi_1 _10452_ (.A1(net578),
    .A2(_00229_),
    .Y(_02915_),
    .B1(_02914_));
 sg13g2_a21oi_2 _10453_ (.B1(_02913_),
    .Y(_02916_),
    .A2(_02915_),
    .A1(net628));
 sg13g2_a21oi_1 _10454_ (.A1(net502),
    .A2(_02916_),
    .Y(_02917_),
    .B1(net350));
 sg13g2_o21ai_1 _10455_ (.B1(_02917_),
    .Y(_02918_),
    .A1(net502),
    .A2(_02911_));
 sg13g2_mux4_1 _10456_ (.S0(net577),
    .A0(_00218_),
    .A1(_00219_),
    .A2(_00220_),
    .A3(_00221_),
    .S1(net631),
    .X(_02919_));
 sg13g2_mux4_1 _10457_ (.S0(net577),
    .A0(_00222_),
    .A1(_00223_),
    .A2(_00224_),
    .A3(_00225_),
    .S1(net630),
    .X(_02920_));
 sg13g2_nand2_1 _10458_ (.Y(_02921_),
    .A(net622),
    .B(_02920_));
 sg13g2_a21oi_1 _10459_ (.A1(net504),
    .A2(_02919_),
    .Y(_02922_),
    .B1(net352));
 sg13g2_a21oi_1 _10460_ (.A1(_02921_),
    .A2(_02922_),
    .Y(_02923_),
    .B1(_02873_));
 sg13g2_a221oi_1 _10461_ (.B2(_02923_),
    .C1(_02881_),
    .B1(_02918_),
    .A1(_02873_),
    .Y(_02924_),
    .A2(_02907_));
 sg13g2_nor3_1 _10462_ (.A(_02856_),
    .B(_02902_),
    .C(_02924_),
    .Y(_02925_));
 sg13g2_or2_1 _10463_ (.X(_02926_),
    .B(_02925_),
    .A(_02857_));
 sg13g2_mux4_1 _10464_ (.S0(net577),
    .A0(_00227_),
    .A1(_00226_),
    .A2(_00225_),
    .A3(_00224_),
    .S1(net629),
    .X(_02927_));
 sg13g2_and2_1 _10465_ (.A(net503),
    .B(_02927_),
    .X(_02928_));
 sg13g2_mux4_1 _10466_ (.S0(net577),
    .A0(_00223_),
    .A1(_00222_),
    .A2(_00221_),
    .A3(_00220_),
    .S1(net630),
    .X(_02929_));
 sg13g2_a21oi_1 _10467_ (.A1(net623),
    .A2(_02929_),
    .Y(_02930_),
    .B1(_02928_));
 sg13g2_mux4_1 _10468_ (.S0(net577),
    .A0(_00219_),
    .A1(_00218_),
    .A2(_00217_),
    .A3(_00216_),
    .S1(net631),
    .X(_02931_));
 sg13g2_nand2_1 _10469_ (.Y(_02932_),
    .A(net504),
    .B(_02931_));
 sg13g2_mux4_1 _10470_ (.S0(net576),
    .A0(_00215_),
    .A1(_00214_),
    .A2(_00213_),
    .A3(_00212_),
    .S1(net627),
    .X(_02933_));
 sg13g2_a21oi_1 _10471_ (.A1(net623),
    .A2(_02933_),
    .Y(_02934_),
    .B1(net349));
 sg13g2_a221oi_1 _10472_ (.B2(_02934_),
    .C1(_02880_),
    .B1(_02932_),
    .A1(net349),
    .Y(_02935_),
    .A2(_02930_));
 sg13g2_mux4_1 _10473_ (.S0(net575),
    .A0(_00208_),
    .A1(_00209_),
    .A2(_00210_),
    .A3(_00211_),
    .S1(net625),
    .X(_02936_));
 sg13g2_mux4_1 _10474_ (.S0(net576),
    .A0(_00212_),
    .A1(_00213_),
    .A2(_00214_),
    .A3(_00215_),
    .S1(net627),
    .X(_02937_));
 sg13g2_nand2_1 _10475_ (.Y(_02938_),
    .A(net621),
    .B(_02937_));
 sg13g2_a21oi_1 _10476_ (.A1(net504),
    .A2(_02936_),
    .Y(_02939_),
    .B1(net351));
 sg13g2_mux4_1 _10477_ (.S0(net577),
    .A0(_00220_),
    .A1(_00221_),
    .A2(_00222_),
    .A3(_00223_),
    .S1(net630),
    .X(_02940_));
 sg13g2_mux4_1 _10478_ (.S0(net576),
    .A0(_00216_),
    .A1(_00217_),
    .A2(_00218_),
    .A3(_00219_),
    .S1(net631),
    .X(_02941_));
 sg13g2_nand2_1 _10479_ (.Y(_02942_),
    .A(net504),
    .B(_02941_));
 sg13g2_a21oi_1 _10480_ (.A1(net623),
    .A2(_02940_),
    .Y(_02943_),
    .B1(net349));
 sg13g2_a221oi_1 _10481_ (.B2(_02943_),
    .C1(_02881_),
    .B1(_02942_),
    .A1(_02938_),
    .Y(_02944_),
    .A2(_02939_));
 sg13g2_nor3_1 _10482_ (.A(_02872_),
    .B(_02935_),
    .C(_02944_),
    .Y(_02945_));
 sg13g2_nand2_1 _10483_ (.Y(_02946_),
    .A(net625),
    .B(_02882_));
 sg13g2_o21ai_1 _10484_ (.B1(_02946_),
    .Y(_02947_),
    .A1(net627),
    .A2(_02896_));
 sg13g2_nor2_1 _10485_ (.A(net625),
    .B(_02883_),
    .Y(_02948_));
 sg13g2_a21oi_1 _10486_ (.A1(net625),
    .A2(_02887_),
    .Y(_02949_),
    .B1(_02948_));
 sg13g2_nand2_1 _10487_ (.Y(_02950_),
    .A(net621),
    .B(_02949_));
 sg13g2_a21oi_1 _10488_ (.A1(net501),
    .A2(_02947_),
    .Y(_02951_),
    .B1(net351));
 sg13g2_nand3_1 _10489_ (.B(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .C(net625),
    .A(\i_tinyqv.cpu.alu_op[3] ),
    .Y(_02952_));
 sg13g2_o21ai_1 _10490_ (.B1(_02952_),
    .Y(_02953_),
    .A1(net625),
    .A2(_02889_));
 sg13g2_nand2b_1 _10491_ (.Y(_02954_),
    .B(net505),
    .A_N(_02953_));
 sg13g2_a21oi_1 _10492_ (.A1(net624),
    .A2(_02846_),
    .Y(_02955_),
    .B1(net350));
 sg13g2_a221oi_1 _10493_ (.B2(_02955_),
    .C1(_02880_),
    .B1(_02954_),
    .A1(_02950_),
    .Y(_02956_),
    .A2(_02951_));
 sg13g2_nand2_1 _10494_ (.Y(_02957_),
    .A(net628),
    .B(_02908_));
 sg13g2_o21ai_1 _10495_ (.B1(_02957_),
    .Y(_02958_),
    .A1(net629),
    .A2(_02915_));
 sg13g2_nand2_1 _10496_ (.Y(_02959_),
    .A(net622),
    .B(_02958_));
 sg13g2_mux4_1 _10497_ (.S0(net578),
    .A0(_00224_),
    .A1(_00225_),
    .A2(_00226_),
    .A3(_00227_),
    .S1(net629),
    .X(_02960_));
 sg13g2_a21oi_1 _10498_ (.A1(net502),
    .A2(_02960_),
    .Y(_02961_),
    .B1(net352));
 sg13g2_nor2_1 _10499_ (.A(net628),
    .B(_02868_),
    .Y(_02962_));
 sg13g2_a21oi_1 _10500_ (.A1(net629),
    .A2(_02859_),
    .Y(_02963_),
    .B1(_02962_));
 sg13g2_and2_1 _10501_ (.A(net623),
    .B(_02963_),
    .X(_02964_));
 sg13g2_nor2_1 _10502_ (.A(net628),
    .B(_02909_),
    .Y(_02965_));
 sg13g2_a21oi_1 _10503_ (.A1(net628),
    .A2(_02867_),
    .Y(_02966_),
    .B1(_02965_));
 sg13g2_a21oi_1 _10504_ (.A1(net503),
    .A2(_02966_),
    .Y(_02967_),
    .B1(_02964_));
 sg13g2_a221oi_1 _10505_ (.B2(net352),
    .C1(_02881_),
    .B1(_02967_),
    .A1(_02959_),
    .Y(_02968_),
    .A2(_02961_));
 sg13g2_nor3_1 _10506_ (.A(_02873_),
    .B(_02956_),
    .C(_02968_),
    .Y(_02969_));
 sg13g2_nor3_1 _10507_ (.A(_02856_),
    .B(_02945_),
    .C(_02969_),
    .Y(_02970_));
 sg13g2_nor2_1 _10508_ (.A(_02857_),
    .B(_02970_),
    .Y(_02971_));
 sg13g2_or2_1 _10509_ (.X(_02972_),
    .B(_02971_),
    .A(net572));
 sg13g2_a21oi_1 _10510_ (.A1(net572),
    .A2(_02926_),
    .Y(_02973_),
    .B1(_02842_));
 sg13g2_and4_1 _10511_ (.A(_01583_),
    .B(net316),
    .C(_02506_),
    .D(_02827_),
    .X(_02974_));
 sg13g2_a21oi_1 _10512_ (.A1(_02972_),
    .A2(_02973_),
    .Y(_02975_),
    .B1(_02974_));
 sg13g2_o21ai_1 _10513_ (.B1(_02975_),
    .Y(_02976_),
    .A1(_02844_),
    .A2(_02845_));
 sg13g2_nand2b_1 _10514_ (.Y(_02977_),
    .B(_02974_),
    .A_N(\i_tinyqv.cpu.i_core.cmp ));
 sg13g2_nand3_1 _10515_ (.B(_02976_),
    .C(_02977_),
    .A(_02162_),
    .Y(_02978_));
 sg13g2_o21ai_1 _10516_ (.B1(_02978_),
    .Y(_02979_),
    .A1(_00206_),
    .A2(_02829_));
 sg13g2_nand2_1 _10517_ (.Y(_02980_),
    .A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .B(_02540_));
 sg13g2_a21oi_2 _10518_ (.B1(_01604_),
    .Y(_02981_),
    .A2(_02980_),
    .A1(_00192_));
 sg13g2_a21o_1 _10519_ (.A2(_02980_),
    .A1(_00192_),
    .B1(_01604_),
    .X(_02982_));
 sg13g2_a22oi_1 _10520_ (.Y(_02983_),
    .B1(net421),
    .B2(_02982_),
    .A2(_01622_),
    .A1(net637));
 sg13g2_inv_1 _10521_ (.Y(_02984_),
    .A(_02983_));
 sg13g2_o21ai_1 _10522_ (.B1(net315),
    .Y(_02985_),
    .A1(\i_tinyqv.cpu.data_ready_latch ),
    .A2(_02983_));
 sg13g2_o21ai_1 _10523_ (.B1(_02985_),
    .Y(_02986_),
    .A1(_00205_),
    .A2(net315));
 sg13g2_nand2_2 _10524_ (.Y(_02987_),
    .A(_02514_),
    .B(_02986_));
 sg13g2_nand2_1 _10525_ (.Y(_02988_),
    .A(\i_tinyqv.cpu.instr_len[2] ),
    .B(\i_tinyqv.cpu.pc[2] ));
 sg13g2_nor2_1 _10526_ (.A(\i_tinyqv.cpu.instr_len[2] ),
    .B(\i_tinyqv.cpu.pc[2] ),
    .Y(_02989_));
 sg13g2_xor2_1 _10527_ (.B(\i_tinyqv.cpu.pc[2] ),
    .A(\i_tinyqv.cpu.instr_len[2] ),
    .X(_02990_));
 sg13g2_nand2_1 _10528_ (.Y(_02991_),
    .A(\i_tinyqv.cpu.instr_len[1] ),
    .B(\i_tinyqv.cpu.pc[1] ));
 sg13g2_o21ai_1 _10529_ (.B1(_02988_),
    .Y(_02992_),
    .A1(_02989_),
    .A2(_02991_));
 sg13g2_nand2_1 _10530_ (.Y(_02993_),
    .A(\i_tinyqv.cpu.instr_data_start[3] ),
    .B(_02992_));
 sg13g2_nor2_1 _10531_ (.A(_00203_),
    .B(_02993_),
    .Y(_02994_));
 sg13g2_and3_1 _10532_ (.X(_02995_),
    .A(\i_tinyqv.cpu.instr_data_start[6] ),
    .B(\i_tinyqv.cpu.instr_data_start[5] ),
    .C(_02994_));
 sg13g2_nand3_1 _10533_ (.B(\i_tinyqv.cpu.instr_data_start[7] ),
    .C(_02995_),
    .A(\i_tinyqv.cpu.instr_data_start[8] ),
    .Y(_02996_));
 sg13g2_nor2_1 _10534_ (.A(_01517_),
    .B(_02996_),
    .Y(_02997_));
 sg13g2_nor3_2 _10535_ (.A(_01516_),
    .B(_01517_),
    .C(_02996_),
    .Y(_02998_));
 sg13g2_and3_1 _10536_ (.X(_02999_),
    .A(\i_tinyqv.cpu.instr_data_start[12] ),
    .B(\i_tinyqv.cpu.instr_data_start[11] ),
    .C(_02998_));
 sg13g2_nand3_1 _10537_ (.B(net614),
    .C(_02999_),
    .A(net613),
    .Y(_03000_));
 sg13g2_nor2_1 _10538_ (.A(_01514_),
    .B(_03000_),
    .Y(_03001_));
 sg13g2_nand3_1 _10539_ (.B(net612),
    .C(_03001_),
    .A(net611),
    .Y(_03002_));
 sg13g2_nor2_1 _10540_ (.A(_01513_),
    .B(_03002_),
    .Y(_03003_));
 sg13g2_nor3_1 _10541_ (.A(_01513_),
    .B(_00207_),
    .C(_03002_),
    .Y(_03004_));
 sg13g2_xnor2_1 _10542_ (.Y(_03005_),
    .A(net610),
    .B(_03004_));
 sg13g2_nand2_1 _10543_ (.Y(_03006_),
    .A(net594),
    .B(_03005_));
 sg13g2_nand2_2 _10544_ (.Y(_03007_),
    .A(net584),
    .B(_00124_));
 sg13g2_xnor2_1 _10545_ (.Y(_03008_),
    .A(net612),
    .B(_03001_));
 sg13g2_a21oi_1 _10546_ (.A1(_01582_),
    .A2(_03008_),
    .Y(_03009_),
    .B1(_03007_));
 sg13g2_a21oi_1 _10547_ (.A1(\i_tinyqv.cpu.instr_data_start[11] ),
    .A2(_02998_),
    .Y(_03010_),
    .B1(\i_tinyqv.cpu.instr_data_start[12] ));
 sg13g2_nor2_1 _10548_ (.A(_02999_),
    .B(_03010_),
    .Y(_03011_));
 sg13g2_a21o_1 _10549_ (.A2(_02995_),
    .A1(\i_tinyqv.cpu.instr_data_start[7] ),
    .B1(\i_tinyqv.cpu.instr_data_start[8] ),
    .X(_03012_));
 sg13g2_and2_1 _10550_ (.A(_02996_),
    .B(_03012_),
    .X(_03013_));
 sg13g2_a22oi_1 _10551_ (.Y(_03014_),
    .B1(_03013_),
    .B2(net465),
    .A2(_03011_),
    .A1(net458));
 sg13g2_nor2_1 _10552_ (.A(net585),
    .B(_03014_),
    .Y(_03015_));
 sg13g2_xor2_1 _10553_ (.B(_02993_),
    .A(_00203_),
    .X(_03016_));
 sg13g2_a221oi_1 _10554_ (.B2(net353),
    .C1(_03015_),
    .B1(_03016_),
    .A1(_03006_),
    .Y(_03017_),
    .A2(_03009_));
 sg13g2_nor2_2 _10555_ (.A(_02505_),
    .B(_02525_),
    .Y(_03018_));
 sg13g2_nand2b_2 _10556_ (.Y(_03019_),
    .B(_02524_),
    .A_N(_02505_));
 sg13g2_nor3_2 _10557_ (.A(\i_tinyqv.cpu.is_jal ),
    .B(\i_tinyqv.cpu.is_jalr ),
    .C(_03019_),
    .Y(_03020_));
 sg13g2_nor2_1 _10558_ (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .Y(_03021_));
 sg13g2_nor3_1 _10559_ (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .Y(_03022_));
 sg13g2_nand2_1 _10560_ (.Y(_03023_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ));
 sg13g2_inv_1 _10561_ (.Y(_03024_),
    .A(_03023_));
 sg13g2_nor3_1 _10562_ (.A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .C(_03023_),
    .Y(_03025_));
 sg13g2_nand3_1 _10563_ (.B(_03022_),
    .C(_03025_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .Y(_03026_));
 sg13g2_nor2_1 _10564_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(net582),
    .Y(_03027_));
 sg13g2_nand3b_1 _10565_ (.B(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .C(_03027_),
    .Y(_03028_),
    .A_N(\i_tinyqv.cpu.i_core.imm_lo[1] ));
 sg13g2_nor3_2 _10566_ (.A(net456),
    .B(_03026_),
    .C(_03028_),
    .Y(_03029_));
 sg13g2_and2_1 _10567_ (.A(_01588_),
    .B(_03022_),
    .X(_03030_));
 sg13g2_nor2_2 _10568_ (.A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .Y(_03031_));
 sg13g2_nand4_1 _10569_ (.B(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .C(_03030_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .Y(_03032_),
    .D(_03031_));
 sg13g2_nor2_2 _10570_ (.A(_03028_),
    .B(_03032_),
    .Y(_03033_));
 sg13g2_nor3_1 _10571_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .Y(_03034_));
 sg13g2_nor2b_1 _10572_ (.A(net582),
    .B_N(_03034_),
    .Y(_03035_));
 sg13g2_nor2b_2 _10573_ (.A(_03032_),
    .B_N(_03035_),
    .Y(_03036_));
 sg13g2_a22oi_1 _10574_ (.Y(_03037_),
    .B1(_03036_),
    .B2(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .A2(_03033_),
    .A1(\i_tinyqv.cpu.i_core.cycle_count[3] ));
 sg13g2_nand3b_1 _10575_ (.B(_03027_),
    .C(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .Y(_03038_),
    .A_N(\i_tinyqv.cpu.i_core.imm_lo[0] ));
 sg13g2_nor2_2 _10576_ (.A(_03032_),
    .B(_03038_),
    .Y(_03039_));
 sg13g2_nor2_2 _10577_ (.A(_03026_),
    .B(_03038_),
    .Y(_03040_));
 sg13g2_nor2_2 _10578_ (.A(_00120_),
    .B(_02169_),
    .Y(_03041_));
 sg13g2_nand2b_2 _10579_ (.Y(_03042_),
    .B(net461),
    .A_N(_00120_));
 sg13g2_and2_1 _10580_ (.A(_03025_),
    .B(_03030_),
    .X(_03043_));
 sg13g2_nand2_1 _10581_ (.Y(_03044_),
    .A(net582),
    .B(_03034_));
 sg13g2_and3_2 _10582_ (.X(_03045_),
    .A(net582),
    .B(_03034_),
    .C(_03043_));
 sg13g2_nor2_2 _10583_ (.A(_03026_),
    .B(_03044_),
    .Y(_03046_));
 sg13g2_inv_1 _10584_ (.Y(_03047_),
    .A(_03046_));
 sg13g2_a22oi_1 _10585_ (.Y(_03048_),
    .B1(_03046_),
    .B2(\i_tinyqv.cpu.i_core.mip[0] ),
    .A2(_03045_),
    .A1(\i_tinyqv.cpu.i_core.mie[0] ));
 sg13g2_nand2b_1 _10586_ (.Y(_03049_),
    .B(_03041_),
    .A_N(_03048_));
 sg13g2_nand2b_1 _10587_ (.Y(_03050_),
    .B(_03043_),
    .A_N(_03028_));
 sg13g2_inv_1 _10588_ (.Y(_03051_),
    .A(_03050_));
 sg13g2_a22oi_1 _10589_ (.Y(_03052_),
    .B1(net316),
    .B2(\i_tinyqv.cpu.i_core.mcause[0] ),
    .A2(net353),
    .A1(\i_tinyqv.cpu.i_core.mcause[4] ));
 sg13g2_inv_1 _10590_ (.Y(_03053_),
    .A(_03052_));
 sg13g2_a22oi_1 _10591_ (.Y(_03054_),
    .B1(_03040_),
    .B2(_03053_),
    .A2(_03029_),
    .A1(\i_tinyqv.cpu.i_core.mepc[0] ));
 sg13g2_a22oi_1 _10592_ (.Y(_03055_),
    .B1(_03051_),
    .B2(net353),
    .A2(_03039_),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.data[0] ));
 sg13g2_nand4_1 _10593_ (.B(_03049_),
    .C(_03054_),
    .A(_03037_),
    .Y(_03056_),
    .D(_03055_));
 sg13g2_a22oi_1 _10594_ (.Y(_03057_),
    .B1(_03020_),
    .B2(_03056_),
    .A2(\i_tinyqv.cpu.is_lui ),
    .A1(net570));
 sg13g2_o21ai_1 _10595_ (.B1(_03057_),
    .Y(_03058_),
    .A1(_02518_),
    .A2(_03017_));
 sg13g2_o21ai_1 _10596_ (.B1(_03058_),
    .Y(_03059_),
    .A1(_02279_),
    .A2(_02519_));
 sg13g2_nor2b_1 _10597_ (.A(net584),
    .B_N(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .Y(_03060_));
 sg13g2_nor3_2 _10598_ (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .B(_02249_),
    .C(_03060_),
    .Y(_03061_));
 sg13g2_or3_2 _10599_ (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .B(_02249_),
    .C(_03060_),
    .X(_03062_));
 sg13g2_a21oi_2 _10600_ (.B1(_02987_),
    .Y(_03063_),
    .A2(_03061_),
    .A1(\i_tinyqv.cpu.i_core.load_top_bit ));
 sg13g2_inv_1 _10601_ (.Y(_03064_),
    .A(_03063_));
 sg13g2_nor3_2 _10602_ (.A(\addr[5] ),
    .B(_02083_),
    .C(net2382),
    .Y(_03065_));
 sg13g2_nor3_2 _10603_ (.A(net632),
    .B(\addr[6] ),
    .C(_02089_),
    .Y(_03066_));
 sg13g2_nor2_2 _10604_ (.A(_01616_),
    .B(_03065_),
    .Y(_03067_));
 sg13g2_and2_2 _10605_ (.A(_02113_),
    .B(_03067_),
    .X(_03068_));
 sg13g2_nand2_2 _10606_ (.Y(_03069_),
    .A(_02113_),
    .B(_03067_));
 sg13g2_and2_1 _10607_ (.A(_02078_),
    .B(_03066_),
    .X(_03070_));
 sg13g2_nand2_2 _10608_ (.Y(_03071_),
    .A(_02078_),
    .B(_03066_));
 sg13g2_and2_1 _10609_ (.A(_01616_),
    .B(_03065_),
    .X(_03072_));
 sg13g2_inv_1 _10610_ (.Y(_03073_),
    .A(_03072_));
 sg13g2_nand2_1 _10611_ (.Y(_03074_),
    .A(\addr[6] ),
    .B(_03072_));
 sg13g2_and2_1 _10612_ (.A(_03066_),
    .B(_03072_),
    .X(_03075_));
 sg13g2_nand2_1 _10613_ (.Y(_03076_),
    .A(_03066_),
    .B(_03072_));
 sg13g2_a22oi_1 _10614_ (.Y(_03077_),
    .B1(net293),
    .B2(uo_out[4]),
    .A2(net294),
    .A1(\i_spi.data[4] ));
 sg13g2_nor3_2 _10615_ (.A(net632),
    .B(_02089_),
    .C(_03074_),
    .Y(_03078_));
 sg13g2_and2_2 _10616_ (.A(\addr[4] ),
    .B(_03065_),
    .X(_03079_));
 sg13g2_and2_1 _10617_ (.A(_03066_),
    .B(_03079_),
    .X(_03080_));
 sg13g2_nand2_1 _10618_ (.Y(_03081_),
    .A(\i_uart_rx.recieved_data[4] ),
    .B(net289));
 sg13g2_and3_2 _10619_ (.X(_03082_),
    .A(net632),
    .B(_02112_),
    .C(_03072_));
 sg13g2_nor2_2 _10620_ (.A(_02091_),
    .B(_03074_),
    .Y(_03083_));
 sg13g2_nor2_2 _10621_ (.A(_02093_),
    .B(_03073_),
    .Y(_03084_));
 sg13g2_a22oi_1 _10622_ (.Y(_03085_),
    .B1(_03084_),
    .B2(net662),
    .A2(net291),
    .A1(\controller1_data[4] ));
 sg13g2_a21o_1 _10623_ (.A2(net287),
    .A1(\controller2_data[4] ),
    .B1(net472),
    .X(_03086_));
 sg13g2_and2_1 _10624_ (.A(_02092_),
    .B(_03067_),
    .X(_03087_));
 sg13g2_a221oi_1 _10625_ (.B2(\i_time.mtime[4] ),
    .C1(_03086_),
    .B1(net221),
    .A1(\i_time.l_mtimecmp.data_out[4] ),
    .Y(_03088_),
    .A2(net298));
 sg13g2_nand4_1 _10626_ (.B(_03081_),
    .C(_03085_),
    .A(_03077_),
    .Y(_03089_),
    .D(_03088_));
 sg13g2_a21o_1 _10627_ (.A2(net307),
    .A1(\gpio_out_sel[4] ),
    .B1(_03089_),
    .X(_03090_));
 sg13g2_nand2_1 _10628_ (.Y(_03091_),
    .A(uo_out[0]),
    .B(net293));
 sg13g2_or3_1 _10629_ (.A(\i_debug_uart_tx.fsm_state[3] ),
    .B(\i_debug_uart_tx.fsm_state[2] ),
    .C(\i_debug_uart_tx.fsm_state[1] ),
    .X(_03092_));
 sg13g2_nor2_2 _10630_ (.A(\i_debug_uart_tx.fsm_state[0] ),
    .B(_03092_),
    .Y(_03093_));
 sg13g2_or2_2 _10631_ (.X(_03094_),
    .B(_03092_),
    .A(\i_debug_uart_tx.fsm_state[0] ));
 sg13g2_nand3_1 _10632_ (.B(_02112_),
    .C(_03094_),
    .A(net632),
    .Y(_03095_));
 sg13g2_nor3_1 _10633_ (.A(\i_uart_tx.fsm_state[3] ),
    .B(\i_uart_tx.fsm_state[2] ),
    .C(\i_uart_tx.fsm_state[1] ),
    .Y(_03096_));
 sg13g2_or3_1 _10634_ (.A(\i_uart_tx.fsm_state[3] ),
    .B(\i_uart_tx.fsm_state[2] ),
    .C(\i_uart_tx.fsm_state[1] ),
    .X(_03097_));
 sg13g2_nor2_2 _10635_ (.A(\i_uart_tx.fsm_state[0] ),
    .B(_03097_),
    .Y(_03098_));
 sg13g2_nand2_2 _10636_ (.Y(_03099_),
    .A(_01568_),
    .B(_03096_));
 sg13g2_a22oi_1 _10637_ (.Y(_03100_),
    .B1(_03084_),
    .B2(net2),
    .A2(net288),
    .A1(\controller2_data[0] ));
 sg13g2_o21ai_1 _10638_ (.B1(_03095_),
    .Y(_03101_),
    .A1(_02093_),
    .A2(_03098_));
 sg13g2_a221oi_1 _10639_ (.B2(_03079_),
    .C1(net592),
    .B1(_03101_),
    .A1(\i_uart_rx.recieved_data[0] ),
    .Y(_03102_),
    .A2(net289));
 sg13g2_nand3_1 _10640_ (.B(_03100_),
    .C(_03102_),
    .A(_03091_),
    .Y(_03103_));
 sg13g2_nor2_2 _10641_ (.A(net299),
    .B(net221),
    .Y(_03104_));
 sg13g2_or2_1 _10642_ (.X(_03105_),
    .B(net222),
    .A(net299));
 sg13g2_a21oi_1 _10643_ (.A1(_01548_),
    .A2(net296),
    .Y(_03106_),
    .B1(_03104_));
 sg13g2_o21ai_1 _10644_ (.B1(_03106_),
    .Y(_03107_),
    .A1(\i_time.l_mtimecmp.data_out[0] ),
    .A2(net296));
 sg13g2_a22oi_1 _10645_ (.Y(_03108_),
    .B1(net292),
    .B2(\controller1_data[0] ),
    .A2(_02094_),
    .A1(net644));
 sg13g2_a22oi_1 _10646_ (.Y(_03109_),
    .B1(net307),
    .B2(\gpio_out_sel[0] ),
    .A2(net294),
    .A1(\i_spi.data[0] ));
 sg13g2_nand3_1 _10647_ (.B(_03108_),
    .C(_03109_),
    .A(_03107_),
    .Y(_03110_));
 sg13g2_o21ai_1 _10648_ (.B1(_03090_),
    .Y(_03111_),
    .A1(_03103_),
    .A2(_03110_));
 sg13g2_or2_1 _10649_ (.X(_03112_),
    .B(_02096_),
    .A(\addr[5] ));
 sg13g2_nor2b_1 _10650_ (.A(net292),
    .B_N(_03112_),
    .Y(_03113_));
 sg13g2_or3_1 _10651_ (.A(net294),
    .B(net293),
    .C(net288),
    .X(_03114_));
 sg13g2_nor4_1 _10652_ (.A(_02094_),
    .B(net290),
    .C(net183),
    .D(_03114_),
    .Y(_03115_));
 sg13g2_and2_2 _10653_ (.A(_03113_),
    .B(_03115_),
    .X(_03116_));
 sg13g2_nand2_1 _10654_ (.Y(_03117_),
    .A(_03113_),
    .B(_03115_));
 sg13g2_a21oi_1 _10655_ (.A1(_03111_),
    .A2(net114),
    .Y(_03118_),
    .B1(net636));
 sg13g2_nor2_1 _10656_ (.A(net592),
    .B(\i_latch_mem.data_out[0] ),
    .Y(_03119_));
 sg13g2_o21ai_1 _10657_ (.B1(net636),
    .Y(_03120_),
    .A1(net472),
    .A2(\i_latch_mem.data_out[4] ));
 sg13g2_o21ai_1 _10658_ (.B1(_02075_),
    .Y(_03121_),
    .A1(_03119_),
    .A2(_03120_));
 sg13g2_nor2_2 _10659_ (.A(_03118_),
    .B(_03121_),
    .Y(_03122_));
 sg13g2_nand2_1 _10660_ (.Y(_03123_),
    .A(_02535_),
    .B(_02981_));
 sg13g2_mux2_1 _10661_ (.A0(\i_tinyqv.cpu.instr_data_in[12] ),
    .A1(\i_tinyqv.cpu.instr_data_in[4] ),
    .S(_03123_),
    .X(_03124_));
 sg13g2_nor2_1 _10662_ (.A(_01661_),
    .B(net117),
    .Y(_03125_));
 sg13g2_a22oi_1 _10663_ (.Y(_03126_),
    .B1(_03125_),
    .B2(_02535_),
    .A2(net108),
    .A1(\i_tinyqv.cpu.instr_data_in[0] ));
 sg13g2_o21ai_1 _10664_ (.B1(net419),
    .Y(_03127_),
    .A1(net591),
    .A2(_03126_));
 sg13g2_a21oi_1 _10665_ (.A1(net595),
    .A2(_03124_),
    .Y(_03128_),
    .B1(_03127_));
 sg13g2_nor4_1 _10666_ (.A(net584),
    .B(net588),
    .C(_03122_),
    .D(_03128_),
    .Y(_03129_));
 sg13g2_nand2_2 _10667_ (.Y(_03130_),
    .A(_02530_),
    .B(_02533_));
 sg13g2_nor2_1 _10668_ (.A(net117),
    .B(_03130_),
    .Y(_03131_));
 sg13g2_or2_1 _10669_ (.X(_03132_),
    .B(_03130_),
    .A(net117));
 sg13g2_nor2_1 _10670_ (.A(\i_time.mtime[8] ),
    .B(net298),
    .Y(_03133_));
 sg13g2_a21oi_1 _10671_ (.A1(_01641_),
    .A2(net298),
    .Y(_03134_),
    .B1(_03133_));
 sg13g2_nand2_1 _10672_ (.Y(_03135_),
    .A(\controller1_data[8] ),
    .B(net291));
 sg13g2_a21oi_1 _10673_ (.A1(_01662_),
    .A2(net105),
    .Y(_03136_),
    .B1(net416));
 sg13g2_o21ai_1 _10674_ (.B1(_03136_),
    .Y(_03137_),
    .A1(\i_tinyqv.mem.qspi_data_buf[12] ),
    .A2(net105));
 sg13g2_a21oi_1 _10675_ (.A1(net634),
    .A2(_01663_),
    .Y(_03138_),
    .B1(net421));
 sg13g2_a21oi_1 _10676_ (.A1(\i_time.mtime[12] ),
    .A2(net222),
    .Y(_03139_),
    .B1(net297));
 sg13g2_a21oi_2 _10677_ (.B1(_03139_),
    .Y(_03140_),
    .A2(net297),
    .A1(_01638_));
 sg13g2_o21ai_1 _10678_ (.B1(_03138_),
    .Y(_03141_),
    .A1(net116),
    .A2(_03140_));
 sg13g2_a21oi_1 _10679_ (.A1(_03137_),
    .A2(_03141_),
    .Y(_03142_),
    .B1(_02171_));
 sg13g2_a21oi_1 _10680_ (.A1(_01661_),
    .A2(net105),
    .Y(_03143_),
    .B1(net415));
 sg13g2_o21ai_1 _10681_ (.B1(_03143_),
    .Y(_03144_),
    .A1(\i_tinyqv.mem.qspi_data_buf[8] ),
    .A2(net105));
 sg13g2_o21ai_1 _10682_ (.B1(net415),
    .Y(_03145_),
    .A1(_01525_),
    .A2(\i_latch_mem.data_out[8] ));
 sg13g2_nand2_1 _10683_ (.Y(_03146_),
    .A(net183),
    .B(_03134_));
 sg13g2_a22oi_1 _10684_ (.Y(_03147_),
    .B1(net288),
    .B2(\controller2_data[8] ),
    .A2(net307),
    .A1(\gpio_out_sel[8] ));
 sg13g2_nand4_1 _10685_ (.B(_03135_),
    .C(_03146_),
    .A(net115),
    .Y(_03148_),
    .D(_03147_));
 sg13g2_nand2b_1 _10686_ (.Y(_03149_),
    .B(_03148_),
    .A_N(_03145_));
 sg13g2_a21oi_1 _10687_ (.A1(_03144_),
    .A2(_03149_),
    .Y(_03150_),
    .B1(net464));
 sg13g2_o21ai_1 _10688_ (.B1(net476),
    .Y(_03151_),
    .A1(_03142_),
    .A2(_03150_));
 sg13g2_a21oi_1 _10689_ (.A1(\i_tinyqv.mem.qspi_data_buf[24] ),
    .A2(net117),
    .Y(_03152_),
    .B1(_03125_));
 sg13g2_o21ai_1 _10690_ (.B1(net591),
    .Y(_03153_),
    .A1(\i_tinyqv.mem.qspi_data_buf[28] ),
    .A2(_02981_));
 sg13g2_a21oi_1 _10691_ (.A1(_01662_),
    .A2(_02981_),
    .Y(_03154_),
    .B1(_03153_));
 sg13g2_o21ai_1 _10692_ (.B1(net418),
    .Y(_03155_),
    .A1(net591),
    .A2(_03152_));
 sg13g2_mux4_1 _10693_ (.S0(net473),
    .A0(\i_time.mtime[28] ),
    .A1(\i_time.mtime[24] ),
    .A2(\i_time.l_mtimecmp.data_out[28] ),
    .A3(\i_time.l_mtimecmp.data_out[24] ),
    .S1(_03068_),
    .X(_03156_));
 sg13g2_a21oi_1 _10694_ (.A1(net590),
    .A2(\i_latch_mem.data_out[28] ),
    .Y(_03157_),
    .B1(net427));
 sg13g2_o21ai_1 _10695_ (.B1(_03157_),
    .Y(_03158_),
    .A1(net590),
    .A2(_01666_));
 sg13g2_a21oi_1 _10696_ (.A1(net183),
    .A2(_03156_),
    .Y(_03159_),
    .B1(net116));
 sg13g2_o21ai_1 _10697_ (.B1(_03158_),
    .Y(_03160_),
    .A1(_03154_),
    .A2(_03155_));
 sg13g2_nor3_1 _10698_ (.A(_01581_),
    .B(_03159_),
    .C(_03160_),
    .Y(_03161_));
 sg13g2_o21ai_1 _10699_ (.B1(net471),
    .Y(_03162_),
    .A1(net427),
    .A2(\i_latch_mem.data_out[20] ));
 sg13g2_a21oi_1 _10700_ (.A1(_01665_),
    .A2(net418),
    .Y(_03163_),
    .B1(_03162_));
 sg13g2_o21ai_1 _10701_ (.B1(net463),
    .Y(_03164_),
    .A1(net427),
    .A2(\i_latch_mem.data_out[16] ));
 sg13g2_a21oi_1 _10702_ (.A1(_01664_),
    .A2(net418),
    .Y(_03165_),
    .B1(_03164_));
 sg13g2_nor2_1 _10703_ (.A(\i_time.l_mtimecmp.data_out[16] ),
    .B(net295),
    .Y(_03166_));
 sg13g2_nor2_1 _10704_ (.A(\i_time.l_mtimecmp.data_out[20] ),
    .B(net296),
    .Y(_03167_));
 sg13g2_a21oi_1 _10705_ (.A1(\i_time.mtime[20] ),
    .A2(net222),
    .Y(_03168_),
    .B1(net300));
 sg13g2_o21ai_1 _10706_ (.B1(net114),
    .Y(_03169_),
    .A1(_03167_),
    .A2(_03168_));
 sg13g2_a21oi_1 _10707_ (.A1(\i_time.mtime[16] ),
    .A2(net220),
    .Y(_03170_),
    .B1(net297));
 sg13g2_o21ai_1 _10708_ (.B1(net114),
    .Y(_03171_),
    .A1(_03166_),
    .A2(_03170_));
 sg13g2_a221oi_1 _10709_ (.B2(_03165_),
    .C1(_03161_),
    .B1(_03171_),
    .A1(_03163_),
    .Y(_03172_),
    .A2(_03169_));
 sg13g2_o21ai_1 _10710_ (.B1(_03151_),
    .Y(_03173_),
    .A1(net476),
    .A2(_03172_));
 sg13g2_o21ai_1 _10711_ (.B1(_03062_),
    .Y(_03174_),
    .A1(_03129_),
    .A2(_03173_));
 sg13g2_a221oi_1 _10712_ (.B2(_03174_),
    .C1(_02826_),
    .B1(_03063_),
    .A1(_02987_),
    .Y(_03175_),
    .A2(_03059_));
 sg13g2_a21o_2 _10713_ (.A2(_02979_),
    .A1(_02826_),
    .B1(_03175_),
    .X(\debug_rd[0] ));
 sg13g2_nor3_1 _10714_ (.A(_02511_),
    .B(_02520_),
    .C(_03018_),
    .Y(_03176_));
 sg13g2_a21oi_1 _10715_ (.A1(_02157_),
    .A2(_02510_),
    .Y(_03177_),
    .B1(_01596_));
 sg13g2_a22oi_1 _10716_ (.Y(_03178_),
    .B1(_03177_),
    .B2(_02830_),
    .A2(_03176_),
    .A1(_02987_));
 sg13g2_and2_2 _10717_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .X(_03179_));
 sg13g2_nand2_1 _10718_ (.Y(_03180_),
    .A(net661),
    .B(_03179_));
 sg13g2_nand4_1 _10719_ (.B(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .C(_03178_),
    .A(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .Y(_03181_),
    .D(_03179_));
 sg13g2_nor2_1 _10720_ (.A(net83),
    .B(_03181_),
    .Y(_03182_));
 sg13g2_a21oi_1 _10721_ (.A1(_01591_),
    .A2(_03181_),
    .Y(_00086_),
    .B1(_03182_));
 sg13g2_mux2_2 _10722_ (.A0(\i_uart_rx.uart_rts ),
    .A1(\gpio_out[1] ),
    .S(\gpio_out_sel[1] ),
    .X(uo_out[1]));
 sg13g2_nand2_1 _10723_ (.Y(_03183_),
    .A(debug_register_data),
    .B(\debug_rd_r[3] ));
 sg13g2_o21ai_1 _10724_ (.B1(_03183_),
    .Y(_03184_),
    .A1(_01554_),
    .A2(debug_register_data));
 sg13g2_mux2_2 _10725_ (.A0(_03184_),
    .A1(\gpio_out[5] ),
    .S(\gpio_out_sel[5] ),
    .X(uo_out[5]));
 sg13g2_nor2_1 _10726_ (.A(_02161_),
    .B(_02974_),
    .Y(_03185_));
 sg13g2_nand2_1 _10727_ (.Y(_03186_),
    .A(net622),
    .B(_02876_));
 sg13g2_a21oi_1 _10728_ (.A1(net502),
    .A2(_02862_),
    .Y(_03187_),
    .B1(net351));
 sg13g2_nand2_1 _10729_ (.Y(_03188_),
    .A(net622),
    .B(_02899_));
 sg13g2_a21oi_1 _10730_ (.A1(net502),
    .A2(_02874_),
    .Y(_03189_),
    .B1(net349));
 sg13g2_a221oi_1 _10731_ (.B2(_03189_),
    .C1(_02880_),
    .B1(_03188_),
    .A1(_03186_),
    .Y(_03190_),
    .A2(_03187_));
 sg13g2_nand2_1 _10732_ (.Y(_03191_),
    .A(net621),
    .B(_02903_));
 sg13g2_a21oi_1 _10733_ (.A1(net501),
    .A2(_02905_),
    .Y(_03192_),
    .B1(net351));
 sg13g2_nand2_1 _10734_ (.Y(_03193_),
    .A(net504),
    .B(_02904_));
 sg13g2_a21oi_1 _10735_ (.A1(net622),
    .A2(_02919_),
    .Y(_03194_),
    .B1(_02865_));
 sg13g2_a221oi_1 _10736_ (.B2(_03194_),
    .C1(_02881_),
    .B1(_03193_),
    .A1(_03191_),
    .Y(_03195_),
    .A2(_03192_));
 sg13g2_nor3_1 _10737_ (.A(_02872_),
    .B(_03190_),
    .C(_03195_),
    .Y(_03196_));
 sg13g2_nand2_1 _10738_ (.Y(_03197_),
    .A(net621),
    .B(_02884_));
 sg13g2_a21oi_1 _10739_ (.A1(net501),
    .A2(_02897_),
    .Y(_03198_),
    .B1(net351));
 sg13g2_nand2_1 _10740_ (.Y(_03199_),
    .A(net501),
    .B(_02891_));
 sg13g2_a22oi_1 _10741_ (.Y(_03200_),
    .B1(_03199_),
    .B2(_02955_),
    .A2(_03198_),
    .A1(_03197_));
 sg13g2_a21oi_1 _10742_ (.A1(net624),
    .A2(_02870_),
    .Y(_03201_),
    .B1(net350));
 sg13g2_o21ai_1 _10743_ (.B1(_03201_),
    .Y(_03202_),
    .A1(net624),
    .A2(_02911_));
 sg13g2_nand2_1 _10744_ (.Y(_03203_),
    .A(net622),
    .B(_02916_));
 sg13g2_a21oi_1 _10745_ (.A1(net502),
    .A2(_02920_),
    .Y(_03204_),
    .B1(net351));
 sg13g2_a21oi_1 _10746_ (.A1(_03203_),
    .A2(_03204_),
    .Y(_03205_),
    .B1(_02881_));
 sg13g2_a221oi_1 _10747_ (.B2(_03205_),
    .C1(_02873_),
    .B1(_03202_),
    .A1(_02881_),
    .Y(_03206_),
    .A2(_03200_));
 sg13g2_nor3_1 _10748_ (.A(_02856_),
    .B(_03196_),
    .C(_03206_),
    .Y(_03207_));
 sg13g2_or2_1 _10749_ (.X(_03208_),
    .B(_03207_),
    .A(_02857_));
 sg13g2_nand2_1 _10750_ (.Y(_03209_),
    .A(net623),
    .B(_02927_));
 sg13g2_a21oi_1 _10751_ (.A1(net503),
    .A2(_02963_),
    .Y(_03210_),
    .B1(net352));
 sg13g2_nand2_1 _10752_ (.Y(_03211_),
    .A(net503),
    .B(_02929_));
 sg13g2_a21oi_1 _10753_ (.A1(net623),
    .A2(_02931_),
    .Y(_03212_),
    .B1(net349));
 sg13g2_a221oi_1 _10754_ (.B2(_03212_),
    .C1(_02872_),
    .B1(_03211_),
    .A1(_03209_),
    .Y(_03213_),
    .A2(_03210_));
 sg13g2_and2_1 _10755_ (.A(net501),
    .B(_02933_),
    .X(_03214_));
 sg13g2_a21oi_1 _10756_ (.A1(net621),
    .A2(_02947_),
    .Y(_03215_),
    .B1(_03214_));
 sg13g2_nand2_1 _10757_ (.Y(_03216_),
    .A(net501),
    .B(_02949_));
 sg13g2_o21ai_1 _10758_ (.B1(_03216_),
    .Y(_03217_),
    .A1(net501),
    .A2(_02953_));
 sg13g2_o21ai_1 _10759_ (.B1(_02872_),
    .Y(_03218_),
    .A1(net350),
    .A2(_03217_));
 sg13g2_a21oi_1 _10760_ (.A1(net350),
    .A2(_03215_),
    .Y(_03219_),
    .B1(_03218_));
 sg13g2_nor3_1 _10761_ (.A(_02880_),
    .B(_03213_),
    .C(_03219_),
    .Y(_03220_));
 sg13g2_mux4_1 _10762_ (.S0(net573),
    .A0(_00236_),
    .A1(_00237_),
    .A2(_00234_),
    .A3(_00235_),
    .S1(net626),
    .X(_03221_));
 sg13g2_mux4_1 _10763_ (.S0(net351),
    .A0(_02936_),
    .A1(_02941_),
    .A2(_03221_),
    .A3(_02937_),
    .S1(net504),
    .X(_03222_));
 sg13g2_nand2_1 _10764_ (.Y(_03223_),
    .A(net622),
    .B(_02966_));
 sg13g2_a21oi_1 _10765_ (.A1(net503),
    .A2(_02958_),
    .Y(_03224_),
    .B1(net349));
 sg13g2_nand2_1 _10766_ (.Y(_03225_),
    .A(_03223_),
    .B(_03224_));
 sg13g2_and2_1 _10767_ (.A(net503),
    .B(_02940_),
    .X(_03226_));
 sg13g2_a21oi_1 _10768_ (.A1(net623),
    .A2(_02960_),
    .Y(_03227_),
    .B1(_03226_));
 sg13g2_a21oi_1 _10769_ (.A1(net349),
    .A2(_03227_),
    .Y(_03228_),
    .B1(_02873_));
 sg13g2_a221oi_1 _10770_ (.B2(_03228_),
    .C1(_02881_),
    .B1(_03225_),
    .A1(_02873_),
    .Y(_03229_),
    .A2(_03222_));
 sg13g2_nor3_1 _10771_ (.A(_02856_),
    .B(_03220_),
    .C(_03229_),
    .Y(_03230_));
 sg13g2_or2_1 _10772_ (.X(_03231_),
    .B(_03230_),
    .A(_02857_));
 sg13g2_mux2_1 _10773_ (.A0(_03208_),
    .A1(_03231_),
    .S(net572),
    .X(_03232_));
 sg13g2_nor2_1 _10774_ (.A(_02842_),
    .B(_03232_),
    .Y(_03233_));
 sg13g2_xnor2_1 _10775_ (.Y(_03234_),
    .A(_02293_),
    .B(_02294_));
 sg13g2_o21ai_1 _10776_ (.B1(net581),
    .Y(_03235_),
    .A1(_02178_),
    .A2(_02223_));
 sg13g2_nand3_1 _10777_ (.B(_02837_),
    .C(_03235_),
    .A(_02496_),
    .Y(_03236_));
 sg13g2_o21ai_1 _10778_ (.B1(_03236_),
    .Y(_03237_),
    .A1(_02833_),
    .A2(_03234_));
 sg13g2_a21oi_1 _10779_ (.A1(_02498_),
    .A2(_02836_),
    .Y(_03238_),
    .B1(_03237_));
 sg13g2_xnor2_1 _10780_ (.Y(_03239_),
    .A(_02559_),
    .B(_02560_));
 sg13g2_o21ai_1 _10781_ (.B1(_02842_),
    .Y(_03240_),
    .A1(net406),
    .A2(_03239_));
 sg13g2_a21oi_1 _10782_ (.A1(net406),
    .A2(_03238_),
    .Y(_03241_),
    .B1(_03240_));
 sg13g2_o21ai_1 _10783_ (.B1(_03185_),
    .Y(_03242_),
    .A1(_03233_),
    .A2(_03241_));
 sg13g2_o21ai_1 _10784_ (.B1(_03242_),
    .Y(_03243_),
    .A1(_00237_),
    .A2(_02829_));
 sg13g2_and3_1 _10785_ (.X(_03244_),
    .A(net610),
    .B(\i_tinyqv.cpu.instr_data_start[19] ),
    .C(_03003_));
 sg13g2_xnor2_1 _10786_ (.Y(_03245_),
    .A(net609),
    .B(_03244_));
 sg13g2_nand2_1 _10787_ (.Y(_03246_),
    .A(net593),
    .B(_03245_));
 sg13g2_a21o_1 _10788_ (.A2(_03001_),
    .A1(net612),
    .B1(net611),
    .X(_03247_));
 sg13g2_nand2_1 _10789_ (.Y(_03248_),
    .A(_03002_),
    .B(_03247_));
 sg13g2_a21oi_1 _10790_ (.A1(_01582_),
    .A2(_03248_),
    .Y(_03249_),
    .B1(_03007_));
 sg13g2_xnor2_1 _10791_ (.Y(_03250_),
    .A(net614),
    .B(_02999_));
 sg13g2_xnor2_1 _10792_ (.Y(_03251_),
    .A(\i_tinyqv.cpu.instr_data_start[5] ),
    .B(_02994_));
 sg13g2_xor2_1 _10793_ (.B(\i_tinyqv.cpu.pc[1] ),
    .A(\i_tinyqv.cpu.instr_len[1] ),
    .X(_03252_));
 sg13g2_o21ai_1 _10794_ (.B1(net474),
    .Y(_03253_),
    .A1(_02169_),
    .A2(_03252_));
 sg13g2_a21oi_1 _10795_ (.A1(net468),
    .A2(_03251_),
    .Y(_03254_),
    .B1(_03253_));
 sg13g2_xnor2_1 _10796_ (.Y(_03255_),
    .A(\i_tinyqv.cpu.instr_data_start[9] ),
    .B(_02996_));
 sg13g2_o21ai_1 _10797_ (.B1(_03254_),
    .Y(_03256_),
    .A1(net464),
    .A2(_03255_));
 sg13g2_a21oi_1 _10798_ (.A1(net458),
    .A2(_03250_),
    .Y(_03257_),
    .B1(_03256_));
 sg13g2_a21oi_2 _10799_ (.B1(_03257_),
    .Y(_03258_),
    .A2(_03249_),
    .A1(_03246_));
 sg13g2_mux2_1 _10800_ (.A0(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .A1(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .S(net313),
    .X(_03259_));
 sg13g2_a22oi_1 _10801_ (.Y(_03260_),
    .B1(_03039_),
    .B2(\i_tinyqv.cpu.i_core.i_instrret.data[1] ),
    .A2(_03036_),
    .A1(\i_tinyqv.cpu.i_core.cycle_count[1] ));
 sg13g2_a22oi_1 _10802_ (.Y(_03261_),
    .B1(_03046_),
    .B2(\i_tinyqv.cpu.i_core.mip[1] ),
    .A2(_03045_),
    .A1(\i_tinyqv.cpu.i_core.mie[1] ));
 sg13g2_nand4_1 _10803_ (.B(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .A(_01588_),
    .Y(_03262_),
    .D(\i_tinyqv.cpu.i_core.imm_lo[4] ));
 sg13g2_nand3_1 _10804_ (.B(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .C(_03024_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .Y(_03263_));
 sg13g2_nor4_1 _10805_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(net582),
    .C(_03262_),
    .D(_03263_),
    .Y(_03264_));
 sg13g2_a22oi_1 _10806_ (.Y(_03265_),
    .B1(_03264_),
    .B2(_03021_),
    .A2(_03040_),
    .A1(\i_tinyqv.cpu.i_core.mcause[1] ));
 sg13g2_o21ai_1 _10807_ (.B1(_03260_),
    .Y(_03266_),
    .A1(net334),
    .A2(_03265_));
 sg13g2_a221oi_1 _10808_ (.B2(_03259_),
    .C1(_03266_),
    .B1(_03033_),
    .A1(\i_tinyqv.cpu.i_core.mepc[1] ),
    .Y(_03267_),
    .A2(_03029_));
 sg13g2_o21ai_1 _10809_ (.B1(_03267_),
    .Y(_03268_),
    .A1(_03042_),
    .A2(_03261_));
 sg13g2_a22oi_1 _10810_ (.Y(_03269_),
    .B1(_03020_),
    .B2(_03268_),
    .A2(\i_tinyqv.cpu.is_lui ),
    .A1(net570));
 sg13g2_o21ai_1 _10811_ (.B1(_03269_),
    .Y(_03270_),
    .A1(_02518_),
    .A2(_03258_));
 sg13g2_o21ai_1 _10812_ (.B1(_03270_),
    .Y(_03271_),
    .A1(_02221_),
    .A2(_02519_));
 sg13g2_and2_1 _10813_ (.A(net592),
    .B(\i_latch_mem.data_out[5] ),
    .X(_03272_));
 sg13g2_a21oi_1 _10814_ (.A1(net472),
    .A2(\i_latch_mem.data_out[1] ),
    .Y(_03273_),
    .B1(_03272_));
 sg13g2_nand2_1 _10815_ (.Y(_03274_),
    .A(\controller1_data[5] ),
    .B(net291));
 sg13g2_nand2_1 _10816_ (.Y(_03275_),
    .A(\i_spi.data[5] ),
    .B(net294));
 sg13g2_a22oi_1 _10817_ (.Y(_03276_),
    .B1(uo_out[5]),
    .B2(net293),
    .A2(net287),
    .A1(\controller2_data[5] ));
 sg13g2_a22oi_1 _10818_ (.Y(_03277_),
    .B1(net307),
    .B2(\gpio_out_sel[5] ),
    .A2(net289),
    .A1(\i_uart_rx.recieved_data[5] ));
 sg13g2_a21oi_1 _10819_ (.A1(net7),
    .A2(_03084_),
    .Y(_03278_),
    .B1(net472));
 sg13g2_a22oi_1 _10820_ (.Y(_03279_),
    .B1(net221),
    .B2(\i_time.mtime[5] ),
    .A2(net298),
    .A1(\i_time.l_mtimecmp.data_out[5] ));
 sg13g2_nand4_1 _10821_ (.B(_03277_),
    .C(_03278_),
    .A(_03275_),
    .Y(_03280_),
    .D(_03279_));
 sg13g2_nand3b_1 _10822_ (.B(_03274_),
    .C(_03276_),
    .Y(_03281_),
    .A_N(_03280_));
 sg13g2_nand2_1 _10823_ (.Y(_03282_),
    .A(\controller2_data[1] ),
    .B(net287));
 sg13g2_nand2_1 _10824_ (.Y(_03283_),
    .A(\i_spi.data[1] ),
    .B(net294));
 sg13g2_nor2b_1 _10825_ (.A(\i_uart_rx.fsm_state[2] ),
    .B_N(\i_uart_rx.fsm_state[3] ),
    .Y(_03284_));
 sg13g2_and2_1 _10826_ (.A(\i_uart_rx.fsm_state[1] ),
    .B(_03284_),
    .X(_03285_));
 sg13g2_nand2_1 _10827_ (.Y(_03286_),
    .A(\i_uart_rx.fsm_state[1] ),
    .B(_03284_));
 sg13g2_and2_2 _10828_ (.A(\i_uart_rx.fsm_state[0] ),
    .B(_03285_),
    .X(_03287_));
 sg13g2_inv_1 _10829_ (.Y(_03288_),
    .A(_03287_));
 sg13g2_nand2_1 _10830_ (.Y(_03289_),
    .A(net3),
    .B(_03084_));
 sg13g2_a22oi_1 _10831_ (.Y(_03290_),
    .B1(uo_out[1]),
    .B2(net293),
    .A2(net221),
    .A1(\i_time.mtime[1] ));
 sg13g2_nand3_1 _10832_ (.B(_03289_),
    .C(_03290_),
    .A(_03282_),
    .Y(_03291_));
 sg13g2_a22oi_1 _10833_ (.Y(_03292_),
    .B1(_03082_),
    .B2(\gpio_out_sel[1] ),
    .A2(net292),
    .A1(\controller1_data[1] ));
 sg13g2_a21oi_1 _10834_ (.A1(\i_time.l_mtimecmp.data_out[1] ),
    .A2(net299),
    .Y(_03293_),
    .B1(net592));
 sg13g2_and2_1 _10835_ (.A(_03079_),
    .B(_03287_),
    .X(_03294_));
 sg13g2_a22oi_1 _10836_ (.Y(_03295_),
    .B1(_03294_),
    .B2(_02092_),
    .A2(net289),
    .A1(\i_uart_rx.recieved_data[1] ));
 sg13g2_nand4_1 _10837_ (.B(_03292_),
    .C(_03293_),
    .A(_03283_),
    .Y(_03296_),
    .D(_03295_));
 sg13g2_o21ai_1 _10838_ (.B1(_03281_),
    .Y(_03297_),
    .A1(_03291_),
    .A2(_03296_));
 sg13g2_a221oi_1 _10839_ (.B2(net115),
    .C1(net588),
    .B1(_03297_),
    .A1(net635),
    .Y(_03298_),
    .A2(_03273_));
 sg13g2_o21ai_1 _10840_ (.B1(net460),
    .Y(_03299_),
    .A1(_01525_),
    .A2(\i_latch_mem.data_out[13] ));
 sg13g2_a21oi_1 _10841_ (.A1(_01538_),
    .A2(net295),
    .Y(_03300_),
    .B1(_03104_));
 sg13g2_o21ai_1 _10842_ (.B1(_03300_),
    .Y(_03301_),
    .A1(\i_time.l_mtimecmp.data_out[13] ),
    .A2(net295));
 sg13g2_a21oi_1 _10843_ (.A1(net115),
    .A2(_03301_),
    .Y(_03302_),
    .B1(_03299_));
 sg13g2_o21ai_1 _10844_ (.B1(net467),
    .Y(_03303_),
    .A1(net427),
    .A2(\i_latch_mem.data_out[9] ));
 sg13g2_nor2_1 _10845_ (.A(\i_time.l_mtimecmp.data_out[9] ),
    .B(net296),
    .Y(_03304_));
 sg13g2_a21oi_1 _10846_ (.A1(_01541_),
    .A2(net296),
    .Y(_03305_),
    .B1(_03304_));
 sg13g2_a22oi_1 _10847_ (.Y(_03306_),
    .B1(net287),
    .B2(\controller2_data[9] ),
    .A2(net291),
    .A1(\controller1_data[9] ));
 sg13g2_inv_1 _10848_ (.Y(_03307_),
    .A(_03306_));
 sg13g2_a221oi_1 _10849_ (.B2(_03305_),
    .C1(_03307_),
    .B1(_03105_),
    .A1(\gpio_out_sel[9] ),
    .Y(_03308_),
    .A2(net307));
 sg13g2_a21oi_1 _10850_ (.A1(net115),
    .A2(_03308_),
    .Y(_03309_),
    .B1(_03303_));
 sg13g2_nor3_2 _10851_ (.A(_03298_),
    .B(_03302_),
    .C(_03309_),
    .Y(_03310_));
 sg13g2_nor2_1 _10852_ (.A(\i_tinyqv.cpu.instr_data_in[13] ),
    .B(net117),
    .Y(_03311_));
 sg13g2_a22oi_1 _10853_ (.Y(_03312_),
    .B1(_03311_),
    .B2(_02535_),
    .A2(net108),
    .A1(_01671_));
 sg13g2_a21oi_1 _10854_ (.A1(_01672_),
    .A2(net105),
    .Y(_03313_),
    .B1(_02171_));
 sg13g2_o21ai_1 _10855_ (.B1(_03313_),
    .Y(_03314_),
    .A1(\i_tinyqv.mem.qspi_data_buf[13] ),
    .A2(net106));
 sg13g2_nor2_1 _10856_ (.A(\i_tinyqv.cpu.instr_data_in[9] ),
    .B(net108),
    .Y(_03315_));
 sg13g2_a21oi_1 _10857_ (.A1(_01669_),
    .A2(net108),
    .Y(_03316_),
    .B1(_03315_));
 sg13g2_a21oi_1 _10858_ (.A1(_01670_),
    .A2(net105),
    .Y(_03317_),
    .B1(net464));
 sg13g2_o21ai_1 _10859_ (.B1(_03317_),
    .Y(_03318_),
    .A1(\i_tinyqv.mem.qspi_data_buf[9] ),
    .A2(net105));
 sg13g2_a21oi_1 _10860_ (.A1(net471),
    .A2(_03312_),
    .Y(_03319_),
    .B1(net416));
 sg13g2_nand2_1 _10861_ (.Y(_03320_),
    .A(_03318_),
    .B(_03319_));
 sg13g2_a21oi_1 _10862_ (.A1(net463),
    .A2(_03316_),
    .Y(_03321_),
    .B1(_03320_));
 sg13g2_a21oi_1 _10863_ (.A1(_03314_),
    .A2(_03321_),
    .Y(_03322_),
    .B1(_03310_));
 sg13g2_o21ai_1 _10864_ (.B1(net591),
    .Y(_03323_),
    .A1(\i_tinyqv.mem.qspi_data_buf[29] ),
    .A2(_02981_));
 sg13g2_o21ai_1 _10865_ (.B1(net419),
    .Y(_03324_),
    .A1(_03311_),
    .A2(_03323_));
 sg13g2_o21ai_1 _10866_ (.B1(net467),
    .Y(_03325_),
    .A1(\i_tinyqv.mem.qspi_data_buf[25] ),
    .A2(_02981_));
 sg13g2_a21oi_1 _10867_ (.A1(_01670_),
    .A2(_02981_),
    .Y(_03326_),
    .B1(_03325_));
 sg13g2_a21oi_1 _10868_ (.A1(net588),
    .A2(_03324_),
    .Y(_03327_),
    .B1(_03326_));
 sg13g2_nor2b_1 _10869_ (.A(net590),
    .B_N(\i_latch_mem.data_out[25] ),
    .Y(_03328_));
 sg13g2_a21oi_1 _10870_ (.A1(net590),
    .A2(\i_latch_mem.data_out[29] ),
    .Y(_03329_),
    .B1(_03328_));
 sg13g2_mux4_1 _10871_ (.S0(net473),
    .A0(\i_time.mtime[29] ),
    .A1(\i_time.mtime[25] ),
    .A2(\i_time.l_mtimecmp.data_out[29] ),
    .A3(\i_time.l_mtimecmp.data_out[25] ),
    .S1(net301),
    .X(_03330_));
 sg13g2_nand2_1 _10872_ (.Y(_03331_),
    .A(net183),
    .B(_03330_));
 sg13g2_a221oi_1 _10873_ (.B2(net115),
    .C1(_03327_),
    .B1(_03331_),
    .A1(net637),
    .Y(_03332_),
    .A2(_03329_));
 sg13g2_nor2_1 _10874_ (.A(\i_time.l_mtimecmp.data_out[21] ),
    .B(net296),
    .Y(_03333_));
 sg13g2_nor2_1 _10875_ (.A(\i_tinyqv.mem.data_from_read[21] ),
    .B(net415),
    .Y(_03334_));
 sg13g2_o21ai_1 _10876_ (.B1(net471),
    .Y(_03335_),
    .A1(net427),
    .A2(\i_latch_mem.data_out[21] ));
 sg13g2_o21ai_1 _10877_ (.B1(net463),
    .Y(_03336_),
    .A1(net427),
    .A2(\i_latch_mem.data_out[17] ));
 sg13g2_a21o_1 _10878_ (.A2(net220),
    .A1(\i_time.mtime[17] ),
    .B1(net297),
    .X(_03337_));
 sg13g2_o21ai_1 _10879_ (.B1(_03337_),
    .Y(_03338_),
    .A1(\i_time.l_mtimecmp.data_out[17] ),
    .A2(net295));
 sg13g2_a221oi_1 _10880_ (.B2(_03338_),
    .C1(_03336_),
    .B1(net115),
    .A1(_01674_),
    .Y(_03339_),
    .A2(net418));
 sg13g2_a21oi_1 _10881_ (.A1(_01533_),
    .A2(net296),
    .Y(_03340_),
    .B1(_03333_));
 sg13g2_a21oi_1 _10882_ (.A1(net183),
    .A2(_03340_),
    .Y(_03341_),
    .B1(net116));
 sg13g2_nor3_1 _10883_ (.A(_03334_),
    .B(_03335_),
    .C(_03341_),
    .Y(_03342_));
 sg13g2_nor4_2 _10884_ (.A(net476),
    .B(_03332_),
    .C(_03339_),
    .Y(_03343_),
    .D(_03342_));
 sg13g2_o21ai_1 _10885_ (.B1(_03062_),
    .Y(_03344_),
    .A1(net584),
    .A2(_03322_));
 sg13g2_o21ai_1 _10886_ (.B1(_03063_),
    .Y(_03345_),
    .A1(_03343_),
    .A2(_03344_));
 sg13g2_nand2b_1 _10887_ (.Y(_03346_),
    .B(_03345_),
    .A_N(_02826_));
 sg13g2_a21oi_1 _10888_ (.A1(_02987_),
    .A2(_03271_),
    .Y(_03347_),
    .B1(_03346_));
 sg13g2_a21o_2 _10889_ (.A2(_03243_),
    .A1(_02826_),
    .B1(_03347_),
    .X(\debug_rd[1] ));
 sg13g2_mux2_1 _10890_ (.A0(net74),
    .A1(net3641),
    .S(_03181_),
    .X(_00087_));
 sg13g2_mux2_1 _10891_ (.A0(\i_spi.spi_dc ),
    .A1(\debug_rd_r[0] ),
    .S(debug_register_data),
    .X(_03348_));
 sg13g2_mux2_2 _10892_ (.A0(_03348_),
    .A1(\gpio_out[2] ),
    .S(\gpio_out_sel[2] ),
    .X(uo_out[2]));
 sg13g2_mux2_1 _10893_ (.A0(debug_uart_txd),
    .A1(\gpio_out[6] ),
    .S(\gpio_out_sel[6] ),
    .X(uo_out[6]));
 sg13g2_nand2b_1 _10894_ (.Y(_03349_),
    .B(_03231_),
    .A_N(net572));
 sg13g2_a21oi_1 _10895_ (.A1(net572),
    .A2(_03208_),
    .Y(_03350_),
    .B1(_02842_));
 sg13g2_or2_1 _10896_ (.X(_03351_),
    .B(_02401_),
    .A(_02295_));
 sg13g2_a21oi_1 _10897_ (.A1(_02295_),
    .A2(_02401_),
    .Y(_03352_),
    .B1(_02833_));
 sg13g2_nand2_1 _10898_ (.Y(_03353_),
    .A(_03351_),
    .B(_03352_));
 sg13g2_nand2b_1 _10899_ (.Y(_03354_),
    .B(_02836_),
    .A_N(_02492_));
 sg13g2_o21ai_1 _10900_ (.B1(\i_tinyqv.cpu.alu_op[0] ),
    .Y(_03355_),
    .A1(_02373_),
    .A2(_02398_));
 sg13g2_nand3_1 _10901_ (.B(_02837_),
    .C(_03355_),
    .A(_02491_),
    .Y(_03356_));
 sg13g2_nand3_1 _10902_ (.B(_03354_),
    .C(_03356_),
    .A(_03353_),
    .Y(_03357_));
 sg13g2_nand2b_1 _10903_ (.Y(_03358_),
    .B(_02831_),
    .A_N(_03357_));
 sg13g2_xnor2_1 _10904_ (.Y(_03359_),
    .A(_02562_),
    .B(_02563_));
 sg13g2_a21oi_1 _10905_ (.A1(_02830_),
    .A2(_03359_),
    .Y(_03360_),
    .B1(_02841_));
 sg13g2_a22oi_1 _10906_ (.Y(_03361_),
    .B1(_03358_),
    .B2(_03360_),
    .A2(_03350_),
    .A1(_03349_));
 sg13g2_nand2b_1 _10907_ (.Y(_03362_),
    .B(_03185_),
    .A_N(_03361_));
 sg13g2_o21ai_1 _10908_ (.B1(_03362_),
    .Y(_03363_),
    .A1(_00235_),
    .A2(_02829_));
 sg13g2_a21oi_1 _10909_ (.A1(_02392_),
    .A2(_02395_),
    .Y(_03364_),
    .B1(_02519_));
 sg13g2_nand3_1 _10910_ (.B(net609),
    .C(_03244_),
    .A(\i_tinyqv.cpu.instr_data_start[22] ),
    .Y(_03365_));
 sg13g2_a21o_1 _10911_ (.A2(_03244_),
    .A1(net609),
    .B1(\i_tinyqv.cpu.instr_data_start[22] ),
    .X(_03366_));
 sg13g2_nand2_1 _10912_ (.Y(_03367_),
    .A(_03365_),
    .B(_03366_));
 sg13g2_xnor2_1 _10913_ (.Y(_03368_),
    .A(\i_tinyqv.cpu.instr_data_start[18] ),
    .B(_03002_));
 sg13g2_a21oi_1 _10914_ (.A1(net593),
    .A2(_03367_),
    .Y(_03369_),
    .B1(_03007_));
 sg13g2_o21ai_1 _10915_ (.B1(_03369_),
    .Y(_03370_),
    .A1(net593),
    .A2(_03368_));
 sg13g2_xnor2_1 _10916_ (.Y(_03371_),
    .A(_02990_),
    .B(_02991_));
 sg13g2_a21o_1 _10917_ (.A2(_02999_),
    .A1(net614),
    .B1(net613),
    .X(_03372_));
 sg13g2_and2_1 _10918_ (.A(_03000_),
    .B(_03372_),
    .X(_03373_));
 sg13g2_a22oi_1 _10919_ (.Y(_03374_),
    .B1(_03373_),
    .B2(net457),
    .A2(_03371_),
    .A1(net461));
 sg13g2_nor2_1 _10920_ (.A(net585),
    .B(_03374_),
    .Y(_03375_));
 sg13g2_xnor2_1 _10921_ (.Y(_03376_),
    .A(_01516_),
    .B(_02997_));
 sg13g2_a21oi_1 _10922_ (.A1(\i_tinyqv.cpu.instr_data_start[5] ),
    .A2(_02994_),
    .Y(_03377_),
    .B1(\i_tinyqv.cpu.instr_data_start[6] ));
 sg13g2_nor2_1 _10923_ (.A(_02995_),
    .B(_03377_),
    .Y(_03378_));
 sg13g2_a221oi_1 _10924_ (.B2(net353),
    .C1(_03375_),
    .B1(_03378_),
    .A1(_02254_),
    .Y(_03379_),
    .A2(_03376_));
 sg13g2_a21oi_1 _10925_ (.A1(_03370_),
    .A2(_03379_),
    .Y(_03380_),
    .B1(_02518_));
 sg13g2_a22oi_1 _10926_ (.Y(_03381_),
    .B1(_03046_),
    .B2(_03287_),
    .A2(_03045_),
    .A1(\i_tinyqv.cpu.i_core.mie[2] ));
 sg13g2_nor2_1 _10927_ (.A(_03042_),
    .B(_03381_),
    .Y(_03382_));
 sg13g2_nand2_1 _10928_ (.Y(_03383_),
    .A(net596),
    .B(net456));
 sg13g2_o21ai_1 _10929_ (.B1(net334),
    .Y(_03384_),
    .A1(_03050_),
    .A2(_03383_));
 sg13g2_a21o_1 _10930_ (.A2(_03040_),
    .A1(\i_tinyqv.cpu.i_core.mcause[2] ),
    .B1(_03051_),
    .X(_03385_));
 sg13g2_a21oi_1 _10931_ (.A1(_03384_),
    .A2(_03385_),
    .Y(_03386_),
    .B1(_03382_));
 sg13g2_and2_1 _10932_ (.A(_03035_),
    .B(_03043_),
    .X(_03387_));
 sg13g2_and2_1 _10933_ (.A(net315),
    .B(_03387_),
    .X(_03388_));
 sg13g2_a22oi_1 _10934_ (.Y(_03389_),
    .B1(_03388_),
    .B2(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .A2(_03029_),
    .A1(\i_tinyqv.cpu.i_core.mepc[2] ));
 sg13g2_nand2_1 _10935_ (.Y(_03390_),
    .A(\i_tinyqv.cpu.i_core.cycle_count[2] ),
    .B(_03036_));
 sg13g2_mux2_1 _10936_ (.A0(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .A1(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .S(net313),
    .X(_03391_));
 sg13g2_a22oi_1 _10937_ (.Y(_03392_),
    .B1(_03391_),
    .B2(_03033_),
    .A2(_03039_),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.data[2] ));
 sg13g2_nand4_1 _10938_ (.B(_03389_),
    .C(_03390_),
    .A(_03386_),
    .Y(_03393_),
    .D(_03392_));
 sg13g2_a221oi_1 _10939_ (.B2(_03393_),
    .C1(_03380_),
    .B1(_03020_),
    .A1(net570),
    .Y(_03394_),
    .A2(\i_tinyqv.cpu.is_lui ));
 sg13g2_or2_1 _10940_ (.X(_03395_),
    .B(_03394_),
    .A(_03364_));
 sg13g2_mux4_1 _10941_ (.S0(net591),
    .A0(\i_tinyqv.cpu.instr_data_in[10] ),
    .A1(\i_tinyqv.cpu.instr_data_in[14] ),
    .A2(\i_tinyqv.cpu.instr_data_in[2] ),
    .A3(\i_tinyqv.cpu.instr_data_in[6] ),
    .S1(net108),
    .X(_03396_));
 sg13g2_nand2_1 _10942_ (.Y(_03397_),
    .A(net293),
    .B(uo_out[6]));
 sg13g2_nand2_1 _10943_ (.Y(_03398_),
    .A(\gpio_out_sel[6] ),
    .B(net307));
 sg13g2_a22oi_1 _10944_ (.Y(_03399_),
    .B1(net289),
    .B2(\i_uart_rx.recieved_data[6] ),
    .A2(net294),
    .A1(\i_spi.data[6] ));
 sg13g2_a21oi_1 _10945_ (.A1(\controller1_data[6] ),
    .A2(net291),
    .Y(_03400_),
    .B1(net472));
 sg13g2_a22oi_1 _10946_ (.Y(_03401_),
    .B1(net287),
    .B2(\controller2_data[6] ),
    .A2(net298),
    .A1(\i_time.l_mtimecmp.data_out[6] ));
 sg13g2_nand4_1 _10947_ (.B(_03399_),
    .C(_03400_),
    .A(_03398_),
    .Y(_03402_),
    .D(_03401_));
 sg13g2_a221oi_1 _10948_ (.B2(\i_time.mtime[6] ),
    .C1(_03402_),
    .B1(net221),
    .A1(net8),
    .Y(_03403_),
    .A2(_03084_));
 sg13g2_nand2_1 _10949_ (.Y(_03404_),
    .A(net293),
    .B(uo_out[2]));
 sg13g2_nand2_1 _10950_ (.Y(_03405_),
    .A(\controller2_data[2] ),
    .B(net287));
 sg13g2_a21oi_1 _10951_ (.A1(\gpio_out_sel[2] ),
    .A2(net307),
    .Y(_03406_),
    .B1(net592));
 sg13g2_o21ai_1 _10952_ (.B1(_03406_),
    .Y(_03407_),
    .A1(_01645_),
    .A2(_03069_));
 sg13g2_a21oi_1 _10953_ (.A1(net4),
    .A2(_03084_),
    .Y(_03408_),
    .B1(_03407_));
 sg13g2_a22oi_1 _10954_ (.Y(_03409_),
    .B1(net289),
    .B2(\i_uart_rx.recieved_data[2] ),
    .A2(net291),
    .A1(\controller1_data[2] ));
 sg13g2_a22oi_1 _10955_ (.Y(_03410_),
    .B1(net221),
    .B2(\i_time.mtime[2] ),
    .A2(net294),
    .A1(\i_spi.data[2] ));
 sg13g2_and4_1 _10956_ (.A(_03404_),
    .B(_03405_),
    .C(_03409_),
    .D(_03410_),
    .X(_03411_));
 sg13g2_a22oi_1 _10957_ (.Y(_03412_),
    .B1(_03408_),
    .B2(_03411_),
    .A2(_03403_),
    .A1(_03397_));
 sg13g2_o21ai_1 _10958_ (.B1(net427),
    .Y(_03413_),
    .A1(net116),
    .A2(_03412_));
 sg13g2_nor2_1 _10959_ (.A(net592),
    .B(\i_latch_mem.data_out[2] ),
    .Y(_03414_));
 sg13g2_o21ai_1 _10960_ (.B1(net634),
    .Y(_03415_),
    .A1(net472),
    .A2(\i_latch_mem.data_out[6] ));
 sg13g2_o21ai_1 _10961_ (.B1(_03413_),
    .Y(_03416_),
    .A1(_03414_),
    .A2(_03415_));
 sg13g2_o21ai_1 _10962_ (.B1(_03416_),
    .Y(_03417_),
    .A1(net415),
    .A2(_03396_));
 sg13g2_nor2_1 _10963_ (.A(\i_tinyqv.cpu.instr_data_in[10] ),
    .B(_03132_),
    .Y(_03418_));
 sg13g2_nor2_1 _10964_ (.A(\i_time.l_mtimecmp.data_out[10] ),
    .B(_03069_),
    .Y(_03419_));
 sg13g2_a22oi_1 _10965_ (.Y(_03420_),
    .B1(net287),
    .B2(\controller2_data[10] ),
    .A2(net291),
    .A1(\controller1_data[10] ));
 sg13g2_o21ai_1 _10966_ (.B1(net419),
    .Y(_03421_),
    .A1(\i_tinyqv.mem.qspi_data_buf[10] ),
    .A2(net106));
 sg13g2_a21oi_1 _10967_ (.A1(net634),
    .A2(_01676_),
    .Y(_03422_),
    .B1(net421));
 sg13g2_a21oi_1 _10968_ (.A1(\i_time.mtime[10] ),
    .A2(net220),
    .Y(_03423_),
    .B1(net298));
 sg13g2_o21ai_1 _10969_ (.B1(_03420_),
    .Y(_03424_),
    .A1(_03419_),
    .A2(_03423_));
 sg13g2_o21ai_1 _10970_ (.B1(_03422_),
    .Y(_03425_),
    .A1(net116),
    .A2(_03424_));
 sg13g2_o21ai_1 _10971_ (.B1(_03425_),
    .Y(_03426_),
    .A1(_03418_),
    .A2(_03421_));
 sg13g2_a21oi_1 _10972_ (.A1(_01675_),
    .A2(net105),
    .Y(_03427_),
    .B1(net415));
 sg13g2_o21ai_1 _10973_ (.B1(_03427_),
    .Y(_03428_),
    .A1(\i_tinyqv.mem.qspi_data_buf[14] ),
    .A2(net106));
 sg13g2_o21ai_1 _10974_ (.B1(net415),
    .Y(_03429_),
    .A1(net427),
    .A2(\i_latch_mem.data_out[14] ));
 sg13g2_a21oi_1 _10975_ (.A1(\i_time.mtime[14] ),
    .A2(net220),
    .Y(_03430_),
    .B1(net297));
 sg13g2_a21oi_2 _10976_ (.B1(_03430_),
    .Y(_03431_),
    .A2(net297),
    .A1(_01636_));
 sg13g2_nor2_1 _10977_ (.A(net116),
    .B(_03431_),
    .Y(_03432_));
 sg13g2_o21ai_1 _10978_ (.B1(_03428_),
    .Y(_03433_),
    .A1(_03429_),
    .A2(_03432_));
 sg13g2_a221oi_1 _10979_ (.B2(net460),
    .C1(net583),
    .B1(_03433_),
    .A1(net467),
    .Y(_03434_),
    .A2(_03426_));
 sg13g2_o21ai_1 _10980_ (.B1(_03434_),
    .Y(_03435_),
    .A1(net588),
    .A2(_03417_));
 sg13g2_mux4_1 _10981_ (.S0(net591),
    .A0(\i_tinyqv.cpu.instr_data_in[10] ),
    .A1(\i_tinyqv.cpu.instr_data_in[14] ),
    .A2(\i_tinyqv.mem.qspi_data_buf[26] ),
    .A3(\i_tinyqv.mem.qspi_data_buf[30] ),
    .S1(net117),
    .X(_03436_));
 sg13g2_nor2_1 _10982_ (.A(net415),
    .B(_03436_),
    .Y(_03437_));
 sg13g2_mux4_1 _10983_ (.S0(net473),
    .A0(\i_time.mtime[30] ),
    .A1(\i_time.mtime[26] ),
    .A2(\i_time.l_mtimecmp.data_out[30] ),
    .A3(\i_time.l_mtimecmp.data_out[26] ),
    .S1(net301),
    .X(_03438_));
 sg13g2_o21ai_1 _10984_ (.B1(net635),
    .Y(_03439_),
    .A1(net590),
    .A2(_01681_));
 sg13g2_a21oi_1 _10985_ (.A1(net590),
    .A2(\i_latch_mem.data_out[30] ),
    .Y(_03440_),
    .B1(_03439_));
 sg13g2_a21oi_1 _10986_ (.A1(net183),
    .A2(_03438_),
    .Y(_03441_),
    .B1(net116));
 sg13g2_nor4_1 _10987_ (.A(_01581_),
    .B(_03437_),
    .C(_03440_),
    .D(_03441_),
    .Y(_03442_));
 sg13g2_a221oi_1 _10988_ (.B2(net418),
    .C1(_02169_),
    .B1(_01678_),
    .A1(net637),
    .Y(_03443_),
    .A2(_01677_));
 sg13g2_a221oi_1 _10989_ (.B2(net418),
    .C1(_02164_),
    .B1(_01680_),
    .A1(net637),
    .Y(_03444_),
    .A2(_01679_));
 sg13g2_nor2_1 _10990_ (.A(\i_time.l_mtimecmp.data_out[22] ),
    .B(net295),
    .Y(_03445_));
 sg13g2_nor2_1 _10991_ (.A(\i_time.l_mtimecmp.data_out[18] ),
    .B(net295),
    .Y(_03446_));
 sg13g2_a21oi_1 _10992_ (.A1(\i_time.mtime[18] ),
    .A2(net220),
    .Y(_03447_),
    .B1(net300));
 sg13g2_o21ai_1 _10993_ (.B1(net114),
    .Y(_03448_),
    .A1(_03446_),
    .A2(_03447_));
 sg13g2_a21oi_1 _10994_ (.A1(\i_time.mtime[22] ),
    .A2(net220),
    .Y(_03449_),
    .B1(net301));
 sg13g2_o21ai_1 _10995_ (.B1(net114),
    .Y(_03450_),
    .A1(_03445_),
    .A2(_03449_));
 sg13g2_a221oi_1 _10996_ (.B2(_03444_),
    .C1(_03442_),
    .B1(_03450_),
    .A1(_03443_),
    .Y(_03451_),
    .A2(_03448_));
 sg13g2_a21oi_1 _10997_ (.A1(net584),
    .A2(_03451_),
    .Y(_03452_),
    .B1(_03061_));
 sg13g2_nand2_2 _10998_ (.Y(_03453_),
    .A(_03435_),
    .B(_03452_));
 sg13g2_a221oi_1 _10999_ (.B2(_03063_),
    .C1(_02826_),
    .B1(_03453_),
    .A1(_02987_),
    .Y(_03454_),
    .A2(_03395_));
 sg13g2_a21o_2 _11000_ (.A2(_03363_),
    .A1(_02826_),
    .B1(_03454_),
    .X(\debug_rd[2] ));
 sg13g2_mux2_1 _11001_ (.A0(net81),
    .A1(net3650),
    .S(_03181_),
    .X(_00088_));
 sg13g2_mux2_1 _11002_ (.A0(\i_spi.data[7] ),
    .A1(\debug_rd_r[1] ),
    .S(debug_register_data),
    .X(_03455_));
 sg13g2_mux2_2 _11003_ (.A0(_03455_),
    .A1(\gpio_out[3] ),
    .S(\gpio_out_sel[3] ),
    .X(uo_out[3]));
 sg13g2_nand2_1 _11004_ (.Y(_03456_),
    .A(\gpio_out_sel[8] ),
    .B(\i_pwm.pwm ));
 sg13g2_xor2_1 _11005_ (.B(\i_tinyqv.cpu.i_core.cmp_out ),
    .A(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .X(_03457_));
 sg13g2_nand4_1 _11006_ (.B(_02505_),
    .C(_02524_),
    .A(_00130_),
    .Y(_03458_),
    .D(_03031_));
 sg13g2_and2_2 _11007_ (.A(_00129_),
    .B(_03458_),
    .X(_03459_));
 sg13g2_nand2_2 _11008_ (.Y(_03460_),
    .A(_00129_),
    .B(_03458_));
 sg13g2_and4_1 _11009_ (.A(_00130_),
    .B(_02505_),
    .C(_02524_),
    .D(_03024_),
    .X(_03461_));
 sg13g2_nand4_1 _11010_ (.B(_02505_),
    .C(_02524_),
    .A(_00130_),
    .Y(_03462_),
    .D(_03024_));
 sg13g2_nand3_1 _11011_ (.B(_03459_),
    .C(net341),
    .A(_02518_),
    .Y(_03463_));
 sg13g2_a21o_1 _11012_ (.A2(_03457_),
    .A1(net414),
    .B1(_03463_),
    .X(_03464_));
 sg13g2_and2_1 _11013_ (.A(net407),
    .B(_03464_),
    .X(_03465_));
 sg13g2_nand2_1 _11014_ (.Y(_03466_),
    .A(net407),
    .B(_03464_));
 sg13g2_nand2_1 _11015_ (.Y(_03467_),
    .A(_00134_),
    .B(net99));
 sg13g2_nand2_1 _11016_ (.Y(_03468_),
    .A(\i_tinyqv.cpu.i_core.mip[0] ),
    .B(\i_tinyqv.cpu.i_core.mie[0] ));
 sg13g2_a22oi_1 _11017_ (.Y(_03469_),
    .B1(\i_tinyqv.cpu.i_core.mie[1] ),
    .B2(\i_tinyqv.cpu.i_core.mip[1] ),
    .A2(\i_tinyqv.cpu.i_core.mie[0] ),
    .A1(\i_tinyqv.cpu.i_core.mip[0] ));
 sg13g2_inv_1 _11018_ (.Y(_03470_),
    .A(_03469_));
 sg13g2_a21oi_1 _11019_ (.A1(\i_tinyqv.cpu.i_core.mie[2] ),
    .A2(_03287_),
    .Y(_03471_),
    .B1(_03470_));
 sg13g2_nor2_1 _11020_ (.A(_00166_),
    .B(_03099_),
    .Y(_03472_));
 sg13g2_nand2_1 _11021_ (.Y(_03473_),
    .A(\i_tinyqv.cpu.i_core.mie[4] ),
    .B(\i_time.timer_interrupt ));
 sg13g2_nor2b_1 _11022_ (.A(_03472_),
    .B_N(_03473_),
    .Y(_03474_));
 sg13g2_a21oi_2 _11023_ (.B1(_01576_),
    .Y(_03475_),
    .A2(_03474_),
    .A1(_03471_));
 sg13g2_nor2_1 _11024_ (.A(net568),
    .B(_00137_),
    .Y(_03476_));
 sg13g2_a21oi_2 _11025_ (.B1(_03476_),
    .Y(_03477_),
    .A2(_03371_),
    .A1(net568));
 sg13g2_a21o_2 _11026_ (.A2(_03371_),
    .A1(net568),
    .B1(_03476_),
    .X(_03478_));
 sg13g2_nor2_1 _11027_ (.A(net568),
    .B(_00136_),
    .Y(_03479_));
 sg13g2_a21oi_2 _11028_ (.B1(_03479_),
    .Y(_03480_),
    .A2(_03252_),
    .A1(net568));
 sg13g2_a21o_2 _11029_ (.A2(_03252_),
    .A1(net568),
    .B1(_03479_),
    .X(_03481_));
 sg13g2_nand2_1 _11030_ (.Y(_03482_),
    .A(_01600_),
    .B(net449));
 sg13g2_mux4_1 _11031_ (.S0(_03480_),
    .A0(\i_tinyqv.cpu.instr_data[1][0] ),
    .A1(\i_tinyqv.cpu.instr_data[0][0] ),
    .A2(\i_tinyqv.cpu.instr_data[3][0] ),
    .A3(\i_tinyqv.cpu.instr_data[2][0] ),
    .S1(_03478_),
    .X(_03483_));
 sg13g2_inv_1 _11032_ (.Y(_03484_),
    .A(_03483_));
 sg13g2_mux4_1 _11033_ (.S0(net438),
    .A0(_00138_),
    .A1(_00139_),
    .A2(_00140_),
    .A3(_00141_),
    .S1(net449),
    .X(_03485_));
 sg13g2_inv_1 _11034_ (.Y(_03486_),
    .A(_03485_));
 sg13g2_nor2_2 _11035_ (.A(_03484_),
    .B(_03485_),
    .Y(_03487_));
 sg13g2_nand2_1 _11036_ (.Y(_03488_),
    .A(_03483_),
    .B(net286));
 sg13g2_xnor2_1 _11037_ (.Y(_03489_),
    .A(\i_tinyqv.cpu.instr_write_offset[1] ),
    .B(net438));
 sg13g2_and2_1 _11038_ (.A(_00131_),
    .B(_03481_),
    .X(_03490_));
 sg13g2_nor2b_1 _11039_ (.A(_00135_),
    .B_N(_02992_),
    .Y(_03491_));
 sg13g2_xnor2_1 _11040_ (.Y(_03492_),
    .A(\i_tinyqv.cpu.instr_write_offset[3] ),
    .B(_03491_));
 sg13g2_a22oi_1 _11041_ (.Y(_03493_),
    .B1(_03490_),
    .B2(_03492_),
    .A2(_03478_),
    .A1(_01597_));
 sg13g2_o21ai_1 _11042_ (.B1(_03492_),
    .Y(_03494_),
    .A1(_01597_),
    .A2(net449));
 sg13g2_a21oi_1 _11043_ (.A1(_03490_),
    .A2(_03494_),
    .Y(_03495_),
    .B1(_03493_));
 sg13g2_a221oi_1 _11044_ (.B2(_03494_),
    .C1(_03495_),
    .B1(_03493_),
    .A1(net219),
    .Y(_03496_),
    .A2(_03489_));
 sg13g2_nand2b_2 _11045_ (.Y(_03497_),
    .B(_00134_),
    .A_N(_03496_));
 sg13g2_a21o_1 _11046_ (.A2(_03475_),
    .A1(_02528_),
    .B1(_03497_),
    .X(_03498_));
 sg13g2_a221oi_1 _11047_ (.B2(_02528_),
    .C1(_03497_),
    .B1(_03475_),
    .A1(net407),
    .Y(_03499_),
    .A2(_03464_));
 sg13g2_or2_1 _11048_ (.X(_03500_),
    .B(\i_tinyqv.cpu.additional_mem_ops[0] ),
    .A(\i_tinyqv.cpu.additional_mem_ops[1] ));
 sg13g2_nor2_2 _11049_ (.A(\i_tinyqv.cpu.additional_mem_ops[2] ),
    .B(_03500_),
    .Y(_03501_));
 sg13g2_inv_4 _11050_ (.A(_03501_),
    .Y(_03502_));
 sg13g2_nand2_2 _11051_ (.Y(_03503_),
    .A(_02529_),
    .B(_03501_));
 sg13g2_nor2_1 _11052_ (.A(net571),
    .B(net313),
    .Y(_03504_));
 sg13g2_a21o_1 _11053_ (.A2(_03501_),
    .A1(_02529_),
    .B1(_03504_),
    .X(_03505_));
 sg13g2_and2_1 _11054_ (.A(_03499_),
    .B(_03505_),
    .X(_03506_));
 sg13g2_nor2_2 _11055_ (.A(_03484_),
    .B(net286),
    .Y(_03507_));
 sg13g2_nand2b_1 _11056_ (.Y(_03508_),
    .B(net440),
    .A_N(_00160_));
 sg13g2_o21ai_1 _11057_ (.B1(_03508_),
    .Y(_03509_),
    .A1(_00158_),
    .A2(net440));
 sg13g2_nand2_1 _11058_ (.Y(_03510_),
    .A(_00161_),
    .B(net440));
 sg13g2_a21oi_1 _11059_ (.A1(_00159_),
    .A2(net450),
    .Y(_03511_),
    .B1(net434));
 sg13g2_a22oi_1 _11060_ (.Y(_03512_),
    .B1(_03510_),
    .B2(_03511_),
    .A2(_03509_),
    .A1(net434));
 sg13g2_nand2b_1 _11061_ (.Y(_03513_),
    .B(net445),
    .A_N(_00156_));
 sg13g2_o21ai_1 _11062_ (.B1(_03513_),
    .Y(_03514_),
    .A1(_00154_),
    .A2(net445));
 sg13g2_nand2_1 _11063_ (.Y(_03515_),
    .A(_00157_),
    .B(net444));
 sg13g2_a21oi_1 _11064_ (.A1(_00155_),
    .A2(net451),
    .Y(_03516_),
    .B1(net436));
 sg13g2_a22oi_1 _11065_ (.Y(_03517_),
    .B1(_03515_),
    .B2(_03516_),
    .A2(_03514_),
    .A1(net436));
 sg13g2_inv_2 _11066_ (.Y(_03518_),
    .A(net210));
 sg13g2_nor2b_2 _11067_ (.A(net210),
    .B_N(net211),
    .Y(_03519_));
 sg13g2_and2_1 _11068_ (.A(_03507_),
    .B(_03519_),
    .X(_03520_));
 sg13g2_nand2_2 _11069_ (.Y(_03521_),
    .A(_03507_),
    .B(_03519_));
 sg13g2_mux4_1 _11070_ (.S0(net438),
    .A0(\i_tinyqv.cpu.instr_data[1][3] ),
    .A1(\i_tinyqv.cpu.instr_data[0][3] ),
    .A2(\i_tinyqv.cpu.instr_data[3][3] ),
    .A3(\i_tinyqv.cpu.instr_data[2][3] ),
    .S1(net448),
    .X(_03522_));
 sg13g2_nand2b_1 _11071_ (.Y(_03523_),
    .B(net447),
    .A_N(_00152_));
 sg13g2_o21ai_1 _11072_ (.B1(_03523_),
    .Y(_03524_),
    .A1(_00150_),
    .A2(net447));
 sg13g2_nand2_1 _11073_ (.Y(_03525_),
    .A(_00153_),
    .B(net447));
 sg13g2_a21oi_1 _11074_ (.A1(_00151_),
    .A2(net451),
    .Y(_03526_),
    .B1(net436));
 sg13g2_a22oi_1 _11075_ (.Y(_03527_),
    .B1(_03525_),
    .B2(_03526_),
    .A2(_03524_),
    .A1(net436));
 sg13g2_inv_2 _11076_ (.Y(_03528_),
    .A(net208));
 sg13g2_nand2b_1 _11077_ (.Y(_03529_),
    .B(net441),
    .A_N(_00148_));
 sg13g2_o21ai_1 _11078_ (.B1(_03529_),
    .Y(_03530_),
    .A1(_00146_),
    .A2(net441));
 sg13g2_nand2_1 _11079_ (.Y(_03531_),
    .A(_00149_),
    .B(net441));
 sg13g2_a21oi_1 _11080_ (.A1(_00147_),
    .A2(net450),
    .Y(_03532_),
    .B1(net436));
 sg13g2_a22oi_1 _11081_ (.Y(_03533_),
    .B1(_03531_),
    .B2(_03532_),
    .A2(_03530_),
    .A1(net436));
 sg13g2_inv_2 _11082_ (.Y(_03534_),
    .A(_03533_));
 sg13g2_nand2_2 _11083_ (.Y(_03535_),
    .A(_03528_),
    .B(_03534_));
 sg13g2_nand2b_1 _11084_ (.Y(_03536_),
    .B(net446),
    .A_N(\i_tinyqv.cpu.instr_data[3][2] ));
 sg13g2_mux4_1 _11085_ (.S0(net438),
    .A0(\i_tinyqv.cpu.instr_data[1][2] ),
    .A1(\i_tinyqv.cpu.instr_data[0][2] ),
    .A2(\i_tinyqv.cpu.instr_data[3][2] ),
    .A3(\i_tinyqv.cpu.instr_data[2][2] ),
    .S1(net446),
    .X(_03537_));
 sg13g2_nand2b_1 _11086_ (.Y(_03538_),
    .B(net446),
    .A_N(_00144_));
 sg13g2_o21ai_1 _11087_ (.B1(_03538_),
    .Y(_03539_),
    .A1(_00142_),
    .A2(net446));
 sg13g2_mux2_1 _11088_ (.A0(_00143_),
    .A1(_00145_),
    .S(net446),
    .X(_03540_));
 sg13g2_nor2_1 _11089_ (.A(net438),
    .B(_03539_),
    .Y(_03541_));
 sg13g2_a21oi_2 _11090_ (.B1(_03541_),
    .Y(_03542_),
    .A2(_03540_),
    .A1(net438));
 sg13g2_nor2_1 _11091_ (.A(_03535_),
    .B(net119),
    .Y(_03543_));
 sg13g2_nand2_1 _11092_ (.Y(_03544_),
    .A(net283),
    .B(_03543_));
 sg13g2_nor2b_2 _11093_ (.A(_03544_),
    .B_N(net332),
    .Y(_03545_));
 sg13g2_nand3_1 _11094_ (.B(net283),
    .C(_03543_),
    .A(net332),
    .Y(_03546_));
 sg13g2_o21ai_1 _11095_ (.B1(_03521_),
    .Y(_03547_),
    .A1(net217),
    .A2(_03546_));
 sg13g2_nand4_1 _11096_ (.B(_03499_),
    .C(_03505_),
    .A(net659),
    .Y(_03548_),
    .D(_03547_));
 sg13g2_nand2_1 _11097_ (.Y(_03549_),
    .A(net211),
    .B(_03517_));
 sg13g2_nand2b_1 _11098_ (.Y(_03550_),
    .B(net439),
    .A_N(_00164_));
 sg13g2_o21ai_1 _11099_ (.B1(_03550_),
    .Y(_03551_),
    .A1(_00162_),
    .A2(net439));
 sg13g2_nand2_1 _11100_ (.Y(_03552_),
    .A(_00165_),
    .B(net439));
 sg13g2_a21oi_1 _11101_ (.A1(_00163_),
    .A2(net450),
    .Y(_03553_),
    .B1(net434));
 sg13g2_a22oi_1 _11102_ (.Y(_03554_),
    .B1(_03552_),
    .B2(_03553_),
    .A2(_03551_),
    .A1(net434));
 sg13g2_or2_2 _11103_ (.X(_03555_),
    .B(_03554_),
    .A(_03483_));
 sg13g2_nor2_2 _11104_ (.A(net333),
    .B(_03555_),
    .Y(_03556_));
 sg13g2_nor3_2 _11105_ (.A(net333),
    .B(net118),
    .C(_03555_),
    .Y(_03557_));
 sg13g2_nor2_2 _11106_ (.A(net332),
    .B(net283),
    .Y(_03558_));
 sg13g2_nand2b_2 _11107_ (.Y(_03559_),
    .B(_03558_),
    .A_N(net119));
 sg13g2_inv_1 _11108_ (.Y(_03560_),
    .A(_03559_));
 sg13g2_nand2_2 _11109_ (.Y(_03561_),
    .A(net208),
    .B(_03533_));
 sg13g2_nor2_2 _11110_ (.A(_03559_),
    .B(_03561_),
    .Y(_03562_));
 sg13g2_and2_1 _11111_ (.A(_03557_),
    .B(_03562_),
    .X(_03563_));
 sg13g2_nand2_2 _11112_ (.Y(_03564_),
    .A(_03557_),
    .B(_03562_));
 sg13g2_nand2b_1 _11113_ (.Y(_03565_),
    .B(net439),
    .A_N(_00181_));
 sg13g2_o21ai_1 _11114_ (.B1(_03565_),
    .Y(_03566_),
    .A1(_00179_),
    .A2(net439));
 sg13g2_nand2_1 _11115_ (.Y(_03567_),
    .A(_00182_),
    .B(net439));
 sg13g2_a21oi_1 _11116_ (.A1(_00180_),
    .A2(net450),
    .Y(_03568_),
    .B1(net434));
 sg13g2_a22oi_1 _11117_ (.Y(_03569_),
    .B1(_03567_),
    .B2(_03568_),
    .A2(_03566_),
    .A1(net434));
 sg13g2_inv_2 _11118_ (.Y(_03570_),
    .A(_03569_));
 sg13g2_nand2b_1 _11119_ (.Y(_03571_),
    .B(net444),
    .A_N(_00177_));
 sg13g2_o21ai_1 _11120_ (.B1(_03571_),
    .Y(_03572_),
    .A1(_00175_),
    .A2(net444));
 sg13g2_nand2_1 _11121_ (.Y(_03573_),
    .A(_00178_),
    .B(net445));
 sg13g2_a21oi_1 _11122_ (.A1(_00176_),
    .A2(net450),
    .Y(_03574_),
    .B1(net437));
 sg13g2_a22oi_1 _11123_ (.Y(_03575_),
    .B1(_03573_),
    .B2(_03574_),
    .A2(_03572_),
    .A1(net437));
 sg13g2_and2_1 _11124_ (.A(_03569_),
    .B(_03575_),
    .X(_03576_));
 sg13g2_nand2b_1 _11125_ (.Y(_03577_),
    .B(net451),
    .A_N(_00183_));
 sg13g2_nand2b_1 _11126_ (.Y(_03578_),
    .B(net447),
    .A_N(_00185_));
 sg13g2_a21oi_1 _11127_ (.A1(_03577_),
    .A2(_03578_),
    .Y(_03579_),
    .B1(net438));
 sg13g2_a21oi_1 _11128_ (.A1(_00186_),
    .A2(net447),
    .Y(_03580_),
    .B1(net436));
 sg13g2_o21ai_1 _11129_ (.B1(_03580_),
    .Y(_03581_),
    .A1(_01603_),
    .A2(net447));
 sg13g2_nor2b_2 _11130_ (.A(_03579_),
    .B_N(_03581_),
    .Y(_03582_));
 sg13g2_nand2b_2 _11131_ (.Y(_03583_),
    .B(_03581_),
    .A_N(_03579_));
 sg13g2_nand2b_1 _11132_ (.Y(_03584_),
    .B(net441),
    .A_N(_00169_));
 sg13g2_o21ai_1 _11133_ (.B1(_03584_),
    .Y(_03585_),
    .A1(_00167_),
    .A2(net442));
 sg13g2_nand2_1 _11134_ (.Y(_03586_),
    .A(_00170_),
    .B(net442));
 sg13g2_a21oi_1 _11135_ (.A1(_00168_),
    .A2(net450),
    .Y(_03587_),
    .B1(net435));
 sg13g2_a22oi_1 _11136_ (.Y(_03588_),
    .B1(_03586_),
    .B2(_03587_),
    .A2(_03585_),
    .A1(net435));
 sg13g2_nand2b_1 _11137_ (.Y(_03589_),
    .B(net444),
    .A_N(_00173_));
 sg13g2_o21ai_1 _11138_ (.B1(_03589_),
    .Y(_03590_),
    .A1(_00171_),
    .A2(net442));
 sg13g2_nand2_1 _11139_ (.Y(_03591_),
    .A(_00174_),
    .B(net441));
 sg13g2_a21oi_1 _11140_ (.A1(_00172_),
    .A2(net450),
    .Y(_03592_),
    .B1(net434));
 sg13g2_a22oi_1 _11141_ (.Y(_03593_),
    .B1(_03591_),
    .B2(_03592_),
    .A2(_03590_),
    .A1(net434));
 sg13g2_nand2_1 _11142_ (.Y(_03594_),
    .A(_03576_),
    .B(net204));
 sg13g2_nor4_2 _11143_ (.A(_03564_),
    .B(net205),
    .C(net282),
    .Y(_03595_),
    .D(_03594_));
 sg13g2_nand4_1 _11144_ (.B(_03499_),
    .C(_03505_),
    .A(net656),
    .Y(_03596_),
    .D(_03595_));
 sg13g2_and3_1 _11145_ (.X(_03597_),
    .A(net656),
    .B(_03506_),
    .C(_03595_));
 sg13g2_nand3_1 _11146_ (.B(_03506_),
    .C(_03595_),
    .A(net658),
    .Y(_03598_));
 sg13g2_nand4_1 _11147_ (.B(_03467_),
    .C(_03548_),
    .A(_00132_),
    .Y(_03599_),
    .D(net86));
 sg13g2_nand3_1 _11148_ (.B(_02992_),
    .C(_03501_),
    .A(_02529_),
    .Y(_03600_));
 sg13g2_nor2b_2 _11149_ (.A(net619),
    .B_N(net620),
    .Y(_03601_));
 sg13g2_nand2_1 _11150_ (.Y(_03602_),
    .A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .B(_03601_));
 sg13g2_nand3_1 _11151_ (.B(\i_tinyqv.mem.q_ctrl.data_ready ),
    .C(_03601_),
    .A(\i_tinyqv.mem.instr_active ),
    .Y(_03603_));
 sg13g2_nor2_2 _11152_ (.A(_00132_),
    .B(_03603_),
    .Y(_03604_));
 sg13g2_nor3_1 _11153_ (.A(_00132_),
    .B(_00131_),
    .C(_03603_),
    .Y(_03605_));
 sg13g2_nand2_1 _11154_ (.Y(_03606_),
    .A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(_03605_));
 sg13g2_xor2_1 _11155_ (.B(_03606_),
    .A(\i_tinyqv.cpu.instr_write_offset[3] ),
    .X(_03607_));
 sg13g2_xnor2_1 _11156_ (.Y(_03608_),
    .A(_03600_),
    .B(_03607_));
 sg13g2_xnor2_1 _11157_ (.Y(_03609_),
    .A(net4094),
    .B(_03604_));
 sg13g2_xnor2_1 _11158_ (.Y(_03610_),
    .A(_00136_),
    .B(_03609_));
 sg13g2_xnor2_1 _11159_ (.Y(_03611_),
    .A(net3978),
    .B(_03605_));
 sg13g2_xnor2_1 _11160_ (.Y(_03612_),
    .A(_00137_),
    .B(_03611_));
 sg13g2_or2_1 _11161_ (.X(_03613_),
    .B(_03612_),
    .A(_03610_));
 sg13g2_nand3_1 _11162_ (.B(_03601_),
    .C(_03603_),
    .A(_01604_),
    .Y(_03614_));
 sg13g2_or3_2 _11163_ (.A(_03608_),
    .B(_03613_),
    .C(_03614_),
    .X(_03615_));
 sg13g2_a21o_1 _11164_ (.A2(_03615_),
    .A1(\i_tinyqv.cpu.instr_fetch_started ),
    .B1(_03599_),
    .X(_03616_));
 sg13g2_o21ai_1 _11165_ (.B1(_03602_),
    .Y(_03617_),
    .A1(_03608_),
    .A2(_03613_));
 sg13g2_a21oi_1 _11166_ (.A1(\i_tinyqv.cpu.data_read_n[1] ),
    .A2(\i_tinyqv.cpu.data_read_n[0] ),
    .Y(_03618_),
    .B1(net417));
 sg13g2_o21ai_1 _11167_ (.B1(net420),
    .Y(_03619_),
    .A1(_02531_),
    .A2(_02532_));
 sg13g2_o21ai_1 _11168_ (.B1(_02534_),
    .Y(_03620_),
    .A1(net417),
    .A2(_02530_));
 sg13g2_a21oi_1 _11169_ (.A1(_03617_),
    .A2(_03620_),
    .Y(_03621_),
    .B1(_01524_));
 sg13g2_nor2b_1 _11170_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .B_N(_00193_),
    .Y(_03622_));
 sg13g2_nor2_2 _11171_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .B(net616),
    .Y(_03623_));
 sg13g2_nor2b_1 _11172_ (.A(net616),
    .B_N(_03622_),
    .Y(_03624_));
 sg13g2_nand2_2 _11173_ (.Y(_03625_),
    .A(_00193_),
    .B(_03623_));
 sg13g2_nand2_2 _11174_ (.Y(_03626_),
    .A(net4057),
    .B(net486));
 sg13g2_inv_1 _11175_ (.Y(_03627_),
    .A(_03626_));
 sg13g2_nor2_2 _11176_ (.A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .B(\i_tinyqv.mem.q_ctrl.data_req ),
    .Y(_03628_));
 sg13g2_nor2_1 _11177_ (.A(debug_data_continue),
    .B(_03628_),
    .Y(_03629_));
 sg13g2_a21oi_1 _11178_ (.A1(_02540_),
    .A2(_03629_),
    .Y(_03630_),
    .B1(net4031));
 sg13g2_or2_1 _11179_ (.X(_03631_),
    .B(_03630_),
    .A(_03627_));
 sg13g2_a21o_2 _11180_ (.A2(_03621_),
    .A1(_03616_),
    .B1(_03631_),
    .X(_03632_));
 sg13g2_a21o_1 _11181_ (.A2(_03615_),
    .A1(net5),
    .B1(net662),
    .X(_03633_));
 sg13g2_a21o_1 _11182_ (.A2(_03632_),
    .A1(_01685_),
    .B1(_03633_),
    .X(_03634_));
 sg13g2_o21ai_1 _11183_ (.B1(net662),
    .Y(_03635_),
    .A1(debug_data_continue),
    .A2(net5));
 sg13g2_a21oi_1 _11184_ (.A1(net5),
    .A2(net336),
    .Y(_03636_),
    .B1(_03635_));
 sg13g2_nor2_1 _11185_ (.A(net7),
    .B(_03636_),
    .Y(_03637_));
 sg13g2_a21oi_1 _11186_ (.A1(net5),
    .A2(net86),
    .Y(_03638_),
    .B1(net662));
 sg13g2_o21ai_1 _11187_ (.B1(_03638_),
    .Y(_03639_),
    .A1(net5),
    .A2(_03178_));
 sg13g2_o21ai_1 _11188_ (.B1(net662),
    .Y(_03640_),
    .A1(_01685_),
    .A2(net99));
 sg13g2_a21oi_1 _11189_ (.A1(_01685_),
    .A2(_03548_),
    .Y(_03641_),
    .B1(_03640_));
 sg13g2_nor2_1 _11190_ (.A(_01673_),
    .B(_03641_),
    .Y(_03642_));
 sg13g2_a221oi_1 _11191_ (.B2(_03642_),
    .C1(net8),
    .B1(_03639_),
    .A1(_03634_),
    .Y(_03643_),
    .A2(_03637_));
 sg13g2_nand2_1 _11192_ (.Y(_03644_),
    .A(_01685_),
    .B(_03599_));
 sg13g2_a21oi_1 _11193_ (.A1(_01487_),
    .A2(net5),
    .Y(_03645_),
    .B1(net662));
 sg13g2_a21oi_1 _11194_ (.A1(_02529_),
    .A2(_03501_),
    .Y(_03646_),
    .B1(_01685_));
 sg13g2_a21oi_1 _11195_ (.A1(_01685_),
    .A2(_03603_),
    .Y(_03647_),
    .B1(_03646_));
 sg13g2_a221oi_1 _11196_ (.B2(net662),
    .C1(_01673_),
    .B1(_03647_),
    .A1(_03644_),
    .Y(_03648_),
    .A2(_03645_));
 sg13g2_a21oi_1 _11197_ (.A1(\i_tinyqv.cpu.data_read_n[1] ),
    .A2(\i_tinyqv.cpu.data_read_n[0] ),
    .Y(_03649_),
    .B1(net420));
 sg13g2_mux4_1 _11198_ (.S0(net6),
    .A0(_02983_),
    .A1(_03649_),
    .A2(_03475_),
    .A3(_02076_),
    .S1(_01685_),
    .X(_03650_));
 sg13g2_o21ai_1 _11199_ (.B1(net8),
    .Y(_03651_),
    .A1(net7),
    .A2(_03650_));
 sg13g2_o21ai_1 _11200_ (.B1(_01688_),
    .Y(_03652_),
    .A1(_03648_),
    .A2(_03651_));
 sg13g2_a21oi_1 _11201_ (.A1(\gpio_out_sel[7] ),
    .A2(_01689_),
    .Y(_03653_),
    .B1(\gpio_out_sel[8] ));
 sg13g2_o21ai_1 _11202_ (.B1(_03653_),
    .Y(_03654_),
    .A1(_03643_),
    .A2(_03652_));
 sg13g2_nand2_2 _11203_ (.Y(uo_out[7]),
    .A(_03456_),
    .B(_03654_));
 sg13g2_a21oi_1 _11204_ (.A1(net638),
    .A2(_01690_),
    .Y(_03655_),
    .B1(net421));
 sg13g2_a21oi_1 _11205_ (.A1(_03456_),
    .A2(_03654_),
    .Y(_03656_),
    .B1(_03076_));
 sg13g2_and2_1 _11206_ (.A(\i_spi.data[7] ),
    .B(net294),
    .X(_03657_));
 sg13g2_a21oi_1 _11207_ (.A1(\i_time.mtime[7] ),
    .A2(net221),
    .Y(_03658_),
    .B1(net299));
 sg13g2_a21oi_1 _11208_ (.A1(_01642_),
    .A2(net298),
    .Y(_03659_),
    .B1(_03658_));
 sg13g2_a221oi_1 _11209_ (.B2(\gpio_out_sel[7] ),
    .C1(_03659_),
    .B1(net307),
    .A1(\i_uart_rx.recieved_data[7] ),
    .Y(_03660_),
    .A2(net289));
 sg13g2_a221oi_1 _11210_ (.B2(net9),
    .C1(_03657_),
    .B1(_03084_),
    .A1(\controller2_data[7] ),
    .Y(_03661_),
    .A2(net288));
 sg13g2_a21oi_1 _11211_ (.A1(\controller1_data[7] ),
    .A2(net292),
    .Y(_03662_),
    .B1(net638));
 sg13g2_nand4_1 _11212_ (.B(_03660_),
    .C(_03661_),
    .A(net114),
    .Y(_03663_),
    .D(_03662_));
 sg13g2_o21ai_1 _11213_ (.B1(_03655_),
    .Y(_03664_),
    .A1(_03656_),
    .A2(_03663_));
 sg13g2_mux2_1 _11214_ (.A0(\i_tinyqv.cpu.instr_data_in[15] ),
    .A1(\i_tinyqv.cpu.instr_data_in[7] ),
    .S(net108),
    .X(_03665_));
 sg13g2_nand2_1 _11215_ (.Y(_03666_),
    .A(net418),
    .B(_03665_));
 sg13g2_a21o_1 _11216_ (.A2(_03666_),
    .A1(_03664_),
    .B1(_02164_),
    .X(_03667_));
 sg13g2_and2_1 _11217_ (.A(\gpio_out_sel[3] ),
    .B(_03082_),
    .X(_03668_));
 sg13g2_nor2_1 _11218_ (.A(_01545_),
    .B(_02113_),
    .Y(_03669_));
 sg13g2_and2_1 _11219_ (.A(\i_uart_rx.recieved_data[3] ),
    .B(net289),
    .X(_03670_));
 sg13g2_a21oi_1 _11220_ (.A1(_01537_),
    .A2(net295),
    .Y(_03671_),
    .B1(_03104_));
 sg13g2_o21ai_1 _11221_ (.B1(_03671_),
    .Y(_03672_),
    .A1(\i_time.l_mtimecmp.data_out[15] ),
    .A2(net295));
 sg13g2_a221oi_1 _11222_ (.B2(_03672_),
    .C1(net421),
    .B1(net114),
    .A1(net634),
    .Y(_03673_),
    .A2(_01693_));
 sg13g2_o21ai_1 _11223_ (.B1(net418),
    .Y(_03674_),
    .A1(\i_tinyqv.mem.qspi_data_buf[15] ),
    .A2(net106));
 sg13g2_a21oi_1 _11224_ (.A1(_01687_),
    .A2(net106),
    .Y(_03675_),
    .B1(_03674_));
 sg13g2_o21ai_1 _11225_ (.B1(net419),
    .Y(_03676_),
    .A1(\i_tinyqv.cpu.instr_data_in[11] ),
    .A2(_03132_));
 sg13g2_a21oi_1 _11226_ (.A1(_01691_),
    .A2(_03132_),
    .Y(_03677_),
    .B1(_03676_));
 sg13g2_a21oi_1 _11227_ (.A1(\i_time.mtime[11] ),
    .A2(net220),
    .Y(_03678_),
    .B1(net297));
 sg13g2_a21oi_1 _11228_ (.A1(_01639_),
    .A2(net297),
    .Y(_03679_),
    .B1(_03678_));
 sg13g2_a221oi_1 _11229_ (.B2(\controller2_data[11] ),
    .C1(_03679_),
    .B1(net288),
    .A1(\controller1_data[11] ),
    .Y(_03680_),
    .A2(net292));
 sg13g2_a221oi_1 _11230_ (.B2(_03680_),
    .C1(net421),
    .B1(net115),
    .A1(net634),
    .Y(_03681_),
    .A2(_01692_));
 sg13g2_o21ai_1 _11231_ (.B1(net467),
    .Y(_03682_),
    .A1(_03677_),
    .A2(_03681_));
 sg13g2_a221oi_1 _11232_ (.B2(uo_out[3]),
    .C1(_03668_),
    .B1(_03075_),
    .A1(\i_spi.data[3] ),
    .Y(_03683_),
    .A2(_03070_));
 sg13g2_nand2_1 _11233_ (.Y(_03684_),
    .A(net5),
    .B(_03084_));
 sg13g2_a22oi_1 _11234_ (.Y(_03685_),
    .B1(net287),
    .B2(\controller2_data[3] ),
    .A2(net291),
    .A1(\controller1_data[3] ));
 sg13g2_a221oi_1 _11235_ (.B2(_03669_),
    .C1(_03670_),
    .B1(net221),
    .A1(\i_time.l_mtimecmp.data_out[3] ),
    .Y(_03686_),
    .A2(net298));
 sg13g2_and4_2 _11236_ (.A(_03683_),
    .B(_03684_),
    .C(_03685_),
    .D(_03686_),
    .X(_03687_));
 sg13g2_a221oi_1 _11237_ (.B2(_03687_),
    .C1(net421),
    .B1(net114),
    .A1(net636),
    .Y(_03688_),
    .A2(_01686_));
 sg13g2_o21ai_1 _11238_ (.B1(net419),
    .Y(_03689_),
    .A1(\i_tinyqv.cpu.instr_data_in[11] ),
    .A2(net108));
 sg13g2_a21oi_1 _11239_ (.A1(_01684_),
    .A2(net108),
    .Y(_03690_),
    .B1(_03689_));
 sg13g2_o21ai_1 _11240_ (.B1(net463),
    .Y(_03691_),
    .A1(_03688_),
    .A2(_03690_));
 sg13g2_o21ai_1 _11241_ (.B1(net460),
    .Y(_03692_),
    .A1(_03673_),
    .A2(_03675_));
 sg13g2_and4_1 _11242_ (.A(net476),
    .B(_03682_),
    .C(_03691_),
    .D(_03692_),
    .X(_03693_));
 sg13g2_mux4_1 _11243_ (.S0(net591),
    .A0(\i_tinyqv.cpu.instr_data_in[11] ),
    .A1(\i_tinyqv.cpu.instr_data_in[15] ),
    .A2(\i_tinyqv.mem.qspi_data_buf[27] ),
    .A3(\i_tinyqv.mem.qspi_data_buf[31] ),
    .S1(net117),
    .X(_03694_));
 sg13g2_nor2_1 _11244_ (.A(net416),
    .B(_03694_),
    .Y(_03695_));
 sg13g2_mux4_1 _11245_ (.S0(net472),
    .A0(\i_time.mtime[31] ),
    .A1(\i_time.mtime[27] ),
    .A2(\i_time.l_mtimecmp.data_out[31] ),
    .A3(\i_time.l_mtimecmp.data_out[27] ),
    .S1(net301),
    .X(_03696_));
 sg13g2_o21ai_1 _11246_ (.B1(net634),
    .Y(_03697_),
    .A1(net592),
    .A2(_01694_));
 sg13g2_a21oi_1 _11247_ (.A1(net590),
    .A2(\i_latch_mem.data_out[31] ),
    .Y(_03698_),
    .B1(_03697_));
 sg13g2_a21oi_1 _11248_ (.A1(net183),
    .A2(_03696_),
    .Y(_03699_),
    .B1(net116));
 sg13g2_nor4_1 _11249_ (.A(_01581_),
    .B(_03695_),
    .C(_03698_),
    .D(_03699_),
    .Y(_03700_));
 sg13g2_nor2_1 _11250_ (.A(\i_tinyqv.mem.data_from_read[19] ),
    .B(net416),
    .Y(_03701_));
 sg13g2_nor2b_1 _11251_ (.A(\i_latch_mem.data_out[19] ),
    .B_N(net634),
    .Y(_03702_));
 sg13g2_nor2_1 _11252_ (.A(\i_tinyqv.mem.data_from_read[23] ),
    .B(net415),
    .Y(_03703_));
 sg13g2_nor2b_1 _11253_ (.A(\i_latch_mem.data_out[23] ),
    .B_N(net634),
    .Y(_03704_));
 sg13g2_mux2_1 _11254_ (.A0(\i_time.mtime[19] ),
    .A1(\i_time.l_mtimecmp.data_out[19] ),
    .S(net300),
    .X(_03705_));
 sg13g2_a21oi_1 _11255_ (.A1(net183),
    .A2(_03705_),
    .Y(_03706_),
    .B1(_03116_));
 sg13g2_nor4_1 _11256_ (.A(_02169_),
    .B(_03701_),
    .C(_03702_),
    .D(_03706_),
    .Y(_03707_));
 sg13g2_a21oi_1 _11257_ (.A1(\i_time.mtime[23] ),
    .A2(net220),
    .Y(_03708_),
    .B1(net301));
 sg13g2_a21oi_1 _11258_ (.A1(_01628_),
    .A2(net301),
    .Y(_03709_),
    .B1(_03708_));
 sg13g2_nor2_1 _11259_ (.A(_03116_),
    .B(_03709_),
    .Y(_03710_));
 sg13g2_nor4_1 _11260_ (.A(_02164_),
    .B(_03703_),
    .C(_03704_),
    .D(_03710_),
    .Y(_03711_));
 sg13g2_nor3_1 _11261_ (.A(_03700_),
    .B(_03707_),
    .C(_03711_),
    .Y(_03712_));
 sg13g2_a22oi_1 _11262_ (.Y(_03713_),
    .B1(_03712_),
    .B2(net583),
    .A2(_03693_),
    .A1(_03667_));
 sg13g2_a21oi_2 _11263_ (.B1(_03064_),
    .Y(_03714_),
    .A2(_03713_),
    .A1(_03062_));
 sg13g2_nor2_1 _11264_ (.A(_02343_),
    .B(_02519_),
    .Y(_03715_));
 sg13g2_xnor2_1 _11265_ (.Y(_03716_),
    .A(_00202_),
    .B(_03365_));
 sg13g2_xnor2_1 _11266_ (.Y(_03717_),
    .A(_00207_),
    .B(_03003_));
 sg13g2_a21oi_1 _11267_ (.A1(net593),
    .A2(_03716_),
    .Y(_03718_),
    .B1(_03007_));
 sg13g2_o21ai_1 _11268_ (.B1(_03718_),
    .Y(_03719_),
    .A1(net593),
    .A2(_03717_));
 sg13g2_xnor2_1 _11269_ (.Y(_03720_),
    .A(_01514_),
    .B(_03000_));
 sg13g2_xnor2_1 _11270_ (.Y(_03721_),
    .A(_01518_),
    .B(_02995_));
 sg13g2_inv_1 _11271_ (.Y(_03722_),
    .A(_03721_));
 sg13g2_xor2_1 _11272_ (.B(_02992_),
    .A(\i_tinyqv.cpu.instr_data_start[3] ),
    .X(_03723_));
 sg13g2_o21ai_1 _11273_ (.B1(net474),
    .Y(_03724_),
    .A1(_02169_),
    .A2(_03723_));
 sg13g2_xnor2_1 _11274_ (.Y(_03725_),
    .A(_00239_),
    .B(_02998_));
 sg13g2_a221oi_1 _11275_ (.B2(net468),
    .C1(_03724_),
    .B1(_03722_),
    .A1(net458),
    .Y(_03726_),
    .A2(_03720_));
 sg13g2_o21ai_1 _11276_ (.B1(_03726_),
    .Y(_03727_),
    .A1(_02166_),
    .A2(_03725_));
 sg13g2_a21oi_1 _11277_ (.A1(_03719_),
    .A2(_03727_),
    .Y(_03728_),
    .B1(_02518_));
 sg13g2_nand2_1 _11278_ (.Y(_03729_),
    .A(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .B(_03387_));
 sg13g2_nor2_1 _11279_ (.A(_00166_),
    .B(_02250_),
    .Y(_03730_));
 sg13g2_a22oi_1 _11280_ (.Y(_03731_),
    .B1(_03730_),
    .B2(_03045_),
    .A2(_03098_),
    .A1(_03046_));
 sg13g2_nand2_1 _11281_ (.Y(_03732_),
    .A(\i_tinyqv.cpu.i_core.mepc[3] ),
    .B(_03029_));
 sg13g2_a22oi_1 _11282_ (.Y(_03733_),
    .B1(net407),
    .B2(\i_tinyqv.cpu.i_core.mcause[5] ),
    .A2(net316),
    .A1(\i_tinyqv.cpu.i_core.mcause[3] ));
 sg13g2_nand2b_1 _11283_ (.Y(_03734_),
    .B(_03040_),
    .A_N(_03733_));
 sg13g2_nand2_1 _11284_ (.Y(_03735_),
    .A(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .B(net313));
 sg13g2_o21ai_1 _11285_ (.B1(_03735_),
    .Y(_03736_),
    .A1(_01578_),
    .A2(net313));
 sg13g2_a22oi_1 _11286_ (.Y(_03737_),
    .B1(_03046_),
    .B2(\i_time.timer_interrupt ),
    .A2(_03045_),
    .A1(\i_tinyqv.cpu.i_core.mie[4] ));
 sg13g2_nand2_1 _11287_ (.Y(_03738_),
    .A(_03729_),
    .B(_03737_));
 sg13g2_nand2_1 _11288_ (.Y(_03739_),
    .A(net353),
    .B(_03738_));
 sg13g2_o21ai_1 _11289_ (.B1(_03732_),
    .Y(_03740_),
    .A1(_03042_),
    .A2(_03731_));
 sg13g2_a221oi_1 _11290_ (.B2(_03033_),
    .C1(_03740_),
    .B1(_03736_),
    .A1(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .Y(_03741_),
    .A2(_03036_));
 sg13g2_a22oi_1 _11291_ (.Y(_03742_),
    .B1(_03388_),
    .B2(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .A2(_03039_),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.data[3] ));
 sg13g2_nand4_1 _11292_ (.B(_03739_),
    .C(_03741_),
    .A(_03734_),
    .Y(_03743_),
    .D(_03742_));
 sg13g2_a221oi_1 _11293_ (.B2(_03743_),
    .C1(_03728_),
    .B1(_03020_),
    .A1(net570),
    .Y(_03744_),
    .A2(\i_tinyqv.cpu.is_lui ));
 sg13g2_o21ai_1 _11294_ (.B1(_02987_),
    .Y(_03745_),
    .A1(_03715_),
    .A2(_03744_));
 sg13g2_nand2b_1 _11295_ (.Y(_03746_),
    .B(_03745_),
    .A_N(_02826_));
 sg13g2_o21ai_1 _11296_ (.B1(_02837_),
    .Y(_03747_),
    .A1(_01595_),
    .A2(_02489_));
 sg13g2_o21ai_1 _11297_ (.B1(_02836_),
    .Y(_03748_),
    .A1(_02318_),
    .A2(_02345_));
 sg13g2_a22oi_1 _11298_ (.Y(_03749_),
    .B1(_03747_),
    .B2(_03748_),
    .A2(_02345_),
    .A1(_02318_));
 sg13g2_nor2_1 _11299_ (.A(_02350_),
    .B(_02400_),
    .Y(_03750_));
 sg13g2_a221oi_1 _11300_ (.B2(_03750_),
    .C1(_02833_),
    .B1(_03351_),
    .A1(_02350_),
    .Y(_03751_),
    .A2(\i_tinyqv.cpu.i_core.cy_out ));
 sg13g2_or2_1 _11301_ (.X(_03752_),
    .B(_03751_),
    .A(_03749_));
 sg13g2_nand2b_1 _11302_ (.Y(_03753_),
    .B(_02576_),
    .A_N(_02564_));
 sg13g2_nor2_1 _11303_ (.A(_02577_),
    .B(net406),
    .Y(_03754_));
 sg13g2_a221oi_1 _11304_ (.B2(_03754_),
    .C1(_02841_),
    .B1(_03753_),
    .A1(net406),
    .Y(_03755_),
    .A2(_03752_));
 sg13g2_a21oi_1 _11305_ (.A1(net572),
    .A2(_02971_),
    .Y(_03756_),
    .B1(_02842_));
 sg13g2_o21ai_1 _11306_ (.B1(_03756_),
    .Y(_03757_),
    .A1(net572),
    .A2(_02926_));
 sg13g2_nand3b_1 _11307_ (.B(_03757_),
    .C(_03185_),
    .Y(_03758_),
    .A_N(_03755_));
 sg13g2_o21ai_1 _11308_ (.B1(_03758_),
    .Y(_03759_),
    .A1(_00209_),
    .A2(_02829_));
 sg13g2_nand2_1 _11309_ (.Y(_03760_),
    .A(_02826_),
    .B(_03759_));
 sg13g2_o21ai_1 _11310_ (.B1(_03760_),
    .Y(\debug_rd[3] ),
    .A1(_03714_),
    .A2(_03746_));
 sg13g2_mux2_1 _11311_ (.A0(net14),
    .A1(net3310),
    .S(_03181_),
    .X(_00089_));
 sg13g2_nor2b_1 _11312_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .Y(_03761_));
 sg13g2_and2_1 _11313_ (.A(_03178_),
    .B(_03761_),
    .X(_03762_));
 sg13g2_nand3_1 _11314_ (.B(net660),
    .C(_03762_),
    .A(net661),
    .Y(_03763_));
 sg13g2_mux2_1 _11315_ (.A0(net84),
    .A1(net3881),
    .S(_03763_),
    .X(_00082_));
 sg13g2_mux2_1 _11316_ (.A0(net75),
    .A1(net3982),
    .S(_03763_),
    .X(_00083_));
 sg13g2_mux2_1 _11317_ (.A0(net82),
    .A1(net3922),
    .S(_03763_),
    .X(_00084_));
 sg13g2_mux2_1 _11318_ (.A0(net15),
    .A1(net4046),
    .S(_03763_),
    .X(_00085_));
 sg13g2_nor2b_1 _11319_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .Y(_03764_));
 sg13g2_and2_1 _11320_ (.A(_03178_),
    .B(_03764_),
    .X(_03765_));
 sg13g2_nand3_1 _11321_ (.B(net660),
    .C(_03765_),
    .A(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .Y(_03766_));
 sg13g2_mux2_1 _11322_ (.A0(net84),
    .A1(net3910),
    .S(_03766_),
    .X(_00078_));
 sg13g2_mux2_1 _11323_ (.A0(net75),
    .A1(net3858),
    .S(_03766_),
    .X(_00079_));
 sg13g2_mux2_1 _11324_ (.A0(net82),
    .A1(net3818),
    .S(_03766_),
    .X(_00080_));
 sg13g2_mux2_1 _11325_ (.A0(net14),
    .A1(net3869),
    .S(_03766_),
    .X(_00081_));
 sg13g2_nor2_2 _11326_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .Y(_03767_));
 sg13g2_nand4_1 _11327_ (.B(net660),
    .C(_03178_),
    .A(net661),
    .Y(_03768_),
    .D(_03767_));
 sg13g2_mux2_1 _11328_ (.A0(net83),
    .A1(net3822),
    .S(_03768_),
    .X(_00074_));
 sg13g2_mux2_1 _11329_ (.A0(net74),
    .A1(net3899),
    .S(_03768_),
    .X(_00075_));
 sg13g2_mux2_1 _11330_ (.A0(net81),
    .A1(net3879),
    .S(_03768_),
    .X(_00076_));
 sg13g2_mux2_1 _11331_ (.A0(net14),
    .A1(net3870),
    .S(_03768_),
    .X(_00077_));
 sg13g2_nand2_1 _11332_ (.Y(_03769_),
    .A(net660),
    .B(_03178_));
 sg13g2_nor2_2 _11333_ (.A(net661),
    .B(_03769_),
    .Y(_03770_));
 sg13g2_nand2_2 _11334_ (.Y(_03771_),
    .A(_03179_),
    .B(_03770_));
 sg13g2_mux2_1 _11335_ (.A0(net83),
    .A1(net3825),
    .S(_03771_),
    .X(_00070_));
 sg13g2_mux2_1 _11336_ (.A0(net74),
    .A1(net3767),
    .S(_03771_),
    .X(_00071_));
 sg13g2_mux2_1 _11337_ (.A0(net81),
    .A1(net3784),
    .S(_03771_),
    .X(_00072_));
 sg13g2_mux2_1 _11338_ (.A0(net14),
    .A1(net3603),
    .S(_03771_),
    .X(_00073_));
 sg13g2_nand2_2 _11339_ (.Y(_03772_),
    .A(_03761_),
    .B(_03770_));
 sg13g2_mux2_1 _11340_ (.A0(net83),
    .A1(net4005),
    .S(_03772_),
    .X(_00066_));
 sg13g2_mux2_1 _11341_ (.A0(net74),
    .A1(net3966),
    .S(_03772_),
    .X(_00067_));
 sg13g2_mux2_1 _11342_ (.A0(net81),
    .A1(net4007),
    .S(_03772_),
    .X(_00068_));
 sg13g2_mux2_1 _11343_ (.A0(net14),
    .A1(net3896),
    .S(_03772_),
    .X(_00069_));
 sg13g2_nand2_2 _11344_ (.Y(_03773_),
    .A(_03764_),
    .B(_03770_));
 sg13g2_mux2_1 _11345_ (.A0(net83),
    .A1(net4016),
    .S(_03773_),
    .X(_00114_));
 sg13g2_mux2_1 _11346_ (.A0(net74),
    .A1(net4041),
    .S(_03773_),
    .X(_00115_));
 sg13g2_mux2_1 _11347_ (.A0(net81),
    .A1(net4059),
    .S(_03773_),
    .X(_00116_));
 sg13g2_mux2_1 _11348_ (.A0(net14),
    .A1(net4090),
    .S(_03773_),
    .X(_00117_));
 sg13g2_nand2_2 _11349_ (.Y(_03774_),
    .A(_03767_),
    .B(_03770_));
 sg13g2_mux2_1 _11350_ (.A0(net84),
    .A1(net3950),
    .S(_03774_),
    .X(_00110_));
 sg13g2_mux2_1 _11351_ (.A0(net75),
    .A1(net3942),
    .S(_03774_),
    .X(_00111_));
 sg13g2_mux2_1 _11352_ (.A0(net82),
    .A1(net3980),
    .S(_03774_),
    .X(_00112_));
 sg13g2_mux2_1 _11353_ (.A0(net15),
    .A1(net4032),
    .S(_03774_),
    .X(_00113_));
 sg13g2_nor2_1 _11354_ (.A(net660),
    .B(_03180_),
    .Y(_03775_));
 sg13g2_nand2_2 _11355_ (.Y(_03776_),
    .A(_03178_),
    .B(_03775_));
 sg13g2_mux2_1 _11356_ (.A0(net84),
    .A1(net3934),
    .S(_03776_),
    .X(_00106_));
 sg13g2_mux2_1 _11357_ (.A0(net75),
    .A1(net3996),
    .S(_03776_),
    .X(_00107_));
 sg13g2_mux2_1 _11358_ (.A0(net82),
    .A1(net4093),
    .S(_03776_),
    .X(_00108_));
 sg13g2_mux2_1 _11359_ (.A0(net15),
    .A1(net4104),
    .S(_03776_),
    .X(_00109_));
 sg13g2_nor2b_1 _11360_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .B_N(net661),
    .Y(_03777_));
 sg13g2_nand2_2 _11361_ (.Y(_03778_),
    .A(_03762_),
    .B(_03777_));
 sg13g2_mux2_1 _11362_ (.A0(net83),
    .A1(net3874),
    .S(_03778_),
    .X(_00102_));
 sg13g2_mux2_1 _11363_ (.A0(net74),
    .A1(net3888),
    .S(_03778_),
    .X(_00103_));
 sg13g2_mux2_1 _11364_ (.A0(net81),
    .A1(net3902),
    .S(_03778_),
    .X(_00104_));
 sg13g2_mux2_1 _11365_ (.A0(net14),
    .A1(net3905),
    .S(_03778_),
    .X(_00105_));
 sg13g2_nand2_2 _11366_ (.Y(_03779_),
    .A(_03765_),
    .B(_03777_));
 sg13g2_mux2_1 _11367_ (.A0(net83),
    .A1(net4021),
    .S(_03779_),
    .X(_00098_));
 sg13g2_mux2_1 _11368_ (.A0(net74),
    .A1(net4092),
    .S(_03779_),
    .X(_00099_));
 sg13g2_mux2_1 _11369_ (.A0(net81),
    .A1(net4039),
    .S(_03779_),
    .X(_00100_));
 sg13g2_mux2_1 _11370_ (.A0(net14),
    .A1(net4073),
    .S(_03779_),
    .X(_00101_));
 sg13g2_nor2_1 _11371_ (.A(net661),
    .B(net660),
    .Y(_03780_));
 sg13g2_nand2_2 _11372_ (.Y(_03781_),
    .A(_03762_),
    .B(_03780_));
 sg13g2_mux2_1 _11373_ (.A0(net84),
    .A1(net3994),
    .S(_03781_),
    .X(_00094_));
 sg13g2_mux2_1 _11374_ (.A0(net75),
    .A1(net4113),
    .S(_03781_),
    .X(_00095_));
 sg13g2_mux2_1 _11375_ (.A0(net82),
    .A1(net4091),
    .S(_03781_),
    .X(_00096_));
 sg13g2_mux2_1 _11376_ (.A0(net15),
    .A1(net4081),
    .S(_03781_),
    .X(_00097_));
 sg13g2_nand2_2 _11377_ (.Y(_03782_),
    .A(_03765_),
    .B(_03780_));
 sg13g2_mux2_1 _11378_ (.A0(net83),
    .A1(net3777),
    .S(_03782_),
    .X(_00090_));
 sg13g2_mux2_1 _11379_ (.A0(net74),
    .A1(net3649),
    .S(_03782_),
    .X(_00091_));
 sg13g2_mux2_1 _11380_ (.A0(net81),
    .A1(net3772),
    .S(_03782_),
    .X(_00092_));
 sg13g2_mux2_1 _11381_ (.A0(net15),
    .A1(net3849),
    .S(_03782_),
    .X(_00093_));
 sg13g2_nand2_2 _11382_ (.Y(_03783_),
    .A(net615),
    .B(net616));
 sg13g2_nor2_2 _11383_ (.A(net4054),
    .B(_03783_),
    .Y(_03784_));
 sg13g2_nand2b_2 _11384_ (.Y(_03785_),
    .B(_01521_),
    .A_N(_03783_));
 sg13g2_a21oi_1 _11385_ (.A1(net618),
    .A2(_01662_),
    .Y(_03786_),
    .B1(_03785_));
 sg13g2_nand2_1 _11386_ (.Y(_03787_),
    .A(net616),
    .B(_03622_));
 sg13g2_nor2_2 _11387_ (.A(_01521_),
    .B(net616),
    .Y(_03788_));
 sg13g2_a21oi_1 _11388_ (.A1(_01520_),
    .A2(_03788_),
    .Y(_03789_),
    .B1(_03784_));
 sg13g2_nand2_1 _11389_ (.Y(_03790_),
    .A(_03787_),
    .B(_03789_));
 sg13g2_inv_1 _11390_ (.Y(_03791_),
    .A(_03790_));
 sg13g2_nor2_1 _11391_ (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .B(_03787_),
    .Y(_03792_));
 sg13g2_nand2_1 _11392_ (.Y(_03793_),
    .A(net515),
    .B(_03792_));
 sg13g2_and2_1 _11393_ (.A(_00193_),
    .B(_03788_),
    .X(_03794_));
 sg13g2_nand2_2 _11394_ (.Y(_03795_),
    .A(_00193_),
    .B(_03788_));
 sg13g2_a21oi_1 _11395_ (.A1(\i_tinyqv.mem.q_ctrl.addr[20] ),
    .A2(_03794_),
    .Y(_03796_),
    .B1(_03786_));
 sg13g2_a21oi_2 _11396_ (.B1(_03791_),
    .Y(uio_out[1]),
    .A2(_03796_),
    .A1(_03793_));
 sg13g2_o21ai_1 _11397_ (.B1(_03784_),
    .Y(_03797_),
    .A1(_01522_),
    .A2(\i_tinyqv.cpu.instr_data_in[13] ));
 sg13g2_a21oi_1 _11398_ (.A1(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .A2(_03794_),
    .Y(_03798_),
    .B1(_03792_));
 sg13g2_nand3_1 _11399_ (.B(_03797_),
    .C(_03798_),
    .A(_03790_),
    .Y(uio_out[2]));
 sg13g2_o21ai_1 _11400_ (.B1(_03784_),
    .Y(_03799_),
    .A1(net515),
    .A2(\i_tinyqv.cpu.instr_data_in[14] ));
 sg13g2_nand3_1 _11401_ (.B(_03790_),
    .C(_03794_),
    .A(\i_tinyqv.mem.q_ctrl.addr[22] ),
    .Y(_03800_));
 sg13g2_nand2_2 _11402_ (.Y(uio_out[4]),
    .A(_03799_),
    .B(_03800_));
 sg13g2_nand2_1 _11403_ (.Y(_03801_),
    .A(net618),
    .B(_01687_));
 sg13g2_a22oi_1 _11404_ (.Y(_03802_),
    .B1(_03801_),
    .B2(_03784_),
    .A2(_03794_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[23] ));
 sg13g2_nand3_1 _11405_ (.B(_03793_),
    .C(_03802_),
    .A(_03790_),
    .Y(uio_out[5]));
 sg13g2_nand2_1 _11406_ (.Y(_03803_),
    .A(_02076_),
    .B(net293));
 sg13g2_nand3_1 _11407_ (.B(net3241),
    .C(net182),
    .A(net528),
    .Y(_03804_));
 sg13g2_o21ai_1 _11408_ (.B1(_03804_),
    .Y(_00000_),
    .A1(_01511_),
    .A2(net182));
 sg13g2_nand3_1 _11409_ (.B(net3325),
    .C(net182),
    .A(net528),
    .Y(_03805_));
 sg13g2_o21ai_1 _11410_ (.B1(_03805_),
    .Y(_00001_),
    .A1(_01510_),
    .A2(net182));
 sg13g2_nand3_1 _11411_ (.B(net3240),
    .C(net181),
    .A(net530),
    .Y(_03806_));
 sg13g2_o21ai_1 _11412_ (.B1(_03806_),
    .Y(_00002_),
    .A1(_01509_),
    .A2(net181));
 sg13g2_nand3_1 _11413_ (.B(net3235),
    .C(net182),
    .A(net527),
    .Y(_03807_));
 sg13g2_o21ai_1 _11414_ (.B1(_03807_),
    .Y(_00003_),
    .A1(_01508_),
    .A2(net182));
 sg13g2_nand3_1 _11415_ (.B(net3213),
    .C(net181),
    .A(net525),
    .Y(_03808_));
 sg13g2_o21ai_1 _11416_ (.B1(_03808_),
    .Y(_00004_),
    .A1(_01507_),
    .A2(net181));
 sg13g2_nand3_1 _11417_ (.B(net3307),
    .C(net181),
    .A(net525),
    .Y(_03809_));
 sg13g2_o21ai_1 _11418_ (.B1(_03809_),
    .Y(_00005_),
    .A1(_01506_),
    .A2(net181));
 sg13g2_nand3_1 _11419_ (.B(net3290),
    .C(net181),
    .A(net529),
    .Y(_03810_));
 sg13g2_o21ai_1 _11420_ (.B1(_03810_),
    .Y(_00006_),
    .A1(_01505_),
    .A2(net181));
 sg13g2_nand3_1 _11421_ (.B(net3136),
    .C(net182),
    .A(net528),
    .Y(_03811_));
 sg13g2_o21ai_1 _11422_ (.B1(_03811_),
    .Y(_00007_),
    .A1(_01504_),
    .A2(net182));
 sg13g2_nand2_1 _11423_ (.Y(_03812_),
    .A(net528),
    .B(net3727));
 sg13g2_nor4_2 _11424_ (.A(_00198_),
    .B(_02077_),
    .C(_02096_),
    .Y(_03813_),
    .D(_03073_));
 sg13g2_nand2_1 _11425_ (.Y(_03814_),
    .A(\data_to_write[0] ),
    .B(net280));
 sg13g2_o21ai_1 _11426_ (.B1(_03814_),
    .Y(_00008_),
    .A1(_03812_),
    .A2(net280));
 sg13g2_nand2_1 _11427_ (.Y(_03815_),
    .A(net529),
    .B(net3556));
 sg13g2_nand2_1 _11428_ (.Y(_03816_),
    .A(net601),
    .B(net281));
 sg13g2_o21ai_1 _11429_ (.B1(_03816_),
    .Y(_00009_),
    .A1(net281),
    .A2(_03815_));
 sg13g2_nand2_1 _11430_ (.Y(_03817_),
    .A(net529),
    .B(net3698));
 sg13g2_nand2_1 _11431_ (.Y(_03818_),
    .A(net600),
    .B(net281));
 sg13g2_o21ai_1 _11432_ (.B1(_03818_),
    .Y(_00010_),
    .A1(net281),
    .A2(_03817_));
 sg13g2_nand2_1 _11433_ (.Y(_03819_),
    .A(net527),
    .B(net3549));
 sg13g2_nand2_1 _11434_ (.Y(_03820_),
    .A(\data_to_write[3] ),
    .B(net279));
 sg13g2_o21ai_1 _11435_ (.B1(_03820_),
    .Y(_00011_),
    .A1(net279),
    .A2(_03819_));
 sg13g2_nand2_1 _11436_ (.Y(_03821_),
    .A(net525),
    .B(net3742));
 sg13g2_nand2_1 _11437_ (.Y(_03822_),
    .A(net599),
    .B(net279));
 sg13g2_o21ai_1 _11438_ (.B1(_03822_),
    .Y(_00012_),
    .A1(net279),
    .A2(_03821_));
 sg13g2_nand2_1 _11439_ (.Y(_03823_),
    .A(net524),
    .B(net3577));
 sg13g2_nand2_1 _11440_ (.Y(_03824_),
    .A(net598),
    .B(net279));
 sg13g2_o21ai_1 _11441_ (.B1(_03824_),
    .Y(_00013_),
    .A1(net279),
    .A2(_03823_));
 sg13g2_nand2_1 _11442_ (.Y(_03825_),
    .A(net525),
    .B(net3566));
 sg13g2_nand2_1 _11443_ (.Y(_03826_),
    .A(net597),
    .B(net279));
 sg13g2_o21ai_1 _11444_ (.B1(_03826_),
    .Y(_00014_),
    .A1(net279),
    .A2(_03825_));
 sg13g2_nor2_1 _11445_ (.A(net521),
    .B(net2),
    .Y(_03827_));
 sg13g2_a21oi_1 _11446_ (.A1(net521),
    .A2(net3877),
    .Y(_03828_),
    .B1(_03827_));
 sg13g2_nand2_1 _11447_ (.Y(_03829_),
    .A(\data_to_write[7] ),
    .B(net281));
 sg13g2_o21ai_1 _11448_ (.B1(_03829_),
    .Y(_00015_),
    .A1(net281),
    .A2(_03828_));
 sg13g2_nand2_1 _11449_ (.Y(_03830_),
    .A(net521),
    .B(net3633));
 sg13g2_nand2_1 _11450_ (.Y(_03831_),
    .A(\data_to_write[8] ),
    .B(net281));
 sg13g2_o21ai_1 _11451_ (.B1(_03831_),
    .Y(_00016_),
    .A1(net281),
    .A2(_03830_));
 sg13g2_nand2_1 _11452_ (.Y(_03832_),
    .A(net529),
    .B(net3808));
 sg13g2_nand2_1 _11453_ (.Y(_03833_),
    .A(\data_to_write[9] ),
    .B(net280));
 sg13g2_o21ai_1 _11454_ (.B1(_03833_),
    .Y(_00017_),
    .A1(net280),
    .A2(_03832_));
 sg13g2_and2_2 _11455_ (.A(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ),
    .B(net1),
    .X(uio_oe[5]));
 sg13g2_mux2_2 _11456_ (.A0(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .A1(\i_pwm.pwm ),
    .S(\gpio_out_sel[9] ),
    .X(uio_out[7]));
 sg13g2_nand2_1 _11457_ (.Y(_03834_),
    .A(\i_tinyqv.mem.q_ctrl.spi_clk_neg ),
    .B(\i_tinyqv.mem.q_ctrl.spi_clk_use_neg ));
 sg13g2_o21ai_1 _11458_ (.B1(_03834_),
    .Y(uio_out[3]),
    .A1(_01523_),
    .A2(\i_tinyqv.mem.q_ctrl.spi_clk_use_neg ));
 sg13g2_nand2b_1 _11459_ (.Y(_03835_),
    .B(_02523_),
    .A_N(_02514_));
 sg13g2_nor2_2 _11460_ (.A(\i_tinyqv.cpu.i_core.cycle[1] ),
    .B(\i_tinyqv.cpu.i_core.cycle[0] ),
    .Y(_03836_));
 sg13g2_and3_2 _11461_ (.X(_03837_),
    .A(net407),
    .B(_03835_),
    .C(_03836_));
 sg13g2_nand3_1 _11462_ (.B(_03835_),
    .C(_03836_),
    .A(net407),
    .Y(_03838_));
 sg13g2_nand2_1 _11463_ (.Y(_03839_),
    .A(\i_tinyqv.cpu.is_load ),
    .B(_03503_));
 sg13g2_nor2_1 _11464_ (.A(net331),
    .B(_03839_),
    .Y(_03840_));
 sg13g2_nand2_1 _11465_ (.Y(_03841_),
    .A(\i_tinyqv.cpu.is_store ),
    .B(_03837_));
 sg13g2_mux2_1 _11466_ (.A0(_03501_),
    .A1(_01610_),
    .S(_03841_),
    .X(_03842_));
 sg13g2_nor3_1 _11467_ (.A(net647),
    .B(_03840_),
    .C(_03842_),
    .Y(_03843_));
 sg13g2_a21o_1 _11468_ (.A2(_03840_),
    .A1(_03502_),
    .B1(_03843_),
    .X(_00064_));
 sg13g2_nand2b_1 _11469_ (.Y(_03844_),
    .B(\i_pwm.pwm_count[2] ),
    .A_N(\i_pwm.l_pwm_level.data_out[2] ));
 sg13g2_a22oi_1 _11470_ (.Y(_03845_),
    .B1(_01618_),
    .B2(\i_pwm.l_pwm_level.data_out[1] ),
    .A2(_01599_),
    .A1(\i_pwm.l_pwm_level.data_out[0] ));
 sg13g2_o21ai_1 _11471_ (.B1(_03844_),
    .Y(_03846_),
    .A1(\i_pwm.l_pwm_level.data_out[1] ),
    .A2(_01618_));
 sg13g2_nand2b_1 _11472_ (.Y(_03847_),
    .B(\i_pwm.l_pwm_level.data_out[2] ),
    .A_N(\i_pwm.pwm_count[2] ));
 sg13g2_o21ai_1 _11473_ (.B1(_03847_),
    .Y(_03848_),
    .A1(_03845_),
    .A2(_03846_));
 sg13g2_a21oi_1 _11474_ (.A1(\i_pwm.l_pwm_level.data_out[3] ),
    .A2(_01619_),
    .Y(_03849_),
    .B1(_03848_));
 sg13g2_a221oi_1 _11475_ (.B2(_01552_),
    .C1(_03849_),
    .B1(\i_pwm.pwm_count[4] ),
    .A1(_01553_),
    .Y(_03850_),
    .A2(\i_pwm.pwm_count[3] ));
 sg13g2_nand2b_1 _11476_ (.Y(_03851_),
    .B(\i_pwm.l_pwm_level.data_out[5] ),
    .A_N(\i_pwm.pwm_count[5] ));
 sg13g2_o21ai_1 _11477_ (.B1(_03851_),
    .Y(_03852_),
    .A1(_01552_),
    .A2(\i_pwm.pwm_count[4] ));
 sg13g2_a22oi_1 _11478_ (.Y(_03853_),
    .B1(\i_pwm.pwm_count[6] ),
    .B2(_01550_),
    .A2(\i_pwm.pwm_count[5] ),
    .A1(_01551_));
 sg13g2_o21ai_1 _11479_ (.B1(_03853_),
    .Y(_03854_),
    .A1(_03850_),
    .A2(_03852_));
 sg13g2_a22oi_1 _11480_ (.Y(_03855_),
    .B1(_01621_),
    .B2(\i_pwm.l_pwm_level.data_out[7] ),
    .A2(_01620_),
    .A1(\i_pwm.l_pwm_level.data_out[6] ));
 sg13g2_a22oi_1 _11481_ (.Y(_00018_),
    .B1(_03854_),
    .B2(_03855_),
    .A2(net3892),
    .A1(_01549_));
 sg13g2_nor2_1 _11482_ (.A(net3398),
    .B(net487),
    .Y(_03856_));
 sg13g2_and2_1 _11483_ (.A(\i_latch_mem.genblk1[15].l_ram.data_out[0] ),
    .B(net242),
    .X(_03857_));
 sg13g2_a22oi_1 _11484_ (.Y(_03858_),
    .B1(net244),
    .B2(\i_latch_mem.genblk1[13].l_ram.data_out[0] ),
    .A2(net245),
    .A1(\i_latch_mem.genblk1[12].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11485_ (.Y(_03859_),
    .B1(_01923_),
    .B2(\i_latch_mem.genblk1[16].l_ram.data_out[0] ),
    .A2(net247),
    .A1(\i_latch_mem.genblk1[10].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11486_ (.Y(_03860_),
    .B1(net243),
    .B2(\i_latch_mem.genblk1[14].l_ram.data_out[0] ),
    .A2(net256),
    .A1(\i_latch_mem.genblk1[4].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11487_ (.Y(_03861_),
    .B1(net228),
    .B2(\i_latch_mem.genblk1[28].l_ram.data_out[0] ),
    .A2(net255),
    .A1(\i_latch_mem.genblk1[5].l_ram.data_out[0] ));
 sg13g2_nand3_1 _11488_ (.B(_03860_),
    .C(_03861_),
    .A(_03858_),
    .Y(_03862_));
 sg13g2_a221oi_1 _11489_ (.B2(\i_latch_mem.genblk1[7].l_ram.data_out[0] ),
    .C1(_03862_),
    .B1(net253),
    .A1(\i_latch_mem.genblk1[6].l_ram.data_out[0] ),
    .Y(_03863_),
    .A2(net254));
 sg13g2_a221oi_1 _11490_ (.B2(\i_latch_mem.genblk1[30].l_ram.data_out[0] ),
    .C1(_03857_),
    .B1(net226),
    .A1(\i_latch_mem.genblk1[22].l_ram.data_out[0] ),
    .Y(_03864_),
    .A2(net234));
 sg13g2_a22oi_1 _11491_ (.Y(_03865_),
    .B1(net235),
    .B2(\i_latch_mem.genblk1[21].l_ram.data_out[0] ),
    .A2(net258),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11492_ (.Y(_03866_),
    .B1(net233),
    .B2(\i_latch_mem.genblk1[23].l_ram.data_out[0] ),
    .A2(net259),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[0] ));
 sg13g2_nand4_1 _11493_ (.B(_03864_),
    .C(_03865_),
    .A(_03863_),
    .Y(_03867_),
    .D(_03866_));
 sg13g2_a22oi_1 _11494_ (.Y(_03868_),
    .B1(net230),
    .B2(\i_latch_mem.genblk1[26].l_ram.data_out[0] ),
    .A2(net238),
    .A1(\i_latch_mem.genblk1[18].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11495_ (.Y(_03869_),
    .B1(net225),
    .B2(\i_latch_mem.genblk1[9].l_ram.data_out[0] ),
    .A2(net246),
    .A1(\i_latch_mem.genblk1[11].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11496_ (.Y(_03870_),
    .B1(net229),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[0] ),
    .A2(net232),
    .A1(\i_latch_mem.genblk1[24].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11497_ (.Y(_03871_),
    .B1(net239),
    .B2(\i_latch_mem.genblk1[17].l_ram.data_out[0] ),
    .A2(net260),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[0] ));
 sg13g2_nand4_1 _11498_ (.B(_03869_),
    .C(_03870_),
    .A(_03868_),
    .Y(_03872_),
    .D(_03871_));
 sg13g2_a221oi_1 _11499_ (.B2(\i_latch_mem.genblk1[20].l_ram.data_out[0] ),
    .C1(net251),
    .B1(net236),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[0] ),
    .Y(_03873_),
    .A2(net252));
 sg13g2_a22oi_1 _11500_ (.Y(_03874_),
    .B1(net227),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[0] ),
    .A2(net257),
    .A1(\i_latch_mem.genblk1[3].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11501_ (.Y(_03875_),
    .B1(net231),
    .B2(\i_latch_mem.genblk1[25].l_ram.data_out[0] ),
    .A2(net237),
    .A1(\i_latch_mem.genblk1[1].l_ram.data_out[0] ));
 sg13g2_nand4_1 _11502_ (.B(_03873_),
    .C(_03874_),
    .A(_03859_),
    .Y(_03876_),
    .D(_03875_));
 sg13g2_nor3_1 _11503_ (.A(_03867_),
    .B(_03872_),
    .C(_03876_),
    .Y(_03877_));
 sg13g2_a21o_2 _11504_ (.A2(net251),
    .A1(_00256_),
    .B1(_03877_),
    .X(_03878_));
 sg13g2_a21oi_1 _11505_ (.A1(net487),
    .A2(_03878_),
    .Y(_00031_),
    .B1(_03856_));
 sg13g2_and2_1 _11506_ (.A(\i_latch_mem.genblk1[15].l_ram.data_out[1] ),
    .B(net242),
    .X(_03879_));
 sg13g2_a22oi_1 _11507_ (.Y(_03880_),
    .B1(net230),
    .B2(\i_latch_mem.genblk1[26].l_ram.data_out[1] ),
    .A2(net232),
    .A1(\i_latch_mem.genblk1[24].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11508_ (.Y(_03881_),
    .B1(net231),
    .B2(\i_latch_mem.genblk1[25].l_ram.data_out[1] ),
    .A2(net252),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11509_ (.Y(_03882_),
    .B1(net256),
    .B2(\i_latch_mem.genblk1[4].l_ram.data_out[1] ),
    .A2(net258),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11510_ (.Y(_03883_),
    .B1(net233),
    .B2(\i_latch_mem.genblk1[23].l_ram.data_out[1] ),
    .A2(net243),
    .A1(\i_latch_mem.genblk1[14].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11511_ (.Y(_03884_),
    .B1(_02063_),
    .B2(\i_latch_mem.genblk1[30].l_ram.data_out[1] ),
    .A2(net234),
    .A1(\i_latch_mem.genblk1[22].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11512_ (.Y(_03885_),
    .B1(net236),
    .B2(\i_latch_mem.genblk1[20].l_ram.data_out[1] ),
    .A2(net253),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[1] ));
 sg13g2_nand3_1 _11513_ (.B(_03884_),
    .C(_03885_),
    .A(_03883_),
    .Y(_03886_));
 sg13g2_a221oi_1 _11514_ (.B2(\i_latch_mem.genblk1[13].l_ram.data_out[1] ),
    .C1(_03886_),
    .B1(net244),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[1] ),
    .Y(_03887_),
    .A2(net259));
 sg13g2_a221oi_1 _11515_ (.B2(\i_latch_mem.genblk1[28].l_ram.data_out[1] ),
    .C1(_03879_),
    .B1(net228),
    .A1(\i_latch_mem.genblk1[12].l_ram.data_out[1] ),
    .Y(_03888_),
    .A2(net245));
 sg13g2_a22oi_1 _11516_ (.Y(_03889_),
    .B1(net254),
    .B2(\i_latch_mem.genblk1[6].l_ram.data_out[1] ),
    .A2(net255),
    .A1(\i_latch_mem.genblk1[5].l_ram.data_out[1] ));
 sg13g2_nand4_1 _11517_ (.B(_03887_),
    .C(_03888_),
    .A(_03882_),
    .Y(_03890_),
    .D(_03889_));
 sg13g2_a22oi_1 _11518_ (.Y(_03891_),
    .B1(net237),
    .B2(\i_latch_mem.genblk1[1].l_ram.data_out[1] ),
    .A2(net238),
    .A1(\i_latch_mem.genblk1[18].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11519_ (.Y(_03892_),
    .B1(net246),
    .B2(\i_latch_mem.genblk1[11].l_ram.data_out[1] ),
    .A2(net257),
    .A1(\i_latch_mem.genblk1[3].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11520_ (.Y(_03893_),
    .B1(net227),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[1] ),
    .A2(net247),
    .A1(\i_latch_mem.genblk1[10].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11521_ (.Y(_03894_),
    .B1(net225),
    .B2(\i_latch_mem.genblk1[9].l_ram.data_out[1] ),
    .A2(_01923_),
    .A1(\i_latch_mem.genblk1[16].l_ram.data_out[1] ));
 sg13g2_nand4_1 _11522_ (.B(_03892_),
    .C(_03893_),
    .A(_03891_),
    .Y(_03895_),
    .D(_03894_));
 sg13g2_a22oi_1 _11523_ (.Y(_03896_),
    .B1(net239),
    .B2(\i_latch_mem.genblk1[17].l_ram.data_out[1] ),
    .A2(net260),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[1] ));
 sg13g2_a221oi_1 _11524_ (.B2(\i_latch_mem.genblk1[27].l_ram.data_out[1] ),
    .C1(net251),
    .B1(net229),
    .A1(\i_latch_mem.genblk1[21].l_ram.data_out[1] ),
    .Y(_03897_),
    .A2(net235));
 sg13g2_nand4_1 _11525_ (.B(_03881_),
    .C(_03896_),
    .A(_03880_),
    .Y(_03898_),
    .D(_03897_));
 sg13g2_nor3_1 _11526_ (.A(_03890_),
    .B(_03895_),
    .C(_03898_),
    .Y(_03899_));
 sg13g2_a21o_1 _11527_ (.A2(net250),
    .A1(_00257_),
    .B1(_03899_),
    .X(_03900_));
 sg13g2_nor2_1 _11528_ (.A(net3371),
    .B(net488),
    .Y(_03901_));
 sg13g2_a21oi_1 _11529_ (.A1(net488),
    .A2(_03900_),
    .Y(_00042_),
    .B1(_03901_));
 sg13g2_a22oi_1 _11530_ (.Y(_03902_),
    .B1(net226),
    .B2(\i_latch_mem.genblk1[30].l_ram.data_out[2] ),
    .A2(net245),
    .A1(\i_latch_mem.genblk1[12].l_ram.data_out[2] ));
 sg13g2_and2_1 _11531_ (.A(\i_latch_mem.genblk1[5].l_ram.data_out[2] ),
    .B(net255),
    .X(_03903_));
 sg13g2_a22oi_1 _11532_ (.Y(_03904_),
    .B1(net229),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[2] ),
    .A2(net231),
    .A1(\i_latch_mem.genblk1[25].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11533_ (.Y(_03905_),
    .B1(net239),
    .B2(\i_latch_mem.genblk1[17].l_ram.data_out[2] ),
    .A2(_01725_),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11534_ (.Y(_03906_),
    .B1(net225),
    .B2(\i_latch_mem.genblk1[9].l_ram.data_out[2] ),
    .A2(_01923_),
    .A1(\i_latch_mem.genblk1[16].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11535_ (.Y(_03907_),
    .B1(net254),
    .B2(\i_latch_mem.genblk1[6].l_ram.data_out[2] ),
    .A2(net258),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11536_ (.Y(_03908_),
    .B1(net233),
    .B2(\i_latch_mem.genblk1[23].l_ram.data_out[2] ),
    .A2(net234),
    .A1(\i_latch_mem.genblk1[22].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11537_ (.Y(_03909_),
    .B1(net235),
    .B2(\i_latch_mem.genblk1[21].l_ram.data_out[2] ),
    .A2(net253),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[2] ));
 sg13g2_nand3_1 _11538_ (.B(_03908_),
    .C(_03909_),
    .A(_03907_),
    .Y(_03910_));
 sg13g2_a221oi_1 _11539_ (.B2(\i_latch_mem.genblk1[28].l_ram.data_out[2] ),
    .C1(_03910_),
    .B1(net228),
    .A1(\i_latch_mem.genblk1[15].l_ram.data_out[2] ),
    .Y(_03911_),
    .A2(net242));
 sg13g2_a221oi_1 _11540_ (.B2(\i_latch_mem.genblk1[4].l_ram.data_out[2] ),
    .C1(_03903_),
    .B1(net256),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[2] ),
    .Y(_03912_),
    .A2(net259));
 sg13g2_a22oi_1 _11541_ (.Y(_03913_),
    .B1(net236),
    .B2(\i_latch_mem.genblk1[20].l_ram.data_out[2] ),
    .A2(net244),
    .A1(\i_latch_mem.genblk1[13].l_ram.data_out[2] ));
 sg13g2_nand4_1 _11542_ (.B(_03911_),
    .C(_03912_),
    .A(_03902_),
    .Y(_03914_),
    .D(_03913_));
 sg13g2_a22oi_1 _11543_ (.Y(_03915_),
    .B1(net227),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[2] ),
    .A2(net237),
    .A1(\i_latch_mem.genblk1[1].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11544_ (.Y(_03916_),
    .B1(net230),
    .B2(\i_latch_mem.genblk1[26].l_ram.data_out[2] ),
    .A2(net238),
    .A1(\i_latch_mem.genblk1[18].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11545_ (.Y(_03917_),
    .B1(net246),
    .B2(\i_latch_mem.genblk1[11].l_ram.data_out[2] ),
    .A2(net247),
    .A1(\i_latch_mem.genblk1[10].l_ram.data_out[2] ));
 sg13g2_nand4_1 _11546_ (.B(_03915_),
    .C(_03916_),
    .A(_03904_),
    .Y(_03918_),
    .D(_03917_));
 sg13g2_a221oi_1 _11547_ (.B2(\i_latch_mem.genblk1[14].l_ram.data_out[2] ),
    .C1(net251),
    .B1(net243),
    .A1(\i_latch_mem.genblk1[3].l_ram.data_out[2] ),
    .Y(_03919_),
    .A2(net257));
 sg13g2_a22oi_1 _11548_ (.Y(_03920_),
    .B1(net232),
    .B2(\i_latch_mem.genblk1[24].l_ram.data_out[2] ),
    .A2(net252),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[2] ));
 sg13g2_nand4_1 _11549_ (.B(_03906_),
    .C(_03919_),
    .A(_03905_),
    .Y(_03921_),
    .D(_03920_));
 sg13g2_nor3_1 _11550_ (.A(_03914_),
    .B(_03918_),
    .C(_03921_),
    .Y(_03922_));
 sg13g2_a21o_1 _11551_ (.A2(net250),
    .A1(_00258_),
    .B1(_03922_),
    .X(_03923_));
 sg13g2_nor2_1 _11552_ (.A(net3368),
    .B(net487),
    .Y(_03924_));
 sg13g2_a21oi_1 _11553_ (.A1(net487),
    .A2(_03923_),
    .Y(_00053_),
    .B1(_03924_));
 sg13g2_and2_1 _11554_ (.A(\i_latch_mem.genblk1[15].l_ram.data_out[3] ),
    .B(net242),
    .X(_03925_));
 sg13g2_a22oi_1 _11555_ (.Y(_03926_),
    .B1(net257),
    .B2(\i_latch_mem.genblk1[3].l_ram.data_out[3] ),
    .A2(net260),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11556_ (.Y(_03927_),
    .B1(net227),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[3] ),
    .A2(net246),
    .A1(\i_latch_mem.genblk1[11].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11557_ (.Y(_03928_),
    .B1(net231),
    .B2(\i_latch_mem.genblk1[25].l_ram.data_out[3] ),
    .A2(net237),
    .A1(\i_latch_mem.genblk1[1].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11558_ (.Y(_03929_),
    .B1(net258),
    .B2(\i_latch_mem.genblk1[31].l_ram.data_out[3] ),
    .A2(net259),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11559_ (.Y(_03930_),
    .B1(net243),
    .B2(\i_latch_mem.genblk1[14].l_ram.data_out[3] ),
    .A2(net254),
    .A1(\i_latch_mem.genblk1[6].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11560_ (.Y(_03931_),
    .B1(net226),
    .B2(\i_latch_mem.genblk1[30].l_ram.data_out[3] ),
    .A2(net235),
    .A1(\i_latch_mem.genblk1[21].l_ram.data_out[3] ));
 sg13g2_nand3_1 _11561_ (.B(_03930_),
    .C(_03931_),
    .A(_03929_),
    .Y(_03932_));
 sg13g2_a221oi_1 _11562_ (.B2(\i_latch_mem.genblk1[23].l_ram.data_out[3] ),
    .C1(_03932_),
    .B1(net233),
    .A1(\i_latch_mem.genblk1[22].l_ram.data_out[3] ),
    .Y(_03933_),
    .A2(net234));
 sg13g2_a221oi_1 _11563_ (.B2(\i_latch_mem.genblk1[20].l_ram.data_out[3] ),
    .C1(_03925_),
    .B1(net236),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[3] ),
    .Y(_03934_),
    .A2(_01831_));
 sg13g2_a22oi_1 _11564_ (.Y(_03935_),
    .B1(net244),
    .B2(\i_latch_mem.genblk1[13].l_ram.data_out[3] ),
    .A2(net255),
    .A1(\i_latch_mem.genblk1[5].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11565_ (.Y(_03936_),
    .B1(net228),
    .B2(\i_latch_mem.genblk1[28].l_ram.data_out[3] ),
    .A2(net245),
    .A1(\i_latch_mem.genblk1[12].l_ram.data_out[3] ));
 sg13g2_nand4_1 _11566_ (.B(_03934_),
    .C(_03935_),
    .A(_03933_),
    .Y(_03937_),
    .D(_03936_));
 sg13g2_a22oi_1 _11567_ (.Y(_03938_),
    .B1(net229),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[3] ),
    .A2(net230),
    .A1(\i_latch_mem.genblk1[26].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11568_ (.Y(_03939_),
    .B1(net232),
    .B2(\i_latch_mem.genblk1[24].l_ram.data_out[3] ),
    .A2(net252),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11569_ (.Y(_03940_),
    .B1(net239),
    .B2(\i_latch_mem.genblk1[17].l_ram.data_out[3] ),
    .A2(net247),
    .A1(\i_latch_mem.genblk1[10].l_ram.data_out[3] ));
 sg13g2_nand4_1 _11570_ (.B(_03938_),
    .C(_03939_),
    .A(_03926_),
    .Y(_03941_),
    .D(_03940_));
 sg13g2_a221oi_1 _11571_ (.B2(\i_latch_mem.genblk1[9].l_ram.data_out[3] ),
    .C1(net251),
    .B1(net225),
    .A1(\i_latch_mem.genblk1[4].l_ram.data_out[3] ),
    .Y(_03942_),
    .A2(net256));
 sg13g2_a22oi_1 _11572_ (.Y(_03943_),
    .B1(net238),
    .B2(\i_latch_mem.genblk1[18].l_ram.data_out[3] ),
    .A2(_01923_),
    .A1(\i_latch_mem.genblk1[16].l_ram.data_out[3] ));
 sg13g2_nand4_1 _11573_ (.B(_03928_),
    .C(_03942_),
    .A(_03927_),
    .Y(_03944_),
    .D(_03943_));
 sg13g2_nor3_2 _11574_ (.A(_03937_),
    .B(_03941_),
    .C(_03944_),
    .Y(_03945_));
 sg13g2_a21o_1 _11575_ (.A2(net250),
    .A1(_00259_),
    .B1(_03945_),
    .X(_03946_));
 sg13g2_nor2_1 _11576_ (.A(net3224),
    .B(net487),
    .Y(_03947_));
 sg13g2_a21oi_1 _11577_ (.A1(net487),
    .A2(_03946_),
    .Y(_00056_),
    .B1(_03947_));
 sg13g2_a22oi_1 _11578_ (.Y(_03948_),
    .B1(net234),
    .B2(\i_latch_mem.genblk1[22].l_ram.data_out[4] ),
    .A2(net244),
    .A1(\i_latch_mem.genblk1[13].l_ram.data_out[4] ));
 sg13g2_and2_1 _11579_ (.A(\i_latch_mem.genblk1[5].l_ram.data_out[4] ),
    .B(net255),
    .X(_03949_));
 sg13g2_a22oi_1 _11580_ (.Y(_03950_),
    .B1(net225),
    .B2(\i_latch_mem.genblk1[9].l_ram.data_out[4] ),
    .A2(_02053_),
    .A1(\i_latch_mem.genblk1[2].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11581_ (.Y(_03951_),
    .B1(net238),
    .B2(\i_latch_mem.genblk1[18].l_ram.data_out[4] ),
    .A2(net247),
    .A1(\i_latch_mem.genblk1[10].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11582_ (.Y(_03952_),
    .B1(net245),
    .B2(\i_latch_mem.genblk1[12].l_ram.data_out[4] ),
    .A2(net256),
    .A1(\i_latch_mem.genblk1[4].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11583_ (.Y(_03953_),
    .B1(net233),
    .B2(\i_latch_mem.genblk1[23].l_ram.data_out[4] ),
    .A2(net243),
    .A1(\i_latch_mem.genblk1[14].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11584_ (.Y(_03954_),
    .B1(net226),
    .B2(\i_latch_mem.genblk1[30].l_ram.data_out[4] ),
    .A2(net236),
    .A1(\i_latch_mem.genblk1[20].l_ram.data_out[4] ));
 sg13g2_nand3_1 _11585_ (.B(_03953_),
    .C(_03954_),
    .A(_03952_),
    .Y(_03955_));
 sg13g2_a221oi_1 _11586_ (.B2(\i_latch_mem.genblk1[28].l_ram.data_out[4] ),
    .C1(_03955_),
    .B1(net228),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[4] ),
    .Y(_03956_),
    .A2(net258));
 sg13g2_a221oi_1 _11587_ (.B2(\i_latch_mem.genblk1[21].l_ram.data_out[4] ),
    .C1(_03949_),
    .B1(net235),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[4] ),
    .Y(_03957_),
    .A2(net253));
 sg13g2_a22oi_1 _11588_ (.Y(_03958_),
    .B1(net242),
    .B2(\i_latch_mem.genblk1[15].l_ram.data_out[4] ),
    .A2(net254),
    .A1(\i_latch_mem.genblk1[6].l_ram.data_out[4] ));
 sg13g2_nand4_1 _11589_ (.B(_03956_),
    .C(_03957_),
    .A(_03948_),
    .Y(_03959_),
    .D(_03958_));
 sg13g2_a22oi_1 _11590_ (.Y(_03960_),
    .B1(net230),
    .B2(\i_latch_mem.genblk1[26].l_ram.data_out[4] ),
    .A2(net252),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11591_ (.Y(_03961_),
    .B1(net231),
    .B2(\i_latch_mem.genblk1[25].l_ram.data_out[4] ),
    .A2(net260),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11592_ (.Y(_03962_),
    .B1(net246),
    .B2(\i_latch_mem.genblk1[11].l_ram.data_out[4] ),
    .A2(net257),
    .A1(\i_latch_mem.genblk1[3].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11593_ (.Y(_03963_),
    .B1(net232),
    .B2(\i_latch_mem.genblk1[24].l_ram.data_out[4] ),
    .A2(net239),
    .A1(\i_latch_mem.genblk1[17].l_ram.data_out[4] ));
 sg13g2_nand4_1 _11594_ (.B(_03961_),
    .C(_03962_),
    .A(_03960_),
    .Y(_03964_),
    .D(_03963_));
 sg13g2_a22oi_1 _11595_ (.Y(_03965_),
    .B1(_02033_),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[4] ),
    .A2(_01953_),
    .A1(\i_latch_mem.genblk1[1].l_ram.data_out[4] ));
 sg13g2_a221oi_1 _11596_ (.B2(\i_latch_mem.genblk1[16].l_ram.data_out[4] ),
    .C1(net250),
    .B1(_01923_),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[4] ),
    .Y(_03966_),
    .A2(net259));
 sg13g2_nand4_1 _11597_ (.B(_03951_),
    .C(_03965_),
    .A(_03950_),
    .Y(_03967_),
    .D(_03966_));
 sg13g2_nor3_1 _11598_ (.A(_03959_),
    .B(_03964_),
    .C(_03967_),
    .Y(_03968_));
 sg13g2_a21o_1 _11599_ (.A2(net250),
    .A1(_00260_),
    .B1(_03968_),
    .X(_03969_));
 sg13g2_nor2_1 _11600_ (.A(net3342),
    .B(net488),
    .Y(_03970_));
 sg13g2_a21oi_1 _11601_ (.A1(net488),
    .A2(_03969_),
    .Y(_00057_),
    .B1(_03970_));
 sg13g2_and2_1 _11602_ (.A(\i_latch_mem.genblk1[13].l_ram.data_out[5] ),
    .B(net244),
    .X(_03971_));
 sg13g2_a22oi_1 _11603_ (.Y(_03972_),
    .B1(net239),
    .B2(\i_latch_mem.genblk1[17].l_ram.data_out[5] ),
    .A2(net260),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11604_ (.Y(_03973_),
    .B1(net225),
    .B2(\i_latch_mem.genblk1[9].l_ram.data_out[5] ),
    .A2(net247),
    .A1(\i_latch_mem.genblk1[10].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11605_ (.Y(_03974_),
    .B1(net228),
    .B2(\i_latch_mem.genblk1[28].l_ram.data_out[5] ),
    .A2(_01993_),
    .A1(\i_latch_mem.genblk1[23].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11606_ (.Y(_03975_),
    .B1(net226),
    .B2(\i_latch_mem.genblk1[30].l_ram.data_out[5] ),
    .A2(_01913_),
    .A1(\i_latch_mem.genblk1[15].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11607_ (.Y(_03976_),
    .B1(_01983_),
    .B2(\i_latch_mem.genblk1[22].l_ram.data_out[5] ),
    .A2(_01777_),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[5] ));
 sg13g2_nand3_1 _11608_ (.B(_03975_),
    .C(_03976_),
    .A(_03974_),
    .Y(_03977_));
 sg13g2_a221oi_1 _11609_ (.B2(\i_latch_mem.genblk1[21].l_ram.data_out[5] ),
    .C1(_03977_),
    .B1(net235),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[5] ),
    .Y(_03978_),
    .A2(net259));
 sg13g2_a221oi_1 _11610_ (.B2(\i_latch_mem.genblk1[20].l_ram.data_out[5] ),
    .C1(_03971_),
    .B1(net236),
    .A1(\i_latch_mem.genblk1[14].l_ram.data_out[5] ),
    .Y(_03979_),
    .A2(net243));
 sg13g2_a22oi_1 _11611_ (.Y(_03980_),
    .B1(net254),
    .B2(\i_latch_mem.genblk1[6].l_ram.data_out[5] ),
    .A2(net256),
    .A1(\i_latch_mem.genblk1[4].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11612_ (.Y(_03981_),
    .B1(net245),
    .B2(\i_latch_mem.genblk1[12].l_ram.data_out[5] ),
    .A2(net253),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[5] ));
 sg13g2_nand4_1 _11613_ (.B(_03979_),
    .C(_03980_),
    .A(_03978_),
    .Y(_03982_),
    .D(_03981_));
 sg13g2_a22oi_1 _11614_ (.Y(_03983_),
    .B1(net227),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[5] ),
    .A2(_01873_),
    .A1(\i_latch_mem.genblk1[11].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11615_ (.Y(_03984_),
    .B1(net229),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[5] ),
    .A2(net257),
    .A1(\i_latch_mem.genblk1[3].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11616_ (.Y(_03985_),
    .B1(net237),
    .B2(\i_latch_mem.genblk1[1].l_ram.data_out[5] ),
    .A2(_01923_),
    .A1(\i_latch_mem.genblk1[16].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11617_ (.Y(_03986_),
    .B1(net231),
    .B2(\i_latch_mem.genblk1[25].l_ram.data_out[5] ),
    .A2(net252),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[5] ));
 sg13g2_nand4_1 _11618_ (.B(_03984_),
    .C(_03985_),
    .A(_03983_),
    .Y(_03987_),
    .D(_03986_));
 sg13g2_a221oi_1 _11619_ (.B2(\i_latch_mem.genblk1[24].l_ram.data_out[5] ),
    .C1(net251),
    .B1(net232),
    .A1(\i_latch_mem.genblk1[5].l_ram.data_out[5] ),
    .Y(_03988_),
    .A2(net255));
 sg13g2_a22oi_1 _11620_ (.Y(_03989_),
    .B1(net230),
    .B2(\i_latch_mem.genblk1[26].l_ram.data_out[5] ),
    .A2(net238),
    .A1(\i_latch_mem.genblk1[18].l_ram.data_out[5] ));
 sg13g2_nand4_1 _11621_ (.B(_03973_),
    .C(_03988_),
    .A(_03972_),
    .Y(_03990_),
    .D(_03989_));
 sg13g2_nor3_2 _11622_ (.A(_03982_),
    .B(_03987_),
    .C(_03990_),
    .Y(_03991_));
 sg13g2_a21o_1 _11623_ (.A2(net250),
    .A1(_00261_),
    .B1(_03991_),
    .X(_03992_));
 sg13g2_nor2_1 _11624_ (.A(net3392),
    .B(net487),
    .Y(_03993_));
 sg13g2_a21oi_1 _11625_ (.A1(net487),
    .A2(_03992_),
    .Y(_00058_),
    .B1(_03993_));
 sg13g2_and2_1 _11626_ (.A(\i_latch_mem.genblk1[13].l_ram.data_out[6] ),
    .B(_01893_),
    .X(_03994_));
 sg13g2_a22oi_1 _11627_ (.Y(_03995_),
    .B1(net225),
    .B2(\i_latch_mem.genblk1[9].l_ram.data_out[6] ),
    .A2(_01923_),
    .A1(\i_latch_mem.genblk1[16].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11628_ (.Y(_03996_),
    .B1(net227),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[6] ),
    .A2(net252),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11629_ (.Y(_03997_),
    .B1(net231),
    .B2(\i_latch_mem.genblk1[25].l_ram.data_out[6] ),
    .A2(net246),
    .A1(\i_latch_mem.genblk1[11].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11630_ (.Y(_03998_),
    .B1(net242),
    .B2(\i_latch_mem.genblk1[15].l_ram.data_out[6] ),
    .A2(net254),
    .A1(\i_latch_mem.genblk1[6].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11631_ (.Y(_03999_),
    .B1(net245),
    .B2(\i_latch_mem.genblk1[12].l_ram.data_out[6] ),
    .A2(net253),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11632_ (.Y(_04000_),
    .B1(_02043_),
    .B2(\i_latch_mem.genblk1[28].l_ram.data_out[6] ),
    .A2(net233),
    .A1(\i_latch_mem.genblk1[23].l_ram.data_out[6] ));
 sg13g2_nand3_1 _11633_ (.B(_03999_),
    .C(_04000_),
    .A(_03998_),
    .Y(_04001_));
 sg13g2_a221oi_1 _11634_ (.B2(\i_latch_mem.genblk1[14].l_ram.data_out[6] ),
    .C1(_04001_),
    .B1(net243),
    .A1(\i_latch_mem.genblk1[4].l_ram.data_out[6] ),
    .Y(_04002_),
    .A2(net256));
 sg13g2_a221oi_1 _11635_ (.B2(\i_latch_mem.genblk1[30].l_ram.data_out[6] ),
    .C1(_03994_),
    .B1(net226),
    .A1(\i_latch_mem.genblk1[22].l_ram.data_out[6] ),
    .Y(_04003_),
    .A2(net234));
 sg13g2_a22oi_1 _11636_ (.Y(_04004_),
    .B1(_01973_),
    .B2(\i_latch_mem.genblk1[21].l_ram.data_out[6] ),
    .A2(net259),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11637_ (.Y(_04005_),
    .B1(net255),
    .B2(\i_latch_mem.genblk1[5].l_ram.data_out[6] ),
    .A2(net258),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[6] ));
 sg13g2_nand4_1 _11638_ (.B(_04003_),
    .C(_04004_),
    .A(_04002_),
    .Y(_04006_),
    .D(_04005_));
 sg13g2_a22oi_1 _11639_ (.Y(_04007_),
    .B1(net229),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[6] ),
    .A2(net238),
    .A1(\i_latch_mem.genblk1[18].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11640_ (.Y(_04008_),
    .B1(net230),
    .B2(\i_latch_mem.genblk1[26].l_ram.data_out[6] ),
    .A2(net232),
    .A1(\i_latch_mem.genblk1[24].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11641_ (.Y(_04009_),
    .B1(net239),
    .B2(\i_latch_mem.genblk1[17].l_ram.data_out[6] ),
    .A2(net260),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[6] ));
 sg13g2_nand4_1 _11642_ (.B(_04007_),
    .C(_04008_),
    .A(_03995_),
    .Y(_04010_),
    .D(_04009_));
 sg13g2_a221oi_1 _11643_ (.B2(\i_latch_mem.genblk1[20].l_ram.data_out[6] ),
    .C1(net251),
    .B1(net236),
    .A1(\i_latch_mem.genblk1[10].l_ram.data_out[6] ),
    .Y(_04011_),
    .A2(net247));
 sg13g2_a22oi_1 _11644_ (.Y(_04012_),
    .B1(net237),
    .B2(\i_latch_mem.genblk1[1].l_ram.data_out[6] ),
    .A2(net257),
    .A1(\i_latch_mem.genblk1[3].l_ram.data_out[6] ));
 sg13g2_nand4_1 _11645_ (.B(_03997_),
    .C(_04011_),
    .A(_03996_),
    .Y(_04013_),
    .D(_04012_));
 sg13g2_nor3_1 _11646_ (.A(_04006_),
    .B(_04010_),
    .C(_04013_),
    .Y(_04014_));
 sg13g2_a21o_1 _11647_ (.A2(net250),
    .A1(_00262_),
    .B1(_04014_),
    .X(_04015_));
 sg13g2_nor2_1 _11648_ (.A(net3326),
    .B(net488),
    .Y(_04016_));
 sg13g2_a21oi_1 _11649_ (.A1(net488),
    .A2(_04015_),
    .Y(_00059_),
    .B1(_04016_));
 sg13g2_nor2_1 _11650_ (.A(net3284),
    .B(net489),
    .Y(_04017_));
 sg13g2_and2_1 _11651_ (.A(\i_latch_mem.genblk1[13].l_ram.data_out[7] ),
    .B(net244),
    .X(_04018_));
 sg13g2_a22oi_1 _11652_ (.Y(_04019_),
    .B1(net227),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[7] ),
    .A2(_01933_),
    .A1(\i_latch_mem.genblk1[17].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11653_ (.Y(_04020_),
    .B1(net237),
    .B2(\i_latch_mem.genblk1[1].l_ram.data_out[7] ),
    .A2(_01943_),
    .A1(\i_latch_mem.genblk1[18].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11654_ (.Y(_04021_),
    .B1(net246),
    .B2(\i_latch_mem.genblk1[11].l_ram.data_out[7] ),
    .A2(net252),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11655_ (.Y(_04022_),
    .B1(net225),
    .B2(\i_latch_mem.genblk1[9].l_ram.data_out[7] ),
    .A2(_02003_),
    .A1(\i_latch_mem.genblk1[24].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11656_ (.Y(_04023_),
    .B1(net229),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[7] ),
    .A2(_02013_),
    .A1(\i_latch_mem.genblk1[25].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11657_ (.Y(_04024_),
    .B1(net226),
    .B2(\i_latch_mem.genblk1[30].l_ram.data_out[7] ),
    .A2(net256),
    .A1(\i_latch_mem.genblk1[4].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11658_ (.Y(_04025_),
    .B1(net254),
    .B2(\i_latch_mem.genblk1[6].l_ram.data_out[7] ),
    .A2(net255),
    .A1(\i_latch_mem.genblk1[5].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11659_ (.Y(_04026_),
    .B1(net235),
    .B2(\i_latch_mem.genblk1[21].l_ram.data_out[7] ),
    .A2(net253),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[7] ));
 sg13g2_nand3_1 _11660_ (.B(_04025_),
    .C(_04026_),
    .A(_04024_),
    .Y(_04027_));
 sg13g2_a221oi_1 _11661_ (.B2(\i_latch_mem.genblk1[22].l_ram.data_out[7] ),
    .C1(_04027_),
    .B1(net234),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[7] ),
    .Y(_04028_),
    .A2(_01767_));
 sg13g2_a221oi_1 _11662_ (.B2(\i_latch_mem.genblk1[23].l_ram.data_out[7] ),
    .C1(_04018_),
    .B1(net233),
    .A1(\i_latch_mem.genblk1[12].l_ram.data_out[7] ),
    .Y(_04029_),
    .A2(_01883_));
 sg13g2_a22oi_1 _11663_ (.Y(_04030_),
    .B1(net228),
    .B2(\i_latch_mem.genblk1[28].l_ram.data_out[7] ),
    .A2(_01903_),
    .A1(\i_latch_mem.genblk1[14].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11664_ (.Y(_04031_),
    .B1(_01963_),
    .B2(\i_latch_mem.genblk1[20].l_ram.data_out[7] ),
    .A2(net242),
    .A1(\i_latch_mem.genblk1[15].l_ram.data_out[7] ));
 sg13g2_nand4_1 _11665_ (.B(_04029_),
    .C(_04030_),
    .A(_04028_),
    .Y(_04032_),
    .D(_04031_));
 sg13g2_a221oi_1 _11666_ (.B2(\i_latch_mem.genblk1[10].l_ram.data_out[7] ),
    .C1(_01853_),
    .B1(net247),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[7] ),
    .Y(_04033_),
    .A2(net258));
 sg13g2_nand4_1 _11667_ (.B(_04021_),
    .C(_04022_),
    .A(_04020_),
    .Y(_04034_),
    .D(_04033_));
 sg13g2_a22oi_1 _11668_ (.Y(_04035_),
    .B1(net230),
    .B2(\i_latch_mem.genblk1[26].l_ram.data_out[7] ),
    .A2(net257),
    .A1(\i_latch_mem.genblk1[3].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11669_ (.Y(_04036_),
    .B1(_01923_),
    .B2(\i_latch_mem.genblk1[16].l_ram.data_out[7] ),
    .A2(net260),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[7] ));
 sg13g2_nand4_1 _11670_ (.B(_04023_),
    .C(_04035_),
    .A(_04019_),
    .Y(_04037_),
    .D(_04036_));
 sg13g2_nor3_1 _11671_ (.A(_04032_),
    .B(_04034_),
    .C(_04037_),
    .Y(_04038_));
 sg13g2_a21o_1 _11672_ (.A2(net250),
    .A1(_00263_),
    .B1(_04038_),
    .X(_04039_));
 sg13g2_a21oi_1 _11673_ (.A1(net489),
    .A2(_04039_),
    .Y(_00060_),
    .B1(_04017_));
 sg13g2_nand2_1 _11674_ (.Y(_04040_),
    .A(net3426),
    .B(net496));
 sg13g2_nor2_2 _11675_ (.A(_00242_),
    .B(net489),
    .Y(_04041_));
 sg13g2_nand2b_1 _11676_ (.Y(_04042_),
    .B(_04041_),
    .A_N(_03878_));
 sg13g2_o21ai_1 _11677_ (.B1(_04040_),
    .Y(_00061_),
    .A1(net492),
    .A2(_04042_));
 sg13g2_nand2_1 _11678_ (.Y(_04043_),
    .A(net3352),
    .B(net496));
 sg13g2_nand2b_1 _11679_ (.Y(_04044_),
    .B(_04041_),
    .A_N(_03900_));
 sg13g2_o21ai_1 _11680_ (.B1(_04043_),
    .Y(_00062_),
    .A1(net492),
    .A2(_04044_));
 sg13g2_nand2_1 _11681_ (.Y(_04045_),
    .A(net3010),
    .B(net496));
 sg13g2_nand2b_1 _11682_ (.Y(_04046_),
    .B(_04041_),
    .A_N(_03923_));
 sg13g2_o21ai_1 _11683_ (.B1(_04045_),
    .Y(_00032_),
    .A1(net491),
    .A2(_04046_));
 sg13g2_nand2_1 _11684_ (.Y(_04047_),
    .A(net3001),
    .B(net496));
 sg13g2_nand2b_1 _11685_ (.Y(_04048_),
    .B(_04041_),
    .A_N(_03946_));
 sg13g2_o21ai_1 _11686_ (.B1(_04047_),
    .Y(_00033_),
    .A1(net493),
    .A2(_04048_));
 sg13g2_nand2_1 _11687_ (.Y(_04049_),
    .A(net3142),
    .B(net496));
 sg13g2_nand2b_1 _11688_ (.Y(_04050_),
    .B(_04041_),
    .A_N(_03969_));
 sg13g2_o21ai_1 _11689_ (.B1(_04049_),
    .Y(_00034_),
    .A1(net494),
    .A2(_04050_));
 sg13g2_nand2_1 _11690_ (.Y(_04051_),
    .A(net3606),
    .B(net496));
 sg13g2_nand2b_1 _11691_ (.Y(_04052_),
    .B(_04041_),
    .A_N(_03992_));
 sg13g2_o21ai_1 _11692_ (.B1(_04051_),
    .Y(_00035_),
    .A1(net491),
    .A2(_04052_));
 sg13g2_nand2_1 _11693_ (.Y(_04053_),
    .A(net3229),
    .B(net496));
 sg13g2_nand2b_1 _11694_ (.Y(_04054_),
    .B(_04041_),
    .A_N(_04015_));
 sg13g2_o21ai_1 _11695_ (.B1(_04053_),
    .Y(_00036_),
    .A1(net494),
    .A2(_04054_));
 sg13g2_nand2_1 _11696_ (.Y(_04055_),
    .A(net3182),
    .B(net496));
 sg13g2_nand2b_1 _11697_ (.Y(_04056_),
    .B(_04041_),
    .A_N(_04039_));
 sg13g2_o21ai_1 _11698_ (.B1(_04055_),
    .Y(_00037_),
    .A1(net494),
    .A2(_04056_));
 sg13g2_nor2_1 _11699_ (.A(net3278),
    .B(net498),
    .Y(_04057_));
 sg13g2_a21oi_1 _11700_ (.A1(net498),
    .A2(_03878_),
    .Y(_00038_),
    .B1(_04057_));
 sg13g2_nor2_1 _11701_ (.A(net3222),
    .B(net497),
    .Y(_04058_));
 sg13g2_a21oi_1 _11702_ (.A1(net497),
    .A2(_03900_),
    .Y(_00039_),
    .B1(_04058_));
 sg13g2_nor2_1 _11703_ (.A(net3482),
    .B(net497),
    .Y(_04059_));
 sg13g2_a21oi_1 _11704_ (.A1(net497),
    .A2(_03923_),
    .Y(_00040_),
    .B1(_04059_));
 sg13g2_nor2_1 _11705_ (.A(net3542),
    .B(net499),
    .Y(_04060_));
 sg13g2_a21oi_1 _11706_ (.A1(net499),
    .A2(_03946_),
    .Y(_00041_),
    .B1(_04060_));
 sg13g2_nor2_1 _11707_ (.A(net3450),
    .B(net497),
    .Y(_04061_));
 sg13g2_a21oi_1 _11708_ (.A1(net497),
    .A2(_03969_),
    .Y(_00043_),
    .B1(_04061_));
 sg13g2_nor2_1 _11709_ (.A(net3522),
    .B(net497),
    .Y(_04062_));
 sg13g2_a21oi_1 _11710_ (.A1(net497),
    .A2(_03992_),
    .Y(_00044_),
    .B1(_04062_));
 sg13g2_nor2_1 _11711_ (.A(net3228),
    .B(net498),
    .Y(_04063_));
 sg13g2_a21oi_1 _11712_ (.A1(net498),
    .A2(_04015_),
    .Y(_00045_),
    .B1(_04063_));
 sg13g2_nor2_1 _11713_ (.A(net3375),
    .B(net499),
    .Y(_04064_));
 sg13g2_a21oi_1 _11714_ (.A1(net499),
    .A2(_04039_),
    .Y(_00046_),
    .B1(_04064_));
 sg13g2_nor2_1 _11715_ (.A(net3220),
    .B(net491),
    .Y(_04065_));
 sg13g2_a21oi_1 _11716_ (.A1(net491),
    .A2(_04042_),
    .Y(_00047_),
    .B1(_04065_));
 sg13g2_nor2_1 _11717_ (.A(net3238),
    .B(net492),
    .Y(_04066_));
 sg13g2_a21oi_1 _11718_ (.A1(net492),
    .A2(_04044_),
    .Y(_00048_),
    .B1(_04066_));
 sg13g2_nor2_1 _11719_ (.A(net3255),
    .B(net491),
    .Y(_04067_));
 sg13g2_a21oi_1 _11720_ (.A1(net491),
    .A2(_04046_),
    .Y(_00049_),
    .B1(_04067_));
 sg13g2_nor2_1 _11721_ (.A(net3288),
    .B(net493),
    .Y(_04068_));
 sg13g2_a21oi_1 _11722_ (.A1(net493),
    .A2(_04048_),
    .Y(_00050_),
    .B1(_04068_));
 sg13g2_nor2_1 _11723_ (.A(net3247),
    .B(net495),
    .Y(_04069_));
 sg13g2_a21oi_1 _11724_ (.A1(net494),
    .A2(_04050_),
    .Y(_00051_),
    .B1(_04069_));
 sg13g2_nor2_1 _11725_ (.A(net3268),
    .B(net491),
    .Y(_04070_));
 sg13g2_a21oi_1 _11726_ (.A1(net491),
    .A2(_04052_),
    .Y(_00052_),
    .B1(_04070_));
 sg13g2_nor2_1 _11727_ (.A(net3257),
    .B(net494),
    .Y(_04071_));
 sg13g2_a21oi_1 _11728_ (.A1(net494),
    .A2(_04054_),
    .Y(_00054_),
    .B1(_04071_));
 sg13g2_nor2_1 _11729_ (.A(net3231),
    .B(net494),
    .Y(_04072_));
 sg13g2_a21oi_1 _11730_ (.A1(net494),
    .A2(_04056_),
    .Y(_00055_),
    .B1(_04072_));
 sg13g2_nor3_1 _11731_ (.A(net3843),
    .B(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .C(net316),
    .Y(_04073_));
 sg13g2_o21ai_1 _11732_ (.B1(net4033),
    .Y(_04074_),
    .A1(net3843),
    .A2(net316));
 sg13g2_nand2_1 _11733_ (.Y(_04075_),
    .A(net653),
    .B(_04074_));
 sg13g2_nor2_1 _11734_ (.A(net3844),
    .B(_04075_),
    .Y(_00592_));
 sg13g2_nor2_2 _11735_ (.A(_01647_),
    .B(_04074_),
    .Y(_04076_));
 sg13g2_a21oi_1 _11736_ (.A1(_01647_),
    .A2(_04074_),
    .Y(_04077_),
    .B1(net510));
 sg13g2_nor2b_1 _11737_ (.A(_04076_),
    .B_N(_04077_),
    .Y(_00593_));
 sg13g2_o21ai_1 _11738_ (.B1(net653),
    .Y(_04078_),
    .A1(net3968),
    .A2(_04076_));
 sg13g2_a21oi_1 _11739_ (.A1(net3968),
    .A2(_04076_),
    .Y(_00594_),
    .B1(_04078_));
 sg13g2_a21oi_1 _11740_ (.A1(\i_tinyqv.cpu.i_core.cycle_count[2] ),
    .A2(_04076_),
    .Y(_04079_),
    .B1(net3915));
 sg13g2_nand3_1 _11741_ (.B(net3915),
    .C(_04076_),
    .A(net3968),
    .Y(_04080_));
 sg13g2_nand2_1 _11742_ (.Y(_04081_),
    .A(net653),
    .B(_04080_));
 sg13g2_nor2_1 _11743_ (.A(net3916),
    .B(_04081_),
    .Y(_00595_));
 sg13g2_nand2_1 _11744_ (.Y(_04082_),
    .A(_00264_),
    .B(net316));
 sg13g2_nand2_1 _11745_ (.Y(_04083_),
    .A(_00265_),
    .B(net334));
 sg13g2_and3_1 _11746_ (.X(_04084_),
    .A(net3644),
    .B(_04082_),
    .C(_04083_));
 sg13g2_and2_1 _11747_ (.A(net3973),
    .B(_04084_),
    .X(_04085_));
 sg13g2_nand2_1 _11748_ (.Y(_04086_),
    .A(net4028),
    .B(_04085_));
 sg13g2_nor3_1 _11749_ (.A(net509),
    .B(_01682_),
    .C(_04086_),
    .Y(_00596_));
 sg13g2_nand2_1 _11750_ (.Y(_04087_),
    .A(net353),
    .B(_03836_));
 sg13g2_nand2_1 _11751_ (.Y(_04088_),
    .A(_02273_),
    .B(_02509_));
 sg13g2_o21ai_1 _11752_ (.B1(_04088_),
    .Y(_04089_),
    .A1(_02280_),
    .A2(_02509_));
 sg13g2_mux2_1 _11753_ (.A0(_04089_),
    .A1(net3770),
    .S(_04087_),
    .X(_00597_));
 sg13g2_nor2_1 _11754_ (.A(net509),
    .B(net3969),
    .Y(_00598_));
 sg13g2_a21oi_1 _11755_ (.A1(_04082_),
    .A2(_04083_),
    .Y(_04090_),
    .B1(net3644));
 sg13g2_nor3_1 _11756_ (.A(net509),
    .B(_04084_),
    .C(net3645),
    .Y(_00599_));
 sg13g2_o21ai_1 _11757_ (.B1(net653),
    .Y(_04091_),
    .A1(net3973),
    .A2(_04084_));
 sg13g2_nor2_1 _11758_ (.A(_04085_),
    .B(_04091_),
    .Y(_00600_));
 sg13g2_o21ai_1 _11759_ (.B1(net653),
    .Y(_04092_),
    .A1(net4028),
    .A2(_04085_));
 sg13g2_nor2b_1 _11760_ (.A(_04092_),
    .B_N(_04086_),
    .Y(_00601_));
 sg13g2_xnor2_1 _11761_ (.Y(_04093_),
    .A(_01682_),
    .B(_04086_));
 sg13g2_nor2_1 _11762_ (.A(net509),
    .B(_04093_),
    .Y(_00602_));
 sg13g2_nand2_1 _11763_ (.Y(_04094_),
    .A(net3292),
    .B(net335));
 sg13g2_nand2_2 _11764_ (.Y(_04095_),
    .A(net315),
    .B(_03836_));
 sg13g2_a22oi_1 _11765_ (.Y(_00603_),
    .B1(_04094_),
    .B2(_02985_),
    .A2(_03836_),
    .A1(net315));
 sg13g2_nand2_1 _11766_ (.Y(_04096_),
    .A(net3768),
    .B(net313));
 sg13g2_nand4_1 _11767_ (.B(_02517_),
    .C(_02527_),
    .A(_02482_),
    .Y(_04097_),
    .D(_02828_));
 sg13g2_a21oi_1 _11768_ (.A1(_04096_),
    .A2(_04097_),
    .Y(_00604_),
    .B1(net511));
 sg13g2_a21oi_1 _11769_ (.A1(\i_tinyqv.cpu.i_core.cycle[0] ),
    .A2(_02482_),
    .Y(_04098_),
    .B1(net3613));
 sg13g2_nor3_1 _11770_ (.A(net511),
    .B(_02528_),
    .C(net3614),
    .Y(_00605_));
 sg13g2_nor2_1 _11771_ (.A(net335),
    .B(_03458_),
    .Y(_04099_));
 sg13g2_nor3_1 _11772_ (.A(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .B(net335),
    .C(_03458_),
    .Y(_04100_));
 sg13g2_a21o_1 _11773_ (.A2(net334),
    .A1(net3395),
    .B1(_04100_),
    .X(_00606_));
 sg13g2_nor2_2 _11774_ (.A(net313),
    .B(_04080_),
    .Y(_04101_));
 sg13g2_o21ai_1 _11775_ (.B1(net653),
    .Y(_04102_),
    .A1(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .A2(_04101_));
 sg13g2_a21oi_1 _11776_ (.A1(_01579_),
    .A2(_04101_),
    .Y(_00607_),
    .B1(_04102_));
 sg13g2_a21oi_1 _11777_ (.A1(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .A2(_04101_),
    .Y(_04103_),
    .B1(net3210));
 sg13g2_nand3_1 _11778_ (.B(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .C(_04101_),
    .A(net3210),
    .Y(_04104_));
 sg13g2_nand2_1 _11779_ (.Y(_04105_),
    .A(net653),
    .B(_04104_));
 sg13g2_nor2_1 _11780_ (.A(net3211),
    .B(_04105_),
    .Y(_00608_));
 sg13g2_o21ai_1 _11781_ (.B1(net653),
    .Y(_04106_),
    .A1(_01578_),
    .A2(_04104_));
 sg13g2_a21oi_1 _11782_ (.A1(_01578_),
    .A2(_04104_),
    .Y(_00609_),
    .B1(_04106_));
 sg13g2_nand2_1 _11783_ (.Y(_04107_),
    .A(net315),
    .B(_03460_));
 sg13g2_nor2_2 _11784_ (.A(net335),
    .B(_03459_),
    .Y(_04108_));
 sg13g2_nand2_1 _11785_ (.Y(_04109_),
    .A(_02396_),
    .B(_04108_));
 sg13g2_nor4_2 _11786_ (.A(net3576),
    .B(_02221_),
    .C(_02343_),
    .Y(_04110_),
    .D(_04109_));
 sg13g2_nand3_1 _11787_ (.B(\i_tinyqv.cpu.i_core.mie[1] ),
    .C(_03468_),
    .A(\i_tinyqv.cpu.i_core.mip[1] ),
    .Y(_04111_));
 sg13g2_a22oi_1 _11788_ (.Y(_04112_),
    .B1(_03471_),
    .B2(_03472_),
    .A2(\i_time.timer_interrupt ),
    .A1(\i_tinyqv.cpu.i_core.mie[4] ));
 sg13g2_nand2_1 _11789_ (.Y(_04113_),
    .A(_04111_),
    .B(_04112_));
 sg13g2_and2_1 _11790_ (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .B(_04108_),
    .X(_04114_));
 sg13g2_a221oi_1 _11791_ (.B2(_04114_),
    .C1(_04110_),
    .B1(_04113_),
    .A1(net3847),
    .Y(_04115_),
    .A2(net180));
 sg13g2_nor2_1 _11792_ (.A(net510),
    .B(net3848),
    .Y(_00610_));
 sg13g2_and3_1 _11793_ (.X(_04116_),
    .A(\i_tinyqv.cpu.i_core.mie[2] ),
    .B(_03287_),
    .C(_03469_));
 sg13g2_nor3_1 _11794_ (.A(_00129_),
    .B(net334),
    .C(_04116_),
    .Y(_04117_));
 sg13g2_o21ai_1 _11795_ (.B1(net655),
    .Y(_04118_),
    .A1(net3598),
    .A2(_04108_));
 sg13g2_a21oi_1 _11796_ (.A1(_04112_),
    .A2(_04117_),
    .Y(_00611_),
    .B1(net3599));
 sg13g2_nor3_1 _11797_ (.A(_00129_),
    .B(net334),
    .C(_03473_),
    .Y(_04119_));
 sg13g2_a21oi_1 _11798_ (.A1(net3520),
    .A2(net180),
    .Y(_04120_),
    .B1(_04119_));
 sg13g2_nor2_1 _11799_ (.A(net510),
    .B(net3521),
    .Y(_00612_));
 sg13g2_a22oi_1 _11800_ (.Y(_04121_),
    .B1(_04110_),
    .B2(_02280_),
    .A2(net180),
    .A1(net3297));
 sg13g2_nor2_1 _11801_ (.A(net510),
    .B(net3298),
    .Y(_00613_));
 sg13g2_a22oi_1 _11802_ (.Y(_04122_),
    .B1(_04114_),
    .B2(_03473_),
    .A2(net180),
    .A1(net3299));
 sg13g2_nor2_1 _11803_ (.A(net513),
    .B(net3300),
    .Y(_00614_));
 sg13g2_a21oi_1 _11804_ (.A1(net3384),
    .A2(_04107_),
    .Y(_04123_),
    .B1(_04114_));
 sg13g2_nor2_1 _11805_ (.A(net513),
    .B(net3385),
    .Y(_00615_));
 sg13g2_or3_2 _11806_ (.A(net648),
    .B(net3395),
    .C(_04100_),
    .X(_04124_));
 sg13g2_nand2_2 _11807_ (.Y(_04125_),
    .A(net585),
    .B(net468));
 sg13g2_nor3_2 _11808_ (.A(_00120_),
    .B(net179),
    .C(_04125_),
    .Y(_04126_));
 sg13g2_nand2_1 _11809_ (.Y(_04127_),
    .A(\i_tinyqv.cpu.i_core.interrupt_req[0] ),
    .B(_04126_));
 sg13g2_o21ai_1 _11810_ (.B1(_04127_),
    .Y(_00616_),
    .A1(_01695_),
    .A2(_04126_));
 sg13g2_mux2_1 _11811_ (.A0(net3275),
    .A1(\i_tinyqv.cpu.i_core.interrupt_req[1] ),
    .S(_04126_),
    .X(_00617_));
 sg13g2_nor2_1 _11812_ (.A(net511),
    .B(_02231_),
    .Y(_04128_));
 sg13g2_nand2_1 _11813_ (.Y(_04129_),
    .A(net659),
    .B(net455));
 sg13g2_nor2_1 _11814_ (.A(_02507_),
    .B(_02525_),
    .Y(_04130_));
 sg13g2_or4_2 _11815_ (.A(\i_tinyqv.cpu.alu_op[1] ),
    .B(_03019_),
    .C(_03026_),
    .D(_03028_),
    .X(_04131_));
 sg13g2_a21oi_1 _11816_ (.A1(_01659_),
    .A2(_04131_),
    .Y(_04132_),
    .B1(_03460_));
 sg13g2_o21ai_1 _11817_ (.B1(_04132_),
    .Y(_04133_),
    .A1(_02248_),
    .A2(_04131_));
 sg13g2_o21ai_1 _11818_ (.B1(_04133_),
    .Y(_04134_),
    .A1(_02255_),
    .A2(_03459_));
 sg13g2_a22oi_1 _11819_ (.Y(_04135_),
    .B1(_04128_),
    .B2(_04134_),
    .A2(net456),
    .A1(net3756));
 sg13g2_inv_1 _11820_ (.Y(_00618_),
    .A(_04135_));
 sg13g2_nand2b_1 _11821_ (.Y(_04136_),
    .B(_02156_),
    .A_N(_04131_));
 sg13g2_a21oi_1 _11822_ (.A1(\i_tinyqv.cpu.i_core.mepc[1] ),
    .A2(_04131_),
    .Y(_04137_),
    .B1(_03460_));
 sg13g2_a221oi_1 _11823_ (.B2(_04137_),
    .C1(_04129_),
    .B1(_04136_),
    .A1(_02176_),
    .Y(_04138_),
    .A2(_03460_));
 sg13g2_a21o_1 _11824_ (.A2(net456),
    .A1(net3871),
    .B1(_04138_),
    .X(_00619_));
 sg13g2_nand2b_1 _11825_ (.Y(_04139_),
    .B(_02365_),
    .A_N(_04131_));
 sg13g2_a21oi_1 _11826_ (.A1(\i_tinyqv.cpu.i_core.mepc[2] ),
    .A2(_04131_),
    .Y(_04140_),
    .B1(_03460_));
 sg13g2_a221oi_1 _11827_ (.B2(_04140_),
    .C1(_04129_),
    .B1(_04139_),
    .A1(_02371_),
    .Y(_04141_),
    .A2(_03460_));
 sg13g2_a21o_1 _11828_ (.A2(_02231_),
    .A1(net3615),
    .B1(_04141_),
    .X(_00620_));
 sg13g2_a21oi_1 _11829_ (.A1(_01683_),
    .A2(_04131_),
    .Y(_04142_),
    .B1(_03460_));
 sg13g2_o21ai_1 _11830_ (.B1(_04142_),
    .Y(_04143_),
    .A1(_02311_),
    .A2(_04131_));
 sg13g2_o21ai_1 _11831_ (.B1(_04143_),
    .Y(_04144_),
    .A1(_02316_),
    .A2(_03459_));
 sg13g2_a22oi_1 _11832_ (.Y(_04145_),
    .B1(_04128_),
    .B2(_04144_),
    .A2(_02231_),
    .A1(net3625));
 sg13g2_inv_1 _11833_ (.Y(_00621_),
    .A(_04145_));
 sg13g2_o21ai_1 _11834_ (.B1(net180),
    .Y(_04146_),
    .A1(net3957),
    .A2(net348));
 sg13g2_nand2b_1 _11835_ (.Y(_00622_),
    .B(_04146_),
    .A_N(net179));
 sg13g2_a21oi_1 _11836_ (.A1(_02308_),
    .A2(_02310_),
    .Y(_04147_),
    .B1(_03019_));
 sg13g2_nor2_1 _11837_ (.A(net340),
    .B(_04147_),
    .Y(_04148_));
 sg13g2_nor2b_1 _11838_ (.A(_04148_),
    .B_N(_03388_),
    .Y(_04149_));
 sg13g2_nor3_1 _11839_ (.A(net348),
    .B(_04108_),
    .C(_04149_),
    .Y(_04150_));
 sg13g2_nand2_1 _11840_ (.Y(_04151_),
    .A(\i_tinyqv.cpu.alu_op[1] ),
    .B(net581));
 sg13g2_nand3_1 _11841_ (.B(_04147_),
    .C(_04151_),
    .A(net180),
    .Y(_04152_));
 sg13g2_nand3_1 _11842_ (.B(net348),
    .C(net180),
    .A(net3863),
    .Y(_04153_));
 sg13g2_a21oi_1 _11843_ (.A1(_04152_),
    .A2(_04153_),
    .Y(_04154_),
    .B1(_04150_));
 sg13g2_a21oi_1 _11844_ (.A1(net3525),
    .A2(_04150_),
    .Y(_04155_),
    .B1(net179));
 sg13g2_nand2b_1 _11845_ (.Y(_00623_),
    .B(_04155_),
    .A_N(_04154_));
 sg13g2_nand3_1 _11846_ (.B(_03387_),
    .C(net341),
    .A(_02250_),
    .Y(_04156_));
 sg13g2_o21ai_1 _11847_ (.B1(net180),
    .Y(_04157_),
    .A1(_04148_),
    .A2(_04156_));
 sg13g2_nand2_1 _11848_ (.Y(_04158_),
    .A(_04152_),
    .B(_04157_));
 sg13g2_a21oi_1 _11849_ (.A1(net3525),
    .A2(_04108_),
    .Y(_04159_),
    .B1(_04158_));
 sg13g2_nor2_1 _11850_ (.A(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .B(_04157_),
    .Y(_04160_));
 sg13g2_nor3_1 _11851_ (.A(net179),
    .B(_04159_),
    .C(_04160_),
    .Y(_00624_));
 sg13g2_and2_1 _11852_ (.A(_02529_),
    .B(_03502_),
    .X(_04161_));
 sg13g2_nand2_1 _11853_ (.Y(_04162_),
    .A(_02529_),
    .B(_03502_));
 sg13g2_nand2b_1 _11854_ (.Y(_04163_),
    .B(net94),
    .A_N(_03505_));
 sg13g2_nor2b_2 _11855_ (.A(_03498_),
    .B_N(_04163_),
    .Y(_04164_));
 sg13g2_nor2_2 _11856_ (.A(net90),
    .B(_04164_),
    .Y(_04165_));
 sg13g2_or2_1 _11857_ (.X(_04166_),
    .B(_04165_),
    .A(net648));
 sg13g2_nand2b_1 _11858_ (.Y(_04167_),
    .B(_03507_),
    .A_N(net207));
 sg13g2_nor2_2 _11859_ (.A(net118),
    .B(_04167_),
    .Y(_04168_));
 sg13g2_or2_1 _11860_ (.X(_04169_),
    .B(_04167_),
    .A(net118));
 sg13g2_nand2_1 _11861_ (.Y(_04170_),
    .A(_03507_),
    .B(net207));
 sg13g2_nand2_2 _11862_ (.Y(_04171_),
    .A(_03484_),
    .B(net207));
 sg13g2_nor2_2 _11863_ (.A(net333),
    .B(_04171_),
    .Y(_04172_));
 sg13g2_nor2_1 _11864_ (.A(net118),
    .B(_04171_),
    .Y(_04173_));
 sg13g2_nand2_1 _11865_ (.Y(_04174_),
    .A(net286),
    .B(_04173_));
 sg13g2_o21ai_1 _11866_ (.B1(_04174_),
    .Y(_04175_),
    .A1(_03518_),
    .A2(_04170_));
 sg13g2_inv_1 _11867_ (.Y(_04176_),
    .A(_04175_));
 sg13g2_nor2_2 _11868_ (.A(net212),
    .B(net210),
    .Y(_04177_));
 sg13g2_nor2b_2 _11869_ (.A(_04170_),
    .B_N(_04177_),
    .Y(_04178_));
 sg13g2_nand3_1 _11870_ (.B(net207),
    .C(_04177_),
    .A(_03507_),
    .Y(_04179_));
 sg13g2_and2_1 _11871_ (.A(_03519_),
    .B(_03556_),
    .X(_04180_));
 sg13g2_nand2_1 _11872_ (.Y(_04181_),
    .A(_03519_),
    .B(_03556_));
 sg13g2_nor3_2 _11873_ (.A(net333),
    .B(net211),
    .C(_04171_),
    .Y(_04182_));
 sg13g2_nor4_1 _11874_ (.A(_04175_),
    .B(_04178_),
    .C(_04180_),
    .D(_04182_),
    .Y(_04183_));
 sg13g2_o21ai_1 _11875_ (.B1(_03557_),
    .Y(_04184_),
    .A1(_03559_),
    .A2(_03561_));
 sg13g2_nand3_1 _11876_ (.B(_04183_),
    .C(_04184_),
    .A(net218),
    .Y(_04185_));
 sg13g2_inv_1 _11877_ (.Y(_04186_),
    .A(_04185_));
 sg13g2_nor2_2 _11878_ (.A(_04168_),
    .B(_04185_),
    .Y(_04187_));
 sg13g2_nor2_1 _11879_ (.A(net282),
    .B(_04187_),
    .Y(_04188_));
 sg13g2_nor2_1 _11880_ (.A(_03557_),
    .B(_04172_),
    .Y(_04189_));
 sg13g2_nand2_1 _11881_ (.Y(_04190_),
    .A(_03507_),
    .B(net211));
 sg13g2_nand3_1 _11882_ (.B(_04189_),
    .C(_04190_),
    .A(_04183_),
    .Y(_04191_));
 sg13g2_nand2_1 _11883_ (.Y(_04192_),
    .A(_03557_),
    .B(net205));
 sg13g2_nand2_2 _11884_ (.Y(_04193_),
    .A(_03519_),
    .B(_04172_));
 sg13g2_a22oi_1 _11885_ (.Y(_04194_),
    .B1(_03563_),
    .B2(net205),
    .A2(net207),
    .A1(_03520_));
 sg13g2_nand2_1 _11886_ (.Y(_04195_),
    .A(_04193_),
    .B(_04194_));
 sg13g2_mux2_1 _11887_ (.A0(net284),
    .A1(_04195_),
    .S(_04191_),
    .X(_04196_));
 sg13g2_a21oi_1 _11888_ (.A1(net216),
    .A2(_04196_),
    .Y(_04197_),
    .B1(_04188_));
 sg13g2_nor2_1 _11889_ (.A(_04161_),
    .B(_04197_),
    .Y(_04198_));
 sg13g2_a21oi_1 _11890_ (.A1(net3035),
    .A2(net90),
    .Y(_04199_),
    .B1(_04198_));
 sg13g2_nand2_1 _11891_ (.Y(_04200_),
    .A(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .B(net64));
 sg13g2_o21ai_1 _11892_ (.B1(_04200_),
    .Y(_00625_),
    .A1(net64),
    .A2(_04199_));
 sg13g2_nand2_1 _11893_ (.Y(_04201_),
    .A(net217),
    .B(_03522_));
 sg13g2_or2_1 _11894_ (.X(_04202_),
    .B(_04201_),
    .A(_04191_));
 sg13g2_o21ai_1 _11895_ (.B1(_04202_),
    .Y(_04203_),
    .A1(net204),
    .A2(_04187_));
 sg13g2_nor3_1 _11896_ (.A(_03179_),
    .B(_03767_),
    .C(net89),
    .Y(_04204_));
 sg13g2_a21oi_1 _11897_ (.A1(net89),
    .A2(_04203_),
    .Y(_04205_),
    .B1(_04204_));
 sg13g2_nand2_1 _11898_ (.Y(_04206_),
    .A(net3638),
    .B(net65));
 sg13g2_o21ai_1 _11899_ (.B1(_04206_),
    .Y(_00626_),
    .A1(net65),
    .A2(_04205_));
 sg13g2_or2_1 _11900_ (.X(_04207_),
    .B(_03179_),
    .A(net661));
 sg13g2_nand3b_1 _11901_ (.B(net120),
    .C(net216),
    .Y(_04208_),
    .A_N(_04191_));
 sg13g2_o21ai_1 _11902_ (.B1(_04208_),
    .Y(_04209_),
    .A1(_03575_),
    .A2(_04187_));
 sg13g2_and3_1 _11903_ (.X(_04210_),
    .A(_03180_),
    .B(net90),
    .C(_04207_));
 sg13g2_a21oi_1 _11904_ (.A1(net89),
    .A2(_04209_),
    .Y(_04211_),
    .B1(_04210_));
 sg13g2_nand2_1 _11905_ (.Y(_04212_),
    .A(net661),
    .B(net65));
 sg13g2_o21ai_1 _11906_ (.B1(_04212_),
    .Y(_00627_),
    .A1(net64),
    .A2(_04211_));
 sg13g2_a21oi_1 _11907_ (.A1(net107),
    .A2(_04191_),
    .Y(_04213_),
    .B1(_03487_));
 sg13g2_a21oi_1 _11908_ (.A1(_04186_),
    .A2(_04193_),
    .Y(_04214_),
    .B1(_03569_));
 sg13g2_nor3_2 _11909_ (.A(net90),
    .B(_04213_),
    .C(_04214_),
    .Y(_04215_));
 sg13g2_xor2_1 _11910_ (.B(_03180_),
    .A(net660),
    .X(_04216_));
 sg13g2_a21oi_1 _11911_ (.A1(net90),
    .A2(_04216_),
    .Y(_04217_),
    .B1(_04215_));
 sg13g2_mux2_1 _11912_ (.A0(_04217_),
    .A1(net660),
    .S(net65),
    .X(_00628_));
 sg13g2_nand2_1 _11913_ (.Y(_04218_),
    .A(net3138),
    .B(\i_uart_tx.cycle_counter[0] ));
 sg13g2_nor2_1 _11914_ (.A(\i_uart_tx.cycle_counter[2] ),
    .B(_04218_),
    .Y(_04219_));
 sg13g2_nand2_1 _11915_ (.Y(_04220_),
    .A(\i_uart_tx.cycle_counter[5] ),
    .B(\i_uart_tx.cycle_counter[3] ));
 sg13g2_nor2_1 _11916_ (.A(\i_uart_tx.cycle_counter[10] ),
    .B(\i_uart_tx.cycle_counter[8] ),
    .Y(_04221_));
 sg13g2_nor4_1 _11917_ (.A(\i_uart_tx.cycle_counter[7] ),
    .B(\i_uart_tx.cycle_counter[6] ),
    .C(\i_uart_tx.cycle_counter[4] ),
    .D(_04220_),
    .Y(_04222_));
 sg13g2_nand4_1 _11918_ (.B(_04219_),
    .C(_04221_),
    .A(\i_uart_tx.cycle_counter[9] ),
    .Y(_04223_),
    .D(_04222_));
 sg13g2_o21ai_1 _11919_ (.B1(net3749),
    .Y(_04224_),
    .A1(\i_uart_tx.fsm_state[2] ),
    .A2(net3983));
 sg13g2_nand3b_1 _11920_ (.B(_04224_),
    .C(_03097_),
    .Y(_04225_),
    .A_N(_04223_));
 sg13g2_and3_1 _11921_ (.X(_04226_),
    .A(_02076_),
    .B(net290),
    .C(_03098_));
 sg13g2_nand3_1 _11922_ (.B(net290),
    .C(_03098_),
    .A(_02076_),
    .Y(_04227_));
 sg13g2_o21ai_1 _11923_ (.B1(net178),
    .Y(_04228_),
    .A1(_01575_),
    .A2(net405));
 sg13g2_a21oi_1 _11924_ (.A1(net3502),
    .A2(net405),
    .Y(_04229_),
    .B1(_04228_));
 sg13g2_o21ai_1 _11925_ (.B1(net537),
    .Y(_04230_),
    .A1(\data_to_write[0] ),
    .A2(net178));
 sg13g2_nor2_1 _11926_ (.A(net3503),
    .B(_04230_),
    .Y(_00629_));
 sg13g2_o21ai_1 _11927_ (.B1(net178),
    .Y(_04231_),
    .A1(_01574_),
    .A2(net405));
 sg13g2_a21oi_1 _11928_ (.A1(net3527),
    .A2(net405),
    .Y(_04232_),
    .B1(_04231_));
 sg13g2_o21ai_1 _11929_ (.B1(net537),
    .Y(_04233_),
    .A1(\data_to_write[1] ),
    .A2(net177));
 sg13g2_nor2_1 _11930_ (.A(_04232_),
    .B(_04233_),
    .Y(_00630_));
 sg13g2_o21ai_1 _11931_ (.B1(net177),
    .Y(_04234_),
    .A1(_01573_),
    .A2(net405));
 sg13g2_a21oi_1 _11932_ (.A1(net3494),
    .A2(net405),
    .Y(_04235_),
    .B1(_04234_));
 sg13g2_o21ai_1 _11933_ (.B1(net535),
    .Y(_04236_),
    .A1(\data_to_write[2] ),
    .A2(net177));
 sg13g2_nor2_1 _11934_ (.A(_04235_),
    .B(_04236_),
    .Y(_00631_));
 sg13g2_o21ai_1 _11935_ (.B1(net178),
    .Y(_04237_),
    .A1(_01572_),
    .A2(net404));
 sg13g2_a21oi_1 _11936_ (.A1(net3472),
    .A2(net404),
    .Y(_04238_),
    .B1(_04237_));
 sg13g2_o21ai_1 _11937_ (.B1(net535),
    .Y(_04239_),
    .A1(\data_to_write[3] ),
    .A2(net178));
 sg13g2_nor2_1 _11938_ (.A(_04238_),
    .B(_04239_),
    .Y(_00632_));
 sg13g2_o21ai_1 _11939_ (.B1(net178),
    .Y(_04240_),
    .A1(_01571_),
    .A2(net404));
 sg13g2_a21oi_1 _11940_ (.A1(net3428),
    .A2(net404),
    .Y(_04241_),
    .B1(_04240_));
 sg13g2_o21ai_1 _11941_ (.B1(net536),
    .Y(_04242_),
    .A1(\data_to_write[4] ),
    .A2(net177));
 sg13g2_nor2_1 _11942_ (.A(net3429),
    .B(_04242_),
    .Y(_00633_));
 sg13g2_o21ai_1 _11943_ (.B1(net177),
    .Y(_04243_),
    .A1(_01570_),
    .A2(net405));
 sg13g2_a21oi_1 _11944_ (.A1(net3514),
    .A2(net404),
    .Y(_04244_),
    .B1(_04243_));
 sg13g2_o21ai_1 _11945_ (.B1(net536),
    .Y(_04245_),
    .A1(net598),
    .A2(net177));
 sg13g2_nor2_1 _11946_ (.A(_04244_),
    .B(_04245_),
    .Y(_00634_));
 sg13g2_o21ai_1 _11947_ (.B1(net177),
    .Y(_04246_),
    .A1(_01569_),
    .A2(net404));
 sg13g2_a21oi_1 _11948_ (.A1(net3452),
    .A2(net404),
    .Y(_04247_),
    .B1(_04246_));
 sg13g2_o21ai_1 _11949_ (.B1(net535),
    .Y(_04248_),
    .A1(\data_to_write[6] ),
    .A2(net177));
 sg13g2_nor2_1 _11950_ (.A(net3453),
    .B(_04248_),
    .Y(_00635_));
 sg13g2_and2_1 _11951_ (.A(\i_uart_tx.data_to_send[7] ),
    .B(net404),
    .X(_04249_));
 sg13g2_o21ai_1 _11952_ (.B1(net535),
    .Y(_04250_),
    .A1(_04226_),
    .A2(_04249_));
 sg13g2_a21oi_1 _11953_ (.A1(net2998),
    .A2(_04226_),
    .Y(_00636_),
    .B1(_04250_));
 sg13g2_nand2b_2 _11954_ (.Y(_04251_),
    .B(_04223_),
    .A_N(net517));
 sg13g2_nand2_1 _11955_ (.Y(_04252_),
    .A(net2833),
    .B(_03099_));
 sg13g2_nand2_1 _11956_ (.Y(_04253_),
    .A(\i_uart_tx.cycle_counter[0] ),
    .B(_03098_));
 sg13g2_a21oi_1 _11957_ (.A1(_04252_),
    .A2(_04253_),
    .Y(_00637_),
    .B1(_04251_));
 sg13g2_a21oi_1 _11958_ (.A1(\i_uart_tx.cycle_counter[0] ),
    .A2(_03099_),
    .Y(_04254_),
    .B1(net3138));
 sg13g2_nor2_1 _11959_ (.A(_03098_),
    .B(_04218_),
    .Y(_04255_));
 sg13g2_nor3_1 _11960_ (.A(net403),
    .B(net3139),
    .C(_04255_),
    .Y(_00638_));
 sg13g2_nor2_1 _11961_ (.A(net3621),
    .B(_04255_),
    .Y(_04256_));
 sg13g2_and2_1 _11962_ (.A(net3621),
    .B(_04255_),
    .X(_04257_));
 sg13g2_nor3_1 _11963_ (.A(_04251_),
    .B(net3622),
    .C(_04257_),
    .Y(_00639_));
 sg13g2_nor2_1 _11964_ (.A(net3594),
    .B(_04257_),
    .Y(_04258_));
 sg13g2_and2_1 _11965_ (.A(net3594),
    .B(_04257_),
    .X(_04259_));
 sg13g2_nor3_1 _11966_ (.A(_04251_),
    .B(net3595),
    .C(_04259_),
    .Y(_00640_));
 sg13g2_nor2_1 _11967_ (.A(net3612),
    .B(_04259_),
    .Y(_04260_));
 sg13g2_and2_1 _11968_ (.A(net3612),
    .B(_04259_),
    .X(_04261_));
 sg13g2_nor3_1 _11969_ (.A(net403),
    .B(_04260_),
    .C(_04261_),
    .Y(_00641_));
 sg13g2_nor2_1 _11970_ (.A(net3608),
    .B(_04261_),
    .Y(_04262_));
 sg13g2_and2_1 _11971_ (.A(net3608),
    .B(_04261_),
    .X(_04263_));
 sg13g2_nor3_1 _11972_ (.A(net403),
    .B(net3609),
    .C(_04263_),
    .Y(_00642_));
 sg13g2_nor2_1 _11973_ (.A(net3601),
    .B(_04263_),
    .Y(_04264_));
 sg13g2_and2_1 _11974_ (.A(net3601),
    .B(_04263_),
    .X(_04265_));
 sg13g2_nor3_1 _11975_ (.A(net403),
    .B(net3602),
    .C(_04265_),
    .Y(_00643_));
 sg13g2_nor2_1 _11976_ (.A(net3516),
    .B(_04265_),
    .Y(_04266_));
 sg13g2_and2_1 _11977_ (.A(net3516),
    .B(_04265_),
    .X(_04267_));
 sg13g2_nor3_1 _11978_ (.A(net403),
    .B(net3517),
    .C(_04267_),
    .Y(_00644_));
 sg13g2_nor2_1 _11979_ (.A(net3581),
    .B(_04267_),
    .Y(_04268_));
 sg13g2_and2_1 _11980_ (.A(net3581),
    .B(_04267_),
    .X(_04269_));
 sg13g2_nor3_1 _11981_ (.A(net403),
    .B(_04268_),
    .C(_04269_),
    .Y(_00645_));
 sg13g2_nor2_1 _11982_ (.A(net3533),
    .B(_04269_),
    .Y(_04270_));
 sg13g2_and2_1 _11983_ (.A(net3533),
    .B(_04269_),
    .X(_04271_));
 sg13g2_nor3_1 _11984_ (.A(net403),
    .B(net3534),
    .C(_04271_),
    .Y(_00646_));
 sg13g2_a21oi_1 _11985_ (.A1(net3806),
    .A2(_04271_),
    .Y(_04272_),
    .B1(net403));
 sg13g2_o21ai_1 _11986_ (.B1(_04272_),
    .Y(_04273_),
    .A1(net3806),
    .A2(_04271_));
 sg13g2_inv_1 _11987_ (.Y(_00647_),
    .A(_04273_));
 sg13g2_nor4_2 _11988_ (.A(_01566_),
    .B(\i_uart_tx.fsm_state[2] ),
    .C(_01567_),
    .Y(_04274_),
    .D(\i_uart_tx.fsm_state[0] ));
 sg13g2_nor4_1 _11989_ (.A(net4062),
    .B(_03096_),
    .C(_04223_),
    .D(_04274_),
    .Y(_04275_));
 sg13g2_a21oi_1 _11990_ (.A1(net4062),
    .A2(_04223_),
    .Y(_04276_),
    .B1(_04275_));
 sg13g2_a21oi_1 _11991_ (.A1(net178),
    .A2(_04276_),
    .Y(_00648_),
    .B1(net398));
 sg13g2_nand2_1 _11992_ (.Y(_04277_),
    .A(_03099_),
    .B(_04223_));
 sg13g2_o21ai_1 _11993_ (.B1(_04277_),
    .Y(_04278_),
    .A1(net4132),
    .A2(_04274_));
 sg13g2_o21ai_1 _11994_ (.B1(net537),
    .Y(_04279_),
    .A1(_01567_),
    .A2(_04278_));
 sg13g2_a21oi_1 _11995_ (.A1(_01567_),
    .A2(_04278_),
    .Y(_00649_),
    .B1(_04279_));
 sg13g2_nor3_1 _11996_ (.A(_01567_),
    .B(_01568_),
    .C(_04223_),
    .Y(_04280_));
 sg13g2_nand3_1 _11997_ (.B(net3983),
    .C(net4132),
    .A(net4000),
    .Y(_04281_));
 sg13g2_nor2_1 _11998_ (.A(_04223_),
    .B(_04281_),
    .Y(_04282_));
 sg13g2_o21ai_1 _11999_ (.B1(net537),
    .Y(_04283_),
    .A1(net4000),
    .A2(_04280_));
 sg13g2_nor2_1 _12000_ (.A(_04282_),
    .B(_04283_),
    .Y(_00650_));
 sg13g2_xnor2_1 _12001_ (.Y(_04284_),
    .A(_01566_),
    .B(_04281_));
 sg13g2_nor2_1 _12002_ (.A(_04274_),
    .B(_04284_),
    .Y(_04285_));
 sg13g2_a22oi_1 _12003_ (.Y(_04286_),
    .B1(_04277_),
    .B2(_04285_),
    .A2(_04223_),
    .A1(net3749));
 sg13g2_nor2_1 _12004_ (.A(net397),
    .B(_04286_),
    .Y(_00651_));
 sg13g2_nor3_1 _12005_ (.A(_01607_),
    .B(\i_uart_rx.cycle_counter[8] ),
    .C(\i_uart_rx.cycle_counter[10] ),
    .Y(_04287_));
 sg13g2_or2_1 _12006_ (.X(_04288_),
    .B(\i_uart_rx.cycle_counter[6] ),
    .A(\i_uart_rx.cycle_counter[7] ));
 sg13g2_and2_1 _12007_ (.A(net3335),
    .B(\i_uart_rx.cycle_counter[1] ),
    .X(_04289_));
 sg13g2_nor3_1 _12008_ (.A(net3903),
    .B(net3642),
    .C(net4051),
    .Y(_04290_));
 sg13g2_o21ai_1 _12009_ (.B1(\i_uart_rx.fsm_state[3] ),
    .Y(_04291_),
    .A1(\i_uart_rx.fsm_state[2] ),
    .A2(\i_uart_rx.fsm_state[1] ));
 sg13g2_nand4_1 _12010_ (.B(\i_uart_rx.cycle_counter[5] ),
    .C(_04287_),
    .A(\i_uart_rx.cycle_counter[3] ),
    .Y(_04292_),
    .D(_04289_));
 sg13g2_nor4_2 _12011_ (.A(\i_uart_rx.cycle_counter[2] ),
    .B(\i_uart_rx.cycle_counter[4] ),
    .C(_04288_),
    .Y(_04293_),
    .D(_04292_));
 sg13g2_inv_1 _12012_ (.Y(_04294_),
    .A(_04293_));
 sg13g2_nand3b_1 _12013_ (.B(_04291_),
    .C(_04293_),
    .Y(_04295_),
    .A_N(_04290_));
 sg13g2_mux2_1 _12014_ (.A0(net3420),
    .A1(\i_uart_rx.recieved_data[0] ),
    .S(_04295_),
    .X(_00652_));
 sg13g2_mux2_1 _12015_ (.A0(net3535),
    .A1(net3420),
    .S(_04295_),
    .X(_00653_));
 sg13g2_mux2_1 _12016_ (.A0(net3587),
    .A1(net3535),
    .S(_04295_),
    .X(_00654_));
 sg13g2_mux2_1 _12017_ (.A0(net3511),
    .A1(\i_uart_rx.recieved_data[3] ),
    .S(_04295_),
    .X(_00655_));
 sg13g2_mux2_1 _12018_ (.A0(net3486),
    .A1(\i_uart_rx.recieved_data[4] ),
    .S(_04295_),
    .X(_00656_));
 sg13g2_mux2_1 _12019_ (.A0(net3505),
    .A1(net3486),
    .S(_04295_),
    .X(_00657_));
 sg13g2_mux2_1 _12020_ (.A0(net3780),
    .A1(net3505),
    .S(_04295_),
    .X(_00658_));
 sg13g2_mux2_1 _12021_ (.A0(net3338),
    .A1(\i_uart_rx.recieved_data[7] ),
    .S(_04295_),
    .X(_00659_));
 sg13g2_a21oi_1 _12022_ (.A1(_03599_),
    .A2(_03619_),
    .Y(_04296_),
    .B1(_03626_));
 sg13g2_a21o_1 _12023_ (.A2(_03619_),
    .A1(_03599_),
    .B1(_03626_),
    .X(_04297_));
 sg13g2_nor2_2 _12024_ (.A(_00199_),
    .B(_03795_),
    .Y(_04298_));
 sg13g2_nor2_1 _12025_ (.A(net72),
    .B(net401),
    .Y(_04299_));
 sg13g2_or2_2 _12026_ (.X(_04300_),
    .B(net401),
    .A(net72));
 sg13g2_nor3_2 _12027_ (.A(_03599_),
    .B(_03620_),
    .C(_03626_),
    .Y(_04301_));
 sg13g2_nor2_2 _12028_ (.A(_01604_),
    .B(_04301_),
    .Y(_04302_));
 sg13g2_nor3_1 _12029_ (.A(_01604_),
    .B(_03619_),
    .C(_03626_),
    .Y(_04303_));
 sg13g2_nand2_2 _12030_ (.Y(_04304_),
    .A(net72),
    .B(_04302_));
 sg13g2_a22oi_1 _12031_ (.Y(_04305_),
    .B1(net276),
    .B2(net2388),
    .A2(net59),
    .A1(net3267));
 sg13g2_inv_1 _12032_ (.Y(_00660_),
    .A(_04305_));
 sg13g2_nand2_1 _12033_ (.Y(_04306_),
    .A(_00120_),
    .B(net457));
 sg13g2_a21oi_1 _12034_ (.A1(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .A2(_04306_),
    .Y(_04307_),
    .B1(\i_tinyqv.cpu.i_core.mem_op[1] ));
 sg13g2_o21ai_1 _12035_ (.B1(_04307_),
    .Y(_04308_),
    .A1(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .A2(net353));
 sg13g2_nor3_1 _12036_ (.A(\i_tinyqv.cpu.i_core.mem_op[2] ),
    .B(_02987_),
    .C(_04308_),
    .Y(_04309_));
 sg13g2_nand2_1 _12037_ (.Y(_04310_),
    .A(_03713_),
    .B(_04309_));
 sg13g2_nand2_1 _12038_ (.Y(_04311_),
    .A(net3388),
    .B(net336));
 sg13g2_o21ai_1 _12039_ (.B1(_04310_),
    .Y(_00661_),
    .A1(_04309_),
    .A2(_04311_));
 sg13g2_nor2b_1 _12040_ (.A(\i_uart_rx.fsm_state[0] ),
    .B_N(_04290_),
    .Y(_04312_));
 sg13g2_or4_2 _12041_ (.A(net517),
    .B(_03287_),
    .C(_04293_),
    .D(_04312_),
    .X(_04313_));
 sg13g2_nor2_1 _12042_ (.A(_01707_),
    .B(net339),
    .Y(_00662_));
 sg13g2_nor2_1 _12043_ (.A(net3335),
    .B(\i_uart_rx.cycle_counter[1] ),
    .Y(_04314_));
 sg13g2_nor3_1 _12044_ (.A(_04289_),
    .B(net339),
    .C(net3336),
    .Y(_00663_));
 sg13g2_and2_1 _12045_ (.A(net3745),
    .B(_04289_),
    .X(_04315_));
 sg13g2_nor2_1 _12046_ (.A(net3745),
    .B(_04289_),
    .Y(_04316_));
 sg13g2_nor3_1 _12047_ (.A(_04313_),
    .B(_04315_),
    .C(net3746),
    .Y(_00664_));
 sg13g2_and2_1 _12048_ (.A(net3610),
    .B(_04315_),
    .X(_04317_));
 sg13g2_nor2_1 _12049_ (.A(net3610),
    .B(_04315_),
    .Y(_04318_));
 sg13g2_nor3_1 _12050_ (.A(net339),
    .B(_04317_),
    .C(net3611),
    .Y(_00665_));
 sg13g2_and2_1 _12051_ (.A(net3744),
    .B(_04317_),
    .X(_04319_));
 sg13g2_nor2_1 _12052_ (.A(net3744),
    .B(_04317_),
    .Y(_04320_));
 sg13g2_nor3_1 _12053_ (.A(net339),
    .B(_04319_),
    .C(_04320_),
    .Y(_00666_));
 sg13g2_and2_1 _12054_ (.A(net3739),
    .B(_04319_),
    .X(_04321_));
 sg13g2_nor2_1 _12055_ (.A(net3739),
    .B(_04319_),
    .Y(_04322_));
 sg13g2_nor3_1 _12056_ (.A(net339),
    .B(_04321_),
    .C(net3740),
    .Y(_00667_));
 sg13g2_nor2_1 _12057_ (.A(net3490),
    .B(_04321_),
    .Y(_04323_));
 sg13g2_and2_1 _12058_ (.A(net3490),
    .B(_04321_),
    .X(_04324_));
 sg13g2_nor3_1 _12059_ (.A(_04313_),
    .B(net3491),
    .C(_04324_),
    .Y(_00668_));
 sg13g2_nor2_1 _12060_ (.A(net3596),
    .B(_04324_),
    .Y(_04325_));
 sg13g2_and2_1 _12061_ (.A(net3596),
    .B(_04324_),
    .X(_04326_));
 sg13g2_nor3_1 _12062_ (.A(_04313_),
    .B(_04325_),
    .C(_04326_),
    .Y(_00669_));
 sg13g2_nor2_1 _12063_ (.A(net3709),
    .B(_04326_),
    .Y(_04327_));
 sg13g2_and2_1 _12064_ (.A(net3709),
    .B(_04326_),
    .X(_04328_));
 sg13g2_nor3_1 _12065_ (.A(net339),
    .B(_04327_),
    .C(_04328_),
    .Y(_00670_));
 sg13g2_nor2_1 _12066_ (.A(net3762),
    .B(_04328_),
    .Y(_04329_));
 sg13g2_and2_1 _12067_ (.A(net3762),
    .B(_04328_),
    .X(_04330_));
 sg13g2_nor3_1 _12068_ (.A(net339),
    .B(_04329_),
    .C(_04330_),
    .Y(_00671_));
 sg13g2_a21oi_1 _12069_ (.A1(net3872),
    .A2(_04330_),
    .Y(_04331_),
    .B1(net339));
 sg13g2_o21ai_1 _12070_ (.B1(_04331_),
    .Y(_04332_),
    .A1(net3872),
    .A2(_04330_));
 sg13g2_inv_1 _12071_ (.Y(_00672_),
    .A(_04332_));
 sg13g2_nor3_1 _12072_ (.A(\i_uart_rx.cycle_counter[3] ),
    .B(_01606_),
    .C(\i_uart_rx.cycle_counter[5] ),
    .Y(_04333_));
 sg13g2_nor3_1 _12073_ (.A(_01605_),
    .B(\i_uart_rx.cycle_counter[1] ),
    .C(_04288_),
    .Y(_04334_));
 sg13g2_nand3_1 _12074_ (.B(_04333_),
    .C(_04334_),
    .A(\i_uart_rx.cycle_counter[4] ),
    .Y(_04335_));
 sg13g2_nor4_2 _12075_ (.A(\i_uart_rx.cycle_counter[9] ),
    .B(_01608_),
    .C(\i_uart_rx.cycle_counter[10] ),
    .Y(_04336_),
    .D(_04335_));
 sg13g2_o21ai_1 _12076_ (.B1(net536),
    .Y(_04337_),
    .A1(\i_uart_rx.bit_sample ),
    .A2(_04336_));
 sg13g2_a21oi_1 _12077_ (.A1(_01565_),
    .A2(_04336_),
    .Y(_00673_),
    .B1(_04337_));
 sg13g2_nand2_1 _12078_ (.Y(_00674_),
    .A(net536),
    .B(_04290_));
 sg13g2_and2_1 _12079_ (.A(_02529_),
    .B(net290),
    .X(_04338_));
 sg13g2_a21oi_2 _12080_ (.B1(_03288_),
    .Y(_04339_),
    .A2(_04338_),
    .A1(\i_tinyqv.cpu.is_load ));
 sg13g2_nor2_1 _12081_ (.A(\i_uart_rx.fsm_state[0] ),
    .B(_03286_),
    .Y(_04340_));
 sg13g2_nor3_1 _12082_ (.A(\i_uart_rx.fsm_state[0] ),
    .B(_00244_),
    .C(_03286_),
    .Y(_04341_));
 sg13g2_nor2_2 _12083_ (.A(_03285_),
    .B(_04312_),
    .Y(_04342_));
 sg13g2_a221oi_1 _12084_ (.B2(_04341_),
    .C1(_04342_),
    .B1(_04336_),
    .A1(_01565_),
    .Y(_04343_),
    .A2(_04312_));
 sg13g2_nor2b_1 _12085_ (.A(_04339_),
    .B_N(_04343_),
    .Y(_04344_));
 sg13g2_nand2_2 _12086_ (.Y(_04345_),
    .A(_04294_),
    .B(_04342_));
 sg13g2_nand3b_1 _12087_ (.B(_04293_),
    .C(_04342_),
    .Y(_04346_),
    .A_N(net3751));
 sg13g2_o21ai_1 _12088_ (.B1(_04346_),
    .Y(_04347_),
    .A1(\i_uart_rx.fsm_state[0] ),
    .A2(_04345_));
 sg13g2_nor3_1 _12089_ (.A(net397),
    .B(_04344_),
    .C(net3752),
    .Y(_00675_));
 sg13g2_nand2_1 _12090_ (.Y(_04348_),
    .A(net4053),
    .B(_04336_));
 sg13g2_a21oi_1 _12091_ (.A1(_04340_),
    .A2(_04348_),
    .Y(_04349_),
    .B1(_04339_));
 sg13g2_inv_1 _12092_ (.Y(_04350_),
    .A(_04349_));
 sg13g2_xor2_1 _12093_ (.B(\i_uart_rx.fsm_state[0] ),
    .A(\i_uart_rx.fsm_state[1] ),
    .X(_04351_));
 sg13g2_a21oi_1 _12094_ (.A1(_03286_),
    .A2(_04351_),
    .Y(_04352_),
    .B1(_04350_));
 sg13g2_o21ai_1 _12095_ (.B1(net536),
    .Y(_04353_),
    .A1(net4051),
    .A2(_04345_));
 sg13g2_a21oi_1 _12096_ (.A1(_04345_),
    .A2(_04352_),
    .Y(_00676_),
    .B1(_04353_));
 sg13g2_nand3_1 _12097_ (.B(\i_uart_rx.fsm_state[0] ),
    .C(_04345_),
    .A(\i_uart_rx.fsm_state[1] ),
    .Y(_04354_));
 sg13g2_nand3_1 _12098_ (.B(\i_uart_rx.fsm_state[1] ),
    .C(\i_uart_rx.fsm_state[0] ),
    .A(\i_uart_rx.fsm_state[2] ),
    .Y(_04355_));
 sg13g2_or2_1 _12099_ (.X(_04356_),
    .B(_04355_),
    .A(_04294_));
 sg13g2_nand3_1 _12100_ (.B(_04342_),
    .C(_04356_),
    .A(net535),
    .Y(_04357_));
 sg13g2_a21oi_1 _12101_ (.A1(_01564_),
    .A2(_04354_),
    .Y(_00677_),
    .B1(_04357_));
 sg13g2_xnor2_1 _12102_ (.Y(_04358_),
    .A(\i_uart_rx.fsm_state[3] ),
    .B(_04355_));
 sg13g2_o21ai_1 _12103_ (.B1(_04342_),
    .Y(_04359_),
    .A1(_04294_),
    .A2(_04358_));
 sg13g2_o21ai_1 _12104_ (.B1(net535),
    .Y(_04360_),
    .A1(net3903),
    .A2(_04345_));
 sg13g2_a21oi_1 _12105_ (.A1(_04349_),
    .A2(_04359_),
    .Y(_00678_),
    .B1(_04360_));
 sg13g2_nand2b_1 _12106_ (.Y(_00679_),
    .B(net536),
    .A_N(net2935));
 sg13g2_nand2b_1 _12107_ (.Y(_00680_),
    .B(net529),
    .A_N(net9));
 sg13g2_nand2_1 _12108_ (.Y(_04361_),
    .A(net617),
    .B(_01523_));
 sg13g2_nor2b_1 _12109_ (.A(_03632_),
    .B_N(_04361_),
    .Y(_04362_));
 sg13g2_nor2_1 _12110_ (.A(net398),
    .B(_03632_),
    .Y(_01305_));
 sg13g2_nor4_1 _12111_ (.A(net398),
    .B(net2837),
    .C(_03632_),
    .D(_04361_),
    .Y(_00681_));
 sg13g2_nor2_2 _12112_ (.A(net99),
    .B(net80),
    .Y(_04363_));
 sg13g2_nand3_1 _12113_ (.B(_03604_),
    .C(net69),
    .A(net656),
    .Y(_04364_));
 sg13g2_a21oi_1 _12114_ (.A1(\i_tinyqv.cpu.instr_write_offset[2] ),
    .A2(\i_tinyqv.cpu.instr_write_offset[1] ),
    .Y(_04365_),
    .B1(_04364_));
 sg13g2_or2_1 _12115_ (.X(_04366_),
    .B(_04365_),
    .A(_04364_));
 sg13g2_nor2_1 _12116_ (.A(\i_tinyqv.cpu.instr_data_in[0] ),
    .B(net19),
    .Y(_04367_));
 sg13g2_a21oi_1 _12117_ (.A1(_03604_),
    .A2(net69),
    .Y(_04368_),
    .B1(net514));
 sg13g2_or2_1 _12118_ (.X(_04369_),
    .B(_04368_),
    .A(_04365_));
 sg13g2_a21oi_1 _12119_ (.A1(_01600_),
    .A2(_04369_),
    .Y(_00682_),
    .B1(_04367_));
 sg13g2_nor2_1 _12120_ (.A(\i_tinyqv.cpu.instr_data_in[1] ),
    .B(net18),
    .Y(_04370_));
 sg13g2_a21oi_1 _12121_ (.A1(_01601_),
    .A2(_04369_),
    .Y(_00683_),
    .B1(_04370_));
 sg13g2_nor3_1 _12122_ (.A(_01597_),
    .B(\i_tinyqv.cpu.instr_write_offset[1] ),
    .C(_04364_),
    .Y(_04371_));
 sg13g2_mux2_1 _12123_ (.A0(net3558),
    .A1(\i_tinyqv.cpu.instr_data_in[2] ),
    .S(net43),
    .X(_00684_));
 sg13g2_nor2_1 _12124_ (.A(net3475),
    .B(net43),
    .Y(_04372_));
 sg13g2_a21oi_1 _12125_ (.A1(_01684_),
    .A2(net44),
    .Y(_00685_),
    .B1(_04372_));
 sg13g2_mux2_1 _12126_ (.A0(net3218),
    .A1(\i_tinyqv.cpu.instr_data_in[4] ),
    .S(net43),
    .X(_00686_));
 sg13g2_nor2_1 _12127_ (.A(net3089),
    .B(net42),
    .Y(_04373_));
 sg13g2_a21oi_1 _12128_ (.A1(_01671_),
    .A2(net42),
    .Y(_00687_),
    .B1(_04373_));
 sg13g2_mux2_1 _12129_ (.A0(net3062),
    .A1(\i_tinyqv.cpu.instr_data_in[6] ),
    .S(net43),
    .X(_00688_));
 sg13g2_mux2_1 _12130_ (.A0(net3073),
    .A1(\i_tinyqv.cpu.instr_data_in[7] ),
    .S(net42),
    .X(_00689_));
 sg13g2_nor2_1 _12131_ (.A(net3106),
    .B(net41),
    .Y(_04374_));
 sg13g2_a21oi_1 _12132_ (.A1(_00245_),
    .A2(net41),
    .Y(_00690_),
    .B1(_04374_));
 sg13g2_nor2_1 _12133_ (.A(net3038),
    .B(net44),
    .Y(_04375_));
 sg13g2_a21oi_1 _12134_ (.A1(_00246_),
    .A2(net44),
    .Y(_00691_),
    .B1(_04375_));
 sg13g2_nor2_1 _12135_ (.A(net3025),
    .B(net41),
    .Y(_04376_));
 sg13g2_a21oi_1 _12136_ (.A1(_00247_),
    .A2(net41),
    .Y(_00692_),
    .B1(_04376_));
 sg13g2_nor2_1 _12137_ (.A(net3043),
    .B(net42),
    .Y(_04377_));
 sg13g2_a21oi_1 _12138_ (.A1(_00248_),
    .A2(net42),
    .Y(_00693_),
    .B1(_04377_));
 sg13g2_nor2_1 _12139_ (.A(net3180),
    .B(net43),
    .Y(_04378_));
 sg13g2_a21oi_1 _12140_ (.A1(_00249_),
    .A2(net43),
    .Y(_00694_),
    .B1(_04378_));
 sg13g2_nor2_1 _12141_ (.A(net3031),
    .B(net42),
    .Y(_04379_));
 sg13g2_a21oi_1 _12142_ (.A1(_00250_),
    .A2(net42),
    .Y(_00695_),
    .B1(_04379_));
 sg13g2_nor2_1 _12143_ (.A(net3023),
    .B(net41),
    .Y(_04380_));
 sg13g2_a21oi_1 _12144_ (.A1(_00251_),
    .A2(net41),
    .Y(_00696_),
    .B1(_04380_));
 sg13g2_nor2_1 _12145_ (.A(net3123),
    .B(net41),
    .Y(_04381_));
 sg13g2_a21oi_1 _12146_ (.A1(_00252_),
    .A2(net41),
    .Y(_00697_),
    .B1(_04381_));
 sg13g2_o21ai_1 _12147_ (.B1(net3794),
    .Y(_04382_),
    .A1(net3723),
    .A2(net3827));
 sg13g2_nor2b_1 _12148_ (.A(\i_debug_uart_tx.cycle_counter[4] ),
    .B_N(\i_debug_uart_tx.cycle_counter[3] ),
    .Y(_04383_));
 sg13g2_and4_1 _12149_ (.A(net3693),
    .B(net3434),
    .C(\i_debug_uart_tx.cycle_counter[0] ),
    .D(_04383_),
    .X(_04384_));
 sg13g2_nand4_1 _12150_ (.B(\i_debug_uart_tx.cycle_counter[1] ),
    .C(\i_debug_uart_tx.cycle_counter[0] ),
    .A(\i_debug_uart_tx.cycle_counter[2] ),
    .Y(_04385_),
    .D(_04383_));
 sg13g2_and2_1 _12151_ (.A(_03092_),
    .B(_04384_),
    .X(_04386_));
 sg13g2_nand2_1 _12152_ (.Y(_04387_),
    .A(_04382_),
    .B(_04386_));
 sg13g2_nand4_1 _12153_ (.B(_02113_),
    .C(_03079_),
    .A(_02076_),
    .Y(_04388_),
    .D(_03093_));
 sg13g2_o21ai_1 _12154_ (.B1(net275),
    .Y(_04389_),
    .A1(_01563_),
    .A2(net400));
 sg13g2_and4_1 _12155_ (.A(_02076_),
    .B(_02113_),
    .C(_03079_),
    .D(_03093_),
    .X(_04390_));
 sg13g2_a21oi_1 _12156_ (.A1(net3478),
    .A2(net400),
    .Y(_04391_),
    .B1(_04389_));
 sg13g2_o21ai_1 _12157_ (.B1(net527),
    .Y(_04392_),
    .A1(\data_to_write[0] ),
    .A2(net275));
 sg13g2_nor2_1 _12158_ (.A(net3479),
    .B(_04392_),
    .Y(_00698_));
 sg13g2_o21ai_1 _12159_ (.B1(net275),
    .Y(_04393_),
    .A1(_01562_),
    .A2(net400));
 sg13g2_a21oi_1 _12160_ (.A1(net3523),
    .A2(net400),
    .Y(_04394_),
    .B1(_04393_));
 sg13g2_o21ai_1 _12161_ (.B1(net527),
    .Y(_04395_),
    .A1(net601),
    .A2(net275));
 sg13g2_nor2_1 _12162_ (.A(_04394_),
    .B(_04395_),
    .Y(_00699_));
 sg13g2_o21ai_1 _12163_ (.B1(net274),
    .Y(_04396_),
    .A1(_01561_),
    .A2(net400));
 sg13g2_a21oi_1 _12164_ (.A1(net3446),
    .A2(net399),
    .Y(_04397_),
    .B1(_04396_));
 sg13g2_o21ai_1 _12165_ (.B1(net527),
    .Y(_04398_),
    .A1(net600),
    .A2(net275));
 sg13g2_nor2_1 _12166_ (.A(net3447),
    .B(_04398_),
    .Y(_00700_));
 sg13g2_o21ai_1 _12167_ (.B1(net275),
    .Y(_04399_),
    .A1(_01560_),
    .A2(net400));
 sg13g2_a21oi_1 _12168_ (.A1(net3555),
    .A2(net400),
    .Y(_04400_),
    .B1(_04399_));
 sg13g2_o21ai_1 _12169_ (.B1(net527),
    .Y(_04401_),
    .A1(\data_to_write[3] ),
    .A2(net274));
 sg13g2_nor2_1 _12170_ (.A(_04400_),
    .B(_04401_),
    .Y(_00701_));
 sg13g2_o21ai_1 _12171_ (.B1(net274),
    .Y(_04402_),
    .A1(_01559_),
    .A2(net399));
 sg13g2_a21oi_1 _12172_ (.A1(net3432),
    .A2(net399),
    .Y(_04403_),
    .B1(_04402_));
 sg13g2_o21ai_1 _12173_ (.B1(net528),
    .Y(_04404_),
    .A1(\data_to_write[4] ),
    .A2(net274));
 sg13g2_nor2_1 _12174_ (.A(_04403_),
    .B(_04404_),
    .Y(_00702_));
 sg13g2_o21ai_1 _12175_ (.B1(net274),
    .Y(_04405_),
    .A1(_01558_),
    .A2(net399));
 sg13g2_a21oi_1 _12176_ (.A1(net3402),
    .A2(net399),
    .Y(_04406_),
    .B1(_04405_));
 sg13g2_o21ai_1 _12177_ (.B1(net527),
    .Y(_04407_),
    .A1(\data_to_write[5] ),
    .A2(net274));
 sg13g2_nor2_1 _12178_ (.A(net3403),
    .B(_04407_),
    .Y(_00703_));
 sg13g2_o21ai_1 _12179_ (.B1(net274),
    .Y(_04408_),
    .A1(_01557_),
    .A2(net399));
 sg13g2_a21oi_1 _12180_ (.A1(net3459),
    .A2(net399),
    .Y(_04409_),
    .B1(_04408_));
 sg13g2_o21ai_1 _12181_ (.B1(net527),
    .Y(_04410_),
    .A1(\data_to_write[6] ),
    .A2(net274));
 sg13g2_nor2_1 _12182_ (.A(_04409_),
    .B(_04410_),
    .Y(_00704_));
 sg13g2_a21oi_1 _12183_ (.A1(net3365),
    .A2(net399),
    .Y(_04411_),
    .B1(_04390_));
 sg13g2_and2_1 _12184_ (.A(net2998),
    .B(_04390_),
    .X(_04412_));
 sg13g2_nor3_1 _12185_ (.A(net397),
    .B(_04411_),
    .C(_04412_),
    .Y(_00705_));
 sg13g2_nor2_1 _12186_ (.A(net2843),
    .B(_03093_),
    .Y(_04413_));
 sg13g2_nand2b_2 _12187_ (.Y(_04414_),
    .B(_04385_),
    .A_N(net516));
 sg13g2_nor2_1 _12188_ (.A(\i_debug_uart_tx.cycle_counter[0] ),
    .B(_03094_),
    .Y(_04415_));
 sg13g2_nor3_1 _12189_ (.A(net2844),
    .B(_04414_),
    .C(_04415_),
    .Y(_00706_));
 sg13g2_a21oi_1 _12190_ (.A1(\i_debug_uart_tx.cycle_counter[0] ),
    .A2(_03094_),
    .Y(_04416_),
    .B1(net3434));
 sg13g2_and3_1 _12191_ (.X(_04417_),
    .A(net3434),
    .B(\i_debug_uart_tx.cycle_counter[0] ),
    .C(_03094_));
 sg13g2_nor3_1 _12192_ (.A(_04414_),
    .B(net3435),
    .C(_04417_),
    .Y(_00707_));
 sg13g2_nor2_1 _12193_ (.A(net3693),
    .B(_04417_),
    .Y(_04418_));
 sg13g2_and2_1 _12194_ (.A(net3693),
    .B(_04417_),
    .X(_04419_));
 sg13g2_nor3_1 _12195_ (.A(_04414_),
    .B(net3694),
    .C(_04419_),
    .Y(_00708_));
 sg13g2_xnor2_1 _12196_ (.Y(_04420_),
    .A(net3651),
    .B(_04419_));
 sg13g2_nor2_1 _12197_ (.A(_04414_),
    .B(net3652),
    .Y(_00709_));
 sg13g2_nand2b_1 _12198_ (.Y(_04421_),
    .B(net2856),
    .A_N(net516));
 sg13g2_a21oi_1 _12199_ (.A1(\i_debug_uart_tx.cycle_counter[3] ),
    .A2(_04419_),
    .Y(_00710_),
    .B1(_04421_));
 sg13g2_nand3_1 _12200_ (.B(_01556_),
    .C(\i_debug_uart_tx.fsm_state[1] ),
    .A(\i_debug_uart_tx.fsm_state[3] ),
    .Y(_04422_));
 sg13g2_nor2b_1 _12201_ (.A(net3852),
    .B_N(_04422_),
    .Y(_04423_));
 sg13g2_a22oi_1 _12202_ (.Y(_04424_),
    .B1(_04386_),
    .B2(_04423_),
    .A2(_04385_),
    .A1(net3852));
 sg13g2_a21oi_1 _12203_ (.A1(_04388_),
    .A2(_04424_),
    .Y(_00711_),
    .B1(net397));
 sg13g2_a21oi_1 _12204_ (.A1(_03094_),
    .A2(_04385_),
    .Y(_04425_),
    .B1(_04423_));
 sg13g2_nor2_1 _12205_ (.A(net3827),
    .B(_04425_),
    .Y(_04426_));
 sg13g2_a21oi_1 _12206_ (.A1(net3827),
    .A2(_04425_),
    .Y(_04427_),
    .B1(net397));
 sg13g2_nor2b_1 _12207_ (.A(_04426_),
    .B_N(_04427_),
    .Y(_00712_));
 sg13g2_nand3_1 _12208_ (.B(\i_debug_uart_tx.fsm_state[0] ),
    .C(_04384_),
    .A(\i_debug_uart_tx.fsm_state[1] ),
    .Y(_04428_));
 sg13g2_nand3_1 _12209_ (.B(\i_debug_uart_tx.fsm_state[1] ),
    .C(\i_debug_uart_tx.fsm_state[0] ),
    .A(net3723),
    .Y(_04429_));
 sg13g2_o21ai_1 _12210_ (.B1(net525),
    .Y(_04430_),
    .A1(_04385_),
    .A2(_04429_));
 sg13g2_a21oi_1 _12211_ (.A1(_01556_),
    .A2(_04428_),
    .Y(_00713_),
    .B1(_04430_));
 sg13g2_xnor2_1 _12212_ (.Y(_04431_),
    .A(\i_debug_uart_tx.fsm_state[3] ),
    .B(_04429_));
 sg13g2_o21ai_1 _12213_ (.B1(_04431_),
    .Y(_04432_),
    .A1(\i_debug_uart_tx.fsm_state[0] ),
    .A2(_04422_));
 sg13g2_a21oi_1 _12214_ (.A1(_03094_),
    .A2(_04385_),
    .Y(_04433_),
    .B1(_04432_));
 sg13g2_a21oi_1 _12215_ (.A1(net3794),
    .A2(_04385_),
    .Y(_04434_),
    .B1(_04433_));
 sg13g2_nor2_1 _12216_ (.A(net397),
    .B(net3795),
    .Y(_00714_));
 sg13g2_nor3_2 _12217_ (.A(net641),
    .B(_02077_),
    .C(_03071_),
    .Y(_04435_));
 sg13g2_and2_1 _12218_ (.A(net524),
    .B(_04435_),
    .X(_04436_));
 sg13g2_mux2_1 _12219_ (.A0(net3259),
    .A1(\data_to_write[8] ),
    .S(_04436_),
    .X(_00715_));
 sg13g2_xor2_1 _12220_ (.B(\i_spi.clock_count[3] ),
    .A(\i_spi.clock_divider[3] ),
    .X(_04437_));
 sg13g2_xor2_1 _12221_ (.B(\i_spi.clock_count[1] ),
    .A(\i_spi.clock_divider[1] ),
    .X(_04438_));
 sg13g2_xor2_1 _12222_ (.B(\i_spi.clock_count[0] ),
    .A(\i_spi.clock_divider[0] ),
    .X(_04439_));
 sg13g2_xor2_1 _12223_ (.B(\i_spi.clock_count[2] ),
    .A(\i_spi.clock_divider[2] ),
    .X(_04440_));
 sg13g2_nor4_2 _12224_ (.A(_04437_),
    .B(_04438_),
    .C(_04439_),
    .Y(_04441_),
    .D(_04440_));
 sg13g2_nand2b_1 _12225_ (.Y(_04442_),
    .B(net641),
    .A_N(_04441_));
 sg13g2_inv_1 _12226_ (.Y(_04443_),
    .A(_04442_));
 sg13g2_o21ai_1 _12227_ (.B1(net526),
    .Y(_04444_),
    .A1(net3658),
    .A2(_04443_));
 sg13g2_a21oi_1 _12228_ (.A1(net641),
    .A2(net3658),
    .Y(_00716_),
    .B1(_04444_));
 sg13g2_nand2_1 _12229_ (.Y(_04445_),
    .A(net646),
    .B(_04441_));
 sg13g2_nand2_2 _12230_ (.Y(_04446_),
    .A(net526),
    .B(_04445_));
 sg13g2_and3_1 _12231_ (.X(_04447_),
    .A(net641),
    .B(net3381),
    .C(net3658));
 sg13g2_a21oi_1 _12232_ (.A1(net641),
    .A2(\i_spi.clock_count[0] ),
    .Y(_04448_),
    .B1(net3381));
 sg13g2_nor3_1 _12233_ (.A(_04446_),
    .B(_04447_),
    .C(net3382),
    .Y(_00717_));
 sg13g2_nand2_1 _12234_ (.Y(_04449_),
    .A(\i_spi.clock_count[2] ),
    .B(_04447_));
 sg13g2_xnor2_1 _12235_ (.Y(_04450_),
    .A(net3793),
    .B(_04447_));
 sg13g2_nor2_1 _12236_ (.A(_04446_),
    .B(_04450_),
    .Y(_00718_));
 sg13g2_xor2_1 _12237_ (.B(_04449_),
    .A(net3765),
    .X(_04451_));
 sg13g2_nor2_1 _12238_ (.A(_04446_),
    .B(net3766),
    .Y(_00719_));
 sg13g2_nor2b_1 _12239_ (.A(_04435_),
    .B_N(_04445_),
    .Y(_04452_));
 sg13g2_nand3_1 _12240_ (.B(net641),
    .C(_04441_),
    .A(_01554_),
    .Y(_04453_));
 sg13g2_a21oi_1 _12241_ (.A1(\i_spi.read_latency ),
    .A2(_01555_),
    .Y(_04454_),
    .B1(_04453_));
 sg13g2_nor3_1 _12242_ (.A(net516),
    .B(_04452_),
    .C(_04454_),
    .Y(_04455_));
 sg13g2_nand2_1 _12243_ (.Y(_04456_),
    .A(net644),
    .B(net4));
 sg13g2_o21ai_1 _12244_ (.B1(_04456_),
    .Y(_04457_),
    .A1(_01511_),
    .A2(net642));
 sg13g2_mux2_1 _12245_ (.A0(net3653),
    .A1(_04457_),
    .S(_04455_),
    .X(_00720_));
 sg13g2_o21ai_1 _12246_ (.B1(_00204_),
    .Y(_04458_),
    .A1(_02077_),
    .A2(_03071_));
 sg13g2_inv_1 _12247_ (.Y(_04459_),
    .A(_04458_));
 sg13g2_o21ai_1 _12248_ (.B1(net526),
    .Y(_04460_),
    .A1(net641),
    .A2(_04459_));
 sg13g2_nor2_1 _12249_ (.A(_04443_),
    .B(_04459_),
    .Y(_04461_));
 sg13g2_nor4_2 _12250_ (.A(net3670),
    .B(\i_spi.bits_remaining[2] ),
    .C(\i_spi.bits_remaining[1] ),
    .Y(_04462_),
    .D(net3461));
 sg13g2_o21ai_1 _12251_ (.B1(net646),
    .Y(_04463_),
    .A1(_01554_),
    .A2(_04462_));
 sg13g2_nand2_1 _12252_ (.Y(_04464_),
    .A(_04461_),
    .B(_04463_));
 sg13g2_nand2_1 _12253_ (.Y(_04465_),
    .A(net3461),
    .B(_04464_));
 sg13g2_or2_1 _12254_ (.X(_04466_),
    .B(_04464_),
    .A(net3461));
 sg13g2_a21oi_1 _12255_ (.A1(_04465_),
    .A2(_04466_),
    .Y(_00721_),
    .B1(_04460_));
 sg13g2_xor2_1 _12256_ (.B(_04466_),
    .A(net3867),
    .X(_04467_));
 sg13g2_nor2_1 _12257_ (.A(_04460_),
    .B(_04467_),
    .Y(_00722_));
 sg13g2_or3_1 _12258_ (.A(net3703),
    .B(\i_spi.bits_remaining[1] ),
    .C(_04466_),
    .X(_04468_));
 sg13g2_o21ai_1 _12259_ (.B1(net3703),
    .Y(_04469_),
    .A1(\i_spi.bits_remaining[1] ),
    .A2(_04466_));
 sg13g2_a21oi_1 _12260_ (.A1(_04468_),
    .A2(net3704),
    .Y(_00723_),
    .B1(_04460_));
 sg13g2_nor2_1 _12261_ (.A(_00204_),
    .B(_04462_),
    .Y(_04470_));
 sg13g2_nor2_1 _12262_ (.A(_04464_),
    .B(_04470_),
    .Y(_04471_));
 sg13g2_a21oi_1 _12263_ (.A1(net3670),
    .A2(_04468_),
    .Y(_04472_),
    .B1(_04471_));
 sg13g2_nor2_1 _12264_ (.A(net397),
    .B(net3671),
    .Y(_00724_));
 sg13g2_nand2_1 _12265_ (.Y(_04473_),
    .A(_01554_),
    .B(_04462_));
 sg13g2_nand2_1 _12266_ (.Y(_04474_),
    .A(net641),
    .B(_04473_));
 sg13g2_nand2_1 _12267_ (.Y(_04475_),
    .A(_04442_),
    .B(_04474_));
 sg13g2_o21ai_1 _12268_ (.B1(net526),
    .Y(_04476_),
    .A1(_04435_),
    .A2(_04475_));
 sg13g2_inv_1 _12269_ (.Y(_00725_),
    .A(_04476_));
 sg13g2_mux2_1 _12270_ (.A0(net3161),
    .A1(\data_to_write[9] ),
    .S(_04436_),
    .X(_00726_));
 sg13g2_nand2b_1 _12271_ (.Y(_04477_),
    .B(_04474_),
    .A_N(_04452_));
 sg13g2_o21ai_1 _12272_ (.B1(net525),
    .Y(_04478_),
    .A1(_01706_),
    .A2(_04473_));
 sg13g2_a22oi_1 _12273_ (.Y(_04479_),
    .B1(_04478_),
    .B2(_04446_),
    .A2(_04477_),
    .A1(net3102));
 sg13g2_inv_1 _12274_ (.Y(_00727_),
    .A(net3103));
 sg13g2_nor2_1 _12275_ (.A(_04453_),
    .B(_04462_),
    .Y(_04480_));
 sg13g2_a21oi_1 _12276_ (.A1(net3333),
    .A2(_04452_),
    .Y(_04481_),
    .B1(_04480_));
 sg13g2_nor2_1 _12277_ (.A(net397),
    .B(net3334),
    .Y(_00728_));
 sg13g2_nand4_1 _12278_ (.B(\i_pwm.pwm_count[4] ),
    .C(\i_pwm.pwm_count[6] ),
    .A(\i_pwm.pwm_count[5] ),
    .Y(_04482_),
    .D(\i_pwm.pwm_count[7] ));
 sg13g2_nand2_1 _12279_ (.Y(_04483_),
    .A(\i_pwm.pwm_count[1] ),
    .B(\i_pwm.pwm_count[2] ));
 sg13g2_nor4_1 _12280_ (.A(\i_pwm.pwm_count[0] ),
    .B(_01619_),
    .C(_04482_),
    .D(_04483_),
    .Y(_04484_));
 sg13g2_or2_2 _12281_ (.X(_04485_),
    .B(_04484_),
    .A(net516));
 sg13g2_nor2_1 _12282_ (.A(_01708_),
    .B(_04485_),
    .Y(_00737_));
 sg13g2_xnor2_1 _12283_ (.Y(_04486_),
    .A(\i_pwm.pwm_count[0] ),
    .B(net3760));
 sg13g2_nor2_1 _12284_ (.A(_04485_),
    .B(net3761),
    .Y(_00738_));
 sg13g2_and3_1 _12285_ (.X(_04487_),
    .A(\i_pwm.pwm_count[0] ),
    .B(\i_pwm.pwm_count[1] ),
    .C(net3584));
 sg13g2_a21oi_1 _12286_ (.A1(\i_pwm.pwm_count[0] ),
    .A2(\i_pwm.pwm_count[1] ),
    .Y(_04488_),
    .B1(net3584));
 sg13g2_nor3_1 _12287_ (.A(_04485_),
    .B(_04487_),
    .C(net3585),
    .Y(_00739_));
 sg13g2_and2_1 _12288_ (.A(net3582),
    .B(_04487_),
    .X(_04489_));
 sg13g2_nor2_1 _12289_ (.A(net3582),
    .B(_04487_),
    .Y(_04490_));
 sg13g2_nor3_1 _12290_ (.A(_04485_),
    .B(_04489_),
    .C(net3583),
    .Y(_00740_));
 sg13g2_nor2_1 _12291_ (.A(net3785),
    .B(_04489_),
    .Y(_04491_));
 sg13g2_and2_1 _12292_ (.A(net3785),
    .B(_04489_),
    .X(_04492_));
 sg13g2_nor3_1 _12293_ (.A(_04485_),
    .B(_04491_),
    .C(_04492_),
    .Y(_00741_));
 sg13g2_nor2_1 _12294_ (.A(net3781),
    .B(_04492_),
    .Y(_04493_));
 sg13g2_and2_1 _12295_ (.A(net3781),
    .B(_04492_),
    .X(_04494_));
 sg13g2_nor3_1 _12296_ (.A(_04485_),
    .B(net3782),
    .C(_04494_),
    .Y(_00742_));
 sg13g2_and2_1 _12297_ (.A(net3807),
    .B(_04494_),
    .X(_04495_));
 sg13g2_nor2_1 _12298_ (.A(net3807),
    .B(_04494_),
    .Y(_04496_));
 sg13g2_nor3_1 _12299_ (.A(_04485_),
    .B(_04495_),
    .C(_04496_),
    .Y(_00743_));
 sg13g2_a21oi_1 _12300_ (.A1(net3892),
    .A2(_04495_),
    .Y(_04497_),
    .B1(_04485_));
 sg13g2_o21ai_1 _12301_ (.B1(_04497_),
    .Y(_04498_),
    .A1(net3892),
    .A2(_04495_));
 sg13g2_inv_1 _12302_ (.Y(_00744_),
    .A(_04498_));
 sg13g2_nor3_2 _12303_ (.A(_01495_),
    .B(\i_tinyqv.cpu.data_write_n[0] ),
    .C(net420),
    .Y(_04499_));
 sg13g2_a21oi_1 _12304_ (.A1(net301),
    .A2(_04499_),
    .Y(_04500_),
    .B1(net517));
 sg13g2_nor2_1 _12305_ (.A(\data_to_write[16] ),
    .B(net167),
    .Y(_04501_));
 sg13g2_a21oi_1 _12306_ (.A1(_01634_),
    .A2(net167),
    .Y(_00753_),
    .B1(_04501_));
 sg13g2_nor2_1 _12307_ (.A(\data_to_write[17] ),
    .B(net167),
    .Y(_04502_));
 sg13g2_a21oi_1 _12308_ (.A1(_01633_),
    .A2(net167),
    .Y(_00754_),
    .B1(_04502_));
 sg13g2_nor2_1 _12309_ (.A(\data_to_write[18] ),
    .B(net167),
    .Y(_04503_));
 sg13g2_a21oi_1 _12310_ (.A1(_01632_),
    .A2(net167),
    .Y(_00755_),
    .B1(_04503_));
 sg13g2_nand2_1 _12311_ (.Y(_04504_),
    .A(net3536),
    .B(net175));
 sg13g2_o21ai_1 _12312_ (.B1(_04504_),
    .Y(_00756_),
    .A1(_01496_),
    .A2(net175));
 sg13g2_nor2_1 _12313_ (.A(\data_to_write[20] ),
    .B(net172),
    .Y(_04505_));
 sg13g2_a21oi_1 _12314_ (.A1(_01631_),
    .A2(net172),
    .Y(_00757_),
    .B1(_04505_));
 sg13g2_nor2_1 _12315_ (.A(\data_to_write[21] ),
    .B(net172),
    .Y(_04506_));
 sg13g2_a21oi_1 _12316_ (.A1(_01630_),
    .A2(net172),
    .Y(_00758_),
    .B1(_04506_));
 sg13g2_nor2_1 _12317_ (.A(\data_to_write[22] ),
    .B(net172),
    .Y(_04507_));
 sg13g2_a21oi_1 _12318_ (.A1(_01629_),
    .A2(net172),
    .Y(_00759_),
    .B1(_04507_));
 sg13g2_nor2_1 _12319_ (.A(\data_to_write[23] ),
    .B(net172),
    .Y(_04508_));
 sg13g2_a21oi_1 _12320_ (.A1(_01628_),
    .A2(net172),
    .Y(_00760_),
    .B1(_04508_));
 sg13g2_nor2_1 _12321_ (.A(\data_to_write[24] ),
    .B(net173),
    .Y(_04509_));
 sg13g2_a21oi_1 _12322_ (.A1(_01627_),
    .A2(net173),
    .Y(_00761_),
    .B1(_04509_));
 sg13g2_nor2_1 _12323_ (.A(\data_to_write[25] ),
    .B(net173),
    .Y(_04510_));
 sg13g2_a21oi_1 _12324_ (.A1(_01626_),
    .A2(net173),
    .Y(_00762_),
    .B1(_04510_));
 sg13g2_mux2_1 _12325_ (.A0(net3792),
    .A1(net3862),
    .S(net174),
    .X(_00763_));
 sg13g2_mux2_1 _12326_ (.A0(\data_to_write[27] ),
    .A1(net3797),
    .S(net174),
    .X(_00764_));
 sg13g2_nor2_1 _12327_ (.A(\data_to_write[28] ),
    .B(net173),
    .Y(_04511_));
 sg13g2_a21oi_1 _12328_ (.A1(_01625_),
    .A2(net173),
    .Y(_00765_),
    .B1(_04511_));
 sg13g2_nor2_1 _12329_ (.A(\data_to_write[29] ),
    .B(net173),
    .Y(_04512_));
 sg13g2_a21oi_1 _12330_ (.A1(_01624_),
    .A2(net173),
    .Y(_00766_),
    .B1(_04512_));
 sg13g2_nor2_1 _12331_ (.A(\data_to_write[30] ),
    .B(net174),
    .Y(_04513_));
 sg13g2_a21oi_1 _12332_ (.A1(_01623_),
    .A2(net174),
    .Y(_00767_),
    .B1(_04513_));
 sg13g2_mux2_1 _12333_ (.A0(\data_to_write[31] ),
    .A1(net3775),
    .S(net174),
    .X(_00768_));
 sg13g2_nand4_1 _12334_ (.B(_02090_),
    .C(_03067_),
    .A(_02088_),
    .Y(_04514_),
    .D(_04499_));
 sg13g2_nand2b_1 _12335_ (.Y(_04515_),
    .B(\i_time.time_pulse ),
    .A_N(net3811));
 sg13g2_o21ai_1 _12336_ (.B1(net3812),
    .Y(_04516_),
    .A1(\i_time.mtime[0] ),
    .A2(\i_time.time_pulse ));
 sg13g2_nand2_1 _12337_ (.Y(_04517_),
    .A(net222),
    .B(_04499_));
 sg13g2_o21ai_1 _12338_ (.B1(net531),
    .Y(_04518_),
    .A1(\data_to_write[0] ),
    .A2(net110));
 sg13g2_a21oi_1 _12339_ (.A1(net269),
    .A2(net3813),
    .Y(_00774_),
    .B1(_04518_));
 sg13g2_nand3_1 _12340_ (.B(net4083),
    .C(\i_time.time_pulse ),
    .A(\i_time.mtime[1] ),
    .Y(_04519_));
 sg13g2_a21o_1 _12341_ (.A2(\i_time.time_pulse ),
    .A1(net4083),
    .B1(\i_time.mtime[1] ),
    .X(_04520_));
 sg13g2_nand2_1 _12342_ (.Y(_04521_),
    .A(_04519_),
    .B(net4084));
 sg13g2_o21ai_1 _12343_ (.B1(net521),
    .Y(_04522_),
    .A1(net601),
    .A2(net269));
 sg13g2_a21oi_1 _12344_ (.A1(net269),
    .A2(_04521_),
    .Y(_00775_),
    .B1(_04522_));
 sg13g2_nor2_2 _12345_ (.A(_01546_),
    .B(_04519_),
    .Y(_04523_));
 sg13g2_xnor2_1 _12346_ (.Y(_04524_),
    .A(_01546_),
    .B(_04519_));
 sg13g2_o21ai_1 _12347_ (.B1(net521),
    .Y(_04525_),
    .A1(net600),
    .A2(net270));
 sg13g2_a21oi_1 _12348_ (.A1(net269),
    .A2(_04524_),
    .Y(_00776_),
    .B1(_04525_));
 sg13g2_xnor2_1 _12349_ (.Y(_04526_),
    .A(net3880),
    .B(_04523_));
 sg13g2_o21ai_1 _12350_ (.B1(net518),
    .Y(_04527_),
    .A1(\data_to_write[3] ),
    .A2(net268));
 sg13g2_a21oi_1 _12351_ (.A1(net268),
    .A2(_04526_),
    .Y(_00777_),
    .B1(_04527_));
 sg13g2_nand3_1 _12352_ (.B(net3880),
    .C(_04523_),
    .A(net4082),
    .Y(_04528_));
 sg13g2_a21o_1 _12353_ (.A2(_04523_),
    .A1(net3880),
    .B1(net4082),
    .X(_04529_));
 sg13g2_nand2_1 _12354_ (.Y(_04530_),
    .A(_04528_),
    .B(_04529_));
 sg13g2_o21ai_1 _12355_ (.B1(net520),
    .Y(_04531_),
    .A1(net599),
    .A2(net268));
 sg13g2_a21oi_1 _12356_ (.A1(net267),
    .A2(_04530_),
    .Y(_00778_),
    .B1(_04531_));
 sg13g2_or2_1 _12357_ (.X(_04532_),
    .B(_04528_),
    .A(_01543_));
 sg13g2_xnor2_1 _12358_ (.Y(_04533_),
    .A(_01543_),
    .B(_04528_));
 sg13g2_o21ai_1 _12359_ (.B1(net518),
    .Y(_04534_),
    .A1(net598),
    .A2(net268));
 sg13g2_a21oi_1 _12360_ (.A1(net267),
    .A2(_04533_),
    .Y(_00779_),
    .B1(_04534_));
 sg13g2_nor2_1 _12361_ (.A(_01542_),
    .B(_04532_),
    .Y(_04535_));
 sg13g2_xnor2_1 _12362_ (.Y(_04536_),
    .A(_01542_),
    .B(_04532_));
 sg13g2_o21ai_1 _12363_ (.B1(net518),
    .Y(_04537_),
    .A1(net597),
    .A2(net267));
 sg13g2_a21oi_1 _12364_ (.A1(net267),
    .A2(_04536_),
    .Y(_00780_),
    .B1(_04537_));
 sg13g2_xnor2_1 _12365_ (.Y(_04538_),
    .A(net4015),
    .B(_04535_));
 sg13g2_o21ai_1 _12366_ (.B1(net518),
    .Y(_04539_),
    .A1(\data_to_write[7] ),
    .A2(net267));
 sg13g2_a21oi_1 _12367_ (.A1(net267),
    .A2(_04538_),
    .Y(_00781_),
    .B1(_04539_));
 sg13g2_nand3_1 _12368_ (.B(\i_time.mtime[7] ),
    .C(_04535_),
    .A(\i_time.mtime[8] ),
    .Y(_04540_));
 sg13g2_a21o_1 _12369_ (.A2(_04535_),
    .A1(net4015),
    .B1(net4080),
    .X(_04541_));
 sg13g2_nand2_1 _12370_ (.Y(_04542_),
    .A(_04540_),
    .B(_04541_));
 sg13g2_o21ai_1 _12371_ (.B1(net518),
    .Y(_04543_),
    .A1(\data_to_write[8] ),
    .A2(net267));
 sg13g2_a21oi_1 _12372_ (.A1(net267),
    .A2(_04542_),
    .Y(_00782_),
    .B1(_04543_));
 sg13g2_nor2_1 _12373_ (.A(_01541_),
    .B(_04540_),
    .Y(_04544_));
 sg13g2_xnor2_1 _12374_ (.Y(_04545_),
    .A(_01541_),
    .B(_04540_));
 sg13g2_o21ai_1 _12375_ (.B1(net521),
    .Y(_04546_),
    .A1(\data_to_write[9] ),
    .A2(net269));
 sg13g2_a21oi_1 _12376_ (.A1(net269),
    .A2(net4108),
    .Y(_00783_),
    .B1(_04546_));
 sg13g2_xnor2_1 _12377_ (.Y(_04547_),
    .A(net3995),
    .B(_04544_));
 sg13g2_o21ai_1 _12378_ (.B1(net521),
    .Y(_04548_),
    .A1(net3889),
    .A2(net269));
 sg13g2_a21oi_1 _12379_ (.A1(net110),
    .A2(_04547_),
    .Y(_00784_),
    .B1(_04548_));
 sg13g2_nand3_1 _12380_ (.B(\i_time.mtime[10] ),
    .C(_04544_),
    .A(\i_time.mtime[11] ),
    .Y(_04549_));
 sg13g2_a21o_1 _12381_ (.A2(_04544_),
    .A1(\i_time.mtime[10] ),
    .B1(net3976),
    .X(_04550_));
 sg13g2_nand2_1 _12382_ (.Y(_04551_),
    .A(_04549_),
    .B(net3977));
 sg13g2_o21ai_1 _12383_ (.B1(net522),
    .Y(_04552_),
    .A1(net3911),
    .A2(net271));
 sg13g2_a21oi_1 _12384_ (.A1(net110),
    .A2(_04551_),
    .Y(_00785_),
    .B1(_04552_));
 sg13g2_nor2_2 _12385_ (.A(_01539_),
    .B(_04549_),
    .Y(_04553_));
 sg13g2_xnor2_1 _12386_ (.Y(_04554_),
    .A(_01539_),
    .B(_04549_));
 sg13g2_o21ai_1 _12387_ (.B1(net521),
    .Y(_04555_),
    .A1(net3800),
    .A2(net269));
 sg13g2_a21oi_1 _12388_ (.A1(net110),
    .A2(net3944),
    .Y(_00786_),
    .B1(_04555_));
 sg13g2_xnor2_1 _12389_ (.Y(_04556_),
    .A(net3954),
    .B(_04553_));
 sg13g2_o21ai_1 _12390_ (.B1(net522),
    .Y(_04557_),
    .A1(net3835),
    .A2(net273));
 sg13g2_a21oi_1 _12391_ (.A1(net113),
    .A2(_04556_),
    .Y(_00787_),
    .B1(_04557_));
 sg13g2_nand3_1 _12392_ (.B(net3954),
    .C(_04553_),
    .A(net4018),
    .Y(_04558_));
 sg13g2_a21o_1 _12393_ (.A2(_04553_),
    .A1(net3954),
    .B1(net4018),
    .X(_04559_));
 sg13g2_nand2_1 _12394_ (.Y(_04560_),
    .A(_04558_),
    .B(_04559_));
 sg13g2_o21ai_1 _12395_ (.B1(net522),
    .Y(_04561_),
    .A1(net3882),
    .A2(net271));
 sg13g2_a21oi_1 _12396_ (.A1(net110),
    .A2(_04560_),
    .Y(_00788_),
    .B1(_04561_));
 sg13g2_nor2_1 _12397_ (.A(_01537_),
    .B(_04558_),
    .Y(_04562_));
 sg13g2_xnor2_1 _12398_ (.Y(_04563_),
    .A(_01537_),
    .B(_04558_));
 sg13g2_o21ai_1 _12399_ (.B1(net522),
    .Y(_04564_),
    .A1(net3873),
    .A2(net271));
 sg13g2_a21oi_1 _12400_ (.A1(net110),
    .A2(net4013),
    .Y(_00789_),
    .B1(_04564_));
 sg13g2_xnor2_1 _12401_ (.Y(_04565_),
    .A(net3984),
    .B(_04562_));
 sg13g2_o21ai_1 _12402_ (.B1(net522),
    .Y(_04566_),
    .A1(net3842),
    .A2(net271));
 sg13g2_a21oi_1 _12403_ (.A1(net110),
    .A2(_04565_),
    .Y(_00790_),
    .B1(_04566_));
 sg13g2_nand3_1 _12404_ (.B(\i_time.mtime[16] ),
    .C(_04562_),
    .A(net4044),
    .Y(_04567_));
 sg13g2_a21o_1 _12405_ (.A2(_04562_),
    .A1(net3984),
    .B1(net4044),
    .X(_04568_));
 sg13g2_nand2_1 _12406_ (.Y(_04569_),
    .A(_04567_),
    .B(_04568_));
 sg13g2_o21ai_1 _12407_ (.B1(net522),
    .Y(_04570_),
    .A1(net3909),
    .A2(net271));
 sg13g2_a21oi_1 _12408_ (.A1(net110),
    .A2(_04569_),
    .Y(_00791_),
    .B1(_04570_));
 sg13g2_nor2_2 _12409_ (.A(_01535_),
    .B(_04567_),
    .Y(_04571_));
 sg13g2_xnor2_1 _12410_ (.Y(_04572_),
    .A(_01535_),
    .B(_04567_));
 sg13g2_o21ai_1 _12411_ (.B1(net522),
    .Y(_04573_),
    .A1(net3920),
    .A2(net273));
 sg13g2_a21oi_1 _12412_ (.A1(net113),
    .A2(_04572_),
    .Y(_00792_),
    .B1(_04573_));
 sg13g2_xnor2_1 _12413_ (.Y(_04574_),
    .A(net3853),
    .B(_04571_));
 sg13g2_o21ai_1 _12414_ (.B1(net532),
    .Y(_04575_),
    .A1(net3771),
    .A2(net273));
 sg13g2_a21oi_1 _12415_ (.A1(net112),
    .A2(_04574_),
    .Y(_00793_),
    .B1(_04575_));
 sg13g2_nand3_1 _12416_ (.B(\i_time.mtime[19] ),
    .C(_04571_),
    .A(\i_time.mtime[20] ),
    .Y(_04576_));
 sg13g2_a21o_1 _12417_ (.A2(_04571_),
    .A1(net3853),
    .B1(net4075),
    .X(_04577_));
 sg13g2_nand2_1 _12418_ (.Y(_04578_),
    .A(_04576_),
    .B(_04577_));
 sg13g2_o21ai_1 _12419_ (.B1(net532),
    .Y(_04579_),
    .A1(net4061),
    .A2(net273));
 sg13g2_a21oi_1 _12420_ (.A1(net112),
    .A2(net4076),
    .Y(_00794_),
    .B1(_04579_));
 sg13g2_nor2_1 _12421_ (.A(_01533_),
    .B(_04576_),
    .Y(_04580_));
 sg13g2_xnor2_1 _12422_ (.Y(_04581_),
    .A(_01533_),
    .B(_04576_));
 sg13g2_o21ai_1 _12423_ (.B1(net532),
    .Y(_04582_),
    .A1(net4050),
    .A2(net273));
 sg13g2_a21oi_1 _12424_ (.A1(net112),
    .A2(net4068),
    .Y(_00795_),
    .B1(_04582_));
 sg13g2_xnor2_1 _12425_ (.Y(_04583_),
    .A(\i_time.mtime[22] ),
    .B(_04580_));
 sg13g2_o21ai_1 _12426_ (.B1(net532),
    .Y(_04584_),
    .A1(net4026),
    .A2(net272));
 sg13g2_a21oi_1 _12427_ (.A1(net111),
    .A2(_04583_),
    .Y(_00796_),
    .B1(_04584_));
 sg13g2_nand3_1 _12428_ (.B(\i_time.mtime[22] ),
    .C(_04580_),
    .A(\i_time.mtime[23] ),
    .Y(_04585_));
 sg13g2_a21o_1 _12429_ (.A2(_04580_),
    .A1(\i_time.mtime[22] ),
    .B1(\i_time.mtime[23] ),
    .X(_04586_));
 sg13g2_nand2_1 _12430_ (.Y(_04587_),
    .A(_04585_),
    .B(_04586_));
 sg13g2_o21ai_1 _12431_ (.B1(net532),
    .Y(_04588_),
    .A1(net4024),
    .A2(net272));
 sg13g2_a21oi_1 _12432_ (.A1(net112),
    .A2(_04587_),
    .Y(_00797_),
    .B1(_04588_));
 sg13g2_nor2_1 _12433_ (.A(_01532_),
    .B(_04585_),
    .Y(_04589_));
 sg13g2_xnor2_1 _12434_ (.Y(_04590_),
    .A(_01532_),
    .B(_04585_));
 sg13g2_o21ai_1 _12435_ (.B1(net532),
    .Y(_04591_),
    .A1(net3926),
    .A2(net272));
 sg13g2_a21oi_1 _12436_ (.A1(net111),
    .A2(net4030),
    .Y(_00798_),
    .B1(_04591_));
 sg13g2_xnor2_1 _12437_ (.Y(_04592_),
    .A(net4008),
    .B(_04589_));
 sg13g2_o21ai_1 _12438_ (.B1(net533),
    .Y(_04593_),
    .A1(net3971),
    .A2(net272));
 sg13g2_a21oi_1 _12439_ (.A1(net111),
    .A2(_04592_),
    .Y(_00799_),
    .B1(_04593_));
 sg13g2_nand3_1 _12440_ (.B(\i_time.mtime[25] ),
    .C(_04589_),
    .A(net3961),
    .Y(_04594_));
 sg13g2_a21o_1 _12441_ (.A2(_04589_),
    .A1(\i_time.mtime[25] ),
    .B1(net3961),
    .X(_04595_));
 sg13g2_nand2_1 _12442_ (.Y(_04596_),
    .A(_04594_),
    .B(net3962));
 sg13g2_o21ai_1 _12443_ (.B1(net532),
    .Y(_04597_),
    .A1(net3792),
    .A2(net272));
 sg13g2_a21oi_1 _12444_ (.A1(net111),
    .A2(_04596_),
    .Y(_00800_),
    .B1(_04597_));
 sg13g2_nor2_1 _12445_ (.A(_01529_),
    .B(_04594_),
    .Y(_04598_));
 sg13g2_xnor2_1 _12446_ (.Y(_04599_),
    .A(_01529_),
    .B(_04594_));
 sg13g2_o21ai_1 _12447_ (.B1(net533),
    .Y(_04600_),
    .A1(net3817),
    .A2(net272));
 sg13g2_a21oi_1 _12448_ (.A1(net111),
    .A2(net3960),
    .Y(_00801_),
    .B1(_04600_));
 sg13g2_xnor2_1 _12449_ (.Y(_04601_),
    .A(net4001),
    .B(_04598_));
 sg13g2_o21ai_1 _12450_ (.B1(net532),
    .Y(_04602_),
    .A1(net3951),
    .A2(net272));
 sg13g2_a21oi_1 _12451_ (.A1(net112),
    .A2(_04601_),
    .Y(_00802_),
    .B1(_04602_));
 sg13g2_nand3_1 _12452_ (.B(\i_time.mtime[28] ),
    .C(_04598_),
    .A(net3997),
    .Y(_04603_));
 sg13g2_a21o_1 _12453_ (.A2(_04598_),
    .A1(\i_time.mtime[28] ),
    .B1(net3997),
    .X(_04604_));
 sg13g2_nand2_1 _12454_ (.Y(_04605_),
    .A(_04603_),
    .B(net3998));
 sg13g2_o21ai_1 _12455_ (.B1(net533),
    .Y(_04606_),
    .A1(net3974),
    .A2(net272));
 sg13g2_a21oi_1 _12456_ (.A1(net111),
    .A2(_04605_),
    .Y(_00803_),
    .B1(_04606_));
 sg13g2_or2_1 _12457_ (.X(_04607_),
    .B(_04603_),
    .A(_01528_));
 sg13g2_xnor2_1 _12458_ (.Y(_04608_),
    .A(_01528_),
    .B(_04603_));
 sg13g2_o21ai_1 _12459_ (.B1(net533),
    .Y(_04609_),
    .A1(net3921),
    .A2(net273));
 sg13g2_a21oi_1 _12460_ (.A1(net111),
    .A2(net3929),
    .Y(_00804_),
    .B1(_04609_));
 sg13g2_xor2_1 _12461_ (.B(_04607_),
    .A(\i_time.mtime[31] ),
    .X(_04610_));
 sg13g2_o21ai_1 _12462_ (.B1(net533),
    .Y(_04611_),
    .A1(net3864),
    .A2(net273));
 sg13g2_a21oi_1 _12463_ (.A1(net111),
    .A2(_04610_),
    .Y(_00805_),
    .B1(_04611_));
 sg13g2_and2_1 _12464_ (.A(net525),
    .B(net662),
    .X(_00806_));
 sg13g2_and2_1 _12465_ (.A(net526),
    .B(net2846),
    .X(_00807_));
 sg13g2_nand2_1 _12466_ (.Y(_04612_),
    .A(net3478),
    .B(_03092_));
 sg13g2_nand4_1 _12467_ (.B(_03094_),
    .C(_04382_),
    .A(net525),
    .Y(_00809_),
    .D(_04612_));
 sg13g2_nand4_1 _12468_ (.B(net3945),
    .C(net637),
    .A(net3859),
    .Y(_04613_),
    .D(_02531_));
 sg13g2_and2_1 _12469_ (.A(net638),
    .B(_02532_),
    .X(_04614_));
 sg13g2_o21ai_1 _12470_ (.B1(_04614_),
    .Y(_04615_),
    .A1(net639),
    .A2(_02531_));
 sg13g2_o21ai_1 _12471_ (.B1(_04615_),
    .Y(_01058_),
    .A1(_01732_),
    .A2(_04613_));
 sg13g2_nor2_1 _12472_ (.A(net3510),
    .B(net545),
    .Y(_04616_));
 sg13g2_a21oi_1 _12473_ (.A1(_00318_),
    .A2(net545),
    .Y(_01059_),
    .B1(_04616_));
 sg13g2_nor2_1 _12474_ (.A(net3417),
    .B(net545),
    .Y(_04617_));
 sg13g2_a21oi_1 _12475_ (.A1(_00319_),
    .A2(net545),
    .Y(_01060_),
    .B1(_04617_));
 sg13g2_nor2_1 _12476_ (.A(net3312),
    .B(net545),
    .Y(_04618_));
 sg13g2_a21oi_1 _12477_ (.A1(_00320_),
    .A2(net544),
    .Y(_01061_),
    .B1(_04618_));
 sg13g2_nor2_1 _12478_ (.A(net3243),
    .B(net545),
    .Y(_04619_));
 sg13g2_a21oi_1 _12479_ (.A1(_00321_),
    .A2(net545),
    .Y(_01062_),
    .B1(_04619_));
 sg13g2_nor2_1 _12480_ (.A(net3504),
    .B(net542),
    .Y(_04620_));
 sg13g2_a21oi_1 _12481_ (.A1(_00322_),
    .A2(net543),
    .Y(_01063_),
    .B1(_04620_));
 sg13g2_nor2_1 _12482_ (.A(net3569),
    .B(net543),
    .Y(_04621_));
 sg13g2_a21oi_1 _12483_ (.A1(_00323_),
    .A2(net543),
    .Y(_01064_),
    .B1(_04621_));
 sg13g2_nor2_1 _12484_ (.A(net3563),
    .B(net542),
    .Y(_04622_));
 sg13g2_a21oi_1 _12485_ (.A1(_00324_),
    .A2(net542),
    .Y(_01065_),
    .B1(_04622_));
 sg13g2_nor2_1 _12486_ (.A(net3733),
    .B(net541),
    .Y(_04623_));
 sg13g2_a21oi_1 _12487_ (.A1(_00325_),
    .A2(net541),
    .Y(_01066_),
    .B1(_04623_));
 sg13g2_nor2_1 _12488_ (.A(net3273),
    .B(net539),
    .Y(_04624_));
 sg13g2_a21oi_1 _12489_ (.A1(_00326_),
    .A2(net539),
    .Y(_01067_),
    .B1(_04624_));
 sg13g2_nor2_1 _12490_ (.A(net3373),
    .B(net539),
    .Y(_04625_));
 sg13g2_a21oi_1 _12491_ (.A1(_00327_),
    .A2(net539),
    .Y(_01068_),
    .B1(_04625_));
 sg13g2_nor2_1 _12492_ (.A(net3281),
    .B(net539),
    .Y(_04626_));
 sg13g2_a21oi_1 _12493_ (.A1(_00328_),
    .A2(net539),
    .Y(_01069_),
    .B1(_04626_));
 sg13g2_nor2_1 _12494_ (.A(net3575),
    .B(net539),
    .Y(_04627_));
 sg13g2_a21oi_1 _12495_ (.A1(_00329_),
    .A2(net539),
    .Y(_01070_),
    .B1(_04627_));
 sg13g2_nor2_1 _12496_ (.A(net3697),
    .B(net542),
    .Y(_04628_));
 sg13g2_a21oi_1 _12497_ (.A1(_00330_),
    .A2(net542),
    .Y(_01071_),
    .B1(_04628_));
 sg13g2_nor2_1 _12498_ (.A(net3485),
    .B(net542),
    .Y(_04629_));
 sg13g2_a21oi_1 _12499_ (.A1(_00331_),
    .A2(net542),
    .Y(_01072_),
    .B1(_04629_));
 sg13g2_nor2_1 _12500_ (.A(net3348),
    .B(net542),
    .Y(_04630_));
 sg13g2_a21oi_1 _12501_ (.A1(_00332_),
    .A2(net543),
    .Y(_01073_),
    .B1(_04630_));
 sg13g2_nor2_1 _12502_ (.A(net3397),
    .B(net544),
    .Y(_04631_));
 sg13g2_a21oi_1 _12503_ (.A1(_00333_),
    .A2(net544),
    .Y(_01074_),
    .B1(_04631_));
 sg13g2_nor2_1 _12504_ (.A(net3477),
    .B(net544),
    .Y(_04632_));
 sg13g2_a21oi_1 _12505_ (.A1(_00334_),
    .A2(net544),
    .Y(_01075_),
    .B1(_04632_));
 sg13g2_nor2_1 _12506_ (.A(net3261),
    .B(net544),
    .Y(_04633_));
 sg13g2_a21oi_1 _12507_ (.A1(_00335_),
    .A2(net544),
    .Y(_01076_),
    .B1(_04633_));
 sg13g2_nor2_1 _12508_ (.A(net3323),
    .B(net540),
    .Y(_04634_));
 sg13g2_a21oi_1 _12509_ (.A1(_00336_),
    .A2(net541),
    .Y(_01077_),
    .B1(_04634_));
 sg13g2_nor2_1 _12510_ (.A(net3741),
    .B(net544),
    .Y(_04635_));
 sg13g2_a21oi_1 _12511_ (.A1(_00337_),
    .A2(net541),
    .Y(_01078_),
    .B1(_04635_));
 sg13g2_nor2_1 _12512_ (.A(net3639),
    .B(net540),
    .Y(_04636_));
 sg13g2_a21oi_1 _12513_ (.A1(_00338_),
    .A2(net540),
    .Y(_01079_),
    .B1(_04636_));
 sg13g2_nor2_1 _12514_ (.A(net3266),
    .B(net540),
    .Y(_04637_));
 sg13g2_a21oi_1 _12515_ (.A1(_00339_),
    .A2(net540),
    .Y(_01080_),
    .B1(_04637_));
 sg13g2_nor2_1 _12516_ (.A(net3283),
    .B(net540),
    .Y(_04638_));
 sg13g2_a21oi_1 _12517_ (.A1(_00340_),
    .A2(net540),
    .Y(_01081_),
    .B1(_04638_));
 sg13g2_mux2_1 _12518_ (.A0(net3493),
    .A1(\i_game.l_data.data_in[23] ),
    .S(net540),
    .X(_01082_));
 sg13g2_nand2_1 _12519_ (.Y(_04639_),
    .A(_02530_),
    .B(_04614_));
 sg13g2_and2_1 _12520_ (.A(_04613_),
    .B(_04639_),
    .X(_04640_));
 sg13g2_nor2_1 _12521_ (.A(_01729_),
    .B(_04614_),
    .Y(_04641_));
 sg13g2_nor2_1 _12522_ (.A(net4095),
    .B(_04641_),
    .Y(_04642_));
 sg13g2_nor2_1 _12523_ (.A(_04640_),
    .B(_04642_),
    .Y(_01083_));
 sg13g2_nor2_1 _12524_ (.A(_02311_),
    .B(net340),
    .Y(_04643_));
 sg13g2_and2_1 _12525_ (.A(_03018_),
    .B(_03045_),
    .X(_04644_));
 sg13g2_nand2_1 _12526_ (.Y(_04645_),
    .A(net353),
    .B(_04644_));
 sg13g2_nor2_1 _12527_ (.A(_04643_),
    .B(_04645_),
    .Y(_04646_));
 sg13g2_a21o_1 _12528_ (.A2(net340),
    .A1(_02311_),
    .B1(_01595_),
    .X(_04647_));
 sg13g2_nor3_1 _12529_ (.A(_04643_),
    .B(_04645_),
    .C(_04647_),
    .Y(_04648_));
 sg13g2_nor2_1 _12530_ (.A(net3759),
    .B(_04646_),
    .Y(_04649_));
 sg13g2_nor3_1 _12531_ (.A(_04124_),
    .B(_04648_),
    .C(_04649_),
    .Y(_01084_));
 sg13g2_nand2_2 _12532_ (.Y(_04650_),
    .A(_03041_),
    .B(_04644_));
 sg13g2_nor2_1 _12533_ (.A(_04643_),
    .B(_04650_),
    .Y(_04651_));
 sg13g2_nor3_1 _12534_ (.A(_04643_),
    .B(_04647_),
    .C(_04650_),
    .Y(_04652_));
 sg13g2_nand2_1 _12535_ (.Y(_04653_),
    .A(_03018_),
    .B(_03041_));
 sg13g2_nor2_1 _12536_ (.A(net3156),
    .B(_04651_),
    .Y(_04654_));
 sg13g2_nor3_1 _12537_ (.A(_04124_),
    .B(_04652_),
    .C(_04654_),
    .Y(_01085_));
 sg13g2_nor2_1 _12538_ (.A(_02365_),
    .B(net340),
    .Y(_04655_));
 sg13g2_o21ai_1 _12539_ (.B1(net4009),
    .Y(_04656_),
    .A1(_04650_),
    .A2(_04655_));
 sg13g2_o21ai_1 _12540_ (.B1(_02365_),
    .Y(_04657_),
    .A1(_01595_),
    .A2(net340));
 sg13g2_o21ai_1 _12541_ (.B1(_04656_),
    .Y(_04658_),
    .A1(_04650_),
    .A2(_04657_));
 sg13g2_nor2b_1 _12542_ (.A(net179),
    .B_N(_04658_),
    .Y(_01086_));
 sg13g2_nor2_1 _12543_ (.A(_02156_),
    .B(_04130_),
    .Y(_04659_));
 sg13g2_or2_1 _12544_ (.X(_04660_),
    .B(net340),
    .A(_02156_));
 sg13g2_o21ai_1 _12545_ (.B1(net3687),
    .Y(_04661_),
    .A1(_04650_),
    .A2(_04659_));
 sg13g2_nor2b_1 _12546_ (.A(_04653_),
    .B_N(_04151_),
    .Y(_04662_));
 sg13g2_and2_1 _12547_ (.A(_02156_),
    .B(_04662_),
    .X(_04663_));
 sg13g2_nand2_1 _12548_ (.Y(_04664_),
    .A(_04644_),
    .B(_04663_));
 sg13g2_a21oi_1 _12549_ (.A1(_04661_),
    .A2(_04664_),
    .Y(_01087_),
    .B1(_04124_));
 sg13g2_nor2_1 _12550_ (.A(_02248_),
    .B(net340),
    .Y(_04665_));
 sg13g2_or2_1 _12551_ (.X(_04666_),
    .B(net340),
    .A(_02248_));
 sg13g2_o21ai_1 _12552_ (.B1(net3659),
    .Y(_04667_),
    .A1(_04650_),
    .A2(_04665_));
 sg13g2_nand3_1 _12553_ (.B(_04644_),
    .C(_04662_),
    .A(_02248_),
    .Y(_04668_));
 sg13g2_a21oi_1 _12554_ (.A1(_04667_),
    .A2(_04668_),
    .Y(_01088_),
    .B1(net179));
 sg13g2_o21ai_1 _12555_ (.B1(_04125_),
    .Y(_04669_),
    .A1(_03047_),
    .A2(_04653_));
 sg13g2_o21ai_1 _12556_ (.B1(_04669_),
    .Y(_04670_),
    .A1(_03042_),
    .A2(_04660_));
 sg13g2_nor2b_1 _12557_ (.A(net3275),
    .B_N(\i_tinyqv.cpu.i_core.interrupt_req[1] ),
    .Y(_04671_));
 sg13g2_o21ai_1 _12558_ (.B1(_03042_),
    .Y(_04672_),
    .A1(net3763),
    .A2(_04671_));
 sg13g2_nor2_1 _12559_ (.A(_04663_),
    .B(_04670_),
    .Y(_04673_));
 sg13g2_a221oi_1 _12560_ (.B2(_04673_),
    .C1(net179),
    .B1(_04672_),
    .A1(_01526_),
    .Y(_01089_),
    .A2(_04670_));
 sg13g2_o21ai_1 _12561_ (.B1(_04669_),
    .Y(_04674_),
    .A1(_03042_),
    .A2(_04666_));
 sg13g2_nor2b_1 _12562_ (.A(net3773),
    .B_N(_04674_),
    .Y(_04675_));
 sg13g2_a21o_1 _12563_ (.A2(_01695_),
    .A1(\i_tinyqv.cpu.i_core.interrupt_req[0] ),
    .B1(net3773),
    .X(_04676_));
 sg13g2_a221oi_1 _12564_ (.B2(_03042_),
    .C1(_04674_),
    .B1(_04676_),
    .A1(_02248_),
    .Y(_04677_),
    .A2(_04662_));
 sg13g2_nor3_1 _12565_ (.A(net179),
    .B(_04675_),
    .C(_04677_),
    .Y(_01090_));
 sg13g2_nand2_1 _12566_ (.Y(_04678_),
    .A(net3502),
    .B(_03097_));
 sg13g2_nand4_1 _12567_ (.B(_03099_),
    .C(_04224_),
    .A(net537),
    .Y(_01091_),
    .D(_04678_));
 sg13g2_a21oi_1 _12568_ (.A1(_03066_),
    .A2(_03067_),
    .Y(_04679_),
    .B1(net516));
 sg13g2_nor2_1 _12569_ (.A(net529),
    .B(net3),
    .Y(_04680_));
 sg13g2_a21oi_1 _12570_ (.A1(_01511_),
    .A2(net529),
    .Y(_04681_),
    .B1(_04680_));
 sg13g2_mux2_1 _12571_ (.A0(_04681_),
    .A1(net4055),
    .S(_04679_),
    .X(_01092_));
 sg13g2_nor2_1 _12572_ (.A(net398),
    .B(_01685_),
    .Y(_01093_));
 sg13g2_and2_1 _12573_ (.A(net536),
    .B(net3099),
    .X(_01094_));
 sg13g2_and2_1 _12574_ (.A(net536),
    .B(net2913),
    .X(_01095_));
 sg13g2_nor3_1 _12575_ (.A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(\i_tinyqv.cpu.instr_write_offset[1] ),
    .C(_04364_),
    .Y(_04682_));
 sg13g2_mux2_1 _12576_ (.A0(net3488),
    .A1(\i_tinyqv.cpu.instr_data_in[2] ),
    .S(net39),
    .X(_01096_));
 sg13g2_nor2_1 _12577_ (.A(net3448),
    .B(net39),
    .Y(_04683_));
 sg13g2_a21oi_1 _12578_ (.A1(_01684_),
    .A2(net40),
    .Y(_01097_),
    .B1(_04683_));
 sg13g2_mux2_1 _12579_ (.A0(net3060),
    .A1(\i_tinyqv.cpu.instr_data_in[4] ),
    .S(net39),
    .X(_01098_));
 sg13g2_nor2_1 _12580_ (.A(net3108),
    .B(net37),
    .Y(_04684_));
 sg13g2_a21oi_1 _12581_ (.A1(_01671_),
    .A2(net37),
    .Y(_01099_),
    .B1(_04684_));
 sg13g2_mux2_1 _12582_ (.A0(net3121),
    .A1(\i_tinyqv.cpu.instr_data_in[6] ),
    .S(net39),
    .X(_01100_));
 sg13g2_mux2_1 _12583_ (.A0(net3070),
    .A1(\i_tinyqv.cpu.instr_data_in[7] ),
    .S(net36),
    .X(_01101_));
 sg13g2_nor2_1 _12584_ (.A(net3176),
    .B(net36),
    .Y(_04685_));
 sg13g2_a21oi_1 _12585_ (.A1(_00245_),
    .A2(net37),
    .Y(_01102_),
    .B1(_04685_));
 sg13g2_nor2_1 _12586_ (.A(net3054),
    .B(net38),
    .Y(_04686_));
 sg13g2_a21oi_1 _12587_ (.A1(_00246_),
    .A2(net38),
    .Y(_01103_),
    .B1(_04686_));
 sg13g2_nor2_1 _12588_ (.A(net3144),
    .B(net36),
    .Y(_04687_));
 sg13g2_a21oi_1 _12589_ (.A1(_00247_),
    .A2(net36),
    .Y(_01104_),
    .B1(_04687_));
 sg13g2_nor2_1 _12590_ (.A(net3097),
    .B(net37),
    .Y(_04688_));
 sg13g2_a21oi_1 _12591_ (.A1(_00248_),
    .A2(net37),
    .Y(_01105_),
    .B1(_04688_));
 sg13g2_nor2_1 _12592_ (.A(net3194),
    .B(net39),
    .Y(_04689_));
 sg13g2_a21oi_1 _12593_ (.A1(_00249_),
    .A2(net39),
    .Y(_01106_),
    .B1(_04689_));
 sg13g2_nor2_1 _12594_ (.A(net3125),
    .B(net37),
    .Y(_04690_));
 sg13g2_a21oi_1 _12595_ (.A1(_00250_),
    .A2(net37),
    .Y(_01107_),
    .B1(_04690_));
 sg13g2_nor2_1 _12596_ (.A(net3066),
    .B(net36),
    .Y(_04691_));
 sg13g2_a21oi_1 _12597_ (.A1(_00251_),
    .A2(net36),
    .Y(_01108_),
    .B1(_04691_));
 sg13g2_nor2_1 _12598_ (.A(net3158),
    .B(net36),
    .Y(_04692_));
 sg13g2_a21oi_1 _12599_ (.A1(_00252_),
    .A2(net36),
    .Y(_01109_),
    .B1(_04692_));
 sg13g2_mux2_1 _12600_ (.A0(\i_tinyqv.cpu.instr_data_in[2] ),
    .A1(net3717),
    .S(net18),
    .X(_01110_));
 sg13g2_nor2_1 _12601_ (.A(\i_tinyqv.cpu.instr_data_in[3] ),
    .B(net18),
    .Y(_04693_));
 sg13g2_a21oi_1 _12602_ (.A1(_01602_),
    .A2(net18),
    .Y(_01111_),
    .B1(_04693_));
 sg13g2_mux2_1 _12603_ (.A0(\i_tinyqv.cpu.instr_data_in[4] ),
    .A1(net3356),
    .S(net18),
    .X(_01112_));
 sg13g2_nand2_1 _12604_ (.Y(_04694_),
    .A(net2899),
    .B(net17));
 sg13g2_o21ai_1 _12605_ (.B1(_04694_),
    .Y(_01113_),
    .A1(_01671_),
    .A2(net17));
 sg13g2_mux2_1 _12606_ (.A0(\i_tinyqv.cpu.instr_data_in[6] ),
    .A1(net3340),
    .S(net18),
    .X(_01114_));
 sg13g2_mux2_1 _12607_ (.A0(\i_tinyqv.cpu.instr_data_in[7] ),
    .A1(net3303),
    .S(net17),
    .X(_01115_));
 sg13g2_nand2_1 _12608_ (.Y(_04695_),
    .A(net2880),
    .B(net19));
 sg13g2_o21ai_1 _12609_ (.B1(_04695_),
    .Y(_01116_),
    .A1(_00245_),
    .A2(net19));
 sg13g2_nand2_1 _12610_ (.Y(_04696_),
    .A(net2910),
    .B(net16));
 sg13g2_o21ai_1 _12611_ (.B1(_04696_),
    .Y(_01117_),
    .A1(_00246_),
    .A2(net16));
 sg13g2_nand2_1 _12612_ (.Y(_04697_),
    .A(net2974),
    .B(net16));
 sg13g2_o21ai_1 _12613_ (.B1(_04697_),
    .Y(_01118_),
    .A1(_00247_),
    .A2(net16));
 sg13g2_nand2_1 _12614_ (.Y(_04698_),
    .A(net2853),
    .B(net17));
 sg13g2_o21ai_1 _12615_ (.B1(_04698_),
    .Y(_01119_),
    .A1(_00248_),
    .A2(net17));
 sg13g2_nand2_1 _12616_ (.Y(_04699_),
    .A(net2897),
    .B(net18));
 sg13g2_o21ai_1 _12617_ (.B1(_04699_),
    .Y(_01120_),
    .A1(_00249_),
    .A2(net18));
 sg13g2_nand2_1 _12618_ (.Y(_04700_),
    .A(net2887),
    .B(net17));
 sg13g2_o21ai_1 _12619_ (.B1(_04700_),
    .Y(_01121_),
    .A1(_00250_),
    .A2(net17));
 sg13g2_nand2_1 _12620_ (.Y(_04701_),
    .A(net2920),
    .B(net16));
 sg13g2_o21ai_1 _12621_ (.B1(_04701_),
    .Y(_01122_),
    .A1(_00251_),
    .A2(net16));
 sg13g2_nand2_1 _12622_ (.Y(_04702_),
    .A(net2950),
    .B(net16));
 sg13g2_o21ai_1 _12623_ (.B1(_04702_),
    .Y(_01123_),
    .A1(_00252_),
    .A2(net16));
 sg13g2_a21oi_1 _12624_ (.A1(_01696_),
    .A2(_04641_),
    .Y(_01124_),
    .B1(_04640_));
 sg13g2_and3_2 _12625_ (.X(_04703_),
    .A(net526),
    .B(_04453_),
    .C(_04461_));
 sg13g2_nand2_1 _12626_ (.Y(_04704_),
    .A(net642),
    .B(net3653));
 sg13g2_o21ai_1 _12627_ (.B1(_04704_),
    .Y(_04705_),
    .A1(_01510_),
    .A2(net643));
 sg13g2_mux2_1 _12628_ (.A0(net3732),
    .A1(_04705_),
    .S(_04703_),
    .X(_01125_));
 sg13g2_nand2_1 _12629_ (.Y(_04706_),
    .A(net643),
    .B(\i_spi.data[1] ));
 sg13g2_o21ai_1 _12630_ (.B1(_04706_),
    .Y(_04707_),
    .A1(_01509_),
    .A2(net642));
 sg13g2_mux2_1 _12631_ (.A0(net3714),
    .A1(_04707_),
    .S(_04703_),
    .X(_01126_));
 sg13g2_nand2_1 _12632_ (.Y(_04708_),
    .A(net642),
    .B(\i_spi.data[2] ));
 sg13g2_o21ai_1 _12633_ (.B1(_04708_),
    .Y(_04709_),
    .A1(_01508_),
    .A2(net642));
 sg13g2_mux2_1 _12634_ (.A0(net3680),
    .A1(_04709_),
    .S(_04703_),
    .X(_01127_));
 sg13g2_nand2_1 _12635_ (.Y(_04710_),
    .A(net642),
    .B(net3680));
 sg13g2_o21ai_1 _12636_ (.B1(_04710_),
    .Y(_04711_),
    .A1(_01507_),
    .A2(net645));
 sg13g2_mux2_1 _12637_ (.A0(net3691),
    .A1(_04711_),
    .S(_04703_),
    .X(_01128_));
 sg13g2_nand2_1 _12638_ (.Y(_04712_),
    .A(net645),
    .B(\i_spi.data[4] ));
 sg13g2_o21ai_1 _12639_ (.B1(_04712_),
    .Y(_04713_),
    .A1(_01506_),
    .A2(net645));
 sg13g2_mux2_1 _12640_ (.A0(net3531),
    .A1(_04713_),
    .S(_04703_),
    .X(_01129_));
 sg13g2_nand2_1 _12641_ (.Y(_04714_),
    .A(net642),
    .B(net3531));
 sg13g2_o21ai_1 _12642_ (.B1(_04714_),
    .Y(_04715_),
    .A1(_01505_),
    .A2(net642));
 sg13g2_mux2_1 _12643_ (.A0(net3816),
    .A1(_04715_),
    .S(_04703_),
    .X(_01130_));
 sg13g2_nand2_1 _12644_ (.Y(_04716_),
    .A(net643),
    .B(\i_spi.data[6] ));
 sg13g2_o21ai_1 _12645_ (.B1(_04716_),
    .Y(_04717_),
    .A1(_01504_),
    .A2(net643));
 sg13g2_mux2_1 _12646_ (.A0(net3285),
    .A1(_04717_),
    .S(_04703_),
    .X(_01131_));
 sg13g2_nor2_2 _12647_ (.A(net347),
    .B(_03838_),
    .Y(_04718_));
 sg13g2_a22oi_1 _12648_ (.Y(_04719_),
    .B1(_04718_),
    .B2(net3840),
    .A2(net331),
    .A1(net3887));
 sg13g2_nor2_1 _12649_ (.A(net508),
    .B(_04719_),
    .Y(_01132_));
 sg13g2_a22oi_1 _12650_ (.Y(_04720_),
    .B1(_04718_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .A2(net331),
    .A1(net3553));
 sg13g2_nor2_1 _12651_ (.A(net508),
    .B(net3554),
    .Y(_01133_));
 sg13g2_a22oi_1 _12652_ (.Y(_04721_),
    .B1(_04718_),
    .B2(net3591),
    .A2(net331),
    .A1(net637));
 sg13g2_nor2_1 _12653_ (.A(net508),
    .B(_04721_),
    .Y(_01134_));
 sg13g2_a22oi_1 _12654_ (.Y(_04722_),
    .B1(_04718_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .A2(_03838_),
    .A1(net3206));
 sg13g2_nor2_1 _12655_ (.A(net508),
    .B(net3207),
    .Y(_01135_));
 sg13g2_nor2_2 _12656_ (.A(net647),
    .B(net331),
    .Y(_04723_));
 sg13g2_nor2_1 _12657_ (.A(net2389),
    .B(net261),
    .Y(_04724_));
 sg13g2_nand2_1 _12658_ (.Y(_04725_),
    .A(_01648_),
    .B(net341));
 sg13g2_o21ai_1 _12659_ (.B1(_04725_),
    .Y(_04726_),
    .A1(\i_tinyqv.cpu.i_core.mepc[0] ),
    .A2(net341));
 sg13g2_a21oi_1 _12660_ (.A1(net261),
    .A2(_04726_),
    .Y(_01136_),
    .B1(_04724_));
 sg13g2_nor2_1 _12661_ (.A(net4011),
    .B(net261),
    .Y(_04727_));
 sg13g2_nand2b_1 _12662_ (.Y(_04728_),
    .B(net341),
    .A_N(\i_tinyqv.cpu.i_core.i_shift.a[5] ));
 sg13g2_o21ai_1 _12663_ (.B1(_04728_),
    .Y(_04729_),
    .A1(\i_tinyqv.cpu.i_core.mepc[1] ),
    .A2(net341));
 sg13g2_a21oi_1 _12664_ (.A1(net261),
    .A2(_04729_),
    .Y(_01137_),
    .B1(_04727_));
 sg13g2_mux2_2 _12665_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[2] ),
    .S(net347),
    .X(_04730_));
 sg13g2_mux2_1 _12666_ (.A0(net4017),
    .A1(_04730_),
    .S(net261),
    .X(_01138_));
 sg13g2_nor2_1 _12667_ (.A(_01683_),
    .B(net341),
    .Y(_04731_));
 sg13g2_a21oi_2 _12668_ (.B1(_04731_),
    .Y(_04732_),
    .A2(net344),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[7] ));
 sg13g2_nor2_1 _12669_ (.A(net4112),
    .B(net261),
    .Y(_04733_));
 sg13g2_a21oi_2 _12670_ (.B1(_04733_),
    .Y(_01139_),
    .A2(_04732_),
    .A1(net261));
 sg13g2_nor2_1 _12671_ (.A(\addr[4] ),
    .B(net261),
    .Y(_04734_));
 sg13g2_nand2b_1 _12672_ (.Y(_04735_),
    .B(net344),
    .A_N(\i_tinyqv.cpu.i_core.i_shift.a[8] ));
 sg13g2_o21ai_1 _12673_ (.B1(_04735_),
    .Y(_04736_),
    .A1(\i_tinyqv.cpu.i_core.mepc[4] ),
    .A2(net341));
 sg13g2_a21oi_1 _12674_ (.A1(_04723_),
    .A2(_04736_),
    .Y(_01140_),
    .B1(_04734_));
 sg13g2_nor2_1 _12675_ (.A(net3987),
    .B(net263),
    .Y(_04737_));
 sg13g2_nand2b_1 _12676_ (.Y(_04738_),
    .B(net343),
    .A_N(\i_tinyqv.cpu.i_core.i_shift.a[9] ));
 sg13g2_o21ai_1 _12677_ (.B1(_04738_),
    .Y(_04739_),
    .A1(\i_tinyqv.cpu.i_core.mepc[5] ),
    .A2(net343));
 sg13g2_a21oi_1 _12678_ (.A1(net263),
    .A2(_04739_),
    .Y(_01141_),
    .B1(_04737_));
 sg13g2_nor2_1 _12679_ (.A(net4088),
    .B(net263),
    .Y(_04740_));
 sg13g2_nand2b_1 _12680_ (.Y(_04741_),
    .B(net343),
    .A_N(\i_tinyqv.cpu.i_core.i_shift.a[10] ));
 sg13g2_o21ai_1 _12681_ (.B1(_04741_),
    .Y(_04742_),
    .A1(\i_tinyqv.cpu.i_core.mepc[6] ),
    .A2(net342));
 sg13g2_a21oi_1 _12682_ (.A1(net263),
    .A2(_04742_),
    .Y(_01142_),
    .B1(_04740_));
 sg13g2_and2_1 _12683_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .B(net343),
    .X(_04743_));
 sg13g2_a21oi_2 _12684_ (.B1(_04743_),
    .Y(_04744_),
    .A2(net347),
    .A1(\i_tinyqv.cpu.i_core.mepc[7] ));
 sg13g2_nor2_1 _12685_ (.A(net3329),
    .B(net263),
    .Y(_04745_));
 sg13g2_a21oi_1 _12686_ (.A1(net263),
    .A2(_04744_),
    .Y(_01143_),
    .B1(_04745_));
 sg13g2_nor2_1 _12687_ (.A(net3507),
    .B(net263),
    .Y(_04746_));
 sg13g2_nand2b_1 _12688_ (.Y(_04747_),
    .B(net343),
    .A_N(\i_tinyqv.cpu.i_core.i_shift.a[12] ));
 sg13g2_o21ai_1 _12689_ (.B1(_04747_),
    .Y(_04748_),
    .A1(net3561),
    .A2(net343));
 sg13g2_a21oi_1 _12690_ (.A1(net263),
    .A2(_04748_),
    .Y(_01144_),
    .B1(_04746_));
 sg13g2_and2_1 _12691_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .B(net342),
    .X(_04749_));
 sg13g2_a21oi_2 _12692_ (.B1(_04749_),
    .Y(_04750_),
    .A2(net346),
    .A1(net3543));
 sg13g2_nor2_1 _12693_ (.A(net3635),
    .B(net264),
    .Y(_04751_));
 sg13g2_a21oi_1 _12694_ (.A1(net264),
    .A2(_04750_),
    .Y(_01145_),
    .B1(_04751_));
 sg13g2_nor2_1 _12695_ (.A(net3716),
    .B(net342),
    .Y(_04752_));
 sg13g2_a21oi_2 _12696_ (.B1(_04752_),
    .Y(_04753_),
    .A2(net342),
    .A1(_01657_));
 sg13g2_mux2_1 _12697_ (.A0(net3712),
    .A1(_04753_),
    .S(net264),
    .X(_01146_));
 sg13g2_mux2_2 _12698_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[15] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[11] ),
    .S(net345),
    .X(_04754_));
 sg13g2_mux2_1 _12699_ (.A0(net3604),
    .A1(_04754_),
    .S(net264),
    .X(_01147_));
 sg13g2_mux2_2 _12700_ (.A0(net3439),
    .A1(\i_tinyqv.cpu.i_core.mepc[12] ),
    .S(net346),
    .X(_04755_));
 sg13g2_nand2_1 _12701_ (.Y(_04756_),
    .A(net265),
    .B(_04755_));
 sg13g2_o21ai_1 _12702_ (.B1(_04756_),
    .Y(_01148_),
    .A1(_01613_),
    .A2(net264));
 sg13g2_nor2_1 _12703_ (.A(net3710),
    .B(net264),
    .Y(_04757_));
 sg13g2_nand2b_1 _12704_ (.Y(_04758_),
    .B(net342),
    .A_N(\i_tinyqv.cpu.i_core.i_shift.a[17] ));
 sg13g2_o21ai_1 _12705_ (.B1(_04758_),
    .Y(_04759_),
    .A1(\i_tinyqv.cpu.i_core.mepc[13] ),
    .A2(net343));
 sg13g2_a21oi_1 _12706_ (.A1(net264),
    .A2(_04759_),
    .Y(_01149_),
    .B1(_04757_));
 sg13g2_mux2_2 _12707_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .A1(net3529),
    .S(net346),
    .X(_04760_));
 sg13g2_mux2_1 _12708_ (.A0(net3803),
    .A1(_04760_),
    .S(net264),
    .X(_01150_));
 sg13g2_and2_1 _12709_ (.A(net3465),
    .B(net342),
    .X(_04761_));
 sg13g2_a21oi_2 _12710_ (.B1(_04761_),
    .Y(_04762_),
    .A2(net345),
    .A1(\i_tinyqv.cpu.i_core.mepc[15] ));
 sg13g2_nor2_1 _12711_ (.A(net3616),
    .B(net265),
    .Y(_04763_));
 sg13g2_a21oi_1 _12712_ (.A1(net265),
    .A2(_04762_),
    .Y(_01151_),
    .B1(_04763_));
 sg13g2_mux2_2 _12713_ (.A0(net3405),
    .A1(net3540),
    .S(net345),
    .X(_04764_));
 sg13g2_mux2_1 _12714_ (.A0(net3570),
    .A1(_04764_),
    .S(net265),
    .X(_01152_));
 sg13g2_nor2_1 _12715_ (.A(net3573),
    .B(net262),
    .Y(_04765_));
 sg13g2_nand2b_1 _12716_ (.Y(_04766_),
    .B(net342),
    .A_N(\i_tinyqv.cpu.i_core.i_shift.a[21] ));
 sg13g2_o21ai_1 _12717_ (.B1(_04766_),
    .Y(_04767_),
    .A1(\i_tinyqv.cpu.i_core.mepc[17] ),
    .A2(net342));
 sg13g2_a21oi_1 _12718_ (.A1(net262),
    .A2(_04767_),
    .Y(_01153_),
    .B1(_04765_));
 sg13g2_mux2_2 _12719_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[18] ),
    .S(net346),
    .X(_04768_));
 sg13g2_mux2_1 _12720_ (.A0(net3319),
    .A1(net3565),
    .S(net266),
    .X(_01154_));
 sg13g2_mux2_2 _12721_ (.A0(net4134),
    .A1(net3425),
    .S(net345),
    .X(_04769_));
 sg13g2_mux2_1 _12722_ (.A0(net3321),
    .A1(_04769_),
    .S(net262),
    .X(_01155_));
 sg13g2_mux2_2 _12723_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[20] ),
    .S(net345),
    .X(_04770_));
 sg13g2_mux2_1 _12724_ (.A0(net3496),
    .A1(_04770_),
    .S(net266),
    .X(_01156_));
 sg13g2_mux2_2 _12725_ (.A0(net3850),
    .A1(\i_tinyqv.cpu.i_core.mepc[21] ),
    .S(net345),
    .X(_04771_));
 sg13g2_nand2_1 _12726_ (.Y(_04772_),
    .A(net262),
    .B(_04771_));
 sg13g2_o21ai_1 _12727_ (.B1(_04772_),
    .Y(_01157_),
    .A1(_01615_),
    .A2(net262));
 sg13g2_mux2_2 _12728_ (.A0(net3538),
    .A1(\i_tinyqv.cpu.i_core.mepc[22] ),
    .S(net345),
    .X(_04773_));
 sg13g2_nand2_1 _12729_ (.Y(_04774_),
    .A(net262),
    .B(_04773_));
 sg13g2_o21ai_1 _12730_ (.B1(_04774_),
    .Y(_01158_),
    .A1(_01614_),
    .A2(net262));
 sg13g2_mux2_2 _12731_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[23] ),
    .S(net345),
    .X(_04775_));
 sg13g2_mux2_1 _12732_ (.A0(net3295),
    .A1(_04775_),
    .S(net262),
    .X(_01159_));
 sg13g2_nor3_1 _12733_ (.A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(_01598_),
    .C(_04364_),
    .Y(_04776_));
 sg13g2_mux2_1 _12734_ (.A0(net3418),
    .A1(\i_tinyqv.cpu.instr_data_in[2] ),
    .S(net35),
    .X(_01160_));
 sg13g2_nor2_1 _12735_ (.A(net3463),
    .B(net33),
    .Y(_04777_));
 sg13g2_a21oi_1 _12736_ (.A1(_01684_),
    .A2(net33),
    .Y(_01161_),
    .B1(_04777_));
 sg13g2_mux2_1 _12737_ (.A0(net3056),
    .A1(\i_tinyqv.cpu.instr_data_in[4] ),
    .S(net35),
    .X(_01162_));
 sg13g2_nor2_1 _12738_ (.A(net3197),
    .B(net31),
    .Y(_04778_));
 sg13g2_a21oi_1 _12739_ (.A1(_01671_),
    .A2(net31),
    .Y(_01163_),
    .B1(_04778_));
 sg13g2_mux2_1 _12740_ (.A0(net3058),
    .A1(\i_tinyqv.cpu.instr_data_in[6] ),
    .S(net35),
    .X(_01164_));
 sg13g2_mux2_1 _12741_ (.A0(net3068),
    .A1(\i_tinyqv.cpu.instr_data_in[7] ),
    .S(net34),
    .X(_01165_));
 sg13g2_nor2_1 _12742_ (.A(net3079),
    .B(net32),
    .Y(_04779_));
 sg13g2_a21oi_1 _12743_ (.A1(_00245_),
    .A2(net32),
    .Y(_01166_),
    .B1(_04779_));
 sg13g2_nor2_1 _12744_ (.A(net3017),
    .B(net32),
    .Y(_04780_));
 sg13g2_a21oi_1 _12745_ (.A1(_00246_),
    .A2(net32),
    .Y(_01167_),
    .B1(_04780_));
 sg13g2_nor2_1 _12746_ (.A(net3128),
    .B(net31),
    .Y(_04781_));
 sg13g2_a21oi_1 _12747_ (.A1(_00247_),
    .A2(net31),
    .Y(_01168_),
    .B1(_04781_));
 sg13g2_nor2_1 _12748_ (.A(net3147),
    .B(net32),
    .Y(_04782_));
 sg13g2_a21oi_1 _12749_ (.A1(_00248_),
    .A2(net32),
    .Y(_01169_),
    .B1(_04782_));
 sg13g2_nor2_1 _12750_ (.A(net3118),
    .B(net35),
    .Y(_04783_));
 sg13g2_a21oi_1 _12751_ (.A1(_00249_),
    .A2(net35),
    .Y(_01170_),
    .B1(_04783_));
 sg13g2_nor2_1 _12752_ (.A(net3033),
    .B(net32),
    .Y(_04784_));
 sg13g2_a21oi_1 _12753_ (.A1(_00250_),
    .A2(net32),
    .Y(_01171_),
    .B1(_04784_));
 sg13g2_nor2_1 _12754_ (.A(net3150),
    .B(net31),
    .Y(_04785_));
 sg13g2_a21oi_1 _12755_ (.A1(_00251_),
    .A2(net31),
    .Y(_01172_),
    .B1(_04785_));
 sg13g2_nor2_1 _12756_ (.A(net3189),
    .B(net31),
    .Y(_04786_));
 sg13g2_a21oi_1 _12757_ (.A1(_00252_),
    .A2(net31),
    .Y(_01173_),
    .B1(_04786_));
 sg13g2_o21ai_1 _12758_ (.B1(_02842_),
    .Y(_04787_),
    .A1(_02828_),
    .A2(net406));
 sg13g2_nand2_1 _12759_ (.Y(_04788_),
    .A(net3737),
    .B(net325));
 sg13g2_o21ai_1 _12760_ (.B1(_04788_),
    .Y(_01174_),
    .A1(_01648_),
    .A2(net325));
 sg13g2_mux2_1 _12761_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .A1(net3923),
    .S(net325),
    .X(_01175_));
 sg13g2_mux2_1 _12762_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .A1(net3918),
    .S(_04787_),
    .X(_01176_));
 sg13g2_mux2_1 _12763_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .A1(net3912),
    .S(net325),
    .X(_01177_));
 sg13g2_nor2_1 _12764_ (.A(net4035),
    .B(net325),
    .Y(_04789_));
 sg13g2_a21oi_1 _12765_ (.A1(_01648_),
    .A2(net325),
    .Y(_01178_),
    .B1(_04789_));
 sg13g2_mux2_1 _12766_ (.A0(net4064),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .S(net326),
    .X(_01179_));
 sg13g2_mux2_1 _12767_ (.A0(net3964),
    .A1(net4066),
    .S(net327),
    .X(_01180_));
 sg13g2_mux2_1 _12768_ (.A0(net4071),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .S(net327),
    .X(_01181_));
 sg13g2_mux2_1 _12769_ (.A0(net4019),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .S(net327),
    .X(_01182_));
 sg13g2_mux2_1 _12770_ (.A0(net4037),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .S(net327),
    .X(_01183_));
 sg13g2_nand2_1 _12771_ (.Y(_04790_),
    .A(net3964),
    .B(net328));
 sg13g2_o21ai_1 _12772_ (.B1(_04790_),
    .Y(_01184_),
    .A1(_01657_),
    .A2(net328));
 sg13g2_mux2_1 _12773_ (.A0(net3952),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .S(net328),
    .X(_01185_));
 sg13g2_mux2_1 _12774_ (.A0(net3439),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .S(net329),
    .X(_01186_));
 sg13g2_mux2_1 _12775_ (.A0(net3684),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .S(net330),
    .X(_01187_));
 sg13g2_nor2_1 _12776_ (.A(net3407),
    .B(net330),
    .Y(_04791_));
 sg13g2_a21oi_1 _12777_ (.A1(_01657_),
    .A2(net330),
    .Y(_01188_),
    .B1(_04791_));
 sg13g2_mux2_1 _12778_ (.A0(net3465),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[15] ),
    .S(net328),
    .X(_01189_));
 sg13g2_mux2_1 _12779_ (.A0(net3405),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .S(net328),
    .X(_01190_));
 sg13g2_mux2_1 _12780_ (.A0(net3668),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .S(net330),
    .X(_01191_));
 sg13g2_mux2_1 _12781_ (.A0(net3629),
    .A1(net3407),
    .S(net328),
    .X(_01192_));
 sg13g2_mux2_1 _12782_ (.A0(net3515),
    .A1(net3465),
    .S(net328),
    .X(_01193_));
 sg13g2_mux2_1 _12783_ (.A0(net3480),
    .A1(net3405),
    .S(net329),
    .X(_01194_));
 sg13g2_mux2_1 _12784_ (.A0(net3672),
    .A1(net3668),
    .S(net328),
    .X(_01195_));
 sg13g2_mux2_1 _12785_ (.A0(net3538),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .S(net327),
    .X(_01196_));
 sg13g2_mux2_1 _12786_ (.A0(net3692),
    .A1(net3515),
    .S(net327),
    .X(_01197_));
 sg13g2_mux2_1 _12787_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .A1(net3480),
    .S(net327),
    .X(_01198_));
 sg13g2_mux2_1 _12788_ (.A0(net3833),
    .A1(net3672),
    .S(net327),
    .X(_01199_));
 sg13g2_mux2_1 _12789_ (.A0(net3591),
    .A1(net3538),
    .S(net326),
    .X(_01200_));
 sg13g2_mux2_1 _12790_ (.A0(net3750),
    .A1(net3692),
    .S(net326),
    .X(_01201_));
 sg13g2_and2_1 _12791_ (.A(net406),
    .B(_03836_),
    .X(_04792_));
 sg13g2_nand2_1 _12792_ (.Y(_04793_),
    .A(net406),
    .B(_03836_));
 sg13g2_nand2_2 _12793_ (.Y(_04794_),
    .A(_02162_),
    .B(_02507_));
 sg13g2_a21o_1 _12794_ (.A2(_04793_),
    .A1(_02388_),
    .B1(_04794_),
    .X(_04795_));
 sg13g2_a21oi_1 _12795_ (.A1(_03357_),
    .A2(_04792_),
    .Y(_04796_),
    .B1(_04795_));
 sg13g2_nand2b_1 _12796_ (.Y(_04797_),
    .B(_04794_),
    .A_N(_02365_));
 sg13g2_nand2b_2 _12797_ (.Y(_04798_),
    .B(_03459_),
    .A_N(net326));
 sg13g2_nand2b_1 _12798_ (.Y(_04799_),
    .B(_04797_),
    .A_N(_04798_));
 sg13g2_a22oi_1 _12799_ (.Y(_04800_),
    .B1(net326),
    .B2(net3591),
    .A2(_04099_),
    .A1(net3957));
 sg13g2_o21ai_1 _12800_ (.B1(_04800_),
    .Y(_01202_),
    .A1(_04796_),
    .A2(_04799_));
 sg13g2_nand2b_1 _12801_ (.Y(_04801_),
    .B(_04792_),
    .A_N(_03752_));
 sg13g2_a21oi_1 _12802_ (.A1(_02337_),
    .A2(_04793_),
    .Y(_04802_),
    .B1(_04794_));
 sg13g2_a22oi_1 _12803_ (.Y(_04803_),
    .B1(_04801_),
    .B2(_04802_),
    .A2(_04794_),
    .A1(_02311_));
 sg13g2_nor3_1 _12804_ (.A(net4042),
    .B(net334),
    .C(net326),
    .Y(_04804_));
 sg13g2_a21oi_1 _12805_ (.A1(net3750),
    .A2(net325),
    .Y(_04805_),
    .B1(_04804_));
 sg13g2_o21ai_1 _12806_ (.B1(_04805_),
    .Y(_01203_),
    .A1(_04798_),
    .A2(_04803_));
 sg13g2_nor3_1 _12807_ (.A(net3897),
    .B(net647),
    .C(net38),
    .Y(_04806_));
 sg13g2_a21oi_1 _12808_ (.A1(_01660_),
    .A2(net38),
    .Y(_01204_),
    .B1(_04806_));
 sg13g2_nor3_1 _12809_ (.A(net3731),
    .B(net647),
    .C(net39),
    .Y(_04807_));
 sg13g2_a21oi_1 _12810_ (.A1(_01669_),
    .A2(net39),
    .Y(_01205_),
    .B1(_04807_));
 sg13g2_nand2_1 _12811_ (.Y(_04808_),
    .A(net3508),
    .B(net455));
 sg13g2_o21ai_1 _12812_ (.B1(_04808_),
    .Y(_01206_),
    .A1(_01659_),
    .A2(net455));
 sg13g2_mux2_1 _12813_ (.A0(net3810),
    .A1(net3700),
    .S(net455),
    .X(_01207_));
 sg13g2_mux2_1 _12814_ (.A0(\i_tinyqv.cpu.i_core.mepc[2] ),
    .A1(net3623),
    .S(net453),
    .X(_01208_));
 sg13g2_nand2_1 _12815_ (.Y(_04809_),
    .A(net3719),
    .B(net455));
 sg13g2_o21ai_1 _12816_ (.B1(_04809_),
    .Y(_01209_),
    .A1(_01683_),
    .A2(net455));
 sg13g2_mux2_1 _12817_ (.A0(net3508),
    .A1(net3546),
    .S(net454),
    .X(_01210_));
 sg13g2_mux2_1 _12818_ (.A0(net3700),
    .A1(net3543),
    .S(net452),
    .X(_01211_));
 sg13g2_mux2_1 _12819_ (.A0(net3623),
    .A1(net3560),
    .S(net453),
    .X(_01212_));
 sg13g2_mux2_1 _12820_ (.A0(\i_tinyqv.cpu.i_core.mepc[7] ),
    .A1(net3627),
    .S(net452),
    .X(_01213_));
 sg13g2_mux2_1 _12821_ (.A0(net3546),
    .A1(\i_tinyqv.cpu.i_core.mepc[12] ),
    .S(net454),
    .X(_01214_));
 sg13g2_mux2_1 _12822_ (.A0(net3543),
    .A1(net3498),
    .S(net452),
    .X(_01215_));
 sg13g2_mux2_1 _12823_ (.A0(net3560),
    .A1(net3529),
    .S(net453),
    .X(_01216_));
 sg13g2_mux2_1 _12824_ (.A0(net3627),
    .A1(net3640),
    .S(net452),
    .X(_01217_));
 sg13g2_mux2_1 _12825_ (.A0(net3574),
    .A1(net3540),
    .S(net454),
    .X(_01218_));
 sg13g2_mux2_1 _12826_ (.A0(net3498),
    .A1(\i_tinyqv.cpu.i_core.mepc[17] ),
    .S(net452),
    .X(_01219_));
 sg13g2_mux2_1 _12827_ (.A0(net3529),
    .A1(\i_tinyqv.cpu.i_core.mepc[18] ),
    .S(net453),
    .X(_01220_));
 sg13g2_mux2_1 _12828_ (.A0(net3640),
    .A1(net3425),
    .S(net452),
    .X(_01221_));
 sg13g2_mux2_1 _12829_ (.A0(net3540),
    .A1(\i_tinyqv.cpu.i_core.mepc[20] ),
    .S(net454),
    .X(_01222_));
 sg13g2_mux2_1 _12830_ (.A0(net3579),
    .A1(\i_tinyqv.cpu.i_core.mepc[21] ),
    .S(net452),
    .X(_01223_));
 sg13g2_mux2_1 _12831_ (.A0(net3564),
    .A1(net3615),
    .S(net452),
    .X(_01224_));
 sg13g2_mux2_1 _12832_ (.A0(net3425),
    .A1(net3625),
    .S(net454),
    .X(_01225_));
 sg13g2_mux2_1 _12833_ (.A0(_04089_),
    .A1(net627),
    .S(_04095_),
    .X(_01226_));
 sg13g2_mux2_1 _12834_ (.A0(_02221_),
    .A1(_02214_),
    .S(_02509_),
    .X(_04810_));
 sg13g2_nor2_1 _12835_ (.A(_04095_),
    .B(_04810_),
    .Y(_04811_));
 sg13g2_a21oi_1 _12836_ (.A1(net505),
    .A2(_04095_),
    .Y(_01227_),
    .B1(_04811_));
 sg13g2_or2_1 _12837_ (.X(_04812_),
    .B(_02509_),
    .A(_02396_));
 sg13g2_a21oi_1 _12838_ (.A1(_02388_),
    .A2(_02509_),
    .Y(_04813_),
    .B1(_04095_));
 sg13g2_a22oi_1 _12839_ (.Y(_01228_),
    .B1(_04812_),
    .B2(_04813_),
    .A2(_04095_),
    .A1(_01668_));
 sg13g2_a21oi_1 _12840_ (.A1(_02337_),
    .A2(_02509_),
    .Y(_04814_),
    .B1(_04095_));
 sg13g2_o21ai_1 _12841_ (.B1(_04814_),
    .Y(_04815_),
    .A1(_02343_),
    .A2(_02509_));
 sg13g2_nand2_1 _12842_ (.Y(_04816_),
    .A(net3673),
    .B(_04095_));
 sg13g2_nand2_1 _12843_ (.Y(_01229_),
    .A(_04815_),
    .B(_04816_));
 sg13g2_nor2_2 _12844_ (.A(net619),
    .B(net620),
    .Y(_04817_));
 sg13g2_nand3_1 _12845_ (.B(_03620_),
    .C(_04817_),
    .A(net117),
    .Y(_04818_));
 sg13g2_xnor2_1 _12846_ (.Y(_04819_),
    .A(net620),
    .B(_02535_));
 sg13g2_xor2_1 _12847_ (.B(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .A(net619),
    .X(_04820_));
 sg13g2_xnor2_1 _12848_ (.Y(_04821_),
    .A(_02534_),
    .B(_04820_));
 sg13g2_and2_1 _12849_ (.A(\i_tinyqv.mem.q_ctrl.data_req ),
    .B(_04821_),
    .X(_04822_));
 sg13g2_a22oi_1 _12850_ (.Y(_04823_),
    .B1(_04819_),
    .B2(_04822_),
    .A2(_04818_),
    .A1(\i_tinyqv.mem.data_stall ));
 sg13g2_a21oi_1 _12851_ (.A1(_02980_),
    .A2(_04823_),
    .Y(_01230_),
    .B1(_01610_));
 sg13g2_o21ai_1 _12852_ (.B1(_02814_),
    .Y(_04824_),
    .A1(_02805_),
    .A2(_02815_));
 sg13g2_nand2_1 _12853_ (.Y(_04825_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .B(net305));
 sg13g2_nor2_1 _12854_ (.A(_02788_),
    .B(_02808_),
    .Y(_04826_));
 sg13g2_a22oi_1 _12855_ (.Y(_04827_),
    .B1(net309),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .A2(net312),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[15] ));
 sg13g2_nor2_1 _12856_ (.A(_04826_),
    .B(_04827_),
    .Y(_04828_));
 sg13g2_o21ai_1 _12857_ (.B1(_02812_),
    .Y(_04829_),
    .A1(_02751_),
    .A2(_02808_));
 sg13g2_nand2_1 _12858_ (.Y(_04830_),
    .A(_04828_),
    .B(_04829_));
 sg13g2_xnor2_1 _12859_ (.Y(_04831_),
    .A(_04828_),
    .B(_04829_));
 sg13g2_xor2_1 _12860_ (.B(_04831_),
    .A(_04825_),
    .X(_04832_));
 sg13g2_nand2_1 _12861_ (.Y(_04833_),
    .A(_04824_),
    .B(_04832_));
 sg13g2_xnor2_1 _12862_ (.Y(_04834_),
    .A(_04824_),
    .B(_04832_));
 sg13g2_a21oi_1 _12863_ (.A1(_02817_),
    .A2(_02820_),
    .Y(_04835_),
    .B1(_04834_));
 sg13g2_nand3_1 _12864_ (.B(_02820_),
    .C(_04834_),
    .A(_02817_),
    .Y(_04836_));
 sg13g2_nand2b_1 _12865_ (.Y(_04837_),
    .B(_04836_),
    .A_N(_04835_));
 sg13g2_a21oi_1 _12866_ (.A1(_02822_),
    .A2(_02824_),
    .Y(_04838_),
    .B1(_04837_));
 sg13g2_nand3_1 _12867_ (.B(_02824_),
    .C(_04837_),
    .A(_02822_),
    .Y(_04839_));
 sg13g2_nor2b_1 _12868_ (.A(_04838_),
    .B_N(_04839_),
    .Y(_01231_));
 sg13g2_o21ai_1 _12869_ (.B1(_04830_),
    .Y(_04840_),
    .A1(_04825_),
    .A2(_04831_));
 sg13g2_nand2_1 _12870_ (.Y(_04841_),
    .A(net4129),
    .B(_04826_));
 sg13g2_a21o_1 _12871_ (.A2(net309),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .B1(_04826_),
    .X(_04842_));
 sg13g2_nand2_1 _12872_ (.Y(_04843_),
    .A(_04841_),
    .B(_04842_));
 sg13g2_nand2_1 _12873_ (.Y(_04844_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[15] ),
    .B(net305));
 sg13g2_xor2_1 _12874_ (.B(_04844_),
    .A(_04843_),
    .X(_04845_));
 sg13g2_xnor2_1 _12875_ (.Y(_04846_),
    .A(_04840_),
    .B(_04845_));
 sg13g2_nor2_1 _12876_ (.A(_04833_),
    .B(_04846_),
    .Y(_04847_));
 sg13g2_xor2_1 _12877_ (.B(_04846_),
    .A(_04833_),
    .X(_04848_));
 sg13g2_nor2_1 _12878_ (.A(_04835_),
    .B(_04838_),
    .Y(_04849_));
 sg13g2_xnor2_1 _12879_ (.Y(_01232_),
    .A(_04848_),
    .B(_04849_));
 sg13g2_o21ai_1 _12880_ (.B1(_04841_),
    .Y(_04850_),
    .A1(_04843_),
    .A2(_04844_));
 sg13g2_nor2_1 _12881_ (.A(_02808_),
    .B(_04850_),
    .Y(_04851_));
 sg13g2_nand3_1 _12882_ (.B(_04845_),
    .C(_04851_),
    .A(_04840_),
    .Y(_04852_));
 sg13g2_a21o_1 _12883_ (.A2(_04845_),
    .A1(_04840_),
    .B1(_04851_),
    .X(_04853_));
 sg13g2_and2_1 _12884_ (.A(_04852_),
    .B(_04853_),
    .X(_04854_));
 sg13g2_nor3_1 _12885_ (.A(_04835_),
    .B(_04838_),
    .C(_04847_),
    .Y(_04855_));
 sg13g2_a21oi_1 _12886_ (.A1(_04833_),
    .A2(_04846_),
    .Y(_04856_),
    .B1(_04855_));
 sg13g2_nand2_1 _12887_ (.Y(_04857_),
    .A(_04854_),
    .B(_04856_));
 sg13g2_xor2_1 _12888_ (.B(_04856_),
    .A(_04854_),
    .X(_01233_));
 sg13g2_nand3b_1 _12889_ (.B(_04852_),
    .C(_04857_),
    .Y(_01234_),
    .A_N(_04850_));
 sg13g2_nand2_1 _12890_ (.Y(_04858_),
    .A(_03130_),
    .B(_04302_));
 sg13g2_o21ai_1 _12891_ (.B1(_02537_),
    .Y(_04859_),
    .A1(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .A2(_02535_));
 sg13g2_nor2_1 _12892_ (.A(_03601_),
    .B(_04859_),
    .Y(_04860_));
 sg13g2_a22oi_1 _12893_ (.Y(_04861_),
    .B1(_04860_),
    .B2(_04302_),
    .A2(_04858_),
    .A1(_03601_));
 sg13g2_nor2b_1 _12894_ (.A(_03628_),
    .B_N(_00196_),
    .Y(_04862_));
 sg13g2_a22oi_1 _12895_ (.Y(_04863_),
    .B1(_04861_),
    .B2(_04862_),
    .A2(_03628_),
    .A1(net3754));
 sg13g2_nor3_1 _12896_ (.A(net517),
    .B(net73),
    .C(net3755),
    .Y(_01235_));
 sg13g2_nor2b_1 _12897_ (.A(_03628_),
    .B_N(_04820_),
    .Y(_04864_));
 sg13g2_a22oi_1 _12898_ (.Y(_04865_),
    .B1(_04861_),
    .B2(_04864_),
    .A2(_03628_),
    .A1(net619));
 sg13g2_nor3_1 _12899_ (.A(net516),
    .B(net73),
    .C(_04865_),
    .Y(_01236_));
 sg13g2_nand2_2 _12900_ (.Y(_04866_),
    .A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .B(_04817_));
 sg13g2_nor2_1 _12901_ (.A(net3886),
    .B(net431),
    .Y(_04867_));
 sg13g2_a21oi_1 _12902_ (.A1(_01660_),
    .A2(net431),
    .Y(_01237_),
    .B1(_04867_));
 sg13g2_nor2_1 _12903_ (.A(net3819),
    .B(net431),
    .Y(_04868_));
 sg13g2_a21oi_1 _12904_ (.A1(_01669_),
    .A2(net431),
    .Y(_01238_),
    .B1(_04868_));
 sg13g2_mux2_1 _12905_ (.A0(net3861),
    .A1(net4085),
    .S(net432),
    .X(_01239_));
 sg13g2_nor2_1 _12906_ (.A(net3937),
    .B(net432),
    .Y(_04869_));
 sg13g2_a21oi_1 _12907_ (.A1(_01684_),
    .A2(net432),
    .Y(_01240_),
    .B1(_04869_));
 sg13g2_nand2_1 _12908_ (.Y(_04870_),
    .A(\i_tinyqv.cpu.instr_data_in[4] ),
    .B(net431));
 sg13g2_o21ai_1 _12909_ (.B1(_04870_),
    .Y(_01241_),
    .A1(_01662_),
    .A2(net431));
 sg13g2_nor2_1 _12910_ (.A(\i_tinyqv.cpu.instr_data_in[13] ),
    .B(net432),
    .Y(_04871_));
 sg13g2_a21oi_1 _12911_ (.A1(_01671_),
    .A2(net431),
    .Y(_01242_),
    .B1(_04871_));
 sg13g2_nand2_1 _12912_ (.Y(_04872_),
    .A(net3947),
    .B(_04866_));
 sg13g2_o21ai_1 _12913_ (.B1(_04872_),
    .Y(_01243_),
    .A1(_01675_),
    .A2(net431));
 sg13g2_nand2_1 _12914_ (.Y(_04873_),
    .A(net3935),
    .B(net432));
 sg13g2_o21ai_1 _12915_ (.B1(_04873_),
    .Y(_01244_),
    .A1(_01687_),
    .A2(net432));
 sg13g2_or2_2 _12916_ (.X(_04874_),
    .B(_04817_),
    .A(_00196_));
 sg13g2_nor2_1 _12917_ (.A(_00245_),
    .B(net429),
    .Y(_04875_));
 sg13g2_nand2_2 _12918_ (.Y(_04876_),
    .A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .B(_04820_));
 sg13g2_nor3_1 _12919_ (.A(_00245_),
    .B(net430),
    .C(_04876_),
    .Y(_04877_));
 sg13g2_a21o_1 _12920_ (.A2(net433),
    .A1(net3416),
    .B1(_04877_),
    .X(_01245_));
 sg13g2_nor2_1 _12921_ (.A(_00246_),
    .B(net429),
    .Y(_04878_));
 sg13g2_nor3_1 _12922_ (.A(_00246_),
    .B(net430),
    .C(_04876_),
    .Y(_04879_));
 sg13g2_a21o_1 _12923_ (.A2(net433),
    .A1(net3415),
    .B1(_04879_),
    .X(_01246_));
 sg13g2_nor2_1 _12924_ (.A(_00247_),
    .B(net429),
    .Y(_04880_));
 sg13g2_nor3_1 _12925_ (.A(_00247_),
    .B(net430),
    .C(_04876_),
    .Y(_04881_));
 sg13g2_a21o_1 _12926_ (.A2(net433),
    .A1(net3399),
    .B1(_04881_),
    .X(_01247_));
 sg13g2_nor2_1 _12927_ (.A(_00248_),
    .B(net429),
    .Y(_04882_));
 sg13g2_nor3_1 _12928_ (.A(_00248_),
    .B(net430),
    .C(_04876_),
    .Y(_04883_));
 sg13g2_a21o_1 _12929_ (.A2(net433),
    .A1(net3366),
    .B1(_04883_),
    .X(_01248_));
 sg13g2_nor2_1 _12930_ (.A(_00249_),
    .B(net429),
    .Y(_04884_));
 sg13g2_nor3_1 _12931_ (.A(_00249_),
    .B(net430),
    .C(_04876_),
    .Y(_04885_));
 sg13g2_a21o_1 _12932_ (.A2(net433),
    .A1(net3351),
    .B1(_04885_),
    .X(_01249_));
 sg13g2_nor2_1 _12933_ (.A(_00250_),
    .B(net429),
    .Y(_04886_));
 sg13g2_nor3_1 _12934_ (.A(_00250_),
    .B(net430),
    .C(_04876_),
    .Y(_04887_));
 sg13g2_a21o_1 _12935_ (.A2(net433),
    .A1(net3358),
    .B1(_04887_),
    .X(_01250_));
 sg13g2_nor2_1 _12936_ (.A(_00251_),
    .B(net429),
    .Y(_04888_));
 sg13g2_nor3_1 _12937_ (.A(_00251_),
    .B(net430),
    .C(_04876_),
    .Y(_04889_));
 sg13g2_a21o_1 _12938_ (.A2(net433),
    .A1(net3412),
    .B1(_04889_),
    .X(_01251_));
 sg13g2_nor2_1 _12939_ (.A(_00252_),
    .B(net429),
    .Y(_04890_));
 sg13g2_nor3_1 _12940_ (.A(_00252_),
    .B(net430),
    .C(_04876_),
    .Y(_04891_));
 sg13g2_a21o_1 _12941_ (.A2(net433),
    .A1(net3410),
    .B1(_04891_),
    .X(_01252_));
 sg13g2_nand3b_1 _12942_ (.B(\i_tinyqv.mem.q_ctrl.data_ready ),
    .C(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .Y(_04892_),
    .A_N(net620));
 sg13g2_nand2_1 _12943_ (.Y(_04893_),
    .A(net3308),
    .B(net485));
 sg13g2_o21ai_1 _12944_ (.B1(_04893_),
    .Y(_01253_),
    .A1(_00245_),
    .A2(net485));
 sg13g2_nand2_1 _12945_ (.Y(_04894_),
    .A(net2988),
    .B(net484));
 sg13g2_o21ai_1 _12946_ (.B1(_04894_),
    .Y(_01254_),
    .A1(_00246_),
    .A2(net484));
 sg13g2_nand2_1 _12947_ (.Y(_04895_),
    .A(net3154),
    .B(net484));
 sg13g2_o21ai_1 _12948_ (.B1(_04895_),
    .Y(_01255_),
    .A1(_00247_),
    .A2(net484));
 sg13g2_nand2_1 _12949_ (.Y(_04896_),
    .A(net3360),
    .B(net484));
 sg13g2_o21ai_1 _12950_ (.B1(_04896_),
    .Y(_01256_),
    .A1(_00248_),
    .A2(net484));
 sg13g2_nand2_1 _12951_ (.Y(_04897_),
    .A(net2996),
    .B(net485));
 sg13g2_o21ai_1 _12952_ (.B1(_04897_),
    .Y(_01257_),
    .A1(_00249_),
    .A2(net485));
 sg13g2_nand2_1 _12953_ (.Y(_04898_),
    .A(net3092),
    .B(net485));
 sg13g2_o21ai_1 _12954_ (.B1(_04898_),
    .Y(_01258_),
    .A1(_00250_),
    .A2(net485));
 sg13g2_nand2_1 _12955_ (.Y(_04899_),
    .A(net3077),
    .B(net484));
 sg13g2_o21ai_1 _12956_ (.B1(_04899_),
    .Y(_01259_),
    .A1(_00251_),
    .A2(net484));
 sg13g2_nand2_1 _12957_ (.Y(_04900_),
    .A(net3331),
    .B(net485));
 sg13g2_o21ai_1 _12958_ (.B1(_04900_),
    .Y(_01260_),
    .A1(_00252_),
    .A2(_04892_));
 sg13g2_nand3_1 _12959_ (.B(net620),
    .C(\i_tinyqv.mem.q_ctrl.data_ready ),
    .A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .Y(_04901_));
 sg13g2_nand2_2 _12960_ (.Y(_04902_),
    .A(net432),
    .B(net483));
 sg13g2_a22oi_1 _12961_ (.Y(_04903_),
    .B1(_04902_),
    .B2(_04875_),
    .A2(net483),
    .A1(net3519));
 sg13g2_inv_1 _12962_ (.Y(_01261_),
    .A(_04903_));
 sg13g2_a22oi_1 _12963_ (.Y(_04904_),
    .B1(_04902_),
    .B2(_04878_),
    .A2(net483),
    .A1(net3455));
 sg13g2_inv_1 _12964_ (.Y(_01262_),
    .A(_04904_));
 sg13g2_a22oi_1 _12965_ (.Y(_04905_),
    .B1(_04902_),
    .B2(_04880_),
    .A2(net483),
    .A1(net3562));
 sg13g2_inv_1 _12966_ (.Y(_01263_),
    .A(_04905_));
 sg13g2_a22oi_1 _12967_ (.Y(_04906_),
    .B1(_04902_),
    .B2(_04882_),
    .A2(net483),
    .A1(net3437));
 sg13g2_inv_1 _12968_ (.Y(_01264_),
    .A(net3438));
 sg13g2_a22oi_1 _12969_ (.Y(_04907_),
    .B1(_04902_),
    .B2(_04884_),
    .A2(net483),
    .A1(net3306));
 sg13g2_inv_1 _12970_ (.Y(_01265_),
    .A(_04907_));
 sg13g2_a22oi_1 _12971_ (.Y(_04908_),
    .B1(_04902_),
    .B2(_04886_),
    .A2(net483),
    .A1(net3390));
 sg13g2_inv_1 _12972_ (.Y(_01266_),
    .A(net3391));
 sg13g2_a22oi_1 _12973_ (.Y(_04909_),
    .B1(_04902_),
    .B2(_04888_),
    .A2(_04901_),
    .A1(net3409));
 sg13g2_inv_1 _12974_ (.Y(_01267_),
    .A(_04909_));
 sg13g2_a22oi_1 _12975_ (.Y(_04910_),
    .B1(_04902_),
    .B2(_04890_),
    .A2(net483),
    .A1(net3363));
 sg13g2_inv_1 _12976_ (.Y(_01268_),
    .A(net3364));
 sg13g2_and2_1 _12977_ (.A(net534),
    .B(_04301_),
    .X(_01269_));
 sg13g2_a21oi_1 _12978_ (.A1(net4031),
    .A2(_03625_),
    .Y(_04911_),
    .B1(_04301_));
 sg13g2_nor2_1 _12979_ (.A(net517),
    .B(_04911_),
    .Y(_04912_));
 sg13g2_and2_1 _12980_ (.A(_03632_),
    .B(_04912_),
    .X(_01270_));
 sg13g2_mux2_1 _12981_ (.A0(net10),
    .A1(net3665),
    .S(net537),
    .X(_01271_));
 sg13g2_mux2_1 _12982_ (.A0(net11),
    .A1(net3829),
    .S(net537),
    .X(_01272_));
 sg13g2_or3_2 _12983_ (.A(net517),
    .B(net2837),
    .C(_04362_),
    .X(_04913_));
 sg13g2_inv_2 _12984_ (.Y(_04914_),
    .A(net30));
 sg13g2_nor2_2 _12985_ (.A(net486),
    .B(_04913_),
    .Y(_04915_));
 sg13g2_nand2b_2 _12986_ (.Y(_04916_),
    .B(_03615_),
    .A_N(\i_tinyqv.mem.data_stall ));
 sg13g2_nor2_1 _12987_ (.A(net3832),
    .B(_04916_),
    .Y(_04917_));
 sg13g2_o21ai_1 _12988_ (.B1(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .Y(_04918_),
    .A1(net3832),
    .A2(_04916_));
 sg13g2_nor3_2 _12989_ (.A(_01520_),
    .B(_01521_),
    .C(net616),
    .Y(_04919_));
 sg13g2_nand2_2 _12990_ (.Y(_04920_),
    .A(net615),
    .B(_03788_));
 sg13g2_nor2_1 _12991_ (.A(_04917_),
    .B(_04920_),
    .Y(_04921_));
 sg13g2_nor2_2 _12992_ (.A(net617),
    .B(_04920_),
    .Y(_04922_));
 sg13g2_a21o_1 _12993_ (.A2(_04922_),
    .A1(net3665),
    .B1(_04921_),
    .X(_04923_));
 sg13g2_nor2_2 _12994_ (.A(_03783_),
    .B(_04916_),
    .Y(_04924_));
 sg13g2_nor3_2 _12995_ (.A(net4056),
    .B(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .C(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .Y(_04925_));
 sg13g2_nand2_2 _12996_ (.Y(_04926_),
    .A(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .B(net616));
 sg13g2_nor2_1 _12997_ (.A(_00193_),
    .B(_04926_),
    .Y(_04927_));
 sg13g2_or2_1 _12998_ (.X(_04928_),
    .B(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .A(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ));
 sg13g2_nor2_1 _12999_ (.A(_03784_),
    .B(_04927_),
    .Y(_04929_));
 sg13g2_nor2_1 _13000_ (.A(_04928_),
    .B(_04929_),
    .Y(_04930_));
 sg13g2_a21oi_1 _13001_ (.A1(_00200_),
    .A2(_03784_),
    .Y(_04931_),
    .B1(_04927_));
 sg13g2_mux2_1 _13002_ (.A0(_04928_),
    .A1(_00199_),
    .S(_04931_),
    .X(_04932_));
 sg13g2_nor2b_1 _13003_ (.A(_04932_),
    .B_N(net547),
    .Y(_04933_));
 sg13g2_o21ai_1 _13004_ (.B1(_04933_),
    .Y(_04934_),
    .A1(_03783_),
    .A2(_04916_));
 sg13g2_nand2_1 _13005_ (.Y(_04935_),
    .A(net615),
    .B(_03623_));
 sg13g2_o21ai_1 _13006_ (.B1(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .Y(_04936_),
    .A1(_01520_),
    .A2(_03788_));
 sg13g2_o21ai_1 _13007_ (.B1(_04936_),
    .Y(_04937_),
    .A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .A2(_04935_));
 sg13g2_a221oi_1 _13008_ (.B2(_04933_),
    .C1(_04919_),
    .B1(_04937_),
    .A1(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .Y(_04938_),
    .A2(_04934_));
 sg13g2_a21oi_1 _13009_ (.A1(_04918_),
    .A2(_04923_),
    .Y(_04939_),
    .B1(_04938_));
 sg13g2_nor2_1 _13010_ (.A(net3900),
    .B(_04915_),
    .Y(_04940_));
 sg13g2_a21oi_1 _13011_ (.A1(_04915_),
    .A2(_04939_),
    .Y(_01273_),
    .B1(_04940_));
 sg13g2_nand2_1 _13012_ (.Y(_04941_),
    .A(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .B(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ));
 sg13g2_nand2_1 _13013_ (.Y(_04942_),
    .A(_04920_),
    .B(net547));
 sg13g2_nand2_1 _13014_ (.Y(_04943_),
    .A(_04920_),
    .B(_04933_));
 sg13g2_nand2b_1 _13015_ (.Y(_04944_),
    .B(_04916_),
    .A_N(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ));
 sg13g2_nand2b_1 _13016_ (.Y(_04945_),
    .B(_04941_),
    .A_N(_04916_));
 sg13g2_nand4_1 _13017_ (.B(net616),
    .C(_04944_),
    .A(net615),
    .Y(_04946_),
    .D(_04945_));
 sg13g2_nor2_1 _13018_ (.A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .B(_04935_),
    .Y(_04947_));
 sg13g2_a21oi_1 _13019_ (.A1(_04935_),
    .A2(_04941_),
    .Y(_04948_),
    .B1(_04947_));
 sg13g2_a21oi_1 _13020_ (.A1(_03783_),
    .A2(_04948_),
    .Y(_04949_),
    .B1(_04943_));
 sg13g2_a22oi_1 _13021_ (.Y(_04950_),
    .B1(_04946_),
    .B2(_04949_),
    .A2(_04943_),
    .A1(_04941_));
 sg13g2_mux2_1 _13022_ (.A0(net3832),
    .A1(_04950_),
    .S(_04915_),
    .X(_01274_));
 sg13g2_nand3_1 _13023_ (.B(_04920_),
    .C(_04932_),
    .A(_03625_),
    .Y(_04951_));
 sg13g2_nand3_1 _13024_ (.B(_03784_),
    .C(net547),
    .A(net617),
    .Y(_04952_));
 sg13g2_nor3_1 _13025_ (.A(net30),
    .B(_04951_),
    .C(_04952_),
    .Y(_01275_));
 sg13g2_nand2_1 _13026_ (.Y(_04953_),
    .A(net3887),
    .B(_04302_));
 sg13g2_nor2_1 _13027_ (.A(_00201_),
    .B(_04953_),
    .Y(_04954_));
 sg13g2_a21oi_1 _13028_ (.A1(_01617_),
    .A2(net3667),
    .Y(_04955_),
    .B1(net70));
 sg13g2_nand3_1 _13029_ (.B(net3666),
    .C(_04302_),
    .A(\addr[24] ),
    .Y(_04956_));
 sg13g2_o21ai_1 _13030_ (.B1(_04955_),
    .Y(_04957_),
    .A1(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ),
    .A2(_04956_));
 sg13g2_and2_1 _13031_ (.A(net486),
    .B(_04957_),
    .X(_04958_));
 sg13g2_inv_1 _13032_ (.Y(_04959_),
    .A(_04958_));
 sg13g2_nand2_1 _13033_ (.Y(_04960_),
    .A(_01523_),
    .B(_04920_));
 sg13g2_a221oi_1 _13034_ (.B2(_04960_),
    .C1(net30),
    .B1(_04959_),
    .A1(_01523_),
    .Y(_01276_),
    .A2(net486));
 sg13g2_nand2_1 _13035_ (.Y(_04961_),
    .A(net547),
    .B(_04926_));
 sg13g2_or4_1 _13036_ (.A(net615),
    .B(_00193_),
    .C(_04932_),
    .D(_04961_),
    .X(_04962_));
 sg13g2_nand3_1 _13037_ (.B(_04951_),
    .C(_04962_),
    .A(_04920_),
    .Y(_04963_));
 sg13g2_nor2_1 _13038_ (.A(_04958_),
    .B(_04963_),
    .Y(_04964_));
 sg13g2_or2_1 _13039_ (.X(_04965_),
    .B(_04963_),
    .A(_04958_));
 sg13g2_nor2_1 _13040_ (.A(net486),
    .B(_04963_),
    .Y(_04966_));
 sg13g2_o21ai_1 _13041_ (.B1(_04914_),
    .Y(_04967_),
    .A1(net3866),
    .A2(_04964_));
 sg13g2_a21oi_1 _13042_ (.A1(net3866),
    .A2(_04966_),
    .Y(_01277_),
    .B1(_04967_));
 sg13g2_a21oi_1 _13043_ (.A1(uio_out[0]),
    .A2(net515),
    .Y(_04968_),
    .B1(_03795_));
 sg13g2_o21ai_1 _13044_ (.B1(_03795_),
    .Y(_04969_),
    .A1(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .A2(_04926_));
 sg13g2_nand2b_1 _13045_ (.Y(_04970_),
    .B(_04969_),
    .A_N(_04968_));
 sg13g2_xor2_1 _13046_ (.B(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .A(net3820),
    .X(_04971_));
 sg13g2_a21oi_1 _13047_ (.A1(net547),
    .A2(_04970_),
    .Y(_04972_),
    .B1(_04971_));
 sg13g2_a22oi_1 _13048_ (.Y(_04973_),
    .B1(_04966_),
    .B2(_04972_),
    .A2(_04965_),
    .A1(net3820));
 sg13g2_nor2_1 _13049_ (.A(net30),
    .B(net3821),
    .Y(_01278_));
 sg13g2_a21oi_2 _13050_ (.B1(_03625_),
    .Y(_04974_),
    .A2(_04302_),
    .A1(\addr[24] ));
 sg13g2_o21ai_1 _13051_ (.B1(net3802),
    .Y(_04975_),
    .A1(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .A2(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ));
 sg13g2_nand2_1 _13052_ (.Y(_04976_),
    .A(_03622_),
    .B(net547));
 sg13g2_a21oi_1 _13053_ (.A1(_04975_),
    .A2(_04976_),
    .Y(_04977_),
    .B1(net486));
 sg13g2_nor3_1 _13054_ (.A(_04965_),
    .B(_04974_),
    .C(_04977_),
    .Y(_04978_));
 sg13g2_o21ai_1 _13055_ (.B1(_04914_),
    .Y(_04979_),
    .A1(net3802),
    .A2(_04964_));
 sg13g2_nor2_1 _13056_ (.A(_04978_),
    .B(_04979_),
    .Y(_01279_));
 sg13g2_a21oi_1 _13057_ (.A1(_01709_),
    .A2(net420),
    .Y(_04980_),
    .B1(_03599_));
 sg13g2_o21ai_1 _13058_ (.B1(_03627_),
    .Y(_04981_),
    .A1(_03618_),
    .A2(_04980_));
 sg13g2_nor2_1 _13059_ (.A(_04953_),
    .B(_04957_),
    .Y(_04982_));
 sg13g2_a22oi_1 _13060_ (.Y(_04983_),
    .B1(_04981_),
    .B2(_04982_),
    .A2(_04957_),
    .A1(net618));
 sg13g2_nor2_1 _13061_ (.A(net30),
    .B(_04983_),
    .Y(_01280_));
 sg13g2_and2_1 _13062_ (.A(net3883),
    .B(_04933_),
    .X(_04984_));
 sg13g2_a22oi_1 _13063_ (.Y(_04985_),
    .B1(_04924_),
    .B2(_04984_),
    .A2(_04922_),
    .A1(_04917_));
 sg13g2_nor3_1 _13064_ (.A(net486),
    .B(net30),
    .C(_04985_),
    .Y(_01281_));
 sg13g2_nor2_1 _13065_ (.A(_04919_),
    .B(net547),
    .Y(_04986_));
 sg13g2_nand2_1 _13066_ (.Y(_04987_),
    .A(_03625_),
    .B(net428));
 sg13g2_o21ai_1 _13067_ (.B1(_04951_),
    .Y(_04988_),
    .A1(_04927_),
    .A2(_04987_));
 sg13g2_or2_1 _13068_ (.X(_04989_),
    .B(_04988_),
    .A(_04921_));
 sg13g2_or2_1 _13069_ (.X(_04990_),
    .B(_04989_),
    .A(_04958_));
 sg13g2_a21oi_1 _13070_ (.A1(_00253_),
    .A2(_03795_),
    .Y(_04991_),
    .B1(_04968_));
 sg13g2_a21oi_1 _13071_ (.A1(net615),
    .A2(\i_tinyqv.mem.q_ctrl.fsm_state[0] ),
    .Y(_04992_),
    .B1(_04991_));
 sg13g2_nor4_1 _13072_ (.A(net486),
    .B(_04924_),
    .C(_04942_),
    .D(_04992_),
    .Y(_04993_));
 sg13g2_nor3_1 _13073_ (.A(_04974_),
    .B(_04990_),
    .C(_04993_),
    .Y(_04994_));
 sg13g2_a21oi_1 _13074_ (.A1(net3686),
    .A2(_04990_),
    .Y(_04995_),
    .B1(_04994_));
 sg13g2_nor2_1 _13075_ (.A(net30),
    .B(_04995_),
    .Y(_01282_));
 sg13g2_o21ai_1 _13076_ (.B1(_03794_),
    .Y(_04996_),
    .A1(uio_out[0]),
    .A2(net617));
 sg13g2_nand3b_1 _13077_ (.B(_04926_),
    .C(_04996_),
    .Y(_04997_),
    .A_N(_03623_));
 sg13g2_a21o_1 _13078_ (.A2(_04997_),
    .A1(_03783_),
    .B1(_04942_),
    .X(_04998_));
 sg13g2_a21oi_1 _13079_ (.A1(net3829),
    .A2(_04922_),
    .Y(_04999_),
    .B1(_04974_));
 sg13g2_o21ai_1 _13080_ (.B1(_04999_),
    .Y(_05000_),
    .A1(_04924_),
    .A2(_04998_));
 sg13g2_o21ai_1 _13081_ (.B1(_04914_),
    .Y(_05001_),
    .A1(_04990_),
    .A2(_05000_));
 sg13g2_a21oi_1 _13082_ (.A1(_01521_),
    .A2(_04990_),
    .Y(_01283_),
    .B1(_05001_));
 sg13g2_nand4_1 _13083_ (.B(_04925_),
    .C(_04926_),
    .A(_01520_),
    .Y(_05002_),
    .D(_04996_));
 sg13g2_nand2_1 _13084_ (.Y(_05003_),
    .A(_04915_),
    .B(_05002_));
 sg13g2_nand3_1 _13085_ (.B(_04914_),
    .C(_04990_),
    .A(net3431),
    .Y(_05004_));
 sg13g2_o21ai_1 _13086_ (.B1(_05004_),
    .Y(_01284_),
    .A1(_04989_),
    .A2(_05003_));
 sg13g2_o21ai_1 _13087_ (.B1(_04914_),
    .Y(_05005_),
    .A1(net3667),
    .A2(_04957_));
 sg13g2_a21o_1 _13088_ (.A2(_04957_),
    .A1(net3369),
    .B1(_05005_),
    .X(_01285_));
 sg13g2_a22oi_1 _13089_ (.Y(_05006_),
    .B1(_04957_),
    .B2(net3990),
    .A2(_04956_),
    .A1(_04955_));
 sg13g2_nand2_1 _13090_ (.Y(_01286_),
    .A(_04914_),
    .B(_05006_));
 sg13g2_a21oi_1 _13091_ (.A1(net4116),
    .A2(_04957_),
    .Y(_05007_),
    .B1(net30));
 sg13g2_nand2b_1 _13092_ (.Y(_01287_),
    .B(_05007_),
    .A_N(_04982_));
 sg13g2_nand2_1 _13093_ (.Y(_05008_),
    .A(_00193_),
    .B(_03783_));
 sg13g2_o21ai_1 _13094_ (.B1(_05008_),
    .Y(_05009_),
    .A1(net615),
    .A2(_04926_));
 sg13g2_or3_1 _13095_ (.A(_00200_),
    .B(_03795_),
    .C(_04942_),
    .X(_05010_));
 sg13g2_nand4_1 _13096_ (.B(_04997_),
    .C(_05009_),
    .A(_04987_),
    .Y(_05011_),
    .D(_05010_));
 sg13g2_nor4_2 _13097_ (.A(_03624_),
    .B(_04919_),
    .C(_04932_),
    .Y(_05012_),
    .D(_05011_));
 sg13g2_nand2b_1 _13098_ (.Y(_05013_),
    .B(net3374),
    .A_N(_05012_));
 sg13g2_a21oi_1 _13099_ (.A1(_04957_),
    .A2(_05013_),
    .Y(_01288_),
    .B1(_04913_));
 sg13g2_nor2_1 _13100_ (.A(_02840_),
    .B(_04793_),
    .Y(_05014_));
 sg13g2_nor2_1 _13101_ (.A(_02273_),
    .B(_04792_),
    .Y(_05015_));
 sg13g2_nor3_1 _13102_ (.A(_04794_),
    .B(_05014_),
    .C(_05015_),
    .Y(_05016_));
 sg13g2_a21oi_1 _13103_ (.A1(_02248_),
    .A2(_04794_),
    .Y(_05017_),
    .B1(_05016_));
 sg13g2_nand2_1 _13104_ (.Y(_05018_),
    .A(net3840),
    .B(net326));
 sg13g2_o21ai_1 _13105_ (.B1(_05018_),
    .Y(_01289_),
    .A1(_04798_),
    .A2(_05017_));
 sg13g2_nand2_1 _13106_ (.Y(_05019_),
    .A(_03238_),
    .B(_04792_));
 sg13g2_nor2_1 _13107_ (.A(_02214_),
    .B(_04792_),
    .Y(_05020_));
 sg13g2_nor2_1 _13108_ (.A(_04794_),
    .B(_05020_),
    .Y(_05021_));
 sg13g2_a22oi_1 _13109_ (.Y(_05022_),
    .B1(_05019_),
    .B2(_05021_),
    .A2(_04794_),
    .A1(_02156_));
 sg13g2_nand2_1 _13110_ (.Y(_05023_),
    .A(net3833),
    .B(net325));
 sg13g2_o21ai_1 _13111_ (.B1(_05023_),
    .Y(_01290_),
    .A1(_04798_),
    .A2(_05022_));
 sg13g2_nand2_1 _13112_ (.Y(_05024_),
    .A(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .B(_04922_));
 sg13g2_nor2_2 _13113_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .B(_05024_),
    .Y(_05025_));
 sg13g2_mux2_1 _13114_ (.A0(net3270),
    .A1(net10),
    .S(_05025_),
    .X(_01291_));
 sg13g2_mux2_1 _13115_ (.A0(net3249),
    .A1(net11),
    .S(_05025_),
    .X(_01292_));
 sg13g2_mux2_1 _13116_ (.A0(net3343),
    .A1(net12),
    .S(_05025_),
    .X(_01293_));
 sg13g2_mux2_1 _13117_ (.A0(net3263),
    .A1(net13),
    .S(_05025_),
    .X(_01294_));
 sg13g2_nand2_1 _13118_ (.Y(_05026_),
    .A(net620),
    .B(\i_tinyqv.mem.q_ctrl.data_req ));
 sg13g2_xor2_1 _13119_ (.B(\i_tinyqv.mem.q_ctrl.data_req ),
    .A(net620),
    .X(_05027_));
 sg13g2_xnor2_1 _13120_ (.Y(_05028_),
    .A(net620),
    .B(\i_tinyqv.mem.q_ctrl.data_req ));
 sg13g2_nand2_1 _13121_ (.Y(_05029_),
    .A(\data_to_write[0] ),
    .B(net480));
 sg13g2_xnor2_1 _13122_ (.Y(_05030_),
    .A(net619),
    .B(_05026_));
 sg13g2_xor2_1 _13123_ (.B(_05026_),
    .A(net619),
    .X(_05031_));
 sg13g2_a21oi_1 _13124_ (.A1(\data_to_write[8] ),
    .A2(net481),
    .Y(_05032_),
    .B1(_05030_));
 sg13g2_nand2_1 _13125_ (.Y(_05033_),
    .A(\data_to_write[16] ),
    .B(net479));
 sg13g2_a21oi_1 _13126_ (.A1(\data_to_write[24] ),
    .A2(net481),
    .Y(_05034_),
    .B1(_05031_));
 sg13g2_a221oi_1 _13127_ (.B2(_05034_),
    .C1(net428),
    .B1(_05033_),
    .A1(_05029_),
    .Y(_05035_),
    .A2(_05032_));
 sg13g2_a21oi_1 _13128_ (.A1(net10),
    .A2(net428),
    .Y(_05036_),
    .B1(net515));
 sg13g2_nand2b_1 _13129_ (.Y(_05037_),
    .B(_05036_),
    .A_N(_05035_));
 sg13g2_nand3b_1 _13130_ (.B(_03785_),
    .C(net428),
    .Y(_05038_),
    .A_N(_00199_));
 sg13g2_a21oi_1 _13131_ (.A1(_01523_),
    .A2(_04920_),
    .Y(_05039_),
    .B1(_01522_));
 sg13g2_a22oi_1 _13132_ (.Y(_05040_),
    .B1(_05038_),
    .B2(_05039_),
    .A2(_04930_),
    .A1(_01522_));
 sg13g2_nor2_2 _13133_ (.A(_03785_),
    .B(_04928_),
    .Y(_05041_));
 sg13g2_or2_1 _13134_ (.X(_05042_),
    .B(_04928_),
    .A(_03785_));
 sg13g2_nand2_1 _13135_ (.Y(_05043_),
    .A(net3270),
    .B(_05042_));
 sg13g2_a21oi_1 _13136_ (.A1(net10),
    .A2(_05041_),
    .Y(_05044_),
    .B1(net617));
 sg13g2_a21oi_2 _13137_ (.B1(net324),
    .Y(_05045_),
    .A2(_05044_),
    .A1(_05043_));
 sg13g2_a22oi_1 _13138_ (.Y(_05046_),
    .B1(_05045_),
    .B2(_05037_),
    .A2(net324),
    .A1(net3886));
 sg13g2_inv_1 _13139_ (.Y(_01295_),
    .A(_05046_));
 sg13g2_nand2_1 _13140_ (.Y(_05047_),
    .A(net601),
    .B(net480));
 sg13g2_a21oi_1 _13141_ (.A1(\data_to_write[9] ),
    .A2(net482),
    .Y(_05048_),
    .B1(_05030_));
 sg13g2_nand2_1 _13142_ (.Y(_05049_),
    .A(\data_to_write[17] ),
    .B(net479));
 sg13g2_a21oi_1 _13143_ (.A1(\data_to_write[25] ),
    .A2(net482),
    .Y(_05050_),
    .B1(_05031_));
 sg13g2_a221oi_1 _13144_ (.B2(_05050_),
    .C1(net428),
    .B1(_05049_),
    .A1(_05047_),
    .Y(_05051_),
    .A2(_05048_));
 sg13g2_a21oi_1 _13145_ (.A1(net11),
    .A2(_04986_),
    .Y(_05052_),
    .B1(net515));
 sg13g2_nand2b_1 _13146_ (.Y(_05053_),
    .B(_05052_),
    .A_N(_05051_));
 sg13g2_nand2_1 _13147_ (.Y(_05054_),
    .A(net3249),
    .B(_05042_));
 sg13g2_a21oi_1 _13148_ (.A1(net11),
    .A2(_05041_),
    .Y(_05055_),
    .B1(net617));
 sg13g2_a21oi_1 _13149_ (.A1(_05054_),
    .A2(_05055_),
    .Y(_05056_),
    .B1(net324));
 sg13g2_a22oi_1 _13150_ (.Y(_05057_),
    .B1(_05053_),
    .B2(_05056_),
    .A2(net324),
    .A1(net3819));
 sg13g2_inv_1 _13151_ (.Y(_01296_),
    .A(_05057_));
 sg13g2_nand2_1 _13152_ (.Y(_05058_),
    .A(net600),
    .B(net480));
 sg13g2_a21oi_1 _13153_ (.A1(\data_to_write[10] ),
    .A2(net482),
    .Y(_05059_),
    .B1(_05030_));
 sg13g2_nand2_1 _13154_ (.Y(_05060_),
    .A(\data_to_write[18] ),
    .B(net480));
 sg13g2_a21oi_1 _13155_ (.A1(\data_to_write[26] ),
    .A2(net482),
    .Y(_05061_),
    .B1(_05031_));
 sg13g2_a221oi_1 _13156_ (.B2(_05061_),
    .C1(net428),
    .B1(_05060_),
    .A1(_05058_),
    .Y(_05062_),
    .A2(_05059_));
 sg13g2_a21oi_1 _13157_ (.A1(net12),
    .A2(net428),
    .Y(_05063_),
    .B1(net515));
 sg13g2_nand2b_1 _13158_ (.Y(_05064_),
    .B(_05063_),
    .A_N(_05062_));
 sg13g2_nand2_1 _13159_ (.Y(_05065_),
    .A(net3343),
    .B(_05042_));
 sg13g2_a21oi_1 _13160_ (.A1(net12),
    .A2(_05041_),
    .Y(_05066_),
    .B1(net617));
 sg13g2_a21oi_1 _13161_ (.A1(_05065_),
    .A2(_05066_),
    .Y(_05067_),
    .B1(net324));
 sg13g2_a22oi_1 _13162_ (.Y(_05068_),
    .B1(_05064_),
    .B2(_05067_),
    .A2(net324),
    .A1(net3861));
 sg13g2_inv_1 _13163_ (.Y(_01297_),
    .A(_05068_));
 sg13g2_nand2_1 _13164_ (.Y(_05069_),
    .A(\data_to_write[11] ),
    .B(net481));
 sg13g2_o21ai_1 _13165_ (.B1(_05069_),
    .Y(_05070_),
    .A1(_01508_),
    .A2(net481));
 sg13g2_nand2_1 _13166_ (.Y(_05071_),
    .A(\data_to_write[19] ),
    .B(net480));
 sg13g2_a21oi_1 _13167_ (.A1(\data_to_write[27] ),
    .A2(net482),
    .Y(_05072_),
    .B1(_05031_));
 sg13g2_a21oi_1 _13168_ (.A1(_05071_),
    .A2(_05072_),
    .Y(_05073_),
    .B1(net428));
 sg13g2_o21ai_1 _13169_ (.B1(_05073_),
    .Y(_05074_),
    .A1(_05030_),
    .A2(_05070_));
 sg13g2_a21oi_1 _13170_ (.A1(net13),
    .A2(_04986_),
    .Y(_05075_),
    .B1(net515));
 sg13g2_and2_1 _13171_ (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .B(_05042_),
    .X(_05076_));
 sg13g2_a21oi_1 _13172_ (.A1(net13),
    .A2(_05041_),
    .Y(_05077_),
    .B1(_05076_));
 sg13g2_a221oi_1 _13173_ (.B2(net515),
    .C1(_05040_),
    .B1(_05077_),
    .A1(_05074_),
    .Y(_05078_),
    .A2(_05075_));
 sg13g2_a21o_1 _13174_ (.A2(net323),
    .A1(net3937),
    .B1(_05078_),
    .X(_01298_));
 sg13g2_o21ai_1 _13175_ (.B1(net617),
    .Y(_05079_),
    .A1(_04919_),
    .A2(net547));
 sg13g2_nand2_1 _13176_ (.Y(_05080_),
    .A(net599),
    .B(net479));
 sg13g2_a21oi_1 _13177_ (.A1(\data_to_write[12] ),
    .A2(net481),
    .Y(_05081_),
    .B1(_05030_));
 sg13g2_mux2_1 _13178_ (.A0(\data_to_write[28] ),
    .A1(\data_to_write[20] ),
    .S(net479),
    .X(_05082_));
 sg13g2_a21oi_1 _13179_ (.A1(_05080_),
    .A2(_05081_),
    .Y(_05083_),
    .B1(_05079_));
 sg13g2_o21ai_1 _13180_ (.B1(_05083_),
    .Y(_05084_),
    .A1(_05031_),
    .A2(_05082_));
 sg13g2_a21oi_1 _13181_ (.A1(net3886),
    .A2(_05079_),
    .Y(_05085_),
    .B1(net324));
 sg13g2_a22oi_1 _13182_ (.Y(_01299_),
    .B1(_05084_),
    .B2(_05085_),
    .A2(net323),
    .A1(_01662_));
 sg13g2_mux2_1 _13183_ (.A0(\data_to_write[29] ),
    .A1(\data_to_write[21] ),
    .S(net480),
    .X(_05086_));
 sg13g2_nand2_1 _13184_ (.Y(_05087_),
    .A(net598),
    .B(net479));
 sg13g2_a21oi_1 _13185_ (.A1(\data_to_write[13] ),
    .A2(net481),
    .Y(_05088_),
    .B1(_05030_));
 sg13g2_a21oi_1 _13186_ (.A1(_05087_),
    .A2(_05088_),
    .Y(_05089_),
    .B1(_05079_));
 sg13g2_o21ai_1 _13187_ (.B1(_05089_),
    .Y(_05090_),
    .A1(_05031_),
    .A2(_05086_));
 sg13g2_a21oi_1 _13188_ (.A1(net3819),
    .A2(_05079_),
    .Y(_05091_),
    .B1(net323));
 sg13g2_a22oi_1 _13189_ (.Y(_01300_),
    .B1(_05090_),
    .B2(_05091_),
    .A2(net323),
    .A1(_01672_));
 sg13g2_mux2_1 _13190_ (.A0(\data_to_write[30] ),
    .A1(\data_to_write[22] ),
    .S(net479),
    .X(_05092_));
 sg13g2_nand2_1 _13191_ (.Y(_05093_),
    .A(net597),
    .B(net480));
 sg13g2_a21oi_1 _13192_ (.A1(\data_to_write[14] ),
    .A2(net481),
    .Y(_05094_),
    .B1(_05030_));
 sg13g2_a21oi_1 _13193_ (.A1(_05093_),
    .A2(_05094_),
    .Y(_05095_),
    .B1(_05079_));
 sg13g2_o21ai_1 _13194_ (.B1(_05095_),
    .Y(_05096_),
    .A1(_05031_),
    .A2(_05092_));
 sg13g2_a21oi_1 _13195_ (.A1(net3861),
    .A2(_05079_),
    .Y(_05097_),
    .B1(net323));
 sg13g2_a22oi_1 _13196_ (.Y(_01301_),
    .B1(_05096_),
    .B2(_05097_),
    .A2(net323),
    .A1(_01675_));
 sg13g2_mux2_1 _13197_ (.A0(\data_to_write[31] ),
    .A1(\data_to_write[23] ),
    .S(net479),
    .X(_05098_));
 sg13g2_nand2_1 _13198_ (.Y(_05099_),
    .A(\data_to_write[7] ),
    .B(net479));
 sg13g2_a21oi_1 _13199_ (.A1(\data_to_write[15] ),
    .A2(net481),
    .Y(_05100_),
    .B1(_05030_));
 sg13g2_a21oi_1 _13200_ (.A1(_05099_),
    .A2(_05100_),
    .Y(_05101_),
    .B1(_05079_));
 sg13g2_o21ai_1 _13201_ (.B1(_05101_),
    .Y(_05102_),
    .A1(_05031_),
    .A2(_05098_));
 sg13g2_a21oi_1 _13202_ (.A1(net3937),
    .A2(_05079_),
    .Y(_05103_),
    .B1(net323));
 sg13g2_a22oi_1 _13203_ (.Y(_01302_),
    .B1(_05102_),
    .B2(_05103_),
    .A2(net323),
    .A1(_01687_));
 sg13g2_nand2b_1 _13204_ (.Y(_01303_),
    .B(net535),
    .A_N(net3369));
 sg13g2_nand2b_1 _13205_ (.Y(_01304_),
    .B(net537),
    .A_N(net3990));
 sg13g2_mux2_1 _13206_ (.A0(net12),
    .A1(net3801),
    .S(net535),
    .X(_01306_));
 sg13g2_nor3_1 _13207_ (.A(net3804),
    .B(net647),
    .C(net44),
    .Y(_05104_));
 sg13g2_a21oi_1 _13208_ (.A1(_01660_),
    .A2(net44),
    .Y(_01307_),
    .B1(_05104_));
 sg13g2_nor3_1 _13209_ (.A(\i_tinyqv.cpu.instr_data[2][1] ),
    .B(net647),
    .C(net43),
    .Y(_05105_));
 sg13g2_a21oi_1 _13210_ (.A1(_01669_),
    .A2(net43),
    .Y(_01308_),
    .B1(_05105_));
 sg13g2_nor3_1 _13211_ (.A(net3875),
    .B(net647),
    .C(net33),
    .Y(_05106_));
 sg13g2_a21oi_1 _13212_ (.A1(_01660_),
    .A2(net33),
    .Y(_01309_),
    .B1(_05106_));
 sg13g2_nor3_1 _13213_ (.A(net3730),
    .B(net647),
    .C(net33),
    .Y(_05107_));
 sg13g2_a21oi_1 _13214_ (.A1(_01669_),
    .A2(net33),
    .Y(_01310_),
    .B1(_05107_));
 sg13g2_nand2_1 _13215_ (.Y(_05108_),
    .A(\i_tinyqv.cpu.pc[1] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[1] ));
 sg13g2_xnor2_1 _13216_ (.Y(_05109_),
    .A(\i_tinyqv.cpu.pc[1] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[1] ));
 sg13g2_mux2_1 _13217_ (.A0(_04729_),
    .A1(_05109_),
    .S(net414),
    .X(_05110_));
 sg13g2_nand3_1 _13218_ (.B(net91),
    .C(net80),
    .A(net2841),
    .Y(_05111_));
 sg13g2_o21ai_1 _13219_ (.B1(_05111_),
    .Y(_05112_),
    .A1(net91),
    .A2(_05110_));
 sg13g2_a21oi_1 _13220_ (.A1(_03609_),
    .A2(net69),
    .Y(_05113_),
    .B1(_05112_));
 sg13g2_nor2_1 _13221_ (.A(net514),
    .B(_05113_),
    .Y(_01311_));
 sg13g2_nand2_1 _13222_ (.Y(_05114_),
    .A(\i_tinyqv.cpu.pc[2] ),
    .B(net582));
 sg13g2_xnor2_1 _13223_ (.Y(_05115_),
    .A(\i_tinyqv.cpu.pc[2] ),
    .B(net582));
 sg13g2_xnor2_1 _13224_ (.Y(_05116_),
    .A(_05108_),
    .B(_05115_));
 sg13g2_nor2_1 _13225_ (.A(net410),
    .B(_05116_),
    .Y(_05117_));
 sg13g2_a21oi_1 _13226_ (.A1(net410),
    .A2(_04730_),
    .Y(_05118_),
    .B1(_05117_));
 sg13g2_nand3_1 _13227_ (.B(net91),
    .C(net80),
    .A(net2842),
    .Y(_05119_));
 sg13g2_o21ai_1 _13228_ (.B1(_05119_),
    .Y(_05120_),
    .A1(net91),
    .A2(_05118_));
 sg13g2_inv_1 _13229_ (.Y(_05121_),
    .A(_05120_));
 sg13g2_a21oi_1 _13230_ (.A1(_03611_),
    .A2(net69),
    .Y(_05122_),
    .B1(_05120_));
 sg13g2_nor2_1 _13231_ (.A(net512),
    .B(_05122_),
    .Y(_01312_));
 sg13g2_nor2_1 _13232_ (.A(net604),
    .B(\i_tinyqv.cpu.instr_write_offset[1] ),
    .Y(_05123_));
 sg13g2_a21oi_2 _13233_ (.B1(_05123_),
    .Y(_05124_),
    .A2(_05109_),
    .A1(net604));
 sg13g2_nor2_1 _13234_ (.A(net70),
    .B(_04302_),
    .Y(_05125_));
 sg13g2_o21ai_1 _13235_ (.B1(net73),
    .Y(_05126_),
    .A1(_01604_),
    .A2(_04301_));
 sg13g2_a22oi_1 _13236_ (.Y(_05127_),
    .B1(_05124_),
    .B2(net58),
    .A2(net276),
    .A1(net2380));
 sg13g2_o21ai_1 _13237_ (.B1(_05127_),
    .Y(_01313_),
    .A1(_01697_),
    .A2(_04300_));
 sg13g2_nand2_1 _13238_ (.Y(_05128_),
    .A(net604),
    .B(_05116_));
 sg13g2_o21ai_1 _13239_ (.B1(_05128_),
    .Y(_05129_),
    .A1(net604),
    .A2(\i_tinyqv.cpu.instr_write_offset[2] ));
 sg13g2_a22oi_1 _13240_ (.Y(_05130_),
    .B1(net276),
    .B2(net633),
    .A2(net59),
    .A1(net3654));
 sg13g2_o21ai_1 _13241_ (.B1(net3655),
    .Y(_01314_),
    .A1(_05126_),
    .A2(_05129_));
 sg13g2_and2_1 _13242_ (.A(\i_tinyqv.cpu.instr_data_start[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .X(_05131_));
 sg13g2_xor2_1 _13243_ (.B(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .A(\i_tinyqv.cpu.instr_data_start[3] ),
    .X(_05132_));
 sg13g2_o21ai_1 _13244_ (.B1(_05114_),
    .Y(_05133_),
    .A1(_05108_),
    .A2(_05115_));
 sg13g2_xor2_1 _13245_ (.B(_05133_),
    .A(_05132_),
    .X(_05134_));
 sg13g2_nand2_2 _13246_ (.Y(_05135_),
    .A(\i_tinyqv.cpu.instr_data_start[3] ),
    .B(\i_tinyqv.cpu.instr_write_offset[3] ));
 sg13g2_nor2_1 _13247_ (.A(\i_tinyqv.cpu.instr_data_start[3] ),
    .B(\i_tinyqv.cpu.instr_write_offset[3] ),
    .Y(_05136_));
 sg13g2_nor2_1 _13248_ (.A(net608),
    .B(_05136_),
    .Y(_05137_));
 sg13g2_a22oi_1 _13249_ (.Y(_05138_),
    .B1(_05135_),
    .B2(_05137_),
    .A2(_05134_),
    .A1(net608));
 sg13g2_a22oi_1 _13250_ (.Y(_05139_),
    .B1(net276),
    .B2(\addr[3] ),
    .A2(net59),
    .A1(net3676));
 sg13g2_o21ai_1 _13251_ (.B1(net3677),
    .Y(_01315_),
    .A1(_05126_),
    .A2(_05138_));
 sg13g2_nand2_1 _13252_ (.Y(_05140_),
    .A(\i_tinyqv.cpu.instr_data_start[4] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[4] ));
 sg13g2_xnor2_1 _13253_ (.Y(_05141_),
    .A(\i_tinyqv.cpu.instr_data_start[4] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[4] ));
 sg13g2_a21oi_1 _13254_ (.A1(_05132_),
    .A2(_05133_),
    .Y(_05142_),
    .B1(_05131_));
 sg13g2_xnor2_1 _13255_ (.Y(_05143_),
    .A(_05141_),
    .B(_05142_));
 sg13g2_nand2_1 _13256_ (.Y(_05144_),
    .A(net608),
    .B(_05143_));
 sg13g2_xnor2_1 _13257_ (.Y(_05145_),
    .A(\i_tinyqv.cpu.instr_data_start[4] ),
    .B(_05135_));
 sg13g2_o21ai_1 _13258_ (.B1(_05144_),
    .Y(_05146_),
    .A1(net608),
    .A2(_05145_));
 sg13g2_a21oi_1 _13259_ (.A1(net3267),
    .A2(net401),
    .Y(_05147_),
    .B1(net73));
 sg13g2_a221oi_1 _13260_ (.B2(_05146_),
    .C1(_05147_),
    .B1(net58),
    .A1(_01616_),
    .Y(_05148_),
    .A2(net276));
 sg13g2_a21o_1 _13261_ (.A2(net59),
    .A1(net3372),
    .B1(_05148_),
    .X(_01316_));
 sg13g2_and2_1 _13262_ (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .X(_05149_));
 sg13g2_xor2_1 _13263_ (.B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .A(\i_tinyqv.cpu.instr_data_start[5] ),
    .X(_05150_));
 sg13g2_o21ai_1 _13264_ (.B1(_05140_),
    .Y(_05151_),
    .A1(_05141_),
    .A2(_05142_));
 sg13g2_xor2_1 _13265_ (.B(_05151_),
    .A(_05150_),
    .X(_05152_));
 sg13g2_nand2_1 _13266_ (.Y(_05153_),
    .A(net608),
    .B(_05152_));
 sg13g2_nor3_2 _13267_ (.A(_01519_),
    .B(_00203_),
    .C(_05135_),
    .Y(_05154_));
 sg13g2_o21ai_1 _13268_ (.B1(_01519_),
    .Y(_05155_),
    .A1(_00203_),
    .A2(_05135_));
 sg13g2_nand2_1 _13269_ (.Y(_05156_),
    .A(net478),
    .B(_05155_));
 sg13g2_o21ai_1 _13270_ (.B1(_05153_),
    .Y(_05157_),
    .A1(_05154_),
    .A2(_05156_));
 sg13g2_nand2_1 _13271_ (.Y(_05158_),
    .A(net56),
    .B(_05157_));
 sg13g2_a221oi_1 _13272_ (.B2(\addr[5] ),
    .C1(net59),
    .B1(net277),
    .A1(net3279),
    .Y(_05159_),
    .A2(net70));
 sg13g2_a22oi_1 _13273_ (.Y(_01317_),
    .B1(_05158_),
    .B2(_05159_),
    .A2(net61),
    .A1(_01698_));
 sg13g2_and2_1 _13274_ (.A(\i_tinyqv.cpu.instr_data_start[6] ),
    .B(_05154_),
    .X(_05160_));
 sg13g2_nand2_1 _13275_ (.Y(_05161_),
    .A(\i_tinyqv.cpu.instr_data_start[6] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[6] ));
 sg13g2_xnor2_1 _13276_ (.Y(_05162_),
    .A(\i_tinyqv.cpu.instr_data_start[6] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[6] ));
 sg13g2_a21oi_2 _13277_ (.B1(_05149_),
    .Y(_05163_),
    .A2(_05151_),
    .A1(_05150_));
 sg13g2_xnor2_1 _13278_ (.Y(_05164_),
    .A(_05162_),
    .B(_05163_));
 sg13g2_nor2_1 _13279_ (.A(net477),
    .B(_05164_),
    .Y(_05165_));
 sg13g2_o21ai_1 _13280_ (.B1(net478),
    .Y(_05166_),
    .A1(\i_tinyqv.cpu.instr_data_start[6] ),
    .A2(_05154_));
 sg13g2_nor2_1 _13281_ (.A(_05160_),
    .B(_05166_),
    .Y(_05167_));
 sg13g2_o21ai_1 _13282_ (.B1(net57),
    .Y(_05168_),
    .A1(_05165_),
    .A2(_05167_));
 sg13g2_a221oi_1 _13283_ (.B2(\addr[6] ),
    .C1(net59),
    .B1(net276),
    .A1(\i_tinyqv.mem.q_ctrl.addr[2] ),
    .Y(_05169_),
    .A2(net70));
 sg13g2_a22oi_1 _13284_ (.Y(_01318_),
    .B1(_05168_),
    .B2(_05169_),
    .A2(net62),
    .A1(_01699_));
 sg13g2_xnor2_1 _13285_ (.Y(_05170_),
    .A(_01518_),
    .B(_05160_));
 sg13g2_nor2_1 _13286_ (.A(net605),
    .B(_05170_),
    .Y(_05171_));
 sg13g2_and2_1 _13287_ (.A(\i_tinyqv.cpu.instr_data_start[7] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .X(_05172_));
 sg13g2_xor2_1 _13288_ (.B(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .A(\i_tinyqv.cpu.instr_data_start[7] ),
    .X(_05173_));
 sg13g2_o21ai_1 _13289_ (.B1(_05161_),
    .Y(_05174_),
    .A1(_05162_),
    .A2(_05163_));
 sg13g2_xnor2_1 _13290_ (.Y(_05175_),
    .A(_05173_),
    .B(_05174_));
 sg13g2_a21oi_1 _13291_ (.A1(net605),
    .A2(_05175_),
    .Y(_05176_),
    .B1(_05171_));
 sg13g2_a22oi_1 _13292_ (.Y(_05177_),
    .B1(net276),
    .B2(net3329),
    .A2(net70),
    .A1(\i_tinyqv.mem.q_ctrl.addr[3] ));
 sg13g2_a22oi_1 _13293_ (.Y(_05178_),
    .B1(net57),
    .B2(_05176_),
    .A2(net62),
    .A1(net3550));
 sg13g2_o21ai_1 _13294_ (.B1(_05178_),
    .Y(_01319_),
    .A1(net62),
    .A2(_05177_));
 sg13g2_nand2b_1 _13295_ (.Y(_05179_),
    .B(net276),
    .A_N(\addr[8] ));
 sg13g2_o21ai_1 _13296_ (.B1(_05179_),
    .Y(_05180_),
    .A1(net3372),
    .A2(net72));
 sg13g2_xnor2_1 _13297_ (.Y(_05181_),
    .A(\i_tinyqv.cpu.instr_data_start[8] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ));
 sg13g2_a21oi_1 _13298_ (.A1(_05173_),
    .A2(_05174_),
    .Y(_05182_),
    .B1(_05172_));
 sg13g2_nor2_1 _13299_ (.A(_05181_),
    .B(_05182_),
    .Y(_05183_));
 sg13g2_xor2_1 _13300_ (.B(_05182_),
    .A(_05181_),
    .X(_05184_));
 sg13g2_a21oi_1 _13301_ (.A1(\i_tinyqv.cpu.instr_data_start[7] ),
    .A2(_05160_),
    .Y(_05185_),
    .B1(\i_tinyqv.cpu.instr_data_start[8] ));
 sg13g2_and3_1 _13302_ (.X(_05186_),
    .A(\i_tinyqv.cpu.instr_data_start[8] ),
    .B(\i_tinyqv.cpu.instr_data_start[7] ),
    .C(_05160_));
 sg13g2_o21ai_1 _13303_ (.B1(net477),
    .Y(_05187_),
    .A1(_05185_),
    .A2(_05186_));
 sg13g2_o21ai_1 _13304_ (.B1(_05187_),
    .Y(_05188_),
    .A1(net477),
    .A2(_05184_));
 sg13g2_nor2_1 _13305_ (.A(net3470),
    .B(_04300_),
    .Y(_05189_));
 sg13g2_a221oi_1 _13306_ (.B2(net56),
    .C1(_05189_),
    .B1(_05188_),
    .A1(_04300_),
    .Y(_01320_),
    .A2(_05180_));
 sg13g2_a21oi_2 _13307_ (.B1(_05183_),
    .Y(_05190_),
    .A2(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .A1(\i_tinyqv.cpu.instr_data_start[8] ));
 sg13g2_nand2_1 _13308_ (.Y(_05191_),
    .A(\i_tinyqv.cpu.instr_data_start[9] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[9] ));
 sg13g2_nor2_1 _13309_ (.A(\i_tinyqv.cpu.instr_data_start[9] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .Y(_05192_));
 sg13g2_xor2_1 _13310_ (.B(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .A(\i_tinyqv.cpu.instr_data_start[9] ),
    .X(_05193_));
 sg13g2_xnor2_1 _13311_ (.Y(_05194_),
    .A(_05190_),
    .B(_05193_));
 sg13g2_and2_1 _13312_ (.A(\i_tinyqv.cpu.instr_data_start[9] ),
    .B(_05186_),
    .X(_05195_));
 sg13g2_o21ai_1 _13313_ (.B1(net477),
    .Y(_05196_),
    .A1(\i_tinyqv.cpu.instr_data_start[9] ),
    .A2(_05186_));
 sg13g2_nor2_1 _13314_ (.A(_05195_),
    .B(_05196_),
    .Y(_05197_));
 sg13g2_a21oi_1 _13315_ (.A1(net605),
    .A2(_05194_),
    .Y(_05198_),
    .B1(_05197_));
 sg13g2_a21oi_1 _13316_ (.A1(\i_tinyqv.mem.q_ctrl.addr[5] ),
    .A2(net402),
    .Y(_05199_),
    .B1(net72));
 sg13g2_a221oi_1 _13317_ (.B2(_05198_),
    .C1(_05199_),
    .B1(net56),
    .A1(_01612_),
    .Y(_05200_),
    .A2(net278));
 sg13g2_a21o_1 _13318_ (.A2(net62),
    .A1(net3346),
    .B1(_05200_),
    .X(_01321_));
 sg13g2_nor2_1 _13319_ (.A(net3712),
    .B(_04304_),
    .Y(_05201_));
 sg13g2_nor2b_1 _13320_ (.A(net402),
    .B_N(\i_tinyqv.mem.q_ctrl.addr[10] ),
    .Y(_05202_));
 sg13g2_a21oi_1 _13321_ (.A1(net3457),
    .A2(net402),
    .Y(_05203_),
    .B1(_05202_));
 sg13g2_o21ai_1 _13322_ (.B1(_05191_),
    .Y(_05204_),
    .A1(_05190_),
    .A2(_05192_));
 sg13g2_and2_1 _13323_ (.A(\i_tinyqv.cpu.instr_data_start[10] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .X(_05205_));
 sg13g2_or2_1 _13324_ (.X(_05206_),
    .B(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .A(\i_tinyqv.cpu.instr_data_start[10] ));
 sg13g2_nand2b_1 _13325_ (.Y(_05207_),
    .B(_05206_),
    .A_N(_05205_));
 sg13g2_xnor2_1 _13326_ (.Y(_05208_),
    .A(_05204_),
    .B(_05207_));
 sg13g2_nor2_1 _13327_ (.A(\i_tinyqv.cpu.instr_data_start[10] ),
    .B(_05195_),
    .Y(_05209_));
 sg13g2_and2_1 _13328_ (.A(\i_tinyqv.cpu.instr_data_start[10] ),
    .B(_05195_),
    .X(_05210_));
 sg13g2_nor3_1 _13329_ (.A(net605),
    .B(_05209_),
    .C(_05210_),
    .Y(_05211_));
 sg13g2_a21oi_1 _13330_ (.A1(net605),
    .A2(_05208_),
    .Y(_05212_),
    .B1(_05211_));
 sg13g2_a221oi_1 _13331_ (.B2(net56),
    .C1(_05201_),
    .B1(_05212_),
    .A1(net71),
    .Y(_01322_),
    .A2(_05203_));
 sg13g2_nand2_1 _13332_ (.Y(_05213_),
    .A(\i_tinyqv.cpu.instr_data_start[11] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[11] ));
 sg13g2_xnor2_1 _13333_ (.Y(_05214_),
    .A(\i_tinyqv.cpu.instr_data_start[11] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[11] ));
 sg13g2_a21oi_1 _13334_ (.A1(_05204_),
    .A2(_05206_),
    .Y(_05215_),
    .B1(_05205_));
 sg13g2_xnor2_1 _13335_ (.Y(_05216_),
    .A(_05214_),
    .B(_05215_));
 sg13g2_nand2_1 _13336_ (.Y(_05217_),
    .A(net606),
    .B(_05216_));
 sg13g2_xnor2_1 _13337_ (.Y(_05218_),
    .A(_00239_),
    .B(_05210_));
 sg13g2_o21ai_1 _13338_ (.B1(_05217_),
    .Y(_05219_),
    .A1(net606),
    .A2(_05218_));
 sg13g2_a22oi_1 _13339_ (.Y(_05220_),
    .B1(net57),
    .B2(_05219_),
    .A2(net71),
    .A1(_01700_));
 sg13g2_o21ai_1 _13340_ (.B1(_05220_),
    .Y(_05221_),
    .A1(\addr[11] ),
    .A2(_04304_));
 sg13g2_nand2_1 _13341_ (.Y(_05222_),
    .A(net3019),
    .B(net61));
 sg13g2_o21ai_1 _13342_ (.B1(_05222_),
    .Y(_01323_),
    .A1(net61),
    .A2(_05221_));
 sg13g2_o21ai_1 _13343_ (.B1(_05213_),
    .Y(_05223_),
    .A1(_05214_),
    .A2(_05215_));
 sg13g2_and2_1 _13344_ (.A(\i_tinyqv.cpu.instr_data_start[12] ),
    .B(\i_tinyqv.cpu.imm[12] ),
    .X(_05224_));
 sg13g2_or2_1 _13345_ (.X(_05225_),
    .B(\i_tinyqv.cpu.imm[12] ),
    .A(\i_tinyqv.cpu.instr_data_start[12] ));
 sg13g2_nand2b_1 _13346_ (.Y(_05226_),
    .B(_05225_),
    .A_N(_05224_));
 sg13g2_xnor2_1 _13347_ (.Y(_05227_),
    .A(_05223_),
    .B(_05226_));
 sg13g2_and3_1 _13348_ (.X(_05228_),
    .A(\i_tinyqv.cpu.instr_data_start[12] ),
    .B(\i_tinyqv.cpu.instr_data_start[11] ),
    .C(_05210_));
 sg13g2_a21oi_1 _13349_ (.A1(\i_tinyqv.cpu.instr_data_start[11] ),
    .A2(_05210_),
    .Y(_05229_),
    .B1(\i_tinyqv.cpu.instr_data_start[12] ));
 sg13g2_nor3_1 _13350_ (.A(net605),
    .B(_05228_),
    .C(_05229_),
    .Y(_05230_));
 sg13g2_a21oi_1 _13351_ (.A1(net606),
    .A2(_05227_),
    .Y(_05231_),
    .B1(_05230_));
 sg13g2_a21oi_1 _13352_ (.A1(\i_tinyqv.mem.q_ctrl.addr[8] ),
    .A2(net402),
    .Y(_05232_),
    .B1(net72));
 sg13g2_a221oi_1 _13353_ (.B2(_05231_),
    .C1(_05232_),
    .B1(net56),
    .A1(_01613_),
    .Y(_05233_),
    .A2(net278));
 sg13g2_a21o_1 _13354_ (.A2(net62),
    .A1(net3441),
    .B1(_05233_),
    .X(_01324_));
 sg13g2_nand2_1 _13355_ (.Y(_05234_),
    .A(net614),
    .B(\i_tinyqv.cpu.imm[13] ));
 sg13g2_xnor2_1 _13356_ (.Y(_05235_),
    .A(net614),
    .B(\i_tinyqv.cpu.imm[13] ));
 sg13g2_a21oi_1 _13357_ (.A1(_05223_),
    .A2(_05225_),
    .Y(_05236_),
    .B1(_05224_));
 sg13g2_xor2_1 _13358_ (.B(_05236_),
    .A(_05235_),
    .X(_05237_));
 sg13g2_and2_1 _13359_ (.A(net614),
    .B(_05228_),
    .X(_05238_));
 sg13g2_o21ai_1 _13360_ (.B1(net477),
    .Y(_05239_),
    .A1(net614),
    .A2(_05228_));
 sg13g2_nor2_1 _13361_ (.A(_05238_),
    .B(_05239_),
    .Y(_05240_));
 sg13g2_a21oi_1 _13362_ (.A1(net605),
    .A2(_05237_),
    .Y(_05241_),
    .B1(_05240_));
 sg13g2_a21o_1 _13363_ (.A2(net402),
    .A1(net3346),
    .B1(net73),
    .X(_05242_));
 sg13g2_o21ai_1 _13364_ (.B1(_05242_),
    .Y(_05243_),
    .A1(\addr[13] ),
    .A2(_04304_));
 sg13g2_nand2_1 _13365_ (.Y(_05244_),
    .A(net3379),
    .B(net61));
 sg13g2_a22oi_1 _13366_ (.Y(_01325_),
    .B1(_05243_),
    .B2(_05244_),
    .A2(_05241_),
    .A1(net56));
 sg13g2_and2_1 _13367_ (.A(net613),
    .B(_05238_),
    .X(_05245_));
 sg13g2_o21ai_1 _13368_ (.B1(net478),
    .Y(_05246_),
    .A1(net613),
    .A2(_05238_));
 sg13g2_nor2_1 _13369_ (.A(_05245_),
    .B(_05246_),
    .Y(_05247_));
 sg13g2_o21ai_1 _13370_ (.B1(_05234_),
    .Y(_05248_),
    .A1(_05235_),
    .A2(_05236_));
 sg13g2_xnor2_1 _13371_ (.Y(_05249_),
    .A(net613),
    .B(\i_tinyqv.cpu.imm[14] ));
 sg13g2_xnor2_1 _13372_ (.Y(_05250_),
    .A(_05248_),
    .B(_05249_));
 sg13g2_a21oi_1 _13373_ (.A1(net605),
    .A2(_05250_),
    .Y(_05251_),
    .B1(_05247_));
 sg13g2_a22oi_1 _13374_ (.Y(_05252_),
    .B1(net278),
    .B2(\addr[14] ),
    .A2(net71),
    .A1(\i_tinyqv.mem.q_ctrl.addr[10] ));
 sg13g2_o21ai_1 _13375_ (.B1(_05252_),
    .Y(_05253_),
    .A1(_05126_),
    .A2(_05251_));
 sg13g2_mux2_1 _13376_ (.A0(net3253),
    .A1(_05253_),
    .S(_04300_),
    .X(_01326_));
 sg13g2_and2_1 _13377_ (.A(\i_tinyqv.cpu.instr_data_start[15] ),
    .B(_05245_),
    .X(_05254_));
 sg13g2_o21ai_1 _13378_ (.B1(net478),
    .Y(_05255_),
    .A1(\i_tinyqv.cpu.instr_data_start[15] ),
    .A2(_05245_));
 sg13g2_nor2_1 _13379_ (.A(_05254_),
    .B(_05255_),
    .Y(_05256_));
 sg13g2_nand2_1 _13380_ (.Y(_05257_),
    .A(\i_tinyqv.cpu.instr_data_start[15] ),
    .B(\i_tinyqv.cpu.imm[15] ));
 sg13g2_xnor2_1 _13381_ (.Y(_05258_),
    .A(\i_tinyqv.cpu.instr_data_start[15] ),
    .B(\i_tinyqv.cpu.imm[15] ));
 sg13g2_a21o_1 _13382_ (.A2(\i_tinyqv.cpu.imm[14] ),
    .A1(net613),
    .B1(_05248_),
    .X(_05259_));
 sg13g2_o21ai_1 _13383_ (.B1(_05259_),
    .Y(_05260_),
    .A1(net613),
    .A2(\i_tinyqv.cpu.imm[14] ));
 sg13g2_xor2_1 _13384_ (.B(_05260_),
    .A(_05258_),
    .X(_05261_));
 sg13g2_a21oi_1 _13385_ (.A1(net607),
    .A2(_05261_),
    .Y(_05262_),
    .B1(_05256_));
 sg13g2_a21oi_1 _13386_ (.A1(net3019),
    .A2(net402),
    .Y(_05263_),
    .B1(net72));
 sg13g2_a21oi_1 _13387_ (.A1(net56),
    .A2(_05262_),
    .Y(_05264_),
    .B1(_05263_));
 sg13g2_o21ai_1 _13388_ (.B1(_05264_),
    .Y(_05265_),
    .A1(\addr[15] ),
    .A2(_04304_));
 sg13g2_o21ai_1 _13389_ (.B1(_05265_),
    .Y(_01327_),
    .A1(_01701_),
    .A2(_04300_));
 sg13g2_a22oi_1 _13390_ (.Y(_05266_),
    .B1(net278),
    .B2(\addr[16] ),
    .A2(net70),
    .A1(net3441));
 sg13g2_xnor2_1 _13391_ (.Y(_05267_),
    .A(\i_tinyqv.cpu.instr_data_start[16] ),
    .B(_05254_));
 sg13g2_o21ai_1 _13392_ (.B1(_05257_),
    .Y(_05268_),
    .A1(_05258_),
    .A2(_05260_));
 sg13g2_xnor2_1 _13393_ (.Y(_05269_),
    .A(net612),
    .B(\i_tinyqv.cpu.imm[16] ));
 sg13g2_xnor2_1 _13394_ (.Y(_05270_),
    .A(_05268_),
    .B(_05269_));
 sg13g2_nor2_1 _13395_ (.A(net477),
    .B(_05270_),
    .Y(_05271_));
 sg13g2_a21oi_1 _13396_ (.A1(net477),
    .A2(_05267_),
    .Y(_05272_),
    .B1(_05271_));
 sg13g2_a22oi_1 _13397_ (.Y(_05273_),
    .B1(net56),
    .B2(_05272_),
    .A2(net61),
    .A1(net3500));
 sg13g2_o21ai_1 _13398_ (.B1(_05273_),
    .Y(_01328_),
    .A1(net61),
    .A2(_05266_));
 sg13g2_a21oi_1 _13399_ (.A1(\i_tinyqv.cpu.instr_data_start[16] ),
    .A2(_05254_),
    .Y(_05274_),
    .B1(net611));
 sg13g2_and3_1 _13400_ (.X(_05275_),
    .A(net611),
    .B(\i_tinyqv.cpu.instr_data_start[16] ),
    .C(_05254_));
 sg13g2_nand2_1 _13401_ (.Y(_05276_),
    .A(net611),
    .B(\i_tinyqv.cpu.imm[17] ));
 sg13g2_nor2_1 _13402_ (.A(net611),
    .B(\i_tinyqv.cpu.imm[17] ),
    .Y(_05277_));
 sg13g2_xor2_1 _13403_ (.B(\i_tinyqv.cpu.imm[17] ),
    .A(net611),
    .X(_05278_));
 sg13g2_a21o_1 _13404_ (.A2(\i_tinyqv.cpu.imm[16] ),
    .A1(net612),
    .B1(_05268_),
    .X(_05279_));
 sg13g2_o21ai_1 _13405_ (.B1(_05279_),
    .Y(_05280_),
    .A1(net612),
    .A2(\i_tinyqv.cpu.imm[16] ));
 sg13g2_xnor2_1 _13406_ (.Y(_05281_),
    .A(_05278_),
    .B(_05280_));
 sg13g2_nor3_1 _13407_ (.A(net607),
    .B(_05274_),
    .C(_05275_),
    .Y(_05282_));
 sg13g2_a21oi_1 _13408_ (.A1(net607),
    .A2(_05281_),
    .Y(_05283_),
    .B1(_05282_));
 sg13g2_or2_1 _13409_ (.X(_05284_),
    .B(_05283_),
    .A(_05126_));
 sg13g2_a221oi_1 _13410_ (.B2(\addr[17] ),
    .C1(net61),
    .B1(net278),
    .A1(net3379),
    .Y(_05285_),
    .A2(net70));
 sg13g2_a22oi_1 _13411_ (.Y(_01329_),
    .B1(_05284_),
    .B2(_05285_),
    .A2(net61),
    .A1(_01702_));
 sg13g2_nand2_1 _13412_ (.Y(_05286_),
    .A(net3319),
    .B(net277));
 sg13g2_and2_1 _13413_ (.A(\i_tinyqv.cpu.instr_data_start[18] ),
    .B(_05275_),
    .X(_05287_));
 sg13g2_xnor2_1 _13414_ (.Y(_05288_),
    .A(_01513_),
    .B(_05275_));
 sg13g2_nor2_1 _13415_ (.A(net603),
    .B(_05288_),
    .Y(_05289_));
 sg13g2_o21ai_1 _13416_ (.B1(_05276_),
    .Y(_05290_),
    .A1(_05277_),
    .A2(_05280_));
 sg13g2_and2_1 _13417_ (.A(\i_tinyqv.cpu.instr_data_start[18] ),
    .B(\i_tinyqv.cpu.imm[18] ),
    .X(_05291_));
 sg13g2_or2_1 _13418_ (.X(_05292_),
    .B(\i_tinyqv.cpu.imm[18] ),
    .A(\i_tinyqv.cpu.instr_data_start[18] ));
 sg13g2_nor2b_1 _13419_ (.A(_05291_),
    .B_N(_05292_),
    .Y(_05293_));
 sg13g2_xnor2_1 _13420_ (.Y(_05294_),
    .A(_05290_),
    .B(_05293_));
 sg13g2_a21oi_1 _13421_ (.A1(net603),
    .A2(_05294_),
    .Y(_05295_),
    .B1(_05289_));
 sg13g2_a221oi_1 _13422_ (.B2(_05295_),
    .C1(net60),
    .B1(net58),
    .A1(net3253),
    .Y(_05296_),
    .A2(net71));
 sg13g2_a22oi_1 _13423_ (.Y(_01330_),
    .B1(_05286_),
    .B2(_05296_),
    .A2(net60),
    .A1(_01703_));
 sg13g2_nand2_1 _13424_ (.Y(_05297_),
    .A(\i_tinyqv.cpu.instr_data_start[19] ),
    .B(\i_tinyqv.cpu.imm[19] ));
 sg13g2_nor2_1 _13425_ (.A(\i_tinyqv.cpu.instr_data_start[19] ),
    .B(\i_tinyqv.cpu.imm[19] ),
    .Y(_05298_));
 sg13g2_xor2_1 _13426_ (.B(\i_tinyqv.cpu.imm[19] ),
    .A(\i_tinyqv.cpu.instr_data_start[19] ),
    .X(_05299_));
 sg13g2_a21oi_1 _13427_ (.A1(_05290_),
    .A2(_05292_),
    .Y(_05300_),
    .B1(_05291_));
 sg13g2_xnor2_1 _13428_ (.Y(_05301_),
    .A(_05299_),
    .B(_05300_));
 sg13g2_nand2_1 _13429_ (.Y(_05302_),
    .A(net602),
    .B(_05301_));
 sg13g2_and2_1 _13430_ (.A(\i_tinyqv.cpu.instr_data_start[19] ),
    .B(_05287_),
    .X(_05303_));
 sg13g2_o21ai_1 _13431_ (.B1(net477),
    .Y(_05304_),
    .A1(\i_tinyqv.cpu.instr_data_start[19] ),
    .A2(_05287_));
 sg13g2_o21ai_1 _13432_ (.B1(_05302_),
    .Y(_05305_),
    .A1(_05303_),
    .A2(_05304_));
 sg13g2_nand2_1 _13433_ (.Y(_05306_),
    .A(net3321),
    .B(net277));
 sg13g2_a221oi_1 _13434_ (.B2(_05305_),
    .C1(net60),
    .B1(net58),
    .A1(\i_tinyqv.mem.q_ctrl.addr[15] ),
    .Y(_05307_),
    .A2(net71));
 sg13g2_a22oi_1 _13435_ (.Y(_01331_),
    .B1(_05306_),
    .B2(_05307_),
    .A2(net60),
    .A1(_01704_));
 sg13g2_o21ai_1 _13436_ (.B1(_05297_),
    .Y(_05308_),
    .A1(_05298_),
    .A2(_05300_));
 sg13g2_and2_1 _13437_ (.A(net610),
    .B(\i_tinyqv.cpu.imm[20] ),
    .X(_05309_));
 sg13g2_or2_1 _13438_ (.X(_05310_),
    .B(\i_tinyqv.cpu.imm[20] ),
    .A(net610));
 sg13g2_nor2b_1 _13439_ (.A(_05309_),
    .B_N(_05310_),
    .Y(_05311_));
 sg13g2_xnor2_1 _13440_ (.Y(_05312_),
    .A(_05308_),
    .B(_05311_));
 sg13g2_nand2b_1 _13441_ (.Y(_05313_),
    .B(_05287_),
    .A_N(_00207_));
 sg13g2_xnor2_1 _13442_ (.Y(_05314_),
    .A(net610),
    .B(_05313_));
 sg13g2_nor2_1 _13443_ (.A(net602),
    .B(_05314_),
    .Y(_05315_));
 sg13g2_a21oi_1 _13444_ (.A1(net603),
    .A2(_05312_),
    .Y(_05316_),
    .B1(_05315_));
 sg13g2_a22oi_1 _13445_ (.Y(_05317_),
    .B1(net277),
    .B2(net3496),
    .A2(net401),
    .A1(net3500));
 sg13g2_a22oi_1 _13446_ (.Y(_05318_),
    .B1(net58),
    .B2(_05316_),
    .A2(net59),
    .A1(net3632));
 sg13g2_nand2_1 _13447_ (.Y(_01332_),
    .A(_05317_),
    .B(_05318_));
 sg13g2_nand2_1 _13448_ (.Y(_05319_),
    .A(net609),
    .B(\i_tinyqv.cpu.imm[21] ));
 sg13g2_nor2_1 _13449_ (.A(net609),
    .B(\i_tinyqv.cpu.imm[21] ),
    .Y(_05320_));
 sg13g2_xor2_1 _13450_ (.B(\i_tinyqv.cpu.imm[21] ),
    .A(net609),
    .X(_05321_));
 sg13g2_a21oi_1 _13451_ (.A1(_05308_),
    .A2(_05310_),
    .Y(_05322_),
    .B1(_05309_));
 sg13g2_xnor2_1 _13452_ (.Y(_05323_),
    .A(_05321_),
    .B(_05322_));
 sg13g2_a21oi_1 _13453_ (.A1(net610),
    .A2(_05303_),
    .Y(_05324_),
    .B1(\i_tinyqv.cpu.instr_data_start[21] ));
 sg13g2_and3_1 _13454_ (.X(_05325_),
    .A(\i_tinyqv.cpu.instr_data_start[21] ),
    .B(\i_tinyqv.cpu.instr_data_start[20] ),
    .C(_05303_));
 sg13g2_nor3_1 _13455_ (.A(net602),
    .B(_05324_),
    .C(_05325_),
    .Y(_05326_));
 sg13g2_a21oi_1 _13456_ (.A1(net602),
    .A2(_05323_),
    .Y(_05327_),
    .B1(_05326_));
 sg13g2_a21oi_1 _13457_ (.A1(\i_tinyqv.mem.q_ctrl.addr[17] ),
    .A2(net401),
    .Y(_05328_),
    .B1(net72));
 sg13g2_a221oi_1 _13458_ (.B2(_05327_),
    .C1(_05328_),
    .B1(net58),
    .A1(_01615_),
    .Y(_05329_),
    .A2(net277));
 sg13g2_a21o_1 _13459_ (.A2(net59),
    .A1(net3393),
    .B1(_05329_),
    .X(_01333_));
 sg13g2_o21ai_1 _13460_ (.B1(_05319_),
    .Y(_05330_),
    .A1(_05320_),
    .A2(_05322_));
 sg13g2_and2_1 _13461_ (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(\i_tinyqv.cpu.imm[22] ),
    .X(_05331_));
 sg13g2_or2_1 _13462_ (.X(_05332_),
    .B(\i_tinyqv.cpu.imm[22] ),
    .A(\i_tinyqv.cpu.instr_data_start[22] ));
 sg13g2_nand2b_1 _13463_ (.Y(_05333_),
    .B(_05332_),
    .A_N(_05331_));
 sg13g2_xnor2_1 _13464_ (.Y(_05334_),
    .A(_05330_),
    .B(_05333_));
 sg13g2_nand2_1 _13465_ (.Y(_05335_),
    .A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(_05325_));
 sg13g2_nor2_1 _13466_ (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(_05325_),
    .Y(_05336_));
 sg13g2_nor2_1 _13467_ (.A(net602),
    .B(_05336_),
    .Y(_05337_));
 sg13g2_a221oi_1 _13468_ (.B2(_05337_),
    .C1(_05126_),
    .B1(_05335_),
    .A1(net602),
    .Y(_05338_),
    .A2(_05334_));
 sg13g2_nor2b_1 _13469_ (.A(net401),
    .B_N(\i_tinyqv.mem.q_ctrl.addr[22] ),
    .Y(_05339_));
 sg13g2_a21oi_1 _13470_ (.A1(net3735),
    .A2(net401),
    .Y(_05340_),
    .B1(_05339_));
 sg13g2_a221oi_1 _13471_ (.B2(net70),
    .C1(_05338_),
    .B1(net3736),
    .A1(_01614_),
    .Y(_01334_),
    .A2(net277));
 sg13g2_xnor2_1 _13472_ (.Y(_05341_),
    .A(_00202_),
    .B(_05335_));
 sg13g2_a21oi_1 _13473_ (.A1(_05330_),
    .A2(_05332_),
    .Y(_05342_),
    .B1(_05331_));
 sg13g2_xor2_1 _13474_ (.B(\i_tinyqv.cpu.imm[23] ),
    .A(\i_tinyqv.cpu.instr_data_start[23] ),
    .X(_05343_));
 sg13g2_xnor2_1 _13475_ (.Y(_05344_),
    .A(_05342_),
    .B(_05343_));
 sg13g2_o21ai_1 _13476_ (.B1(net58),
    .Y(_05345_),
    .A1(net602),
    .A2(_05341_));
 sg13g2_a21oi_1 _13477_ (.A1(net602),
    .A2(_05344_),
    .Y(_05346_),
    .B1(_05345_));
 sg13g2_a22oi_1 _13478_ (.Y(_05347_),
    .B1(net277),
    .B2(net3666),
    .A2(net401),
    .A1(_01704_));
 sg13g2_o21ai_1 _13479_ (.B1(_05347_),
    .Y(_05348_),
    .A1(net3706),
    .A2(_04300_));
 sg13g2_nor2_1 _13480_ (.A(_05346_),
    .B(net3707),
    .Y(_01335_));
 sg13g2_and2_1 _13481_ (.A(_03503_),
    .B(net69),
    .X(_05349_));
 sg13g2_nand2_1 _13482_ (.Y(_05350_),
    .A(_03503_),
    .B(net69));
 sg13g2_a21oi_1 _13483_ (.A1(_03252_),
    .A2(net69),
    .Y(_05351_),
    .B1(_05112_));
 sg13g2_o21ai_1 _13484_ (.B1(net656),
    .Y(_05352_),
    .A1(net4052),
    .A2(net50));
 sg13g2_a21oi_1 _13485_ (.A1(net50),
    .A2(_05351_),
    .Y(_01336_),
    .B1(_05352_));
 sg13g2_o21ai_1 _13486_ (.B1(net69),
    .Y(_05353_),
    .A1(_03371_),
    .A2(_03503_));
 sg13g2_o21ai_1 _13487_ (.B1(net656),
    .Y(_05354_),
    .A1(net4077),
    .A2(net50));
 sg13g2_a21oi_1 _13488_ (.A1(_05121_),
    .A2(_05353_),
    .Y(_01337_),
    .B1(_05354_));
 sg13g2_nand2_1 _13489_ (.Y(_05355_),
    .A(net3251),
    .B(net171));
 sg13g2_o21ai_1 _13490_ (.B1(_05355_),
    .Y(_01338_),
    .A1(_01511_),
    .A2(net171));
 sg13g2_nor2_1 _13491_ (.A(net601),
    .B(net169),
    .Y(_05356_));
 sg13g2_a21oi_1 _13492_ (.A1(_01646_),
    .A2(net171),
    .Y(_01339_),
    .B1(_05356_));
 sg13g2_nor2_1 _13493_ (.A(net600),
    .B(net169),
    .Y(_05357_));
 sg13g2_a21oi_1 _13494_ (.A1(_01645_),
    .A2(net170),
    .Y(_01340_),
    .B1(_05357_));
 sg13g2_nand2_1 _13495_ (.Y(_05358_),
    .A(net3506),
    .B(net169));
 sg13g2_o21ai_1 _13496_ (.B1(_05358_),
    .Y(_01341_),
    .A1(_01508_),
    .A2(net169));
 sg13g2_nor2_1 _13497_ (.A(net599),
    .B(net169),
    .Y(_05359_));
 sg13g2_a21oi_1 _13498_ (.A1(_01644_),
    .A2(net169),
    .Y(_01342_),
    .B1(_05359_));
 sg13g2_nand2_1 _13499_ (.Y(_05360_),
    .A(net3376),
    .B(net169));
 sg13g2_o21ai_1 _13500_ (.B1(_05360_),
    .Y(_01343_),
    .A1(_01506_),
    .A2(net169));
 sg13g2_nor2_1 _13501_ (.A(net597),
    .B(net170),
    .Y(_05361_));
 sg13g2_a21oi_1 _13502_ (.A1(_01643_),
    .A2(net170),
    .Y(_01344_),
    .B1(_05361_));
 sg13g2_nor2_1 _13503_ (.A(\data_to_write[7] ),
    .B(net170),
    .Y(_05362_));
 sg13g2_a21oi_1 _13504_ (.A1(_01642_),
    .A2(net170),
    .Y(_01345_),
    .B1(_05362_));
 sg13g2_nor2_1 _13505_ (.A(\data_to_write[8] ),
    .B(net168),
    .Y(_05363_));
 sg13g2_a21oi_1 _13506_ (.A1(_01641_),
    .A2(net168),
    .Y(_01346_),
    .B1(_05363_));
 sg13g2_mux2_1 _13507_ (.A0(\data_to_write[9] ),
    .A1(net3830),
    .S(net170),
    .X(_01347_));
 sg13g2_mux2_1 _13508_ (.A0(\data_to_write[10] ),
    .A1(net3778),
    .S(net170),
    .X(_01348_));
 sg13g2_mux2_1 _13509_ (.A0(\data_to_write[11] ),
    .A1(net3747),
    .S(net168),
    .X(_01349_));
 sg13g2_nor2_1 _13510_ (.A(net3800),
    .B(net171),
    .Y(_05364_));
 sg13g2_a21oi_1 _13511_ (.A1(_01638_),
    .A2(net167),
    .Y(_01350_),
    .B1(_05364_));
 sg13g2_nor2_1 _13512_ (.A(\data_to_write[13] ),
    .B(net167),
    .Y(_05365_));
 sg13g2_a21oi_1 _13513_ (.A1(_01637_),
    .A2(net176),
    .Y(_01351_),
    .B1(_05365_));
 sg13g2_nor2_1 _13514_ (.A(\data_to_write[14] ),
    .B(net168),
    .Y(_05366_));
 sg13g2_a21oi_1 _13515_ (.A1(_01636_),
    .A2(net168),
    .Y(_01352_),
    .B1(_05366_));
 sg13g2_nor2_1 _13516_ (.A(\data_to_write[15] ),
    .B(net168),
    .Y(_05367_));
 sg13g2_a21oi_1 _13517_ (.A1(_01635_),
    .A2(net168),
    .Y(_01353_),
    .B1(_05367_));
 sg13g2_nand2_1 _13518_ (.Y(_05368_),
    .A(net85),
    .B(_03723_));
 sg13g2_nand2_1 _13519_ (.Y(_05369_),
    .A(net2826),
    .B(net78));
 sg13g2_nand3_1 _13520_ (.B(_05368_),
    .C(_05369_),
    .A(net91),
    .Y(_05370_));
 sg13g2_nor2_1 _13521_ (.A(net414),
    .B(_04732_),
    .Y(_05371_));
 sg13g2_a21oi_1 _13522_ (.A1(net414),
    .A2(_05134_),
    .Y(_05372_),
    .B1(_05371_));
 sg13g2_a21oi_1 _13523_ (.A1(net95),
    .A2(_05372_),
    .Y(_05373_),
    .B1(net51));
 sg13g2_a22oi_1 _13524_ (.Y(_05374_),
    .B1(_05370_),
    .B2(_05373_),
    .A2(net51),
    .A1(net4111));
 sg13g2_nor2_1 _13525_ (.A(net512),
    .B(_05374_),
    .Y(_01354_));
 sg13g2_mux2_1 _13526_ (.A0(_03016_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .S(net78),
    .X(_05375_));
 sg13g2_mux2_1 _13527_ (.A0(_04736_),
    .A1(_05143_),
    .S(net414),
    .X(_05376_));
 sg13g2_a21oi_1 _13528_ (.A1(net95),
    .A2(_05376_),
    .Y(_05377_),
    .B1(net51));
 sg13g2_o21ai_1 _13529_ (.B1(_05377_),
    .Y(_05378_),
    .A1(net95),
    .A2(_05375_));
 sg13g2_nand2_1 _13530_ (.Y(_05379_),
    .A(net3895),
    .B(net51));
 sg13g2_a21oi_1 _13531_ (.A1(_05378_),
    .A2(_05379_),
    .Y(_01355_),
    .B1(net512));
 sg13g2_nor2_2 _13532_ (.A(net411),
    .B(_04739_),
    .Y(_05380_));
 sg13g2_a21oi_1 _13533_ (.A1(net414),
    .A2(_05152_),
    .Y(_05381_),
    .B1(_05380_));
 sg13g2_nor2_1 _13534_ (.A(net3981),
    .B(net50),
    .Y(_05382_));
 sg13g2_nand2_1 _13535_ (.Y(_05383_),
    .A(net2798),
    .B(net78));
 sg13g2_o21ai_1 _13536_ (.B1(_05383_),
    .Y(_05384_),
    .A1(_03251_),
    .A2(net78));
 sg13g2_o21ai_1 _13537_ (.B1(net50),
    .Y(_05385_),
    .A1(net91),
    .A2(_05381_));
 sg13g2_a21oi_1 _13538_ (.A1(net94),
    .A2(_05384_),
    .Y(_05386_),
    .B1(_05385_));
 sg13g2_nor3_1 _13539_ (.A(net512),
    .B(_05382_),
    .C(_05386_),
    .Y(_01356_));
 sg13g2_mux2_1 _13540_ (.A0(_03378_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .S(net78),
    .X(_05387_));
 sg13g2_mux2_1 _13541_ (.A0(_04742_),
    .A1(_05164_),
    .S(net412),
    .X(_05388_));
 sg13g2_a21oi_1 _13542_ (.A1(net95),
    .A2(_05388_),
    .Y(_05389_),
    .B1(net54));
 sg13g2_o21ai_1 _13543_ (.B1(_05389_),
    .Y(_05390_),
    .A1(net98),
    .A2(_05387_));
 sg13g2_nand2_1 _13544_ (.Y(_05391_),
    .A(net3967),
    .B(net54));
 sg13g2_a21oi_1 _13545_ (.A1(_05390_),
    .A2(_05391_),
    .Y(_01357_),
    .B1(net511));
 sg13g2_mux2_1 _13546_ (.A0(_04744_),
    .A1(_05175_),
    .S(net413),
    .X(_05392_));
 sg13g2_a21oi_1 _13547_ (.A1(net85),
    .A2(_03721_),
    .Y(_05393_),
    .B1(net95));
 sg13g2_nand2_1 _13548_ (.Y(_05394_),
    .A(net2809),
    .B(net78));
 sg13g2_a22oi_1 _13549_ (.Y(_05395_),
    .B1(_05393_),
    .B2(_05394_),
    .A2(_05392_),
    .A1(net98));
 sg13g2_o21ai_1 _13550_ (.B1(net659),
    .Y(_05396_),
    .A1(net54),
    .A2(_05395_));
 sg13g2_a21oi_1 _13551_ (.A1(_01518_),
    .A2(net54),
    .Y(_01358_),
    .B1(_05396_));
 sg13g2_a21oi_1 _13552_ (.A1(_03013_),
    .A2(net85),
    .Y(_05397_),
    .B1(net97));
 sg13g2_nand2_1 _13553_ (.Y(_05398_),
    .A(net2817),
    .B(net79));
 sg13g2_nor2_1 _13554_ (.A(net413),
    .B(_04748_),
    .Y(_05399_));
 sg13g2_a21oi_1 _13555_ (.A1(net412),
    .A2(_05184_),
    .Y(_05400_),
    .B1(_05399_));
 sg13g2_a221oi_1 _13556_ (.B2(net97),
    .C1(net53),
    .B1(_05400_),
    .A1(_05397_),
    .Y(_05401_),
    .A2(_05398_));
 sg13g2_a21oi_1 _13557_ (.A1(net3986),
    .A2(net55),
    .Y(_05402_),
    .B1(_05401_));
 sg13g2_nor2_1 _13558_ (.A(net511),
    .B(_05402_),
    .Y(_01359_));
 sg13g2_a21oi_1 _13559_ (.A1(_03255_),
    .A2(net85),
    .Y(_05403_),
    .B1(net95));
 sg13g2_nand2_1 _13560_ (.Y(_05404_),
    .A(net2793),
    .B(net78));
 sg13g2_nor2_1 _13561_ (.A(net413),
    .B(_04750_),
    .Y(_05405_));
 sg13g2_a21oi_2 _13562_ (.B1(_05405_),
    .Y(_05406_),
    .A2(_05194_),
    .A1(net412));
 sg13g2_a22oi_1 _13563_ (.Y(_05407_),
    .B1(_05406_),
    .B2(net95),
    .A2(_05404_),
    .A1(_05403_));
 sg13g2_o21ai_1 _13564_ (.B1(net659),
    .Y(_05408_),
    .A1(net54),
    .A2(_05407_));
 sg13g2_a21oi_1 _13565_ (.A1(_01517_),
    .A2(net54),
    .Y(_01360_),
    .B1(_05408_));
 sg13g2_a21oi_1 _13566_ (.A1(_03376_),
    .A2(net86),
    .Y(_05409_),
    .B1(net97));
 sg13g2_nand2_1 _13567_ (.Y(_05410_),
    .A(net2806),
    .B(net79));
 sg13g2_nand2_1 _13568_ (.Y(_05411_),
    .A(net412),
    .B(_05208_));
 sg13g2_a21oi_1 _13569_ (.A1(net409),
    .A2(_04753_),
    .Y(_05412_),
    .B1(net93));
 sg13g2_a22oi_1 _13570_ (.Y(_05413_),
    .B1(_05411_),
    .B2(_05412_),
    .A2(_05410_),
    .A1(_05409_));
 sg13g2_o21ai_1 _13571_ (.B1(net659),
    .Y(_05414_),
    .A1(net54),
    .A2(_05413_));
 sg13g2_a21oi_1 _13572_ (.A1(_01516_),
    .A2(net53),
    .Y(_01361_),
    .B1(_05414_));
 sg13g2_a21oi_1 _13573_ (.A1(net85),
    .A2(_03725_),
    .Y(_05415_),
    .B1(net97));
 sg13g2_nand2_1 _13574_ (.Y(_05416_),
    .A(net2797),
    .B(net79));
 sg13g2_nor2_1 _13575_ (.A(net409),
    .B(_05216_),
    .Y(_05417_));
 sg13g2_a21oi_1 _13576_ (.A1(net408),
    .A2(_04754_),
    .Y(_05418_),
    .B1(_05417_));
 sg13g2_a221oi_1 _13577_ (.B2(net96),
    .C1(net53),
    .B1(_05418_),
    .A1(_05415_),
    .Y(_05419_),
    .A2(_05416_));
 sg13g2_a21oi_1 _13578_ (.A1(net3979),
    .A2(net55),
    .Y(_05420_),
    .B1(_05419_));
 sg13g2_nor2_1 _13579_ (.A(net512),
    .B(_05420_),
    .Y(_01362_));
 sg13g2_a21oi_1 _13580_ (.A1(_03011_),
    .A2(net85),
    .Y(_05421_),
    .B1(net96));
 sg13g2_nand2_1 _13581_ (.Y(_05422_),
    .A(net2799),
    .B(net79));
 sg13g2_nand2_1 _13582_ (.Y(_05423_),
    .A(net412),
    .B(_05227_));
 sg13g2_a21oi_1 _13583_ (.A1(net409),
    .A2(_04755_),
    .Y(_05424_),
    .B1(net93));
 sg13g2_a22oi_1 _13584_ (.Y(_05425_),
    .B1(_05423_),
    .B2(_05424_),
    .A2(_05422_),
    .A1(_05421_));
 sg13g2_o21ai_1 _13585_ (.B1(net659),
    .Y(_05426_),
    .A1(net53),
    .A2(_05425_));
 sg13g2_a21oi_1 _13586_ (.A1(_01515_),
    .A2(net53),
    .Y(_01363_),
    .B1(_05426_));
 sg13g2_nand2_1 _13587_ (.Y(_05427_),
    .A(net412),
    .B(_05237_));
 sg13g2_o21ai_1 _13588_ (.B1(_05427_),
    .Y(_05428_),
    .A1(net412),
    .A2(_04759_));
 sg13g2_nand2_1 _13589_ (.Y(_05429_),
    .A(net2821),
    .B(net78));
 sg13g2_o21ai_1 _13590_ (.B1(_05429_),
    .Y(_05430_),
    .A1(_03250_),
    .A2(net79));
 sg13g2_nand2_1 _13591_ (.Y(_05431_),
    .A(net93),
    .B(_05430_));
 sg13g2_a21oi_1 _13592_ (.A1(net97),
    .A2(_05428_),
    .Y(_05432_),
    .B1(net53));
 sg13g2_o21ai_1 _13593_ (.B1(net658),
    .Y(_05433_),
    .A1(net3734),
    .A2(net49));
 sg13g2_a21oi_1 _13594_ (.A1(_05431_),
    .A2(_05432_),
    .Y(_01364_),
    .B1(_05433_));
 sg13g2_a21oi_1 _13595_ (.A1(_03373_),
    .A2(net77),
    .Y(_05434_),
    .B1(net96));
 sg13g2_nand2_1 _13596_ (.Y(_05435_),
    .A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .B(net79));
 sg13g2_nand2_1 _13597_ (.Y(_05436_),
    .A(net412),
    .B(_05250_));
 sg13g2_a21oi_1 _13598_ (.A1(net409),
    .A2(_04760_),
    .Y(_05437_),
    .B1(net93));
 sg13g2_a221oi_1 _13599_ (.B2(_05437_),
    .C1(net53),
    .B1(_05436_),
    .A1(_05434_),
    .Y(_05438_),
    .A2(_05435_));
 sg13g2_a21o_1 _13600_ (.A2(net53),
    .A1(net4014),
    .B1(_05438_),
    .X(_05439_));
 sg13g2_and2_1 _13601_ (.A(net657),
    .B(_05439_),
    .X(_01365_));
 sg13g2_nor2_1 _13602_ (.A(net409),
    .B(_05261_),
    .Y(_05440_));
 sg13g2_a21oi_1 _13603_ (.A1(net408),
    .A2(_04762_),
    .Y(_05441_),
    .B1(_05440_));
 sg13g2_a21oi_1 _13604_ (.A1(net96),
    .A2(_05441_),
    .Y(_05442_),
    .B1(net51));
 sg13g2_a21oi_1 _13605_ (.A1(net85),
    .A2(_03720_),
    .Y(_05443_),
    .B1(net95));
 sg13g2_o21ai_1 _13606_ (.B1(_05443_),
    .Y(_05444_),
    .A1(net2824),
    .A2(net77));
 sg13g2_a221oi_1 _13607_ (.B2(_05444_),
    .C1(net512),
    .B1(_05442_),
    .A1(_01514_),
    .Y(_01366_),
    .A2(net52));
 sg13g2_a21oi_1 _13608_ (.A1(_03008_),
    .A2(net85),
    .Y(_05445_),
    .B1(net96));
 sg13g2_o21ai_1 _13609_ (.B1(_05445_),
    .Y(_05446_),
    .A1(net2816),
    .A2(net76));
 sg13g2_mux2_1 _13610_ (.A0(_04764_),
    .A1(_05270_),
    .S(net413),
    .X(_05447_));
 sg13g2_a21oi_1 _13611_ (.A1(net96),
    .A2(_05447_),
    .Y(_05448_),
    .B1(net52));
 sg13g2_o21ai_1 _13612_ (.B1(net657),
    .Y(_05449_),
    .A1(net612),
    .A2(net50));
 sg13g2_a21oi_1 _13613_ (.A1(_05446_),
    .A2(_05448_),
    .Y(_01367_),
    .B1(_05449_));
 sg13g2_a21oi_1 _13614_ (.A1(net411),
    .A2(_05281_),
    .Y(_05450_),
    .B1(net92));
 sg13g2_o21ai_1 _13615_ (.B1(_05450_),
    .Y(_05451_),
    .A1(net413),
    .A2(_04767_));
 sg13g2_nor2_1 _13616_ (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .B(net76),
    .Y(_05452_));
 sg13g2_a21oi_1 _13617_ (.A1(_03248_),
    .A2(net76),
    .Y(_05453_),
    .B1(_05452_));
 sg13g2_o21ai_1 _13618_ (.B1(_05451_),
    .Y(_05454_),
    .A1(net96),
    .A2(_05453_));
 sg13g2_o21ai_1 _13619_ (.B1(net657),
    .Y(_05455_),
    .A1(net3826),
    .A2(net49));
 sg13g2_a21oi_1 _13620_ (.A1(net49),
    .A2(_05454_),
    .Y(_01368_),
    .B1(_05455_));
 sg13g2_a21oi_1 _13621_ (.A1(net408),
    .A2(_04768_),
    .Y(_05456_),
    .B1(net92));
 sg13g2_o21ai_1 _13622_ (.B1(_05456_),
    .Y(_05457_),
    .A1(net408),
    .A2(_05294_));
 sg13g2_nand2_1 _13623_ (.Y(_05458_),
    .A(_03368_),
    .B(net86));
 sg13g2_a21oi_1 _13624_ (.A1(net2808),
    .A2(net79),
    .Y(_05459_),
    .B1(net96));
 sg13g2_a21oi_1 _13625_ (.A1(_05458_),
    .A2(_05459_),
    .Y(_05460_),
    .B1(net52));
 sg13g2_a22oi_1 _13626_ (.Y(_05461_),
    .B1(_05457_),
    .B2(_05460_),
    .A2(net51),
    .A1(net3931));
 sg13g2_nor2_1 _13627_ (.A(net512),
    .B(_05461_),
    .Y(_01369_));
 sg13g2_nor2_1 _13628_ (.A(net411),
    .B(_04769_),
    .Y(_05462_));
 sg13g2_nor2_1 _13629_ (.A(net92),
    .B(_05462_),
    .Y(_05463_));
 sg13g2_o21ai_1 _13630_ (.B1(_05463_),
    .Y(_05464_),
    .A1(net408),
    .A2(_05301_));
 sg13g2_mux2_1 _13631_ (.A0(_03717_),
    .A1(net2810),
    .S(net80),
    .X(_05465_));
 sg13g2_a21oi_1 _13632_ (.A1(net92),
    .A2(_05465_),
    .Y(_05466_),
    .B1(net52));
 sg13g2_o21ai_1 _13633_ (.B1(net657),
    .Y(_05467_),
    .A1(net4043),
    .A2(net49));
 sg13g2_a21oi_1 _13634_ (.A1(_05464_),
    .A2(_05466_),
    .Y(_01370_),
    .B1(_05467_));
 sg13g2_o21ai_1 _13635_ (.B1(net99),
    .Y(_05468_),
    .A1(net411),
    .A2(_04770_));
 sg13g2_a21oi_1 _13636_ (.A1(net411),
    .A2(_05312_),
    .Y(_05469_),
    .B1(_05468_));
 sg13g2_o21ai_1 _13637_ (.B1(net93),
    .Y(_05470_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .A2(net77));
 sg13g2_a21oi_1 _13638_ (.A1(_03005_),
    .A2(net77),
    .Y(_05471_),
    .B1(_05470_));
 sg13g2_nor3_1 _13639_ (.A(net52),
    .B(_05469_),
    .C(_05471_),
    .Y(_05472_));
 sg13g2_o21ai_1 _13640_ (.B1(net657),
    .Y(_05473_),
    .A1(net610),
    .A2(net49));
 sg13g2_nor2_1 _13641_ (.A(_05472_),
    .B(_05473_),
    .Y(_01371_));
 sg13g2_nor2_1 _13642_ (.A(net411),
    .B(_04771_),
    .Y(_05474_));
 sg13g2_nor2_1 _13643_ (.A(net92),
    .B(_05474_),
    .Y(_05475_));
 sg13g2_o21ai_1 _13644_ (.B1(_05475_),
    .Y(_05476_),
    .A1(net408),
    .A2(_05323_));
 sg13g2_o21ai_1 _13645_ (.B1(net91),
    .Y(_05477_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .A2(net86));
 sg13g2_a21oi_1 _13646_ (.A1(_03245_),
    .A2(net76),
    .Y(_05478_),
    .B1(_05477_));
 sg13g2_nor2_1 _13647_ (.A(net51),
    .B(_05478_),
    .Y(_05479_));
 sg13g2_o21ai_1 _13648_ (.B1(net657),
    .Y(_05480_),
    .A1(net609),
    .A2(net49));
 sg13g2_a21oi_1 _13649_ (.A1(_05476_),
    .A2(_05479_),
    .Y(_01372_),
    .B1(_05480_));
 sg13g2_nor2_1 _13650_ (.A(net411),
    .B(_04773_),
    .Y(_05481_));
 sg13g2_nor2_1 _13651_ (.A(net92),
    .B(_05481_),
    .Y(_05482_));
 sg13g2_o21ai_1 _13652_ (.B1(_05482_),
    .Y(_05483_),
    .A1(net408),
    .A2(_05334_));
 sg13g2_o21ai_1 _13653_ (.B1(net92),
    .Y(_05484_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .A2(net76));
 sg13g2_a21oi_1 _13654_ (.A1(_03367_),
    .A2(net76),
    .Y(_05485_),
    .B1(_05484_));
 sg13g2_nor2_1 _13655_ (.A(net52),
    .B(_05485_),
    .Y(_05486_));
 sg13g2_o21ai_1 _13656_ (.B1(net657),
    .Y(_05487_),
    .A1(net4047),
    .A2(net49));
 sg13g2_a21oi_1 _13657_ (.A1(_05483_),
    .A2(_05486_),
    .Y(_01373_),
    .B1(_05487_));
 sg13g2_nor2_1 _13658_ (.A(net411),
    .B(_04775_),
    .Y(_05488_));
 sg13g2_nor2_1 _13659_ (.A(net92),
    .B(_05488_),
    .Y(_05489_));
 sg13g2_o21ai_1 _13660_ (.B1(_05489_),
    .Y(_05490_),
    .A1(net408),
    .A2(_05344_));
 sg13g2_o21ai_1 _13661_ (.B1(net91),
    .Y(_05491_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .A2(net76));
 sg13g2_a21oi_1 _13662_ (.A1(net76),
    .A2(_03716_),
    .Y(_05492_),
    .B1(_05491_));
 sg13g2_nor2_1 _13663_ (.A(net51),
    .B(_05492_),
    .Y(_05493_));
 sg13g2_o21ai_1 _13664_ (.B1(net657),
    .Y(_05494_),
    .A1(net3851),
    .A2(net49));
 sg13g2_a21oi_1 _13665_ (.A1(_05490_),
    .A2(_05493_),
    .Y(_01374_),
    .B1(_05494_));
 sg13g2_nand2_1 _13666_ (.Y(_05495_),
    .A(_03548_),
    .B(_04363_));
 sg13g2_a21oi_1 _13667_ (.A1(_01611_),
    .A2(net3836),
    .Y(_05496_),
    .B1(_05495_));
 sg13g2_a21oi_1 _13668_ (.A1(net604),
    .A2(net99),
    .Y(_05497_),
    .B1(net3837));
 sg13g2_nor4_1 _13669_ (.A(\i_tinyqv.cpu.instr_fetch_running ),
    .B(\i_tinyqv.cpu.instr_fetch_started ),
    .C(net3836),
    .D(_05495_),
    .Y(_05498_));
 sg13g2_nor3_1 _13670_ (.A(net508),
    .B(net3838),
    .C(_05498_),
    .Y(_01375_));
 sg13g2_o21ai_1 _13671_ (.B1(net656),
    .Y(_05499_),
    .A1(net604),
    .A2(net407));
 sg13g2_a21oi_1 _13672_ (.A1(net407),
    .A2(_03548_),
    .Y(_01376_),
    .B1(_05499_));
 sg13g2_nor2_2 _13673_ (.A(net336),
    .B(_02522_),
    .Y(_05500_));
 sg13g2_nand2_1 _13674_ (.Y(_05501_),
    .A(_00266_),
    .B(_05500_));
 sg13g2_a21oi_2 _13675_ (.B1(_03061_),
    .Y(_05502_),
    .A2(_02272_),
    .A1(_02269_));
 sg13g2_inv_1 _13676_ (.Y(_05503_),
    .A(_05502_));
 sg13g2_a22oi_1 _13677_ (.Y(_05504_),
    .B1(_05502_),
    .B2(_05500_),
    .A2(_05501_),
    .A1(\data_to_write[0] ));
 sg13g2_nor2_1 _13678_ (.A(net506),
    .B(_05504_),
    .Y(_01377_));
 sg13g2_and2_2 _13679_ (.A(_02214_),
    .B(_03062_),
    .X(_05505_));
 sg13g2_inv_1 _13680_ (.Y(_05506_),
    .A(_05505_));
 sg13g2_a22oi_1 _13681_ (.Y(_05507_),
    .B1(_05505_),
    .B2(_05500_),
    .A2(_05501_),
    .A1(net601));
 sg13g2_nor2_1 _13682_ (.A(net507),
    .B(_05507_),
    .Y(_01378_));
 sg13g2_and2_2 _13683_ (.A(_02388_),
    .B(_03062_),
    .X(_05508_));
 sg13g2_inv_1 _13684_ (.Y(_05509_),
    .A(_05508_));
 sg13g2_a22oi_1 _13685_ (.Y(_05510_),
    .B1(_05508_),
    .B2(_05500_),
    .A2(_05501_),
    .A1(net600));
 sg13g2_nor2_1 _13686_ (.A(net507),
    .B(_05510_),
    .Y(_01379_));
 sg13g2_nor2_2 _13687_ (.A(_02337_),
    .B(_03061_),
    .Y(_05511_));
 sg13g2_inv_1 _13688_ (.Y(_05512_),
    .A(_05511_));
 sg13g2_a22oi_1 _13689_ (.Y(_05513_),
    .B1(_05511_),
    .B2(_05500_),
    .A2(_05501_),
    .A1(\data_to_write[3] ));
 sg13g2_nor2_1 _13690_ (.A(net506),
    .B(_05513_),
    .Y(_01380_));
 sg13g2_xnor2_1 _13691_ (.Y(_05514_),
    .A(net583),
    .B(net463));
 sg13g2_and2_2 _13692_ (.A(_02521_),
    .B(_05514_),
    .X(_05515_));
 sg13g2_inv_1 _13693_ (.Y(_05516_),
    .A(_05515_));
 sg13g2_nor2_2 _13694_ (.A(net471),
    .B(net467),
    .Y(_05517_));
 sg13g2_nor3_2 _13695_ (.A(_00266_),
    .B(_05516_),
    .C(_05517_),
    .Y(_05518_));
 sg13g2_nand2_1 _13696_ (.Y(_05519_),
    .A(net336),
    .B(_05502_));
 sg13g2_o21ai_1 _13697_ (.B1(net649),
    .Y(_05520_),
    .A1(net599),
    .A2(_05518_));
 sg13g2_a21oi_1 _13698_ (.A1(_05518_),
    .A2(_05519_),
    .Y(_01381_),
    .B1(_05520_));
 sg13g2_nand2_1 _13699_ (.Y(_05521_),
    .A(net336),
    .B(_05505_));
 sg13g2_o21ai_1 _13700_ (.B1(net649),
    .Y(_05522_),
    .A1(net598),
    .A2(_05518_));
 sg13g2_a21oi_1 _13701_ (.A1(_05518_),
    .A2(_05521_),
    .Y(_01382_),
    .B1(_05522_));
 sg13g2_nand2_1 _13702_ (.Y(_05523_),
    .A(net336),
    .B(_05508_));
 sg13g2_o21ai_1 _13703_ (.B1(net651),
    .Y(_05524_),
    .A1(net597),
    .A2(_05518_));
 sg13g2_a21oi_1 _13704_ (.A1(_05518_),
    .A2(_05523_),
    .Y(_01383_),
    .B1(_05524_));
 sg13g2_nand2_1 _13705_ (.Y(_05525_),
    .A(net336),
    .B(_05511_));
 sg13g2_o21ai_1 _13706_ (.B1(net649),
    .Y(_05526_),
    .A1(\data_to_write[7] ),
    .A2(_05518_));
 sg13g2_a21oi_1 _13707_ (.A1(_05518_),
    .A2(_05525_),
    .Y(_01384_),
    .B1(_05526_));
 sg13g2_nand2_2 _13708_ (.Y(_05527_),
    .A(_02254_),
    .B(_02521_));
 sg13g2_nor2_1 _13709_ (.A(net464),
    .B(_05503_),
    .Y(_05528_));
 sg13g2_a22oi_1 _13710_ (.Y(_05529_),
    .B1(_05528_),
    .B2(_05515_),
    .A2(_05527_),
    .A1(\data_to_write[8] ));
 sg13g2_nor2_1 _13711_ (.A(net506),
    .B(_05529_),
    .Y(_01385_));
 sg13g2_nor2_1 _13712_ (.A(net464),
    .B(_05506_),
    .Y(_05530_));
 sg13g2_a22oi_1 _13713_ (.Y(_05531_),
    .B1(_05530_),
    .B2(_05515_),
    .A2(_05527_),
    .A1(net4120));
 sg13g2_nor2_1 _13714_ (.A(net506),
    .B(_05531_),
    .Y(_01386_));
 sg13g2_nor2_1 _13715_ (.A(net464),
    .B(_05509_),
    .Y(_05532_));
 sg13g2_a22oi_1 _13716_ (.Y(_05533_),
    .B1(_05532_),
    .B2(_05515_),
    .A2(_05527_),
    .A1(net3889));
 sg13g2_nor2_1 _13717_ (.A(net507),
    .B(_05533_),
    .Y(_01387_));
 sg13g2_nor2_1 _13718_ (.A(net464),
    .B(_05512_),
    .Y(_05534_));
 sg13g2_a22oi_1 _13719_ (.Y(_05535_),
    .B1(_05534_),
    .B2(_05515_),
    .A2(_05527_),
    .A1(net3911));
 sg13g2_nor2_1 _13720_ (.A(net506),
    .B(_05535_),
    .Y(_01388_));
 sg13g2_nor4_2 _13721_ (.A(_00266_),
    .B(net471),
    .C(net467),
    .Y(_05536_),
    .D(_02249_));
 sg13g2_nand2_2 _13722_ (.Y(_05537_),
    .A(_05515_),
    .B(_05536_));
 sg13g2_o21ai_1 _13723_ (.B1(net649),
    .Y(_05538_),
    .A1(_05502_),
    .A2(_05537_));
 sg13g2_a21oi_1 _13724_ (.A1(_01503_),
    .A2(_05537_),
    .Y(_01389_),
    .B1(_05538_));
 sg13g2_o21ai_1 _13725_ (.B1(net650),
    .Y(_05539_),
    .A1(_05505_),
    .A2(_05537_));
 sg13g2_a21oi_1 _13726_ (.A1(_01502_),
    .A2(_05537_),
    .Y(_01390_),
    .B1(_05539_));
 sg13g2_o21ai_1 _13727_ (.B1(net650),
    .Y(_05540_),
    .A1(_05508_),
    .A2(_05537_));
 sg13g2_a21oi_1 _13728_ (.A1(_01501_),
    .A2(_05537_),
    .Y(_01391_),
    .B1(_05540_));
 sg13g2_o21ai_1 _13729_ (.B1(net650),
    .Y(_05541_),
    .A1(_05511_),
    .A2(_05537_));
 sg13g2_a21oi_1 _13730_ (.A1(_01500_),
    .A2(_05537_),
    .Y(_01392_),
    .B1(_05541_));
 sg13g2_nand3_1 _13731_ (.B(net463),
    .C(_02521_),
    .A(net583),
    .Y(_05542_));
 sg13g2_o21ai_1 _13732_ (.B1(net650),
    .Y(_05543_),
    .A1(_05502_),
    .A2(_05542_));
 sg13g2_a21oi_1 _13733_ (.A1(_01499_),
    .A2(_05542_),
    .Y(_01393_),
    .B1(_05543_));
 sg13g2_o21ai_1 _13734_ (.B1(net650),
    .Y(_05544_),
    .A1(_05505_),
    .A2(_05542_));
 sg13g2_a21oi_1 _13735_ (.A1(_01498_),
    .A2(_05542_),
    .Y(_01394_),
    .B1(_05544_));
 sg13g2_o21ai_1 _13736_ (.B1(net650),
    .Y(_05545_),
    .A1(_05508_),
    .A2(_05542_));
 sg13g2_a21oi_1 _13737_ (.A1(_01497_),
    .A2(_05542_),
    .Y(_01395_),
    .B1(_05545_));
 sg13g2_o21ai_1 _13738_ (.B1(net650),
    .Y(_05546_),
    .A1(_05511_),
    .A2(_05542_));
 sg13g2_a21oi_1 _13739_ (.A1(_01496_),
    .A2(_05542_),
    .Y(_01396_),
    .B1(_05546_));
 sg13g2_nor2_2 _13740_ (.A(_02522_),
    .B(_05514_),
    .Y(_05547_));
 sg13g2_nor4_2 _13741_ (.A(_00266_),
    .B(_02522_),
    .C(_05514_),
    .Y(_05548_),
    .D(_05517_));
 sg13g2_o21ai_1 _13742_ (.B1(net649),
    .Y(_05549_),
    .A1(net4061),
    .A2(_05548_));
 sg13g2_a21oi_1 _13743_ (.A1(_05519_),
    .A2(_05548_),
    .Y(_01397_),
    .B1(_05549_));
 sg13g2_o21ai_1 _13744_ (.B1(net649),
    .Y(_05550_),
    .A1(net4050),
    .A2(_05548_));
 sg13g2_a21oi_1 _13745_ (.A1(_05521_),
    .A2(_05548_),
    .Y(_01398_),
    .B1(_05550_));
 sg13g2_o21ai_1 _13746_ (.B1(net651),
    .Y(_05551_),
    .A1(net4026),
    .A2(_05548_));
 sg13g2_a21oi_1 _13747_ (.A1(_05523_),
    .A2(_05548_),
    .Y(_01399_),
    .B1(_05551_));
 sg13g2_o21ai_1 _13748_ (.B1(net649),
    .Y(_05552_),
    .A1(net4024),
    .A2(_05548_));
 sg13g2_a21oi_1 _13749_ (.A1(_05525_),
    .A2(_05548_),
    .Y(_01400_),
    .B1(_05552_));
 sg13g2_nand3_1 _13750_ (.B(net467),
    .C(_02521_),
    .A(net583),
    .Y(_05553_));
 sg13g2_a22oi_1 _13751_ (.Y(_05554_),
    .B1(_05553_),
    .B2(net3926),
    .A2(_05547_),
    .A1(_05528_));
 sg13g2_nor2_1 _13752_ (.A(net506),
    .B(_05554_),
    .Y(_01401_));
 sg13g2_a22oi_1 _13753_ (.Y(_05555_),
    .B1(_05553_),
    .B2(net3971),
    .A2(_05547_),
    .A1(_05530_));
 sg13g2_nor2_1 _13754_ (.A(net506),
    .B(_05555_),
    .Y(_01402_));
 sg13g2_a22oi_1 _13755_ (.Y(_05556_),
    .B1(_05553_),
    .B2(net3792),
    .A2(_05547_),
    .A1(_05532_));
 sg13g2_nor2_1 _13756_ (.A(net507),
    .B(_05556_),
    .Y(_01403_));
 sg13g2_a22oi_1 _13757_ (.Y(_05557_),
    .B1(_05553_),
    .B2(net3817),
    .A2(_05547_),
    .A1(_05534_));
 sg13g2_nor2_1 _13758_ (.A(net506),
    .B(_05557_),
    .Y(_01404_));
 sg13g2_and2_2 _13759_ (.A(_05536_),
    .B(_05547_),
    .X(_05558_));
 sg13g2_o21ai_1 _13760_ (.B1(net649),
    .Y(_05559_),
    .A1(net3951),
    .A2(_05558_));
 sg13g2_a21oi_1 _13761_ (.A1(_05503_),
    .A2(_05558_),
    .Y(_01405_),
    .B1(_05559_));
 sg13g2_o21ai_1 _13762_ (.B1(net651),
    .Y(_05560_),
    .A1(net3974),
    .A2(_05558_));
 sg13g2_a21oi_1 _13763_ (.A1(_05506_),
    .A2(_05558_),
    .Y(_01406_),
    .B1(_05560_));
 sg13g2_o21ai_1 _13764_ (.B1(net651),
    .Y(_05561_),
    .A1(net3921),
    .A2(_05558_));
 sg13g2_a21oi_1 _13765_ (.A1(_05509_),
    .A2(_05558_),
    .Y(_01407_),
    .B1(_05561_));
 sg13g2_o21ai_1 _13766_ (.B1(net651),
    .Y(_05562_),
    .A1(net3864),
    .A2(_05558_));
 sg13g2_a21oi_1 _13767_ (.A1(_05512_),
    .A2(_05558_),
    .Y(_01408_),
    .B1(_05562_));
 sg13g2_nand2_1 _13768_ (.Y(_05563_),
    .A(_02984_),
    .B(_03841_));
 sg13g2_nor2_1 _13769_ (.A(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .B(net331),
    .Y(_05564_));
 sg13g2_nand2_1 _13770_ (.Y(_05565_),
    .A(\i_tinyqv.cpu.is_store ),
    .B(_05564_));
 sg13g2_o21ai_1 _13771_ (.B1(_05565_),
    .Y(_05566_),
    .A1(net4048),
    .A2(_05563_));
 sg13g2_nand2_1 _13772_ (.Y(_01409_),
    .A(net652),
    .B(_05566_));
 sg13g2_nor2_1 _13773_ (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .B(net331),
    .Y(_05567_));
 sg13g2_nand2_1 _13774_ (.Y(_05568_),
    .A(\i_tinyqv.cpu.is_store ),
    .B(_05567_));
 sg13g2_o21ai_1 _13775_ (.B1(_05568_),
    .Y(_05569_),
    .A1(net3945),
    .A2(_05563_));
 sg13g2_nand2_1 _13776_ (.Y(_01410_),
    .A(net652),
    .B(_05569_));
 sg13g2_a21oi_1 _13777_ (.A1(net3178),
    .A2(_02983_),
    .Y(_05570_),
    .B1(_03839_));
 sg13g2_nor2_1 _13778_ (.A(net3846),
    .B(_03837_),
    .Y(_05571_));
 sg13g2_o21ai_1 _13779_ (.B1(_05570_),
    .Y(_01411_),
    .A1(_05564_),
    .A2(_05571_));
 sg13g2_nor2_1 _13780_ (.A(net3859),
    .B(_03837_),
    .Y(_05572_));
 sg13g2_o21ai_1 _13781_ (.B1(_05570_),
    .Y(_01412_),
    .A1(_05567_),
    .A2(_05572_));
 sg13g2_a221oi_1 _13782_ (.B2(\i_tinyqv.cpu.is_store ),
    .C1(net314),
    .B1(_03837_),
    .A1(_01709_),
    .Y(_05573_),
    .A2(_02984_));
 sg13g2_a21oi_1 _13783_ (.A1(net3790),
    .A2(net314),
    .Y(_05574_),
    .B1(_05573_));
 sg13g2_nand2_1 _13784_ (.Y(_01413_),
    .A(net652),
    .B(_05574_));
 sg13g2_a21oi_1 _13785_ (.A1(_01494_),
    .A2(net331),
    .Y(_01414_),
    .B1(_03839_));
 sg13g2_and2_1 _13786_ (.A(net652),
    .B(net3856),
    .X(_01415_));
 sg13g2_nor2_1 _13787_ (.A(net508),
    .B(_05517_),
    .Y(_01416_));
 sg13g2_nand2_1 _13788_ (.Y(_05575_),
    .A(net655),
    .B(_03383_));
 sg13g2_a21oi_1 _13789_ (.A1(net474),
    .A2(_02171_),
    .Y(_01417_),
    .B1(_05575_));
 sg13g2_nand2_1 _13790_ (.Y(_05576_),
    .A(net3049),
    .B(net334));
 sg13g2_a21oi_1 _13791_ (.A1(_02985_),
    .A2(_05576_),
    .Y(_01418_),
    .B1(net511));
 sg13g2_nand2_1 _13792_ (.Y(_05577_),
    .A(net3823),
    .B(_03837_));
 sg13g2_o21ai_1 _13793_ (.B1(_05577_),
    .Y(_05578_),
    .A1(net3823),
    .A2(_02983_));
 sg13g2_nor3_1 _13794_ (.A(net648),
    .B(net315),
    .C(_05578_),
    .Y(_01419_));
 sg13g2_nand2_1 _13795_ (.Y(_05579_),
    .A(net88),
    .B(_04163_));
 sg13g2_nor2_2 _13796_ (.A(_03498_),
    .B(_05579_),
    .Y(_05580_));
 sg13g2_nand2_2 _13797_ (.Y(_05581_),
    .A(net88),
    .B(_04164_));
 sg13g2_nor2_2 _13798_ (.A(net218),
    .B(net66),
    .Y(_05582_));
 sg13g2_and2_1 _13799_ (.A(net118),
    .B(_04172_),
    .X(_05583_));
 sg13g2_nor4_2 _13800_ (.A(_03483_),
    .B(net286),
    .C(net212),
    .Y(_05584_),
    .D(_03518_));
 sg13g2_a21oi_2 _13801_ (.B1(_05583_),
    .Y(_05585_),
    .A2(_05584_),
    .A1(net207));
 sg13g2_nor3_2 _13802_ (.A(net286),
    .B(net118),
    .C(_03555_),
    .Y(_05586_));
 sg13g2_nand2b_1 _13803_ (.Y(_05587_),
    .B(net444),
    .A_N(_00189_));
 sg13g2_o21ai_1 _13804_ (.B1(_05587_),
    .Y(_05588_),
    .A1(_00187_),
    .A2(net444));
 sg13g2_nand2_1 _13805_ (.Y(_05589_),
    .A(_00190_),
    .B(net444));
 sg13g2_a21oi_1 _13806_ (.A1(_00188_),
    .A2(net450),
    .Y(_05590_),
    .B1(net435));
 sg13g2_a22oi_1 _13807_ (.Y(_05591_),
    .B1(_05589_),
    .B2(_05590_),
    .A2(_05588_),
    .A1(net435));
 sg13g2_inv_2 _13808_ (.Y(_05592_),
    .A(_05591_));
 sg13g2_a22oi_1 _13809_ (.Y(_05593_),
    .B1(_05586_),
    .B2(_05591_),
    .A2(_03562_),
    .A1(_03487_));
 sg13g2_and2_1 _13810_ (.A(_05580_),
    .B(_05585_),
    .X(_05594_));
 sg13g2_a221oi_1 _13811_ (.B2(_05594_),
    .C1(net511),
    .B1(_05593_),
    .A1(_01493_),
    .Y(_01420_),
    .A2(net67));
 sg13g2_nand3_1 _13812_ (.B(net119),
    .C(_03558_),
    .A(net285),
    .Y(_05595_));
 sg13g2_nor2_1 _13813_ (.A(_03561_),
    .B(_05595_),
    .Y(_05596_));
 sg13g2_nand3b_1 _13814_ (.B(net282),
    .C(_03576_),
    .Y(_05597_),
    .A_N(net204));
 sg13g2_nor2_1 _13815_ (.A(_04179_),
    .B(_05597_),
    .Y(_05598_));
 sg13g2_or2_1 _13816_ (.X(_05599_),
    .B(_05597_),
    .A(_04179_));
 sg13g2_nor2_2 _13817_ (.A(_03569_),
    .B(_05591_),
    .Y(_05600_));
 sg13g2_and2_1 _13818_ (.A(net206),
    .B(_05600_),
    .X(_05601_));
 sg13g2_nand2_1 _13819_ (.Y(_05602_),
    .A(net206),
    .B(_05600_));
 sg13g2_o21ai_1 _13820_ (.B1(_05599_),
    .Y(_05603_),
    .A1(_04169_),
    .A2(_05601_));
 sg13g2_nor4_1 _13821_ (.A(_04173_),
    .B(_04175_),
    .C(_05596_),
    .D(_05603_),
    .Y(_05604_));
 sg13g2_o21ai_1 _13822_ (.B1(net654),
    .Y(_05605_),
    .A1(net4004),
    .A2(net68));
 sg13g2_a21oi_1 _13823_ (.A1(net68),
    .A2(_05604_),
    .Y(_01421_),
    .B1(_05605_));
 sg13g2_nand3b_1 _13824_ (.B(net283),
    .C(net119),
    .Y(_05606_),
    .A_N(net332));
 sg13g2_nor2_1 _13825_ (.A(_03528_),
    .B(_05606_),
    .Y(_05607_));
 sg13g2_or2_1 _13826_ (.X(_05608_),
    .B(_05606_),
    .A(_03528_));
 sg13g2_nor2_1 _13827_ (.A(_03561_),
    .B(_05606_),
    .Y(_05609_));
 sg13g2_a22oi_1 _13828_ (.Y(_05610_),
    .B1(_05582_),
    .B2(_05609_),
    .A2(net66),
    .A1(net3949));
 sg13g2_nor2_1 _13829_ (.A(net509),
    .B(_05610_),
    .Y(_01422_));
 sg13g2_nand2_1 _13830_ (.Y(_05611_),
    .A(_05586_),
    .B(_05592_));
 sg13g2_or2_2 _13831_ (.X(_05612_),
    .B(_03555_),
    .A(net212));
 sg13g2_nand4_1 _13832_ (.B(net68),
    .C(_05611_),
    .A(net216),
    .Y(_05613_),
    .D(_05612_));
 sg13g2_o21ai_1 _13833_ (.B1(_05613_),
    .Y(_05614_),
    .A1(\i_tinyqv.cpu.is_store ),
    .A2(net68));
 sg13g2_nor2_1 _13834_ (.A(_03533_),
    .B(_03559_),
    .Y(_05615_));
 sg13g2_nand2_1 _13835_ (.Y(_05616_),
    .A(net208),
    .B(_05615_));
 sg13g2_a21oi_1 _13836_ (.A1(_05582_),
    .A2(_05616_),
    .Y(_05617_),
    .B1(net509));
 sg13g2_nor2b_1 _13837_ (.A(_05614_),
    .B_N(_05617_),
    .Y(_01423_));
 sg13g2_a21oi_1 _13838_ (.A1(_04168_),
    .A2(_05601_),
    .Y(_05618_),
    .B1(_04180_));
 sg13g2_nand3_1 _13839_ (.B(_04184_),
    .C(_05618_),
    .A(net218),
    .Y(_05619_));
 sg13g2_nand4_1 _13840_ (.B(_03534_),
    .C(net119),
    .A(net208),
    .Y(_05620_),
    .D(_03558_));
 sg13g2_o21ai_1 _13841_ (.B1(net654),
    .Y(_05621_),
    .A1(net66),
    .A2(_05619_));
 sg13g2_a221oi_1 _13842_ (.B2(_05620_),
    .C1(_05621_),
    .B1(_05582_),
    .A1(_01492_),
    .Y(_01424_),
    .A2(net66));
 sg13g2_nor2_1 _13843_ (.A(net3991),
    .B(net68),
    .Y(_05622_));
 sg13g2_nand2_1 _13844_ (.Y(_05623_),
    .A(_04178_),
    .B(_05597_));
 sg13g2_inv_1 _13845_ (.Y(_05624_),
    .A(_05623_));
 sg13g2_nor3_1 _13846_ (.A(net213),
    .B(_03533_),
    .C(net103),
    .Y(_05625_));
 sg13g2_nor3_1 _13847_ (.A(net67),
    .B(_05624_),
    .C(_05625_),
    .Y(_05626_));
 sg13g2_nor3_1 _13848_ (.A(net510),
    .B(_05622_),
    .C(_05626_),
    .Y(_01425_));
 sg13g2_nor2_1 _13849_ (.A(_03535_),
    .B(_03559_),
    .Y(_05627_));
 sg13g2_or2_2 _13850_ (.X(_05628_),
    .B(_04167_),
    .A(net211));
 sg13g2_nor2_1 _13851_ (.A(net66),
    .B(_05628_),
    .Y(_05629_));
 sg13g2_a221oi_1 _13852_ (.B2(net100),
    .C1(_05629_),
    .B1(_05582_),
    .A1(net4105),
    .Y(_05630_),
    .A2(net66));
 sg13g2_nor2_1 _13853_ (.A(net509),
    .B(_05630_),
    .Y(_01426_));
 sg13g2_nor2_1 _13854_ (.A(net332),
    .B(_03544_),
    .Y(_05631_));
 sg13g2_and4_1 _13855_ (.A(_03576_),
    .B(net282),
    .C(net204),
    .D(_05591_),
    .X(_05632_));
 sg13g2_nor3_1 _13856_ (.A(_03564_),
    .B(net66),
    .C(_05632_),
    .Y(_05633_));
 sg13g2_a221oi_1 _13857_ (.B2(_05631_),
    .C1(_05633_),
    .B1(_05582_),
    .A1(net4097),
    .Y(_05634_),
    .A2(net66));
 sg13g2_nor2_1 _13858_ (.A(net509),
    .B(_05634_),
    .Y(_01427_));
 sg13g2_o21ai_1 _13859_ (.B1(net659),
    .Y(_05635_),
    .A1(_03547_),
    .A2(net67));
 sg13g2_a21oi_1 _13860_ (.A1(_01490_),
    .A2(net67),
    .Y(_01428_),
    .B1(_05635_));
 sg13g2_nand2_1 _13861_ (.Y(_05636_),
    .A(net107),
    .B(_04176_));
 sg13g2_nand2_1 _13862_ (.Y(_05637_),
    .A(_03521_),
    .B(net109));
 sg13g2_or2_1 _13863_ (.X(_05638_),
    .B(_05637_),
    .A(_05636_));
 sg13g2_or2_1 _13864_ (.X(_05639_),
    .B(_05586_),
    .A(_05584_));
 sg13g2_nor3_2 _13865_ (.A(net286),
    .B(_03549_),
    .C(_04171_),
    .Y(_05640_));
 sg13g2_nor2_2 _13866_ (.A(net333),
    .B(_05612_),
    .Y(_05641_));
 sg13g2_nor2_1 _13867_ (.A(net210),
    .B(_05612_),
    .Y(_05642_));
 sg13g2_nor3_2 _13868_ (.A(net286),
    .B(net210),
    .C(_05612_),
    .Y(_05643_));
 sg13g2_nand2_2 _13869_ (.Y(_05644_),
    .A(net333),
    .B(_05642_));
 sg13g2_nor3_2 _13870_ (.A(_05640_),
    .B(_05641_),
    .C(_05643_),
    .Y(_05645_));
 sg13g2_nand3b_1 _13871_ (.B(_05645_),
    .C(_04179_),
    .Y(_05646_),
    .A_N(_05638_));
 sg13g2_nor4_1 _13872_ (.A(_03557_),
    .B(_04172_),
    .C(_05639_),
    .D(_05646_),
    .Y(_05647_));
 sg13g2_nor2_1 _13873_ (.A(_03535_),
    .B(_05595_),
    .Y(_05648_));
 sg13g2_a221oi_1 _13874_ (.B2(net333),
    .C1(_05648_),
    .B1(_05647_),
    .A1(_03563_),
    .Y(_05649_),
    .A2(_05632_));
 sg13g2_o21ai_1 _13875_ (.B1(net654),
    .Y(_05650_),
    .A1(net3972),
    .A2(net68));
 sg13g2_a21oi_1 _13876_ (.A1(net68),
    .A2(_05649_),
    .Y(_01429_),
    .B1(_05650_));
 sg13g2_o21ai_1 _13877_ (.B1(net656),
    .Y(_05651_),
    .A1(net219),
    .A2(net67));
 sg13g2_a21oi_1 _13878_ (.A1(_01489_),
    .A2(net67),
    .Y(_01430_),
    .B1(_05651_));
 sg13g2_a21o_1 _13879_ (.A2(net67),
    .A1(net3783),
    .B1(_05651_),
    .X(_01431_));
 sg13g2_nor2_2 _13880_ (.A(net648),
    .B(net67),
    .Y(_05652_));
 sg13g2_nand2b_1 _13881_ (.Y(_05653_),
    .B(net68),
    .A_N(net648));
 sg13g2_nor2_2 _13882_ (.A(net214),
    .B(net104),
    .Y(_05654_));
 sg13g2_nand2_2 _13883_ (.Y(_05655_),
    .A(net285),
    .B(net102));
 sg13g2_nor2_2 _13884_ (.A(net441),
    .B(net436),
    .Y(_05656_));
 sg13g2_nor2_2 _13885_ (.A(net451),
    .B(net438),
    .Y(_05657_));
 sg13g2_or2_1 _13886_ (.X(_05658_),
    .B(net337),
    .A(net321));
 sg13g2_o21ai_1 _13887_ (.B1(_03538_),
    .Y(_05659_),
    .A1(_00145_),
    .A2(net446));
 sg13g2_a22oi_1 _13888_ (.Y(_05660_),
    .B1(net338),
    .B2(_00143_),
    .A2(net322),
    .A1(_00142_));
 sg13g2_o21ai_1 _13889_ (.B1(_05660_),
    .Y(_05661_),
    .A1(net203),
    .A2(_05659_));
 sg13g2_or3_1 _13890_ (.A(_03545_),
    .B(net101),
    .C(_05661_),
    .X(_05662_));
 sg13g2_o21ai_1 _13891_ (.B1(_05662_),
    .Y(_05663_),
    .A1(net282),
    .A2(_05616_));
 sg13g2_nor2_1 _13892_ (.A(net206),
    .B(net107),
    .Y(_05664_));
 sg13g2_nand2_1 _13893_ (.Y(_05665_),
    .A(net205),
    .B(_05600_));
 sg13g2_nor2_2 _13894_ (.A(net107),
    .B(_05665_),
    .Y(_05666_));
 sg13g2_nand2_1 _13895_ (.Y(_05667_),
    .A(_05600_),
    .B(_05664_));
 sg13g2_nor2_1 _13896_ (.A(net208),
    .B(_03570_),
    .Y(_05668_));
 sg13g2_a221oi_1 _13897_ (.B2(_05586_),
    .C1(_05666_),
    .B1(_05668_),
    .A1(_03557_),
    .Y(_05669_),
    .A2(_05632_));
 sg13g2_a22oi_1 _13898_ (.Y(_05670_),
    .B1(_05654_),
    .B2(_05663_),
    .A2(_05636_),
    .A1(net283));
 sg13g2_a21oi_1 _13899_ (.A1(_05669_),
    .A2(_05670_),
    .Y(_05671_),
    .B1(net45));
 sg13g2_a21o_1 _13900_ (.A2(net46),
    .A1(net3908),
    .B1(_05671_),
    .X(_01432_));
 sg13g2_o21ai_1 _13901_ (.B1(_03529_),
    .Y(_05672_),
    .A1(_00149_),
    .A2(net441));
 sg13g2_a22oi_1 _13902_ (.Y(_05673_),
    .B1(net337),
    .B2(_00147_),
    .A2(net321),
    .A1(_00146_));
 sg13g2_o21ai_1 _13903_ (.B1(_05673_),
    .Y(_05674_),
    .A1(net202),
    .A2(_05672_));
 sg13g2_nor2b_1 _13904_ (.A(net101),
    .B_N(_05674_),
    .Y(_05675_));
 sg13g2_a21oi_1 _13905_ (.A1(net204),
    .A2(net101),
    .Y(_05676_),
    .B1(_05675_));
 sg13g2_a22oi_1 _13906_ (.Y(_05677_),
    .B1(_05638_),
    .B2(net332),
    .A2(_05586_),
    .A1(_03534_));
 sg13g2_nand3b_1 _13907_ (.B(_05667_),
    .C(_05677_),
    .Y(_05678_),
    .A_N(_05647_));
 sg13g2_a22oi_1 _13908_ (.Y(_05679_),
    .B1(_05678_),
    .B2(net215),
    .A2(_05676_),
    .A1(_05654_));
 sg13g2_nor2_1 _13909_ (.A(net4069),
    .B(net22),
    .Y(_05680_));
 sg13g2_a21oi_1 _13910_ (.A1(net22),
    .A2(_05679_),
    .Y(_01433_),
    .B1(_05680_));
 sg13g2_o21ai_1 _13911_ (.B1(_05638_),
    .Y(_05681_),
    .A1(net119),
    .A2(_05666_));
 sg13g2_o21ai_1 _13912_ (.B1(_03523_),
    .Y(_05682_),
    .A1(_00153_),
    .A2(net447));
 sg13g2_a22oi_1 _13913_ (.Y(_05683_),
    .B1(net338),
    .B2(_00151_),
    .A2(net322),
    .A1(_00150_));
 sg13g2_o21ai_1 _13914_ (.B1(_05683_),
    .Y(_05684_),
    .A1(net203),
    .A2(_05682_));
 sg13g2_o21ai_1 _13915_ (.B1(_05684_),
    .Y(_05685_),
    .A1(_03533_),
    .A2(_03559_));
 sg13g2_a21oi_1 _13916_ (.A1(_03575_),
    .A2(net101),
    .Y(_05686_),
    .B1(_05655_));
 sg13g2_nor2_1 _13917_ (.A(_05584_),
    .B(_05640_),
    .Y(_05687_));
 sg13g2_nand2b_1 _13918_ (.Y(_05688_),
    .B(_05641_),
    .A_N(_03575_));
 sg13g2_nand3_1 _13919_ (.B(net119),
    .C(_04182_),
    .A(net215),
    .Y(_05689_));
 sg13g2_o21ai_1 _13920_ (.B1(_05688_),
    .Y(_05690_),
    .A1(net209),
    .A2(_05687_));
 sg13g2_a21oi_1 _13921_ (.A1(_05685_),
    .A2(_05686_),
    .Y(_05691_),
    .B1(_05690_));
 sg13g2_nand4_1 _13922_ (.B(_05681_),
    .C(_05689_),
    .A(net20),
    .Y(_05692_),
    .D(_05691_));
 sg13g2_o21ai_1 _13923_ (.B1(_05692_),
    .Y(_05693_),
    .A1(net3796),
    .A2(net28));
 sg13g2_inv_1 _13924_ (.Y(_01434_),
    .A(_05693_));
 sg13g2_nor2_2 _13925_ (.A(_03520_),
    .B(_05640_),
    .Y(_05694_));
 sg13g2_nor2_1 _13926_ (.A(_04182_),
    .B(_05636_),
    .Y(_05695_));
 sg13g2_a21oi_1 _13927_ (.A1(_05694_),
    .A2(_05695_),
    .Y(_05696_),
    .B1(_03533_));
 sg13g2_nand2b_1 _13928_ (.Y(_05697_),
    .B(net109),
    .A_N(_05584_));
 sg13g2_nor2_1 _13929_ (.A(_05641_),
    .B(_05697_),
    .Y(_05698_));
 sg13g2_nand2_1 _13930_ (.Y(_05699_),
    .A(net101),
    .B(_05654_));
 sg13g2_a21oi_1 _13931_ (.A1(_05698_),
    .A2(_05699_),
    .Y(_05700_),
    .B1(_03569_));
 sg13g2_o21ai_1 _13932_ (.B1(_03584_),
    .Y(_05701_),
    .A1(_00170_),
    .A2(net442));
 sg13g2_a22oi_1 _13933_ (.Y(_05702_),
    .B1(net337),
    .B2(_00168_),
    .A2(net321),
    .A1(_00167_));
 sg13g2_o21ai_1 _13934_ (.B1(_05702_),
    .Y(_05703_),
    .A1(net202),
    .A2(_05701_));
 sg13g2_nor2_2 _13935_ (.A(net213),
    .B(_05703_),
    .Y(_05704_));
 sg13g2_nor4_1 _13936_ (.A(net215),
    .B(net104),
    .C(net101),
    .D(_05703_),
    .Y(_05705_));
 sg13g2_nor4_2 _13937_ (.A(_05666_),
    .B(_05696_),
    .C(_05700_),
    .Y(_05706_),
    .D(_05705_));
 sg13g2_nor2_1 _13938_ (.A(net4034),
    .B(net23),
    .Y(_05707_));
 sg13g2_a21oi_1 _13939_ (.A1(net23),
    .A2(_05706_),
    .Y(_01435_),
    .B1(_05707_));
 sg13g2_a221oi_1 _13940_ (.B2(_03528_),
    .C1(_05636_),
    .B1(_05598_),
    .A1(net118),
    .Y(_05708_),
    .A2(_04172_));
 sg13g2_a21oi_1 _13941_ (.A1(net209),
    .A2(_05667_),
    .Y(_05709_),
    .B1(_05708_));
 sg13g2_nand3_1 _13942_ (.B(_05694_),
    .C(_05698_),
    .A(_05644_),
    .Y(_05710_));
 sg13g2_o21ai_1 _13943_ (.B1(_03589_),
    .Y(_05711_),
    .A1(_00174_),
    .A2(net441));
 sg13g2_a22oi_1 _13944_ (.Y(_05712_),
    .B1(net337),
    .B2(_00172_),
    .A2(net321),
    .A1(_00171_));
 sg13g2_o21ai_1 _13945_ (.B1(_05712_),
    .Y(_05713_),
    .A1(net202),
    .A2(_05711_));
 sg13g2_nand2_1 _13946_ (.Y(_05714_),
    .A(_05592_),
    .B(net101));
 sg13g2_o21ai_1 _13947_ (.B1(_05714_),
    .Y(_05715_),
    .A1(net101),
    .A2(_05713_));
 sg13g2_a221oi_1 _13948_ (.B2(_05654_),
    .C1(_05709_),
    .B1(_05715_),
    .A1(_05592_),
    .Y(_05716_),
    .A2(_05710_));
 sg13g2_nor2_1 _13949_ (.A(net3985),
    .B(net23),
    .Y(_05717_));
 sg13g2_a21oi_1 _13950_ (.A1(net23),
    .A2(_05716_),
    .Y(_01436_),
    .B1(_05717_));
 sg13g2_nand3b_1 _13951_ (.B(_05687_),
    .C(_05695_),
    .Y(_05718_),
    .A_N(_05641_));
 sg13g2_o21ai_1 _13952_ (.B1(_03571_),
    .Y(_05719_),
    .A1(_00178_),
    .A2(net445));
 sg13g2_a22oi_1 _13953_ (.Y(_05720_),
    .B1(net337),
    .B2(_00176_),
    .A2(net321),
    .A1(_00175_));
 sg13g2_o21ai_1 _13954_ (.B1(_05720_),
    .Y(_05721_),
    .A1(net203),
    .A2(_05719_));
 sg13g2_nor2_1 _13955_ (.A(net215),
    .B(_05721_),
    .Y(_05722_));
 sg13g2_nand2_1 _13956_ (.Y(_05723_),
    .A(_04193_),
    .B(_05599_));
 sg13g2_o21ai_1 _13957_ (.B1(net283),
    .Y(_05724_),
    .A1(_05637_),
    .A2(_05723_));
 sg13g2_o21ai_1 _13958_ (.B1(_05724_),
    .Y(_05725_),
    .A1(_03569_),
    .A2(_05644_));
 sg13g2_a221oi_1 _13959_ (.B2(net102),
    .C1(_05725_),
    .B1(_05722_),
    .A1(net205),
    .Y(_05726_),
    .A2(_05718_));
 sg13g2_nor2_1 _13960_ (.A(net3956),
    .B(net23),
    .Y(_05727_));
 sg13g2_a21oi_1 _13961_ (.A1(net26),
    .A2(_05726_),
    .Y(_01437_),
    .B1(_05727_));
 sg13g2_o21ai_1 _13962_ (.B1(_03534_),
    .Y(_05728_),
    .A1(_05697_),
    .A2(_05723_));
 sg13g2_a21oi_1 _13963_ (.A1(net107),
    .A2(_04176_),
    .Y(_05729_),
    .B1(net206));
 sg13g2_a21oi_1 _13964_ (.A1(_03521_),
    .A2(_05645_),
    .Y(_05730_),
    .B1(net282));
 sg13g2_o21ai_1 _13965_ (.B1(_03565_),
    .Y(_05731_),
    .A1(_00182_),
    .A2(net439));
 sg13g2_a22oi_1 _13966_ (.Y(_05732_),
    .B1(net337),
    .B2(_00180_),
    .A2(net321),
    .A1(_00179_));
 sg13g2_o21ai_1 _13967_ (.B1(_05732_),
    .Y(_05733_),
    .A1(net202),
    .A2(_05731_));
 sg13g2_nor2_1 _13968_ (.A(net213),
    .B(_05733_),
    .Y(_05734_));
 sg13g2_a21oi_1 _13969_ (.A1(net103),
    .A2(_05734_),
    .Y(_05735_),
    .B1(_05729_));
 sg13g2_a21oi_1 _13970_ (.A1(net284),
    .A2(_04182_),
    .Y(_05736_),
    .B1(_05730_));
 sg13g2_and4_1 _13971_ (.A(net21),
    .B(_05728_),
    .C(_05735_),
    .D(_05736_),
    .X(_05737_));
 sg13g2_a21oi_1 _13972_ (.A1(_01588_),
    .A2(net46),
    .Y(_01438_),
    .B1(_05737_));
 sg13g2_a21oi_1 _13973_ (.A1(_03521_),
    .A2(net109),
    .Y(_05738_),
    .B1(net208));
 sg13g2_o21ai_1 _13974_ (.B1(_05587_),
    .Y(_05739_),
    .A1(_00190_),
    .A2(net444));
 sg13g2_a22oi_1 _13975_ (.Y(_05740_),
    .B1(net338),
    .B2(_00188_),
    .A2(net322),
    .A1(_00187_));
 sg13g2_o21ai_1 _13976_ (.B1(_05740_),
    .Y(_05741_),
    .A1(net202),
    .A2(_05739_));
 sg13g2_nor2_1 _13977_ (.A(_05655_),
    .B(_05741_),
    .Y(_05742_));
 sg13g2_o21ai_1 _13978_ (.B1(net332),
    .Y(_05743_),
    .A1(_05583_),
    .A2(_05598_));
 sg13g2_o21ai_1 _13979_ (.B1(_05743_),
    .Y(_05744_),
    .A1(net204),
    .A2(_05645_));
 sg13g2_nor4_2 _13980_ (.A(_05729_),
    .B(_05738_),
    .C(_05742_),
    .Y(_05745_),
    .D(_05744_));
 sg13g2_nor2_1 _13981_ (.A(net4023),
    .B(net27),
    .Y(_05746_));
 sg13g2_a21oi_1 _13982_ (.A1(net27),
    .A2(_05745_),
    .Y(_01439_),
    .B1(_05746_));
 sg13g2_nand2_1 _13983_ (.Y(_05747_),
    .A(net120),
    .B(_05723_));
 sg13g2_a21oi_1 _13984_ (.A1(_05644_),
    .A2(_05694_),
    .Y(_05748_),
    .B1(_03575_));
 sg13g2_a21oi_1 _13985_ (.A1(_04176_),
    .A2(net109),
    .Y(_05749_),
    .B1(net206));
 sg13g2_o21ai_1 _13986_ (.B1(_03578_),
    .Y(_05750_),
    .A1(_00186_),
    .A2(net446));
 sg13g2_a22oi_1 _13987_ (.Y(_05751_),
    .B1(net338),
    .B2(_00184_),
    .A2(net322),
    .A1(_00183_));
 sg13g2_o21ai_1 _13988_ (.B1(_05751_),
    .Y(_05752_),
    .A1(net203),
    .A2(_05750_));
 sg13g2_nand2_1 _13989_ (.Y(_05753_),
    .A(_05600_),
    .B(_05606_));
 sg13g2_nand2_1 _13990_ (.Y(_05754_),
    .A(_05664_),
    .B(_05753_));
 sg13g2_nand2_1 _13991_ (.Y(_05755_),
    .A(net332),
    .B(_05664_));
 sg13g2_nand2_1 _13992_ (.Y(_05756_),
    .A(_05754_),
    .B(_05755_));
 sg13g2_o21ai_1 _13993_ (.B1(_05747_),
    .Y(_05757_),
    .A1(_05655_),
    .A2(_05752_));
 sg13g2_nor4_2 _13994_ (.A(_05748_),
    .B(_05749_),
    .C(_05756_),
    .Y(_05758_),
    .D(_05757_));
 sg13g2_nor2_1 _13995_ (.A(net4074),
    .B(net27),
    .Y(_05759_));
 sg13g2_a21oi_1 _13996_ (.A1(net27),
    .A2(_05758_),
    .Y(_01440_),
    .B1(_05759_));
 sg13g2_nor2_1 _13997_ (.A(net206),
    .B(_04193_),
    .Y(_05760_));
 sg13g2_nor2_1 _13998_ (.A(_05749_),
    .B(_05760_),
    .Y(_05761_));
 sg13g2_o21ai_1 _13999_ (.B1(net205),
    .Y(_05762_),
    .A1(_05598_),
    .A2(_05643_));
 sg13g2_nand4_1 _14000_ (.B(_05755_),
    .C(_05761_),
    .A(_05754_),
    .Y(_05763_),
    .D(_05762_));
 sg13g2_o21ai_1 _14001_ (.B1(_03513_),
    .Y(_05764_),
    .A1(_00157_),
    .A2(net445));
 sg13g2_a22oi_1 _14002_ (.Y(_05765_),
    .B1(net338),
    .B2(_00155_),
    .A2(net322),
    .A1(_00154_));
 sg13g2_o21ai_1 _14003_ (.B1(_05765_),
    .Y(_05766_),
    .A1(net202),
    .A2(_05764_));
 sg13g2_nor2_1 _14004_ (.A(net213),
    .B(_05766_),
    .Y(_05767_));
 sg13g2_nand2_1 _14005_ (.Y(_05768_),
    .A(net102),
    .B(_05767_));
 sg13g2_o21ai_1 _14006_ (.B1(_05768_),
    .Y(_05769_),
    .A1(_03569_),
    .A2(_05694_));
 sg13g2_nor3_2 _14007_ (.A(net45),
    .B(_05763_),
    .C(_05769_),
    .Y(_05770_));
 sg13g2_a21oi_1 _14008_ (.A1(_01589_),
    .A2(net47),
    .Y(_01441_),
    .B1(_05770_));
 sg13g2_o21ai_1 _14009_ (.B1(_03508_),
    .Y(_05771_),
    .A1(_00161_),
    .A2(net440));
 sg13g2_a22oi_1 _14010_ (.Y(_05772_),
    .B1(net337),
    .B2(_00159_),
    .A2(net321),
    .A1(_00158_));
 sg13g2_o21ai_1 _14011_ (.B1(_05772_),
    .Y(_05773_),
    .A1(net202),
    .A2(_05771_));
 sg13g2_nor2_1 _14012_ (.A(net215),
    .B(_05773_),
    .Y(_05774_));
 sg13g2_a21oi_1 _14013_ (.A1(net102),
    .A2(_05774_),
    .Y(_05775_),
    .B1(_05763_));
 sg13g2_o21ai_1 _14014_ (.B1(_05775_),
    .Y(_05776_),
    .A1(_03521_),
    .A2(net204));
 sg13g2_mux2_1 _14015_ (.A0(net4089),
    .A1(_05776_),
    .S(net21),
    .X(_01442_));
 sg13g2_nand2_1 _14016_ (.Y(_05777_),
    .A(_03520_),
    .B(net205));
 sg13g2_nand2b_1 _14017_ (.Y(_05778_),
    .B(_05777_),
    .A_N(_05763_));
 sg13g2_nor2_1 _14018_ (.A(_03546_),
    .B(_05661_),
    .Y(_05779_));
 sg13g2_o21ai_1 _14019_ (.B1(_03550_),
    .Y(_05780_),
    .A1(_00165_),
    .A2(net439));
 sg13g2_a22oi_1 _14020_ (.Y(_05781_),
    .B1(net337),
    .B2(_00163_),
    .A2(net321),
    .A1(_00162_));
 sg13g2_o21ai_1 _14021_ (.B1(_05781_),
    .Y(_05782_),
    .A1(net202),
    .A2(_05780_));
 sg13g2_nor2_1 _14022_ (.A(_03545_),
    .B(_05782_),
    .Y(_05783_));
 sg13g2_nor3_1 _14023_ (.A(net100),
    .B(_05779_),
    .C(_05783_),
    .Y(_05784_));
 sg13g2_a21oi_1 _14024_ (.A1(net282),
    .A2(net100),
    .Y(_05785_),
    .B1(_05784_));
 sg13g2_a21oi_1 _14025_ (.A1(_05654_),
    .A2(_05785_),
    .Y(_05786_),
    .B1(_05778_));
 sg13g2_nor2_1 _14026_ (.A(net4106),
    .B(net27),
    .Y(_05787_));
 sg13g2_a21oi_1 _14027_ (.A1(net27),
    .A2(_05786_),
    .Y(_01443_),
    .B1(_05787_));
 sg13g2_nand2_1 _14028_ (.Y(_05788_),
    .A(_05654_),
    .B(_05783_));
 sg13g2_nand2b_1 _14029_ (.Y(_05789_),
    .B(_05788_),
    .A_N(_05778_));
 sg13g2_nor2_1 _14030_ (.A(_03545_),
    .B(net104),
    .Y(_05790_));
 sg13g2_nand2_2 _14031_ (.Y(_05791_),
    .A(_03546_),
    .B(net103));
 sg13g2_nor2_1 _14032_ (.A(net217),
    .B(_03582_),
    .Y(_05792_));
 sg13g2_a221oi_1 _14033_ (.B2(_05792_),
    .C1(_05789_),
    .B1(_05791_),
    .A1(net283),
    .Y(_05793_),
    .A2(_05624_));
 sg13g2_nor2_1 _14034_ (.A(net3955),
    .B(net27),
    .Y(_05794_));
 sg13g2_a21oi_1 _14035_ (.A1(net27),
    .A2(_05793_),
    .Y(_01444_),
    .B1(_05794_));
 sg13g2_nor3_1 _14036_ (.A(net217),
    .B(_03517_),
    .C(_05790_),
    .Y(_05795_));
 sg13g2_nor2_1 _14037_ (.A(_04201_),
    .B(_05623_),
    .Y(_05796_));
 sg13g2_nor4_2 _14038_ (.A(net47),
    .B(_05789_),
    .C(_05795_),
    .Y(_05797_),
    .D(_05796_));
 sg13g2_a21oi_1 _14039_ (.A1(_01590_),
    .A2(net47),
    .Y(_01445_),
    .B1(_05797_));
 sg13g2_nand2b_1 _14040_ (.Y(_05798_),
    .B(_05791_),
    .A_N(net211));
 sg13g2_a21oi_1 _14041_ (.A1(net102),
    .A2(_05783_),
    .Y(_05799_),
    .B1(net214));
 sg13g2_nand2_1 _14042_ (.Y(_05800_),
    .A(net119),
    .B(_05624_));
 sg13g2_nor2_1 _14043_ (.A(net285),
    .B(_05778_),
    .Y(_05801_));
 sg13g2_a221oi_1 _14044_ (.B2(_05801_),
    .C1(net45),
    .B1(_05800_),
    .A1(_05798_),
    .Y(_05802_),
    .A2(_05799_));
 sg13g2_a21o_1 _14045_ (.A2(net46),
    .A1(net4063),
    .B1(_05802_),
    .X(_01446_));
 sg13g2_o21ai_1 _14046_ (.B1(_05799_),
    .Y(_05803_),
    .A1(net207),
    .A2(_05790_));
 sg13g2_o21ai_1 _14047_ (.B1(_05801_),
    .Y(_05804_),
    .A1(_03533_),
    .A2(_05623_));
 sg13g2_nand3_1 _14048_ (.B(_05803_),
    .C(_05804_),
    .A(net20),
    .Y(_05805_));
 sg13g2_o21ai_1 _14049_ (.B1(_05805_),
    .Y(_01447_),
    .A1(_01586_),
    .A2(net23));
 sg13g2_o21ai_1 _14050_ (.B1(_03482_),
    .Y(_05806_),
    .A1(\i_tinyqv.cpu.instr_data[2][0] ),
    .A2(net449));
 sg13g2_a22oi_1 _14051_ (.Y(_05807_),
    .B1(net338),
    .B2(\i_tinyqv.cpu.instr_data[0][0] ),
    .A2(net322),
    .A1(\i_tinyqv.cpu.instr_data[1][0] ));
 sg13g2_o21ai_1 _14052_ (.B1(_05807_),
    .Y(_05808_),
    .A1(net203),
    .A2(_05806_));
 sg13g2_nand2_1 _14053_ (.Y(_05809_),
    .A(_05791_),
    .B(_05808_));
 sg13g2_nand3_1 _14054_ (.B(_05761_),
    .C(_05777_),
    .A(_05754_),
    .Y(_05810_));
 sg13g2_a221oi_1 _14055_ (.B2(_05624_),
    .C1(_05810_),
    .B1(_03528_),
    .A1(_03483_),
    .Y(_05811_),
    .A2(_03486_));
 sg13g2_a221oi_1 _14056_ (.B2(_05762_),
    .C1(net45),
    .B1(_05811_),
    .A1(_05799_),
    .Y(_05812_),
    .A2(_05809_));
 sg13g2_a21o_1 _14057_ (.A2(net46),
    .A1(net4045),
    .B1(_05812_),
    .X(_01448_));
 sg13g2_a21oi_1 _14058_ (.A1(_04179_),
    .A2(_05644_),
    .Y(_05813_),
    .B1(_03582_));
 sg13g2_nor2_1 _14059_ (.A(_05810_),
    .B(_05813_),
    .Y(_05814_));
 sg13g2_nand2_1 _14060_ (.Y(_05815_),
    .A(_05788_),
    .B(_05814_));
 sg13g2_a22oi_1 _14061_ (.Y(_05816_),
    .B1(_03481_),
    .B2(\i_tinyqv.cpu.instr_data[2][1] ),
    .A2(net449),
    .A1(\i_tinyqv.cpu.instr_data[3][1] ));
 sg13g2_a22oi_1 _14062_ (.Y(_05817_),
    .B1(_05657_),
    .B2(\i_tinyqv.cpu.instr_data[0][1] ),
    .A2(_05656_),
    .A1(\i_tinyqv.cpu.instr_data[1][1] ));
 sg13g2_o21ai_1 _14063_ (.B1(_05817_),
    .Y(_05818_),
    .A1(_05657_),
    .A2(_05816_));
 sg13g2_nand2_1 _14064_ (.Y(_05819_),
    .A(net285),
    .B(_05818_));
 sg13g2_inv_1 _14065_ (.Y(_05820_),
    .A(_05819_));
 sg13g2_a21oi_1 _14066_ (.A1(_05791_),
    .A2(_05820_),
    .Y(_05821_),
    .B1(_05815_));
 sg13g2_nor2_1 _14067_ (.A(net3975),
    .B(net25),
    .Y(_05822_));
 sg13g2_a21oi_1 _14068_ (.A1(net24),
    .A2(_05821_),
    .Y(_01449_),
    .B1(_05822_));
 sg13g2_o21ai_1 _14069_ (.B1(_03536_),
    .Y(_05823_),
    .A1(\i_tinyqv.cpu.instr_data[2][2] ),
    .A2(net446));
 sg13g2_a22oi_1 _14070_ (.Y(_05824_),
    .B1(net338),
    .B2(\i_tinyqv.cpu.instr_data[0][2] ),
    .A2(net322),
    .A1(\i_tinyqv.cpu.instr_data[1][2] ));
 sg13g2_o21ai_1 _14071_ (.B1(_05824_),
    .Y(_05825_),
    .A1(net203),
    .A2(_05823_));
 sg13g2_nand2_2 _14072_ (.Y(_05826_),
    .A(net285),
    .B(_05825_));
 sg13g2_inv_1 _14073_ (.Y(_05827_),
    .A(_05826_));
 sg13g2_a21oi_1 _14074_ (.A1(_05791_),
    .A2(_05827_),
    .Y(_05828_),
    .B1(_05815_));
 sg13g2_nor2_1 _14075_ (.A(net3941),
    .B(net20),
    .Y(_05829_));
 sg13g2_a21oi_1 _14076_ (.A1(net20),
    .A2(_05828_),
    .Y(_01450_),
    .B1(_05829_));
 sg13g2_a21oi_1 _14077_ (.A1(_01602_),
    .A2(net448),
    .Y(_05830_),
    .B1(net203));
 sg13g2_o21ai_1 _14078_ (.B1(_05830_),
    .Y(_05831_),
    .A1(\i_tinyqv.cpu.instr_data[2][3] ),
    .A2(net448));
 sg13g2_a22oi_1 _14079_ (.Y(_05832_),
    .B1(_05657_),
    .B2(\i_tinyqv.cpu.instr_data[0][3] ),
    .A2(_05656_),
    .A1(\i_tinyqv.cpu.instr_data[1][3] ));
 sg13g2_a21oi_1 _14080_ (.A1(_05831_),
    .A2(_05832_),
    .Y(_05833_),
    .B1(net213));
 sg13g2_a21oi_1 _14081_ (.A1(_05791_),
    .A2(_05833_),
    .Y(_05834_),
    .B1(_05815_));
 sg13g2_nor2_1 _14082_ (.A(net3992),
    .B(net20),
    .Y(_05835_));
 sg13g2_a21oi_1 _14083_ (.A1(net20),
    .A2(_05834_),
    .Y(_01451_),
    .B1(_05835_));
 sg13g2_o21ai_1 _14084_ (.B1(_05814_),
    .Y(_05836_),
    .A1(_05655_),
    .A2(_05782_));
 sg13g2_or2_1 _14085_ (.X(_05837_),
    .B(_05661_),
    .A(net214));
 sg13g2_nor2_1 _14086_ (.A(net103),
    .B(_05837_),
    .Y(_05838_));
 sg13g2_nor3_1 _14087_ (.A(net45),
    .B(net87),
    .C(_05838_),
    .Y(_05839_));
 sg13g2_a21oi_1 _14088_ (.A1(_01592_),
    .A2(net46),
    .Y(_01452_),
    .B1(_05839_));
 sg13g2_nor2_2 _14089_ (.A(net215),
    .B(_05674_),
    .Y(_05840_));
 sg13g2_a21oi_1 _14090_ (.A1(net104),
    .A2(_05840_),
    .Y(_05841_),
    .B1(net87));
 sg13g2_nor2_1 _14091_ (.A(net3988),
    .B(net24),
    .Y(_05842_));
 sg13g2_a21oi_1 _14092_ (.A1(net24),
    .A2(_05841_),
    .Y(_01453_),
    .B1(_05842_));
 sg13g2_nor2_2 _14093_ (.A(net215),
    .B(_05684_),
    .Y(_05843_));
 sg13g2_a21oi_1 _14094_ (.A1(net104),
    .A2(_05843_),
    .Y(_05844_),
    .B1(net87));
 sg13g2_nor2_1 _14095_ (.A(net3890),
    .B(net24),
    .Y(_05845_));
 sg13g2_a21oi_1 _14096_ (.A1(net24),
    .A2(_05844_),
    .Y(_01454_),
    .B1(_05845_));
 sg13g2_a21oi_1 _14097_ (.A1(net104),
    .A2(_05704_),
    .Y(_05846_),
    .B1(_05836_));
 sg13g2_nor2_1 _14098_ (.A(net3841),
    .B(net24),
    .Y(_05847_));
 sg13g2_a21oi_1 _14099_ (.A1(net24),
    .A2(_05846_),
    .Y(_01455_),
    .B1(_05847_));
 sg13g2_nor3_1 _14100_ (.A(net213),
    .B(net102),
    .C(_05713_),
    .Y(_05848_));
 sg13g2_nor3_1 _14101_ (.A(net45),
    .B(net87),
    .C(_05848_),
    .Y(_05849_));
 sg13g2_a21oi_1 _14102_ (.A1(_01593_),
    .A2(net46),
    .Y(_01456_),
    .B1(_05849_));
 sg13g2_a21oi_1 _14103_ (.A1(net104),
    .A2(_05722_),
    .Y(_05850_),
    .B1(_05836_));
 sg13g2_nor2_1 _14104_ (.A(net3492),
    .B(net22),
    .Y(_05851_));
 sg13g2_a21oi_1 _14105_ (.A1(net23),
    .A2(_05850_),
    .Y(_01457_),
    .B1(_05851_));
 sg13g2_a21oi_1 _14106_ (.A1(net104),
    .A2(_05734_),
    .Y(_05852_),
    .B1(net87));
 sg13g2_nor2_1 _14107_ (.A(net3620),
    .B(net20),
    .Y(_05853_));
 sg13g2_a21oi_1 _14108_ (.A1(net21),
    .A2(_05852_),
    .Y(_01458_),
    .B1(_05853_));
 sg13g2_nor3_1 _14109_ (.A(net213),
    .B(net102),
    .C(_05741_),
    .Y(_05854_));
 sg13g2_nor3_1 _14110_ (.A(net45),
    .B(net87),
    .C(_05854_),
    .Y(_05855_));
 sg13g2_a21oi_1 _14111_ (.A1(_01587_),
    .A2(net46),
    .Y(_01459_),
    .B1(_05855_));
 sg13g2_nor3_1 _14112_ (.A(net213),
    .B(net102),
    .C(_05752_),
    .Y(_05856_));
 sg13g2_nor3_1 _14113_ (.A(net45),
    .B(_05836_),
    .C(_05856_),
    .Y(_05857_));
 sg13g2_a21oi_1 _14114_ (.A1(_01594_),
    .A2(net46),
    .Y(_01460_),
    .B1(_05857_));
 sg13g2_a21oi_1 _14115_ (.A1(_05607_),
    .A2(_05767_),
    .Y(_05858_),
    .B1(net87));
 sg13g2_nor2_1 _14116_ (.A(net3370),
    .B(net22),
    .Y(_05859_));
 sg13g2_a21oi_1 _14117_ (.A1(net22),
    .A2(_05858_),
    .Y(_01461_),
    .B1(_05859_));
 sg13g2_a21oi_1 _14118_ (.A1(_05607_),
    .A2(_05774_),
    .Y(_05860_),
    .B1(net87));
 sg13g2_nor2_1 _14119_ (.A(net3443),
    .B(net22),
    .Y(_05861_));
 sg13g2_a21oi_1 _14120_ (.A1(net20),
    .A2(_05860_),
    .Y(_01462_),
    .B1(_05861_));
 sg13g2_o21ai_1 _14121_ (.B1(_05814_),
    .Y(_05862_),
    .A1(net214),
    .A2(_05782_));
 sg13g2_mux2_1 _14122_ (.A0(net3313),
    .A1(_05862_),
    .S(net25),
    .X(_01463_));
 sg13g2_nor2_2 _14123_ (.A(_05620_),
    .B(_05733_),
    .Y(_05863_));
 sg13g2_nor2_1 _14124_ (.A(net100),
    .B(_05863_),
    .Y(_05864_));
 sg13g2_o21ai_1 _14125_ (.B1(net210),
    .Y(_05865_),
    .A1(_05627_),
    .A2(_05863_));
 sg13g2_a221oi_1 _14126_ (.B2(net208),
    .C1(net218),
    .B1(_03560_),
    .A1(net283),
    .Y(_05866_),
    .A2(_03543_));
 sg13g2_nand2b_1 _14127_ (.Y(_05867_),
    .B(_05866_),
    .A_N(_05609_));
 sg13g2_a21oi_1 _14128_ (.A1(net206),
    .A2(_05864_),
    .Y(_05868_),
    .B1(_05867_));
 sg13g2_o21ai_1 _14129_ (.B1(_04168_),
    .Y(_05869_),
    .A1(_05606_),
    .A2(_05665_));
 sg13g2_a21oi_1 _14130_ (.A1(_03535_),
    .A2(_05601_),
    .Y(_05870_),
    .B1(_05869_));
 sg13g2_a221oi_1 _14131_ (.B2(_05868_),
    .C1(_05870_),
    .B1(_05865_),
    .A1(net286),
    .Y(_05871_),
    .A2(_04173_));
 sg13g2_nor2_1 _14132_ (.A(net3891),
    .B(net29),
    .Y(_05872_));
 sg13g2_a21oi_1 _14133_ (.A1(net29),
    .A2(_05871_),
    .Y(_01464_),
    .B1(_05872_));
 sg13g2_a221oi_1 _14134_ (.B2(net210),
    .C1(_05867_),
    .B1(_05864_),
    .A1(net211),
    .Y(_05873_),
    .A2(net100));
 sg13g2_o21ai_1 _14135_ (.B1(_05592_),
    .Y(_05874_),
    .A1(_03528_),
    .A2(_05602_));
 sg13g2_o21ai_1 _14136_ (.B1(_04181_),
    .Y(_05875_),
    .A1(_05869_),
    .A2(_05874_));
 sg13g2_o21ai_1 _14137_ (.B1(net21),
    .Y(_05876_),
    .A1(_05873_),
    .A2(_05875_));
 sg13g2_o21ai_1 _14138_ (.B1(_05876_),
    .Y(_01465_),
    .A1(_01584_),
    .A2(net29));
 sg13g2_mux2_1 _14139_ (.A0(net211),
    .A1(_05741_),
    .S(_05863_),
    .X(_05877_));
 sg13g2_inv_1 _14140_ (.Y(_05878_),
    .A(_05877_));
 sg13g2_nor2_1 _14141_ (.A(net100),
    .B(_05867_),
    .Y(_05879_));
 sg13g2_nor2_1 _14142_ (.A(_03561_),
    .B(_05602_),
    .Y(_05880_));
 sg13g2_a21oi_1 _14143_ (.A1(net100),
    .A2(_05878_),
    .Y(_05881_),
    .B1(_05867_));
 sg13g2_o21ai_1 _14144_ (.B1(_05881_),
    .Y(_05882_),
    .A1(net100),
    .A2(_05878_));
 sg13g2_o21ai_1 _14145_ (.B1(_05882_),
    .Y(_05883_),
    .A1(net107),
    .A2(_05880_));
 sg13g2_nor2b_2 _14146_ (.A(_05883_),
    .B_N(_05628_),
    .Y(_05884_));
 sg13g2_nor2_1 _14147_ (.A(net574),
    .B(net29),
    .Y(_05885_));
 sg13g2_a21oi_1 _14148_ (.A1(net29),
    .A2(_05884_),
    .Y(_01466_),
    .B1(_05885_));
 sg13g2_a21oi_1 _14149_ (.A1(net210),
    .A2(net205),
    .Y(_05886_),
    .B1(_03534_));
 sg13g2_nor2_1 _14150_ (.A(_05773_),
    .B(_05886_),
    .Y(_05887_));
 sg13g2_o21ai_1 _14151_ (.B1(_05879_),
    .Y(_05888_),
    .A1(_05863_),
    .A2(_05887_));
 sg13g2_a21oi_1 _14152_ (.A1(_03570_),
    .A2(_05591_),
    .Y(_05889_),
    .B1(_05880_));
 sg13g2_o21ai_1 _14153_ (.B1(_05888_),
    .Y(_05890_),
    .A1(net107),
    .A2(_05889_));
 sg13g2_o21ai_1 _14154_ (.B1(net21),
    .Y(_05891_),
    .A1(_04180_),
    .A2(_05890_));
 sg13g2_o21ai_1 _14155_ (.B1(_05891_),
    .Y(_01467_),
    .A1(_01583_),
    .A2(net29));
 sg13g2_nand3_1 _14156_ (.B(net209),
    .C(_03560_),
    .A(_03518_),
    .Y(_05892_));
 sg13g2_nand2_1 _14157_ (.Y(_05893_),
    .A(_05585_),
    .B(_05612_));
 sg13g2_nor2b_1 _14158_ (.A(_05893_),
    .B_N(net109),
    .Y(_05894_));
 sg13g2_nand2_1 _14159_ (.Y(_05895_),
    .A(_03570_),
    .B(_05894_));
 sg13g2_o21ai_1 _14160_ (.B1(_05895_),
    .Y(_05896_),
    .A1(_03517_),
    .A2(net109));
 sg13g2_a22oi_1 _14161_ (.Y(_05897_),
    .B1(_05896_),
    .B2(net217),
    .A2(_05892_),
    .A1(_05792_));
 sg13g2_nor2_1 _14162_ (.A(net4006),
    .B(net25),
    .Y(_05898_));
 sg13g2_a21oi_1 _14163_ (.A1(net25),
    .A2(_05897_),
    .Y(_01468_),
    .B1(_05898_));
 sg13g2_a21oi_2 _14164_ (.B1(_05893_),
    .Y(_05899_),
    .A2(_03518_),
    .A1(net285));
 sg13g2_nor2_1 _14165_ (.A(net3958),
    .B(net24),
    .Y(_05900_));
 sg13g2_a21oi_1 _14166_ (.A1(net25),
    .A2(_05899_),
    .Y(_01469_),
    .B1(_05900_));
 sg13g2_a221oi_1 _14167_ (.B2(_03570_),
    .C1(_05592_),
    .B1(_03528_),
    .A1(_03483_),
    .Y(_05901_),
    .A2(_03486_));
 sg13g2_nor2_1 _14168_ (.A(net217),
    .B(net212),
    .Y(_05902_));
 sg13g2_nand4_1 _14169_ (.B(net206),
    .C(_04177_),
    .A(net208),
    .Y(_05903_),
    .D(_05615_));
 sg13g2_nand2b_1 _14170_ (.Y(_05904_),
    .B(_03583_),
    .A_N(_05892_));
 sg13g2_and2_1 _14171_ (.A(_05903_),
    .B(_05904_),
    .X(_05905_));
 sg13g2_a22oi_1 _14172_ (.Y(_05906_),
    .B1(_05902_),
    .B2(_05905_),
    .A2(_05901_),
    .A1(_05894_));
 sg13g2_nor2_1 _14173_ (.A(net3513),
    .B(net22),
    .Y(_05907_));
 sg13g2_a21oi_1 _14174_ (.A1(net22),
    .A2(_05906_),
    .Y(_01470_),
    .B1(_05907_));
 sg13g2_nand3b_1 _14175_ (.B(net109),
    .C(net107),
    .Y(_05908_),
    .A_N(_05639_));
 sg13g2_o21ai_1 _14176_ (.B1(_04192_),
    .Y(_05909_),
    .A1(net118),
    .A2(_04170_));
 sg13g2_nand3_1 _14177_ (.B(_04174_),
    .C(_04181_),
    .A(_03564_),
    .Y(_05910_));
 sg13g2_nor3_2 _14178_ (.A(_05908_),
    .B(_05909_),
    .C(_05910_),
    .Y(_05911_));
 sg13g2_nor2_1 _14179_ (.A(_03588_),
    .B(_05911_),
    .Y(_05912_));
 sg13g2_nor2_1 _14180_ (.A(net216),
    .B(net207),
    .Y(_05913_));
 sg13g2_nand2_1 _14181_ (.Y(_05914_),
    .A(_04193_),
    .B(_05644_));
 sg13g2_nor4_1 _14182_ (.A(net48),
    .B(_05912_),
    .C(_05913_),
    .D(_05914_),
    .Y(_05915_));
 sg13g2_a21oi_1 _14183_ (.A1(_01585_),
    .A2(net48),
    .Y(_01471_),
    .B1(_05915_));
 sg13g2_nor3_1 _14184_ (.A(net333),
    .B(net212),
    .C(_03518_),
    .Y(_05916_));
 sg13g2_nor4_1 _14185_ (.A(net285),
    .B(_04178_),
    .C(_05640_),
    .D(_05916_),
    .Y(_05917_));
 sg13g2_nor2b_1 _14186_ (.A(_05914_),
    .B_N(_05917_),
    .Y(_05918_));
 sg13g2_o21ai_1 _14187_ (.B1(_05918_),
    .Y(_05919_),
    .A1(net204),
    .A2(_05911_));
 sg13g2_o21ai_1 _14188_ (.B1(_05919_),
    .Y(_05920_),
    .A1(net216),
    .A2(_05808_));
 sg13g2_nand2_1 _14189_ (.Y(_05921_),
    .A(net3906),
    .B(net48));
 sg13g2_o21ai_1 _14190_ (.B1(_05921_),
    .Y(_01472_),
    .A1(net48),
    .A2(_05920_));
 sg13g2_nand2_1 _14191_ (.Y(_05922_),
    .A(_03486_),
    .B(_04177_));
 sg13g2_o21ai_1 _14192_ (.B1(_05922_),
    .Y(_05923_),
    .A1(_03575_),
    .A2(_05911_));
 sg13g2_a21oi_1 _14193_ (.A1(net217),
    .A2(_05923_),
    .Y(_05924_),
    .B1(_05820_));
 sg13g2_nor2_1 _14194_ (.A(net3930),
    .B(_05652_),
    .Y(_05925_));
 sg13g2_a21oi_1 _14195_ (.A1(net29),
    .A2(_05924_),
    .Y(_01473_),
    .B1(_05925_));
 sg13g2_o21ai_1 _14196_ (.B1(net218),
    .Y(_05926_),
    .A1(_03570_),
    .A2(_05908_));
 sg13g2_o21ai_1 _14197_ (.B1(_05826_),
    .Y(_05927_),
    .A1(_05911_),
    .A2(_05926_));
 sg13g2_mux2_1 _14198_ (.A0(net4022),
    .A1(_05927_),
    .S(net29),
    .X(_01474_));
 sg13g2_and2_1 _14199_ (.A(net216),
    .B(net109),
    .X(_05928_));
 sg13g2_o21ai_1 _14200_ (.B1(_05928_),
    .Y(_05929_),
    .A1(net284),
    .A2(_05643_));
 sg13g2_xor2_1 _14201_ (.B(\i_tinyqv.cpu.mem_op_increment_reg ),
    .A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .X(_05930_));
 sg13g2_nand3_1 _14202_ (.B(_05837_),
    .C(_05929_),
    .A(net88),
    .Y(_05931_));
 sg13g2_o21ai_1 _14203_ (.B1(_05931_),
    .Y(_05932_),
    .A1(net88),
    .A2(_05930_));
 sg13g2_nand2_1 _14204_ (.Y(_05933_),
    .A(net3999),
    .B(net64));
 sg13g2_o21ai_1 _14205_ (.B1(_05933_),
    .Y(_01475_),
    .A1(net64),
    .A2(_05932_));
 sg13g2_nand2_1 _14206_ (.Y(_05934_),
    .A(\i_tinyqv.cpu.mem_op_increment_reg ),
    .B(net557));
 sg13g2_a21o_1 _14207_ (.A2(\i_tinyqv.cpu.mem_op_increment_reg ),
    .A1(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .B1(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .X(_05935_));
 sg13g2_nand2_1 _14208_ (.Y(_05936_),
    .A(_05934_),
    .B(_05935_));
 sg13g2_and2_1 _14209_ (.A(_05628_),
    .B(_05644_),
    .X(_05937_));
 sg13g2_nor2b_1 _14210_ (.A(_04201_),
    .B_N(_05937_),
    .Y(_05938_));
 sg13g2_o21ai_1 _14211_ (.B1(net88),
    .Y(_05939_),
    .A1(_05840_),
    .A2(_05938_));
 sg13g2_o21ai_1 _14212_ (.B1(_05939_),
    .Y(_05940_),
    .A1(net89),
    .A2(_05936_));
 sg13g2_mux2_1 _14213_ (.A0(_05940_),
    .A1(net4003),
    .S(net64),
    .X(_01476_));
 sg13g2_nand3_1 _14214_ (.B(\i_tinyqv.cpu.mem_op_increment_reg ),
    .C(net557),
    .A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .Y(_05941_));
 sg13g2_xor2_1 _14215_ (.B(_05934_),
    .A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .X(_05942_));
 sg13g2_and3_1 _14216_ (.X(_05943_),
    .A(net216),
    .B(net120),
    .C(_05937_));
 sg13g2_o21ai_1 _14217_ (.B1(net88),
    .Y(_05944_),
    .A1(_05843_),
    .A2(_05943_));
 sg13g2_o21ai_1 _14218_ (.B1(_05944_),
    .Y(_05945_),
    .A1(net89),
    .A2(_05942_));
 sg13g2_mux2_1 _14219_ (.A0(_05945_),
    .A1(net4096),
    .S(net64),
    .X(_01477_));
 sg13g2_o21ai_1 _14220_ (.B1(_03533_),
    .Y(_05946_),
    .A1(_03556_),
    .A2(_05642_));
 sg13g2_a21oi_2 _14221_ (.B1(_05704_),
    .Y(_05947_),
    .A2(_05946_),
    .A1(_05928_));
 sg13g2_xnor2_1 _14222_ (.Y(_05948_),
    .A(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .B(_05941_));
 sg13g2_nand2_1 _14223_ (.Y(_05949_),
    .A(net90),
    .B(_05948_));
 sg13g2_o21ai_1 _14224_ (.B1(_05949_),
    .Y(_05950_),
    .A1(_04161_),
    .A2(_05947_));
 sg13g2_mux2_1 _14225_ (.A0(_05950_),
    .A1(net4070),
    .S(net64),
    .X(_01478_));
 sg13g2_o21ai_1 _14226_ (.B1(net216),
    .Y(_05951_),
    .A1(net282),
    .A2(_04193_));
 sg13g2_a21oi_1 _14227_ (.A1(net284),
    .A2(_05643_),
    .Y(_05952_),
    .B1(_05951_));
 sg13g2_a21oi_1 _14228_ (.A1(net285),
    .A2(_05905_),
    .Y(_05953_),
    .B1(_05952_));
 sg13g2_mux2_1 _14229_ (.A0(_00254_),
    .A1(_05953_),
    .S(net88),
    .X(_05954_));
 sg13g2_o21ai_1 _14230_ (.B1(net655),
    .Y(_05955_),
    .A1(_04165_),
    .A2(_05954_));
 sg13g2_a21oi_1 _14231_ (.A1(_01488_),
    .A2(_04165_),
    .Y(_01479_),
    .B1(_05955_));
 sg13g2_nor2b_1 _14232_ (.A(_05905_),
    .B_N(_05902_),
    .Y(_05956_));
 sg13g2_a21oi_1 _14233_ (.A1(_03522_),
    .A2(_05643_),
    .Y(_05957_),
    .B1(_05956_));
 sg13g2_o21ai_1 _14234_ (.B1(_05957_),
    .Y(_05958_),
    .A1(_03593_),
    .A2(_04193_));
 sg13g2_xor2_1 _14235_ (.B(net3444),
    .A(net3524),
    .X(_05959_));
 sg13g2_a21oi_1 _14236_ (.A1(net90),
    .A2(_05959_),
    .Y(_05960_),
    .B1(_04165_));
 sg13g2_o21ai_1 _14237_ (.B1(_05960_),
    .Y(_05961_),
    .A1(net90),
    .A2(_05958_));
 sg13g2_nand2_1 _14238_ (.Y(_05962_),
    .A(net3524),
    .B(_04165_));
 sg13g2_a21oi_1 _14239_ (.A1(_05961_),
    .A2(_05962_),
    .Y(_01480_),
    .B1(net510));
 sg13g2_nand2_1 _14240_ (.Y(_05963_),
    .A(net120),
    .B(_05643_));
 sg13g2_o21ai_1 _14241_ (.B1(_05963_),
    .Y(_05964_),
    .A1(_03575_),
    .A2(_04193_));
 sg13g2_a21o_1 _14242_ (.A2(_03500_),
    .A1(_02529_),
    .B1(_04165_),
    .X(_05965_));
 sg13g2_a22oi_1 _14243_ (.Y(_05966_),
    .B1(_05965_),
    .B2(net3217),
    .A2(_05964_),
    .A1(_05580_));
 sg13g2_nor2_1 _14244_ (.A(net510),
    .B(_05966_),
    .Y(_01481_));
 sg13g2_nor2_1 _14245_ (.A(net648),
    .B(_05903_),
    .Y(_05967_));
 sg13g2_a22oi_1 _14246_ (.Y(_01482_),
    .B1(_05967_),
    .B2(_05582_),
    .A2(net48),
    .A1(_01705_));
 sg13g2_nand3_1 _14247_ (.B(_03475_),
    .C(net88),
    .A(_02528_),
    .Y(_05968_));
 sg13g2_nand2_1 _14248_ (.Y(_05969_),
    .A(net3576),
    .B(_05579_));
 sg13g2_a21oi_1 _14249_ (.A1(_05968_),
    .A2(_05969_),
    .Y(_01483_),
    .B1(net511));
 sg13g2_nand2_1 _14250_ (.Y(_05970_),
    .A(_05579_),
    .B(_05968_));
 sg13g2_nand2b_1 _14251_ (.Y(_05971_),
    .B(_03499_),
    .A_N(_03595_));
 sg13g2_o21ai_1 _14252_ (.B1(net658),
    .Y(_05972_),
    .A1(net571),
    .A2(_05970_));
 sg13g2_a21oi_1 _14253_ (.A1(_05970_),
    .A2(_05971_),
    .Y(_01484_),
    .B1(_05972_));
 sg13g2_nor2b_1 _14254_ (.A(net2828),
    .B_N(_01095_),
    .Y(_01485_));
 sg13g2_nor4_1 _14255_ (.A(net648),
    .B(net99),
    .C(net80),
    .D(_03608_),
    .Y(_01486_));
 sg13g2_inv_1 _14257__3 (.Y(net2110),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _14258__4 (.Y(net2111),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _14259__5 (.Y(net2112),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _14260__6 (.Y(net2113),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _14261__7 (.Y(net2114),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _14262__8 (.Y(net2115),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _14263__9 (.Y(net2116),
    .A(clknet_leaf_32_clk));
 sg13g2_inv_1 _14264__10 (.Y(net2117),
    .A(clknet_leaf_32_clk));
 sg13g2_inv_1 _14265__11 (.Y(net2118),
    .A(clknet_leaf_32_clk));
 sg13g2_inv_1 _14266__12 (.Y(net2119),
    .A(clknet_leaf_32_clk));
 sg13g2_inv_1 _14267__13 (.Y(net2120),
    .A(clknet_leaf_32_clk));
 sg13g2_inv_1 _14268__14 (.Y(net2121),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 _14269__15 (.Y(net2122),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _14270__16 (.Y(net2123),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _14271__17 (.Y(net2124),
    .A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 _14272__18 (.Y(net2125),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _14273__19 (.Y(net2126),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _14274__20 (.Y(net2127),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _14275__21 (.Y(net2128),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _14276__22 (.Y(net2129),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _14277__23 (.Y(net2130),
    .A(clknet_leaf_25_clk));
 sg13g2_inv_1 _14278__24 (.Y(net2131),
    .A(clknet_leaf_24_clk));
 sg13g2_inv_1 _14279__25 (.Y(net2132),
    .A(clknet_leaf_35_clk));
 sg13g2_inv_1 _14280__26 (.Y(net2133),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _14281__27 (.Y(net2134),
    .A(clknet_leaf_27_clk));
 sg13g2_inv_1 _14282__28 (.Y(net2135),
    .A(clknet_leaf_24_clk));
 sg13g2_inv_1 _14283__29 (.Y(net2136),
    .A(clknet_leaf_24_clk));
 sg13g2_inv_1 _14284__30 (.Y(net2137),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _14285__31 (.Y(net2138),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _14286__32 (.Y(net2139),
    .A(clknet_leaf_30_clk));
 sg13g2_inv_1 _14287__33 (.Y(net2140),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _14288__34 (.Y(net2141),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 _14289__35 (.Y(net2142),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 _14290__36 (.Y(net2143),
    .A(clknet_leaf_8_clk));
 sg13g2_inv_1 _14291__37 (.Y(net2144),
    .A(clknet_leaf_7_clk));
 sg13g2_inv_1 _14292__38 (.Y(net2145),
    .A(clknet_leaf_3_clk));
 sg13g2_inv_1 _14293__39 (.Y(net2146),
    .A(clknet_leaf_36_clk));
 sg13g2_inv_1 _14294__40 (.Y(net2147),
    .A(clknet_leaf_36_clk));
 sg13g2_inv_1 _14295__41 (.Y(net2148),
    .A(clknet_leaf_35_clk));
 sg13g2_inv_1 _14296__42 (.Y(net2149),
    .A(clknet_leaf_36_clk));
 sg13g2_inv_1 _14297__43 (.Y(net2150),
    .A(clknet_leaf_26_clk));
 sg13g2_inv_1 _14298__44 (.Y(net2151),
    .A(clknet_leaf_24_clk));
 sg13g2_inv_1 _14299__45 (.Y(net2152),
    .A(clknet_leaf_26_clk));
 sg13g2_inv_1 _14300__46 (.Y(net2153),
    .A(clknet_leaf_25_clk));
 sg13g2_inv_1 _14301__47 (.Y(net2154),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _14302__48 (.Y(net2155),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _14303__49 (.Y(net2156),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 _14304__50 (.Y(net2157),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _14305__51 (.Y(net2158),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _14306__52 (.Y(net2159),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _14307__53 (.Y(net2160),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 _14308__54 (.Y(net2161),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _14309__55 (.Y(net2162),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _14310__56 (.Y(net2163),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _14311__57 (.Y(net2164),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _14312__58 (.Y(net2165),
    .A(clknet_leaf_7_clk));
 sg13g2_inv_1 _14313__59 (.Y(net2166),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _14314__60 (.Y(net2167),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _14315__61 (.Y(net2168),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _14316__62 (.Y(net2169),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _14317__63 (.Y(net2170),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _14318__64 (.Y(net2171),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _14319__65 (.Y(net2172),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _14320__66 (.Y(net2173),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _14321__67 (.Y(net2174),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _14322__68 (.Y(net2175),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _14323__69 (.Y(net2176),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _14324__70 (.Y(net2177),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _14325__71 (.Y(net2178),
    .A(clknet_leaf_4_clk));
 sg13g2_inv_1 _14326__72 (.Y(net2179),
    .A(clknet_leaf_0_clk));
 sg13g2_inv_1 _14327__73 (.Y(net2180),
    .A(clknet_leaf_0_clk));
 sg13g2_inv_1 _14328__74 (.Y(net2181),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _14329__75 (.Y(net2182),
    .A(clknet_leaf_0_clk));
 sg13g2_inv_1 _14330__76 (.Y(net2183),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _14331__77 (.Y(net2184),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _14332__78 (.Y(net2185),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _14333__79 (.Y(net2186),
    .A(clknet_leaf_22_clk));
 sg13g2_inv_1 _14334__80 (.Y(net2187),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _14335__81 (.Y(net2188),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _14336__82 (.Y(net2189),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _14337__83 (.Y(net2190),
    .A(clknet_leaf_22_clk));
 sg13g2_inv_1 _14338__84 (.Y(net2191),
    .A(clknet_leaf_24_clk));
 sg13g2_inv_1 _14339__85 (.Y(net2192),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _14340__86 (.Y(net2193),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _14341__87 (.Y(net2194),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _14342__88 (.Y(net2195),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _14343__89 (.Y(net2196),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _14344__90 (.Y(net2197),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _14345__91 (.Y(net2198),
    .A(clknet_leaf_22_clk));
 sg13g2_inv_1 _14346__92 (.Y(net2199),
    .A(clknet_leaf_22_clk));
 sg13g2_inv_1 _14347__93 (.Y(net2200),
    .A(clknet_leaf_24_clk));
 sg13g2_inv_1 _14348__94 (.Y(net2201),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _14349__95 (.Y(net2202),
    .A(clknet_leaf_22_clk));
 sg13g2_inv_1 _14350__96 (.Y(net2203),
    .A(clknet_leaf_0_clk));
 sg13g2_inv_1 _14351__97 (.Y(net2204),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _14352__98 (.Y(net2205),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _14353__99 (.Y(net2206),
    .A(clknet_leaf_0_clk));
 sg13g2_inv_1 _14354__100 (.Y(net2207),
    .A(clknet_leaf_22_clk));
 sg13g2_inv_1 _14355__101 (.Y(net2208),
    .A(clknet_leaf_22_clk));
 sg13g2_inv_1 _14356__102 (.Y(net2209),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _14357__103 (.Y(net2210),
    .A(clknet_leaf_2_clk));
 sg13g2_inv_1 _14358__104 (.Y(net2211),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _14359__105 (.Y(net2212),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _14360__106 (.Y(net2213),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _14361__107 (.Y(net2214),
    .A(clknet_leaf_0_clk));
 sg13g2_inv_1 _14362__108 (.Y(net2215),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _14363__109 (.Y(net2216),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 _14364__110 (.Y(net2217),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _14365__111 (.Y(net2218),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _14366__112 (.Y(net2219),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _14367__113 (.Y(net2220),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _14368__114 (.Y(net2221),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _14369__115 (.Y(net2222),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _14370__116 (.Y(net2223),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _14371__117 (.Y(net2224),
    .A(clknet_leaf_7_clk));
 sg13g2_inv_1 _14372__118 (.Y(net2225),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 _14373__119 (.Y(net2226),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 _14374__120 (.Y(net2227),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _14375__121 (.Y(net2228),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 _14376__122 (.Y(net2229),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 _14377__123 (.Y(net2230),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 _14378__124 (.Y(net2231),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _14379__125 (.Y(net2232),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 _14380__126 (.Y(net2233),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _14381__127 (.Y(net2234),
    .A(clknet_leaf_3_clk));
 sg13g2_inv_1 _14382__128 (.Y(net2235),
    .A(clknet_leaf_4_clk));
 sg13g2_inv_1 _14383__129 (.Y(net2236),
    .A(clknet_leaf_3_clk));
 sg13g2_inv_1 _14384__130 (.Y(net2237),
    .A(clknet_leaf_3_clk));
 sg13g2_inv_1 _14385__131 (.Y(net2238),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _14386__132 (.Y(net2239),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _14387__133 (.Y(net2240),
    .A(clknet_leaf_4_clk));
 sg13g2_inv_1 _14388__134 (.Y(net2241),
    .A(clknet_leaf_3_clk));
 sg13g2_inv_1 _14389__135 (.Y(net2242),
    .A(clknet_leaf_31_clk));
 sg13g2_inv_1 _14390__136 (.Y(net2243),
    .A(clknet_leaf_30_clk));
 sg13g2_inv_1 _14391__137 (.Y(net2244),
    .A(clknet_leaf_31_clk));
 sg13g2_inv_1 _14392__138 (.Y(net2245),
    .A(clknet_leaf_30_clk));
 sg13g2_inv_1 _14393__139 (.Y(net2246),
    .A(clknet_leaf_31_clk));
 sg13g2_inv_1 _14394__140 (.Y(net2247),
    .A(clknet_leaf_30_clk));
 sg13g2_inv_1 _14395__141 (.Y(net2248),
    .A(clknet_leaf_30_clk));
 sg13g2_inv_1 _14396__142 (.Y(net2249),
    .A(clknet_leaf_30_clk));
 sg13g2_inv_1 _14397__143 (.Y(net2250),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _14398__144 (.Y(net2251),
    .A(clknet_leaf_36_clk));
 sg13g2_inv_1 _14399__145 (.Y(net2252),
    .A(clknet_leaf_35_clk));
 sg13g2_inv_1 _14400__146 (.Y(net2253),
    .A(clknet_leaf_36_clk));
 sg13g2_inv_1 _14401__147 (.Y(net2254),
    .A(clknet_leaf_35_clk));
 sg13g2_inv_1 _14402__148 (.Y(net2255),
    .A(clknet_leaf_24_clk));
 sg13g2_inv_1 _14403__149 (.Y(net2256),
    .A(clknet_leaf_36_clk));
 sg13g2_inv_1 _14404__150 (.Y(net2257),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _14405__151 (.Y(net2258),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 _14406__152 (.Y(net2259),
    .A(clknet_leaf_25_clk));
 sg13g2_inv_1 _14407__153 (.Y(net2260),
    .A(clknet_leaf_2_clk));
 sg13g2_inv_1 _14408__154 (.Y(net2261),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _14409__155 (.Y(net2262),
    .A(clknet_leaf_27_clk));
 sg13g2_inv_1 _14410__156 (.Y(net2263),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 _14411__157 (.Y(net2264),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _14412__158 (.Y(net2265),
    .A(clknet_leaf_26_clk));
 sg13g2_inv_1 _14413__159 (.Y(net2266),
    .A(clknet_leaf_36_clk));
 sg13g2_inv_1 _14414__160 (.Y(net2267),
    .A(clknet_leaf_27_clk));
 sg13g2_inv_1 _14415__161 (.Y(net2268),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 _14416__162 (.Y(net2269),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 _14417__163 (.Y(net2270),
    .A(clknet_leaf_25_clk));
 sg13g2_inv_1 _14418__164 (.Y(net2271),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 _14419__165 (.Y(net2272),
    .A(clknet_leaf_25_clk));
 sg13g2_inv_1 _14420__166 (.Y(net2273),
    .A(clknet_leaf_26_clk));
 sg13g2_inv_1 _14421__167 (.Y(net2274),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 _14422__168 (.Y(net2275),
    .A(clknet_leaf_35_clk));
 sg13g2_inv_1 _14423__169 (.Y(net2276),
    .A(clknet_leaf_26_clk));
 sg13g2_inv_1 _14424__170 (.Y(net2277),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 _14425__171 (.Y(net2278),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _14426__172 (.Y(net2279),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 _14427__173 (.Y(net2280),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 _14428__174 (.Y(net2281),
    .A(clknet_leaf_26_clk));
 sg13g2_inv_1 _14429__175 (.Y(net2282),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _14430__176 (.Y(net2283),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _14431__177 (.Y(net2284),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _14432__178 (.Y(net2285),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _14433__179 (.Y(net2286),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _14434__180 (.Y(net2287),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _14435__181 (.Y(net2288),
    .A(clknet_leaf_8_clk));
 sg13g2_inv_1 _14436__182 (.Y(net2289),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _14437__183 (.Y(net2290),
    .A(clknet_leaf_32_clk));
 sg13g2_inv_1 _14438__184 (.Y(net2291),
    .A(clknet_leaf_31_clk));
 sg13g2_inv_1 _14439__185 (.Y(net2292),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _14440__186 (.Y(net2293),
    .A(clknet_leaf_2_clk));
 sg13g2_inv_1 _14441__187 (.Y(net2294),
    .A(clknet_leaf_30_clk));
 sg13g2_inv_1 _14442__188 (.Y(net2295),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 _14443__189 (.Y(net2296),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 _14444__190 (.Y(net2297),
    .A(clknet_leaf_31_clk));
 sg13g2_inv_1 _14445__191 (.Y(net2298),
    .A(clknet_leaf_31_clk));
 sg13g2_inv_1 _14446__192 (.Y(net2299),
    .A(clknet_leaf_29_clk));
 sg13g2_inv_1 _14447__193 (.Y(net2300),
    .A(clknet_leaf_29_clk));
 sg13g2_inv_1 _14448__194 (.Y(net2301),
    .A(clknet_leaf_29_clk));
 sg13g2_inv_1 _14449__195 (.Y(net2302),
    .A(clknet_leaf_29_clk));
 sg13g2_inv_1 _14450__196 (.Y(net2303),
    .A(clknet_leaf_28_clk));
 sg13g2_inv_1 _14451__197 (.Y(net2304),
    .A(clknet_leaf_30_clk));
 sg13g2_inv_1 _14452__198 (.Y(net2305),
    .A(clknet_leaf_29_clk));
 sg13g2_inv_1 _14453__199 (.Y(net2306),
    .A(clknet_leaf_2_clk));
 sg13g2_inv_1 _14454__200 (.Y(net2307),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _14455__201 (.Y(net2308),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _14456__202 (.Y(net2309),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _14457__203 (.Y(net2310),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _14458__204 (.Y(net2311),
    .A(clknet_leaf_7_clk));
 sg13g2_inv_1 _14459__205 (.Y(net2312),
    .A(clknet_leaf_7_clk));
 sg13g2_inv_1 _14460__206 (.Y(net2313),
    .A(clknet_leaf_3_clk));
 sg13g2_inv_1 _14461__207 (.Y(net2314),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 _14462__208 (.Y(net2315),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _14463__209 (.Y(net2316),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _14464__210 (.Y(net2317),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 _14465__211 (.Y(net2318),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _14466__212 (.Y(net2319),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _14467__213 (.Y(net2320),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 _14468__214 (.Y(net2321),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _14469__215 (.Y(net2322),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 _14470__216 (.Y(net2323),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _14471__217 (.Y(net2324),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 _14472__218 (.Y(net2325),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _14473__219 (.Y(net2326),
    .A(clknet_leaf_35_clk));
 sg13g2_inv_1 _14474__220 (.Y(net2327),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 _14475__221 (.Y(net2328),
    .A(clknet_leaf_36_clk));
 sg13g2_inv_1 _14476__222 (.Y(net2329),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 _14477__223 (.Y(net2330),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 _14478__224 (.Y(net2331),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 _14479__225 (.Y(net2332),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 _14480__226 (.Y(net2333),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 _14481__227 (.Y(net2334),
    .A(clknet_leaf_0_clk));
 sg13g2_inv_1 _14482__228 (.Y(net2335),
    .A(clknet_leaf_0_clk));
 sg13g2_inv_1 _14483__229 (.Y(net2336),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _14484__230 (.Y(net2337),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 _14485__231 (.Y(net2338),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 _14486__232 (.Y(net2339),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _14487__233 (.Y(net2340),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _14488__234 (.Y(net2341),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _14489__235 (.Y(net2342),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _14490__236 (.Y(net2343),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 _14491__237 (.Y(net2344),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _14492__238 (.Y(net2345),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _14493__239 (.Y(net2346),
    .A(clknet_leaf_2_clk));
 sg13g2_inv_1 _14494__240 (.Y(net2347),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _14495__241 (.Y(net2348),
    .A(clknet_leaf_2_clk));
 sg13g2_inv_1 _14496__242 (.Y(net2349),
    .A(clknet_leaf_2_clk));
 sg13g2_inv_1 _14497__243 (.Y(net2350),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _14498__244 (.Y(net2351),
    .A(clknet_leaf_8_clk));
 sg13g2_inv_1 _14499__245 (.Y(net2352),
    .A(clknet_leaf_8_clk));
 sg13g2_inv_1 _14500__246 (.Y(net2353),
    .A(clknet_leaf_7_clk));
 sg13g2_inv_1 _14501__247 (.Y(net2354),
    .A(clknet_leaf_28_clk));
 sg13g2_inv_1 _14502__248 (.Y(net2355),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _14503__249 (.Y(net2356),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _14504__250 (.Y(net2357),
    .A(clknet_leaf_28_clk));
 sg13g2_inv_1 _14505__251 (.Y(net2358),
    .A(clknet_leaf_27_clk));
 sg13g2_inv_1 _14506__252 (.Y(net2359),
    .A(clknet_leaf_22_clk));
 sg13g2_inv_1 _14507__253 (.Y(net2360),
    .A(clknet_leaf_27_clk));
 sg13g2_inv_1 _14508__254 (.Y(net2361),
    .A(clknet_leaf_27_clk));
 sg13g2_inv_1 _14509__255 (.Y(net2362),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _14510__256 (.Y(net2363),
    .A(clknet_leaf_28_clk));
 sg13g2_inv_1 _14511__257 (.Y(net2364),
    .A(clknet_leaf_28_clk));
 sg13g2_inv_1 _14512__258 (.Y(net2365),
    .A(clknet_leaf_28_clk));
 sg13g2_inv_1 _14513__259 (.Y(net2366),
    .A(clknet_leaf_27_clk));
 sg13g2_inv_1 _14514__260 (.Y(net2367),
    .A(clknet_leaf_28_clk));
 sg13g2_inv_1 _14515__261 (.Y(net2368),
    .A(clknet_leaf_28_clk));
 sg13g2_inv_1 _14516__262 (.Y(net2369),
    .A(clknet_leaf_27_clk));
 sg13g2_inv_1 _14517__263 (.Y(net2370),
    .A(clknet_leaf_4_clk));
 sg13g2_inv_1 _14518__264 (.Y(net2371),
    .A(clknet_leaf_4_clk));
 sg13g2_inv_1 _14519__265 (.Y(net2372),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _14520__266 (.Y(net2373),
    .A(clknet_leaf_2_clk));
 sg13g2_inv_1 _14521__267 (.Y(net2374),
    .A(clknet_leaf_4_clk));
 sg13g2_inv_1 _14522__268 (.Y(net2375),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _14523__269 (.Y(net2376),
    .A(clknet_leaf_4_clk));
 sg13g2_inv_1 _14524__270 (.Y(net2377),
    .A(clknet_leaf_3_clk));
 sg13g2_inv_1 _14525__271 (.Y(net2378),
    .A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 _14526__272 (.Y(net2379),
    .A(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_dfrbp_1 _14527_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net2097),
    .D(net2724),
    .Q_N(_06723_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[0] ));
 sg13g2_dfrbp_1 _14528_ (.CLK(clknet_leaf_119_clk_regs),
    .RESET_B(net2098),
    .D(net2777),
    .Q_N(_06724_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[1] ));
 sg13g2_dfrbp_1 _14529_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net2099),
    .D(net2399),
    .Q_N(_06725_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[2] ));
 sg13g2_dfrbp_1 _14530_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net2100),
    .D(net2534),
    .Q_N(_06726_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[3] ));
 sg13g2_dfrbp_1 _14531_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net2101),
    .D(net2583),
    .Q_N(_06727_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ));
 sg13g2_dfrbp_1 _14532_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net2102),
    .D(net2710),
    .Q_N(_06728_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ));
 sg13g2_dfrbp_1 _14533_ (.CLK(clknet_leaf_119_clk_regs),
    .RESET_B(net2103),
    .D(net2538),
    .Q_N(_06729_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ));
 sg13g2_dfrbp_1 _14534_ (.CLK(clknet_leaf_119_clk_regs),
    .RESET_B(net2104),
    .D(net2618),
    .Q_N(_06730_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ));
 sg13g2_dfrbp_1 _14535_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net2105),
    .D(net2784),
    .Q_N(_06731_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ));
 sg13g2_dfrbp_1 _14536_ (.CLK(clknet_leaf_127_clk_regs),
    .RESET_B(net2106),
    .D(net2476),
    .Q_N(_06732_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ));
 sg13g2_dfrbp_1 _14537_ (.CLK(clknet_leaf_119_clk_regs),
    .RESET_B(net2107),
    .D(net2594),
    .Q_N(_06733_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ));
 sg13g2_dfrbp_1 _14538_ (.CLK(clknet_leaf_119_clk_regs),
    .RESET_B(net663),
    .D(net2708),
    .Q_N(_06734_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ));
 sg13g2_dfrbp_1 _14539_ (.CLK(clknet_leaf_123_clk_regs),
    .RESET_B(net664),
    .D(net2493),
    .Q_N(_06735_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ));
 sg13g2_dfrbp_1 _14540_ (.CLK(clknet_leaf_127_clk_regs),
    .RESET_B(net665),
    .D(net2704),
    .Q_N(_06736_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ));
 sg13g2_dfrbp_1 _14541_ (.CLK(clknet_leaf_119_clk_regs),
    .RESET_B(net666),
    .D(net2433),
    .Q_N(_06737_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ));
 sg13g2_dfrbp_1 _14542_ (.CLK(clknet_leaf_119_clk_regs),
    .RESET_B(net667),
    .D(net2718),
    .Q_N(_06738_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ));
 sg13g2_dfrbp_1 _14543_ (.CLK(clknet_leaf_123_clk_regs),
    .RESET_B(net668),
    .D(net2674),
    .Q_N(_06739_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ));
 sg13g2_dfrbp_1 _14544_ (.CLK(clknet_leaf_127_clk_regs),
    .RESET_B(net669),
    .D(net2641),
    .Q_N(_06740_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ));
 sg13g2_dfrbp_1 _14545_ (.CLK(clknet_leaf_119_clk_regs),
    .RESET_B(net670),
    .D(net2757),
    .Q_N(_06741_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ));
 sg13g2_dfrbp_1 _14546_ (.CLK(clknet_leaf_126_clk_regs),
    .RESET_B(net671),
    .D(net2658),
    .Q_N(_06742_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ));
 sg13g2_dfrbp_1 _14547_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net672),
    .D(net2547),
    .Q_N(_06743_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ));
 sg13g2_dfrbp_1 _14548_ (.CLK(clknet_leaf_127_clk_regs),
    .RESET_B(net673),
    .D(net2650),
    .Q_N(_06744_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ));
 sg13g2_dfrbp_1 _14549_ (.CLK(clknet_leaf_126_clk_regs),
    .RESET_B(net674),
    .D(net2612),
    .Q_N(_06745_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ));
 sg13g2_dfrbp_1 _14550_ (.CLK(clknet_leaf_126_clk_regs),
    .RESET_B(net675),
    .D(net2545),
    .Q_N(_06746_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ));
 sg13g2_dfrbp_1 _14551_ (.CLK(clknet_leaf_123_clk_regs),
    .RESET_B(net676),
    .D(net2596),
    .Q_N(_06747_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ));
 sg13g2_dfrbp_1 _14552_ (.CLK(clknet_leaf_127_clk_regs),
    .RESET_B(net677),
    .D(net2521),
    .Q_N(_06748_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ));
 sg13g2_dfrbp_1 _14553_ (.CLK(clknet_leaf_126_clk_regs),
    .RESET_B(net683),
    .D(net2445),
    .Q_N(_06749_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ));
 sg13g2_dfrbp_1 _14554_ (.CLK(clknet_leaf_126_clk_regs),
    .RESET_B(net2096),
    .D(net2443),
    .Q_N(_06722_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ));
 sg13g2_dfrbp_1 _14555_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net1565),
    .D(net3845),
    .Q_N(_06721_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ));
 sg13g2_dfrbp_1 _14556_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net1564),
    .D(_00593_),
    .Q_N(_06720_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ));
 sg13g2_dfrbp_1 _14557_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net1563),
    .D(_00594_),
    .Q_N(_06719_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ));
 sg13g2_dfrbp_1 _14558_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net1562),
    .D(_00595_),
    .Q_N(_06718_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ));
 sg13g2_dfrbp_1 _14559_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net684),
    .D(net3885),
    .Q_N(_00265_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.cy ));
 sg13g2_dfrbp_1 _14560_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net685),
    .D(net2813),
    .Q_N(_06750_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[0] ));
 sg13g2_dfrbp_1 _14561_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net686),
    .D(net2825),
    .Q_N(_06751_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[1] ));
 sg13g2_dfrbp_1 _14562_ (.CLK(clknet_leaf_127_clk_regs),
    .RESET_B(net687),
    .D(net2807),
    .Q_N(_06752_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[2] ));
 sg13g2_dfrbp_1 _14563_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net688),
    .D(net2472),
    .Q_N(_06753_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[3] ));
 sg13g2_dfrbp_1 _14564_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net689),
    .D(net2764),
    .Q_N(_06754_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ));
 sg13g2_dfrbp_1 _14565_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net690),
    .D(net2478),
    .Q_N(_06755_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ));
 sg13g2_dfrbp_1 _14566_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net691),
    .D(net2567),
    .Q_N(_06756_),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ));
 sg13g2_dfrbp_1 _14567_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net692),
    .D(net2570),
    .Q_N(_06757_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ));
 sg13g2_dfrbp_1 _14568_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net693),
    .D(net2750),
    .Q_N(_06758_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ));
 sg13g2_dfrbp_1 _14569_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net694),
    .D(net2667),
    .Q_N(_06759_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ));
 sg13g2_dfrbp_1 _14570_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net695),
    .D(net2497),
    .Q_N(_06760_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ));
 sg13g2_dfrbp_1 _14571_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net696),
    .D(net2574),
    .Q_N(_06761_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ));
 sg13g2_dfrbp_1 _14572_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net697),
    .D(net2556),
    .Q_N(_06762_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ));
 sg13g2_dfrbp_1 _14573_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net698),
    .D(net2522),
    .Q_N(_06763_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ));
 sg13g2_dfrbp_1 _14574_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net699),
    .D(net2716),
    .Q_N(_06764_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ));
 sg13g2_dfrbp_1 _14575_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net700),
    .D(net2722),
    .Q_N(_06765_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ));
 sg13g2_dfrbp_1 _14576_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net701),
    .D(net2730),
    .Q_N(_06766_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ));
 sg13g2_dfrbp_1 _14577_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net702),
    .D(net2701),
    .Q_N(_06767_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ));
 sg13g2_dfrbp_1 _14578_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net703),
    .D(net2616),
    .Q_N(_06768_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ));
 sg13g2_dfrbp_1 _14579_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net704),
    .D(net2484),
    .Q_N(_06769_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ));
 sg13g2_dfrbp_1 _14580_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net705),
    .D(net2744),
    .Q_N(_06770_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ));
 sg13g2_dfrbp_1 _14581_ (.CLK(clknet_leaf_126_clk_regs),
    .RESET_B(net706),
    .D(net2765),
    .Q_N(_06771_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ));
 sg13g2_dfrbp_1 _14582_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net707),
    .D(net2715),
    .Q_N(_06772_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ));
 sg13g2_dfrbp_1 _14583_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net708),
    .D(net2615),
    .Q_N(_06773_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ));
 sg13g2_dfrbp_1 _14584_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net709),
    .D(net2516),
    .Q_N(_06774_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ));
 sg13g2_dfrbp_1 _14585_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net710),
    .D(net2491),
    .Q_N(_06775_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ));
 sg13g2_dfrbp_1 _14586_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net717),
    .D(net2697),
    .Q_N(_06776_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ));
 sg13g2_dfrbp_1 _14587_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net1561),
    .D(net2711),
    .Q_N(_06717_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ));
 sg13g2_dfrbp_1 _14588_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net1560),
    .D(_00597_),
    .Q_N(_06716_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[4] ));
 sg13g2_dfrbp_1 _14589_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net1559),
    .D(_00598_),
    .Q_N(_06715_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.cy ));
 sg13g2_dfrbp_1 _14590_ (.CLK(clknet_leaf_123_clk_regs),
    .RESET_B(net1558),
    .D(net3646),
    .Q_N(_06714_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ));
 sg13g2_dfrbp_1 _14591_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net1557),
    .D(_00600_),
    .Q_N(_06713_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ));
 sg13g2_dfrbp_1 _14592_ (.CLK(clknet_leaf_126_clk_regs),
    .RESET_B(net1556),
    .D(_00601_),
    .Q_N(_06712_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ));
 sg13g2_dfrbp_1 _14593_ (.CLK(clknet_leaf_126_clk_regs),
    .RESET_B(net718),
    .D(_00602_),
    .Q_N(_06777_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ));
 sg13g2_dfrbp_1 _14594_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net719),
    .D(net2760),
    .Q_N(_06778_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ));
 sg13g2_dfrbp_1 _14595_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net720),
    .D(net2624),
    .Q_N(_00127_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ));
 sg13g2_dfrbp_1 _14596_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net721),
    .D(net2394),
    .Q_N(_00126_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ));
 sg13g2_dfrbp_1 _14597_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net722),
    .D(net2460),
    .Q_N(_00123_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ));
 sg13g2_dfrbp_1 _14598_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net723),
    .D(net2573),
    .Q_N(_06779_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 _14599_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net724),
    .D(net2467),
    .Q_N(_06780_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 _14600_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net725),
    .D(net2677),
    .Q_N(_06781_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 _14601_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net726),
    .D(net2587),
    .Q_N(_06782_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 _14602_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net727),
    .D(net2699),
    .Q_N(_06783_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 _14603_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net728),
    .D(net2627),
    .Q_N(_06784_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 _14604_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net729),
    .D(net2693),
    .Q_N(_06785_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 _14605_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net730),
    .D(net2703),
    .Q_N(_06786_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 _14606_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net731),
    .D(net2449),
    .Q_N(_06787_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 _14607_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net732),
    .D(net2510),
    .Q_N(_06788_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 _14608_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net733),
    .D(net2588),
    .Q_N(_06789_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 _14609_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net734),
    .D(net2660),
    .Q_N(_06790_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 _14610_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net735),
    .D(net2638),
    .Q_N(_06791_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 _14611_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net736),
    .D(net2620),
    .Q_N(_06792_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 _14612_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net737),
    .D(net2561),
    .Q_N(_06793_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 _14613_ (.CLK(clknet_leaf_121_clk_regs),
    .RESET_B(net738),
    .D(net2815),
    .Q_N(_06794_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 _14614_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net739),
    .D(net2670),
    .Q_N(_06795_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 _14615_ (.CLK(clknet_leaf_122_clk_regs),
    .RESET_B(net740),
    .D(net2779),
    .Q_N(_06796_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 _14616_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net741),
    .D(net2621),
    .Q_N(_06797_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 _14617_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net742),
    .D(net2513),
    .Q_N(_06798_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 _14618_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net743),
    .D(net2754),
    .Q_N(_06799_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 _14619_ (.CLK(clknet_leaf_123_clk_regs),
    .RESET_B(net744),
    .D(net2492),
    .Q_N(_06800_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 _14620_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net745),
    .D(net2663),
    .Q_N(_06801_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 _14621_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net746),
    .D(net2404),
    .Q_N(_06802_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 _14622_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net747),
    .D(net3589),
    .Q_N(_06803_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 _14623_ (.CLK(clknet_leaf_123_clk_regs),
    .RESET_B(net748),
    .D(_00087_),
    .Q_N(_06804_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 _14624_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net749),
    .D(_00088_),
    .Q_N(_06805_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 _14625_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net750),
    .D(_00089_),
    .Q_N(_06806_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 _14626_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net751),
    .D(net2625),
    .Q_N(_06807_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ));
 sg13g2_dfrbp_1 _14627_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net752),
    .D(net2734),
    .Q_N(_06808_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ));
 sg13g2_dfrbp_1 _14628_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net753),
    .D(net2520),
    .Q_N(_06809_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ));
 sg13g2_dfrbp_1 _14629_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net754),
    .D(net2606),
    .Q_N(_06810_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ));
 sg13g2_dfrbp_1 _14630_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net755),
    .D(net2422),
    .Q_N(_06811_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 _14631_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net756),
    .D(net2740),
    .Q_N(_06812_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 _14632_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net757),
    .D(net2712),
    .Q_N(_06813_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 _14633_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net758),
    .D(net2640),
    .Q_N(_06814_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 _14634_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net759),
    .D(net2598),
    .Q_N(_06815_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 _14635_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net760),
    .D(net2792),
    .Q_N(_06816_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 _14636_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net761),
    .D(net2662),
    .Q_N(_06817_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 _14637_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net762),
    .D(net2482),
    .Q_N(_06818_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 _14638_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net763),
    .D(net2565),
    .Q_N(_06819_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 _14639_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net764),
    .D(net2503),
    .Q_N(_06820_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 _14640_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net765),
    .D(net2508),
    .Q_N(_06821_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 _14641_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net766),
    .D(net2564),
    .Q_N(_06822_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 _14642_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net767),
    .D(net2589),
    .Q_N(_06823_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 _14643_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net768),
    .D(net2398),
    .Q_N(_06824_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 _14644_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net769),
    .D(net2487),
    .Q_N(_06825_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 _14645_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net770),
    .D(net2633),
    .Q_N(_06826_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 _14646_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net771),
    .D(net2733),
    .Q_N(_06827_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 _14647_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net772),
    .D(net2786),
    .Q_N(_06828_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 _14648_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net773),
    .D(net2785),
    .Q_N(_06829_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 _14649_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net774),
    .D(net2480),
    .Q_N(_06830_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 _14650_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net775),
    .D(net2553),
    .Q_N(_06831_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 _14651_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net776),
    .D(net2393),
    .Q_N(_06832_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 _14652_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net777),
    .D(net2540),
    .Q_N(_06833_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 _14653_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net778),
    .D(net2794),
    .Q_N(_06834_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 _14654_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net779),
    .D(_00082_),
    .Q_N(_06835_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 _14655_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net780),
    .D(_00083_),
    .Q_N(_06836_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 _14656_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net781),
    .D(_00084_),
    .Q_N(_06837_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 _14657_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net782),
    .D(_00085_),
    .Q_N(_06838_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 _14658_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net783),
    .D(net2632),
    .Q_N(_06839_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ));
 sg13g2_dfrbp_1 _14659_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net784),
    .D(net2713),
    .Q_N(_06840_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ));
 sg13g2_dfrbp_1 _14660_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net785),
    .D(net2523),
    .Q_N(_06841_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ));
 sg13g2_dfrbp_1 _14661_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net786),
    .D(net2767),
    .Q_N(_06842_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ));
 sg13g2_dfrbp_1 _14662_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net787),
    .D(net2557),
    .Q_N(_06843_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 _14663_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net788),
    .D(net2576),
    .Q_N(_06844_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 _14664_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net789),
    .D(net2529),
    .Q_N(_06845_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 _14665_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net790),
    .D(net2411),
    .Q_N(_06846_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 _14666_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net791),
    .D(net2698),
    .Q_N(_06847_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 _14667_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net792),
    .D(net2692),
    .Q_N(_06848_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 _14668_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net793),
    .D(net2423),
    .Q_N(_06849_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 _14669_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net794),
    .D(net2438),
    .Q_N(_06850_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 _14670_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net795),
    .D(net2469),
    .Q_N(_06851_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 _14671_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net796),
    .D(net2577),
    .Q_N(_06852_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 _14672_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net797),
    .D(net2763),
    .Q_N(_06853_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 _14673_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net798),
    .D(net2751),
    .Q_N(_06854_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 _14674_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net799),
    .D(net2611),
    .Q_N(_06855_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 _14675_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net800),
    .D(net2601),
    .Q_N(_06856_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 _14676_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net801),
    .D(net2549),
    .Q_N(_06857_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 _14677_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net802),
    .D(net2431),
    .Q_N(_06858_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 _14678_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net803),
    .D(net2439),
    .Q_N(_06859_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 _14679_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net804),
    .D(net2626),
    .Q_N(_06860_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 _14680_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net805),
    .D(net2473),
    .Q_N(_06861_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 _14681_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net806),
    .D(net2731),
    .Q_N(_06862_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 _14682_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net807),
    .D(net2434),
    .Q_N(_06863_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 _14683_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net808),
    .D(net2408),
    .Q_N(_06864_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 _14684_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net809),
    .D(net2474),
    .Q_N(_06865_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 _14685_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net810),
    .D(net2599),
    .Q_N(_06866_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 _14686_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net811),
    .D(_00078_),
    .Q_N(_06867_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 _14687_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net812),
    .D(_00079_),
    .Q_N(_06868_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 _14688_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net813),
    .D(_00080_),
    .Q_N(_06869_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 _14689_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net814),
    .D(_00081_),
    .Q_N(_06870_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 _14690_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net815),
    .D(net2689),
    .Q_N(_06871_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ));
 sg13g2_dfrbp_1 _14691_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net816),
    .D(net2459),
    .Q_N(_06872_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ));
 sg13g2_dfrbp_1 _14692_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net817),
    .D(net2688),
    .Q_N(_06873_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ));
 sg13g2_dfrbp_1 _14693_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net818),
    .D(net2748),
    .Q_N(_06874_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ));
 sg13g2_dfrbp_1 _14694_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net819),
    .D(net2500),
    .Q_N(_06875_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 _14695_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net820),
    .D(net2406),
    .Q_N(_06876_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 _14696_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net821),
    .D(net2546),
    .Q_N(_06877_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 _14697_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net822),
    .D(net2395),
    .Q_N(_06878_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 _14698_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net823),
    .D(net2686),
    .Q_N(_06879_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 _14699_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net824),
    .D(net2672),
    .Q_N(_06880_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 _14700_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net825),
    .D(net2560),
    .Q_N(_06881_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 _14701_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net826),
    .D(net2762),
    .Q_N(_06882_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 _14702_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net827),
    .D(net2592),
    .Q_N(_06883_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 _14703_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net828),
    .D(net2481),
    .Q_N(_06884_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 _14704_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net829),
    .D(net2723),
    .Q_N(_06885_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 _14705_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net830),
    .D(net2629),
    .Q_N(_06886_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 _14706_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net831),
    .D(net2669),
    .Q_N(_06887_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 _14707_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net832),
    .D(net2466),
    .Q_N(_06888_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 _14708_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net833),
    .D(net2544),
    .Q_N(_06889_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 _14709_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net834),
    .D(net2691),
    .Q_N(_06890_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 _14710_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net835),
    .D(net2485),
    .Q_N(_06891_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 _14711_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net836),
    .D(net2820),
    .Q_N(_06892_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 _14712_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net837),
    .D(net2495),
    .Q_N(_06893_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 _14713_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net838),
    .D(net2648),
    .Q_N(_06894_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 _14714_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net839),
    .D(net2471),
    .Q_N(_06895_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 _14715_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net840),
    .D(net2695),
    .Q_N(_06896_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 _14716_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net841),
    .D(net2496),
    .Q_N(_06897_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 _14717_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net842),
    .D(net2668),
    .Q_N(_06898_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 _14718_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net843),
    .D(_00074_),
    .Q_N(_06899_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 _14719_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net844),
    .D(_00075_),
    .Q_N(_06900_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 _14720_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net845),
    .D(_00076_),
    .Q_N(_06901_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 _14721_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net846),
    .D(_00077_),
    .Q_N(_06902_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 _14722_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net847),
    .D(net2653),
    .Q_N(_06903_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ));
 sg13g2_dfrbp_1 _14723_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net848),
    .D(net2707),
    .Q_N(_06904_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ));
 sg13g2_dfrbp_1 _14724_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net849),
    .D(net2652),
    .Q_N(_06905_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ));
 sg13g2_dfrbp_1 _14725_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net850),
    .D(net2543),
    .Q_N(_06906_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ));
 sg13g2_dfrbp_1 _14726_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net851),
    .D(net2426),
    .Q_N(_06907_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 _14727_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net852),
    .D(net2412),
    .Q_N(_06908_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 _14728_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net853),
    .D(net2518),
    .Q_N(_06909_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 _14729_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net854),
    .D(net2468),
    .Q_N(_06910_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 _14730_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net855),
    .D(net2608),
    .Q_N(_06911_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 _14731_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net856),
    .D(net2591),
    .Q_N(_06912_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 _14732_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net857),
    .D(net2645),
    .Q_N(_06913_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 _14733_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net858),
    .D(net2421),
    .Q_N(_06914_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 _14734_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net859),
    .D(net2607),
    .Q_N(_06915_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 _14735_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net860),
    .D(net2427),
    .Q_N(_06916_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 _14736_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net861),
    .D(net2729),
    .Q_N(_06917_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 _14737_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net862),
    .D(net2541),
    .Q_N(_06918_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 _14738_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net863),
    .D(net2732),
    .Q_N(_06919_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 _14739_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net864),
    .D(net2542),
    .Q_N(_06920_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 _14740_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net865),
    .D(net2428),
    .Q_N(_06921_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 _14741_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net866),
    .D(net2535),
    .Q_N(_06922_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 _14742_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net867),
    .D(net2597),
    .Q_N(_06923_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 _14743_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net868),
    .D(net2582),
    .Q_N(_06924_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 _14744_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net869),
    .D(net2634),
    .Q_N(_06925_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 _14745_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net870),
    .D(net2782),
    .Q_N(_06926_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 _14746_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net871),
    .D(net2605),
    .Q_N(_06927_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 _14747_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net872),
    .D(net2788),
    .Q_N(_06928_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 _14748_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net873),
    .D(net2635),
    .Q_N(_06929_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 _14749_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net874),
    .D(net2819),
    .Q_N(_06930_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 _14750_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net875),
    .D(_00070_),
    .Q_N(_06931_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 _14751_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net876),
    .D(_00071_),
    .Q_N(_06932_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 _14752_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net877),
    .D(_00072_),
    .Q_N(_06933_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 _14753_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net878),
    .D(_00073_),
    .Q_N(_06934_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 _14754_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net879),
    .D(net2679),
    .Q_N(_06935_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ));
 sg13g2_dfrbp_1 _14755_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net880),
    .D(net2700),
    .Q_N(_06936_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ));
 sg13g2_dfrbp_1 _14756_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net881),
    .D(net2569),
    .Q_N(_06937_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ));
 sg13g2_dfrbp_1 _14757_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net882),
    .D(net2814),
    .Q_N(_06938_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ));
 sg13g2_dfrbp_1 _14758_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net883),
    .D(net2507),
    .Q_N(_06939_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 _14759_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net884),
    .D(net2403),
    .Q_N(_06940_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 _14760_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net885),
    .D(net2578),
    .Q_N(_06941_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 _14761_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net886),
    .D(net2571),
    .Q_N(_06942_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 _14762_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net887),
    .D(net2551),
    .Q_N(_06943_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 _14763_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net888),
    .D(net2639),
    .Q_N(_06944_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 _14764_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net889),
    .D(net2409),
    .Q_N(_06945_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 _14765_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net890),
    .D(net2572),
    .Q_N(_06946_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 _14766_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net891),
    .D(net2690),
    .Q_N(_06947_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 _14767_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net892),
    .D(net2477),
    .Q_N(_06948_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 _14768_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net893),
    .D(net2738),
    .Q_N(_06949_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 _14769_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net894),
    .D(net2656),
    .Q_N(_06950_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 _14770_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net895),
    .D(net2486),
    .Q_N(_06951_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 _14771_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net896),
    .D(net2665),
    .Q_N(_06952_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 _14772_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net897),
    .D(net2425),
    .Q_N(_06953_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 _14773_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net898),
    .D(net2489),
    .Q_N(_06954_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 _14774_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net899),
    .D(net2511),
    .Q_N(_06955_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 _14775_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net900),
    .D(net2526),
    .Q_N(_06956_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 _14776_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net901),
    .D(net2558),
    .Q_N(_06957_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 _14777_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net902),
    .D(net2405),
    .Q_N(_06958_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 _14778_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net903),
    .D(net2396),
    .Q_N(_06959_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 _14779_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net904),
    .D(net2462),
    .Q_N(_06960_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 _14780_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net905),
    .D(net2397),
    .Q_N(_06961_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 _14781_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net906),
    .D(net2696),
    .Q_N(_06962_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 _14782_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net907),
    .D(_00066_),
    .Q_N(_06963_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 _14783_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net908),
    .D(_00067_),
    .Q_N(_06964_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 _14784_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net909),
    .D(_00068_),
    .Q_N(_06965_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 _14785_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net910),
    .D(_00069_),
    .Q_N(_06966_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 _14786_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net911),
    .D(net2609),
    .Q_N(_06967_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ));
 sg13g2_dfrbp_1 _14787_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net912),
    .D(net2530),
    .Q_N(_06968_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ));
 sg13g2_dfrbp_1 _14788_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net913),
    .D(net2617),
    .Q_N(_06969_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ));
 sg13g2_dfrbp_1 _14789_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net914),
    .D(net2647),
    .Q_N(_06970_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ));
 sg13g2_dfrbp_1 _14790_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net915),
    .D(net2502),
    .Q_N(_06971_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 _14791_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net916),
    .D(net2604),
    .Q_N(_06972_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 _14792_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net917),
    .D(net2475),
    .Q_N(_06973_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 _14793_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net918),
    .D(net2407),
    .Q_N(_06974_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 _14794_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net919),
    .D(net2504),
    .Q_N(_06975_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 _14795_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net920),
    .D(net2675),
    .Q_N(_06976_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 _14796_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net921),
    .D(net2429),
    .Q_N(_06977_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 _14797_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net922),
    .D(net2671),
    .Q_N(_06978_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 _14798_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net923),
    .D(net2415),
    .Q_N(_06979_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 _14799_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net924),
    .D(net2401),
    .Q_N(_06980_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 _14800_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net925),
    .D(net2651),
    .Q_N(_06981_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 _14801_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net926),
    .D(net2458),
    .Q_N(_06982_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 _14802_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net927),
    .D(net2600),
    .Q_N(_06983_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 _14803_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net928),
    .D(net2446),
    .Q_N(_06984_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 _14804_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net929),
    .D(net2437),
    .Q_N(_06985_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 _14805_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net930),
    .D(net2555),
    .Q_N(_06986_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 _14806_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net931),
    .D(net2451),
    .Q_N(_06987_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 _14807_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net932),
    .D(net2532),
    .Q_N(_06988_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 _14808_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net933),
    .D(net2676),
    .Q_N(_06989_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 _14809_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net934),
    .D(net2524),
    .Q_N(_06990_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 _14810_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net935),
    .D(net2450),
    .Q_N(_06991_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 _14811_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net936),
    .D(net2435),
    .Q_N(_06992_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 _14812_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net937),
    .D(net2657),
    .Q_N(_06993_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 _14813_ (.CLK(clknet_leaf_127_clk_regs),
    .RESET_B(net938),
    .D(net2739),
    .Q_N(_06994_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 _14814_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net939),
    .D(_00114_),
    .Q_N(_06995_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 _14815_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net940),
    .D(_00115_),
    .Q_N(_06996_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 _14816_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net941),
    .D(_00116_),
    .Q_N(_06997_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 _14817_ (.CLK(clknet_leaf_127_clk_regs),
    .RESET_B(net942),
    .D(_00117_),
    .Q_N(_06998_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 _14818_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net943),
    .D(net2681),
    .Q_N(_06999_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ));
 sg13g2_dfrbp_1 _14819_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net944),
    .D(net2702),
    .Q_N(_07000_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ));
 sg13g2_dfrbp_1 _14820_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net945),
    .D(net2766),
    .Q_N(_07001_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ));
 sg13g2_dfrbp_1 _14821_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net946),
    .D(net2623),
    .Q_N(_07002_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ));
 sg13g2_dfrbp_1 _14822_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net947),
    .D(net2430),
    .Q_N(_07003_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 _14823_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net948),
    .D(net2593),
    .Q_N(_07004_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 _14824_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net949),
    .D(net2800),
    .Q_N(_07005_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 _14825_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net950),
    .D(net2483),
    .Q_N(_07006_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 _14826_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net951),
    .D(net2575),
    .Q_N(_07007_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 _14827_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net952),
    .D(net2631),
    .Q_N(_07008_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 _14828_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net953),
    .D(net2683),
    .Q_N(_07009_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 _14829_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net954),
    .D(net2579),
    .Q_N(_07010_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 _14830_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net955),
    .D(net2636),
    .Q_N(_07011_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 _14831_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net956),
    .D(net2726),
    .Q_N(_07012_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 _14832_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net957),
    .D(net2501),
    .Q_N(_07013_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 _14833_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net958),
    .D(net2655),
    .Q_N(_07014_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 _14834_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net959),
    .D(net2756),
    .Q_N(_07015_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 _14835_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net960),
    .D(net2773),
    .Q_N(_07016_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 _14836_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net961),
    .D(net2610),
    .Q_N(_07017_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 _14837_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net962),
    .D(net2479),
    .Q_N(_07018_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 _14838_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net963),
    .D(net2562),
    .Q_N(_07019_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 _14839_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net964),
    .D(net2539),
    .Q_N(_07020_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 _14840_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net965),
    .D(net2536),
    .Q_N(_07021_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 _14841_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net966),
    .D(net2791),
    .Q_N(_07022_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 _14842_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net967),
    .D(net2661),
    .Q_N(_07023_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 _14843_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net968),
    .D(net2488),
    .Q_N(_07024_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 _14844_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net969),
    .D(net2603),
    .Q_N(_07025_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 _14845_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net970),
    .D(net2568),
    .Q_N(_07026_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 _14846_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net971),
    .D(_00110_),
    .Q_N(_07027_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 _14847_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net972),
    .D(_00111_),
    .Q_N(_07028_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 _14848_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net973),
    .D(_00112_),
    .Q_N(_07029_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 _14849_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net974),
    .D(_00113_),
    .Q_N(_07030_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 _14850_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net975),
    .D(net2761),
    .Q_N(_07031_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ));
 sg13g2_dfrbp_1 _14851_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net976),
    .D(net2747),
    .Q_N(_07032_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ));
 sg13g2_dfrbp_1 _14852_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net977),
    .D(net2737),
    .Q_N(_07033_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ));
 sg13g2_dfrbp_1 _14853_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net978),
    .D(net2682),
    .Q_N(_07034_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ));
 sg13g2_dfrbp_1 _14854_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net979),
    .D(net2418),
    .Q_N(_07035_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 _14855_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net980),
    .D(net2554),
    .Q_N(_07036_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 _14856_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net981),
    .D(net2392),
    .Q_N(_07037_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 _14857_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net982),
    .D(net2512),
    .Q_N(_07038_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 _14858_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net983),
    .D(net2768),
    .Q_N(_07039_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 _14859_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net984),
    .D(net2461),
    .Q_N(_07040_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 _14860_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net985),
    .D(net2613),
    .Q_N(_07041_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 _14861_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net986),
    .D(net2390),
    .Q_N(_07042_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 _14862_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net987),
    .D(net2509),
    .Q_N(_07043_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 _14863_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net988),
    .D(net2465),
    .Q_N(_07044_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 _14864_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net989),
    .D(net2440),
    .Q_N(_07045_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 _14865_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net990),
    .D(net2727),
    .Q_N(_07046_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 _14866_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net991),
    .D(net2498),
    .Q_N(_07047_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 _14867_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net992),
    .D(net2559),
    .Q_N(_07048_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 _14868_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net993),
    .D(net2566),
    .Q_N(_07049_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 _14869_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net994),
    .D(net2514),
    .Q_N(_07050_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 _14870_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net995),
    .D(net2666),
    .Q_N(_07051_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 _14871_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net996),
    .D(net2781),
    .Q_N(_07052_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 _14872_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net997),
    .D(net2805),
    .Q_N(_07053_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 _14873_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net998),
    .D(net2441),
    .Q_N(_07054_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 _14874_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net999),
    .D(net2758),
    .Q_N(_07055_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 _14875_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net1000),
    .D(net2448),
    .Q_N(_07056_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 _14876_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net1001),
    .D(net2494),
    .Q_N(_07057_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 _14877_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net1002),
    .D(net2728),
    .Q_N(_07058_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 _14878_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net1003),
    .D(_00106_),
    .Q_N(_07059_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 _14879_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net1004),
    .D(_00107_),
    .Q_N(_07060_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 _14880_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net1005),
    .D(_00108_),
    .Q_N(_07061_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 _14881_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net1006),
    .D(_00109_),
    .Q_N(_07062_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 _14882_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net1007),
    .D(net2687),
    .Q_N(_07063_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ));
 sg13g2_dfrbp_1 _14883_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net1008),
    .D(net2595),
    .Q_N(_07064_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ));
 sg13g2_dfrbp_1 _14884_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net1009),
    .D(net2432),
    .Q_N(_07065_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ));
 sg13g2_dfrbp_1 _14885_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net1010),
    .D(net2725),
    .Q_N(_07066_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ));
 sg13g2_dfrbp_1 _14886_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net1011),
    .D(net2499),
    .Q_N(_07067_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 _14887_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net1012),
    .D(net2519),
    .Q_N(_07068_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 _14888_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net1013),
    .D(net2563),
    .Q_N(_07069_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 _14889_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net1014),
    .D(net2552),
    .Q_N(_07070_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 _14890_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net1015),
    .D(net2759),
    .Q_N(_07071_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 _14891_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net1016),
    .D(net2646),
    .Q_N(_07072_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 _14892_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net1017),
    .D(net2664),
    .Q_N(_07073_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 _14893_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net1018),
    .D(net2719),
    .Q_N(_07074_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 _14894_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net1019),
    .D(net2463),
    .Q_N(_07075_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 _14895_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net1020),
    .D(net2736),
    .Q_N(_07076_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 _14896_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net1021),
    .D(net2528),
    .Q_N(_07077_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 _14897_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net1022),
    .D(net2643),
    .Q_N(_07078_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 _14898_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net1023),
    .D(net2452),
    .Q_N(_07079_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 _14899_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net1024),
    .D(net2424),
    .Q_N(_07080_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 _14900_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net1025),
    .D(net2457),
    .Q_N(_07081_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 _14901_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net1026),
    .D(net2416),
    .Q_N(_07082_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 _14902_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net1027),
    .D(net2454),
    .Q_N(_07083_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 _14903_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net1028),
    .D(net2453),
    .Q_N(_07084_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 _14904_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net1029),
    .D(net2742),
    .Q_N(_07085_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 _14905_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net1030),
    .D(net2455),
    .Q_N(_07086_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 _14906_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net1031),
    .D(net2776),
    .Q_N(_07087_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 _14907_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net1032),
    .D(net2680),
    .Q_N(_07088_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 _14908_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net1033),
    .D(net2746),
    .Q_N(_07089_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 _14909_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net1034),
    .D(net2778),
    .Q_N(_07090_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 _14910_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net1035),
    .D(_00102_),
    .Q_N(_07091_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 _14911_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net1036),
    .D(_00103_),
    .Q_N(_07092_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 _14912_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net1037),
    .D(_00104_),
    .Q_N(_07093_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 _14913_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net1038),
    .D(_00105_),
    .Q_N(_07094_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 _14914_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net1039),
    .D(net2654),
    .Q_N(_07095_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ));
 sg13g2_dfrbp_1 _14915_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net1040),
    .D(net2721),
    .Q_N(_07096_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ));
 sg13g2_dfrbp_1 _14916_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net1041),
    .D(net2741),
    .Q_N(_07097_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ));
 sg13g2_dfrbp_1 _14917_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net1042),
    .D(net2442),
    .Q_N(_07098_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ));
 sg13g2_dfrbp_1 _14918_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net1043),
    .D(net2602),
    .Q_N(_07099_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 _14919_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net1044),
    .D(net2753),
    .Q_N(_07100_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 _14920_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net1045),
    .D(net2630),
    .Q_N(_07101_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 _14921_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1046),
    .D(net2622),
    .Q_N(_07102_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 _14922_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net1047),
    .D(net2402),
    .Q_N(_07103_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 _14923_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net1048),
    .D(net2419),
    .Q_N(_07104_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 _14924_ (.CLK(clknet_leaf_113_clk_regs),
    .RESET_B(net1049),
    .D(net2515),
    .Q_N(_07105_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 _14925_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1050),
    .D(net2444),
    .Q_N(_07106_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 _14926_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net1051),
    .D(net2706),
    .Q_N(_07107_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 _14927_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1052),
    .D(net2447),
    .Q_N(_07108_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 _14928_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net1053),
    .D(net2410),
    .Q_N(_07109_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 _14929_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1054),
    .D(net2537),
    .Q_N(_07110_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 _14930_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net1055),
    .D(net2649),
    .Q_N(_07111_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 _14931_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1056),
    .D(net2586),
    .Q_N(_07112_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 _14932_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net1057),
    .D(net2550),
    .Q_N(_07113_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 _14933_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net1058),
    .D(net2585),
    .Q_N(_07114_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 _14934_ (.CLK(clknet_leaf_118_clk_regs),
    .RESET_B(net1059),
    .D(net2795),
    .Q_N(_07115_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 _14935_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1060),
    .D(net2659),
    .Q_N(_07116_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 _14936_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net1061),
    .D(net2531),
    .Q_N(_07117_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 _14937_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net1062),
    .D(net2637),
    .Q_N(_07118_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 _14938_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net1063),
    .D(net2464),
    .Q_N(_07119_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 _14939_ (.CLK(clknet_leaf_114_clk_regs),
    .RESET_B(net1064),
    .D(net2400),
    .Q_N(_07120_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 _14940_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net1065),
    .D(net2413),
    .Q_N(_07121_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 _14941_ (.CLK(clknet_leaf_115_clk_regs),
    .RESET_B(net1066),
    .D(net2414),
    .Q_N(_07122_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 _14942_ (.CLK(clknet_leaf_120_clk_regs),
    .RESET_B(net1067),
    .D(_00098_),
    .Q_N(_07123_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 _14943_ (.CLK(clknet_leaf_117_clk_regs),
    .RESET_B(net1068),
    .D(_00099_),
    .Q_N(_07124_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 _14944_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net1069),
    .D(_00100_),
    .Q_N(_07125_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 _14945_ (.CLK(clknet_leaf_116_clk_regs),
    .RESET_B(net1070),
    .D(_00101_),
    .Q_N(_07126_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 _14946_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net1071),
    .D(net2770),
    .Q_N(_07127_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ));
 sg13g2_dfrbp_1 _14947_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net1072),
    .D(net2743),
    .Q_N(_07128_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ));
 sg13g2_dfrbp_1 _14948_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net1073),
    .D(net2769),
    .Q_N(_07129_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ));
 sg13g2_dfrbp_1 _14949_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net1074),
    .D(net2709),
    .Q_N(_07130_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ));
 sg13g2_dfrbp_1 _14950_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net1075),
    .D(net2517),
    .Q_N(_07131_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 _14951_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net1076),
    .D(net2685),
    .Q_N(_07132_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 _14952_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net1077),
    .D(net2505),
    .Q_N(_07133_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 _14953_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net1078),
    .D(net2644),
    .Q_N(_07134_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 _14954_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net1079),
    .D(net2694),
    .Q_N(_07135_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 _14955_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net1080),
    .D(net2506),
    .Q_N(_07136_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 _14956_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net1081),
    .D(net2456),
    .Q_N(_07137_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 _14957_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net1082),
    .D(net2580),
    .Q_N(_07138_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 _14958_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net1083),
    .D(net2783),
    .Q_N(_07139_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 _14959_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net1084),
    .D(net2417),
    .Q_N(_07140_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 _14960_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net1085),
    .D(net2420),
    .Q_N(_07141_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 _14961_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net1086),
    .D(net2391),
    .Q_N(_07142_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 _14962_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net1087),
    .D(net2590),
    .Q_N(_07143_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 _14963_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net1088),
    .D(net2436),
    .Q_N(_07144_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 _14964_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net1089),
    .D(net2752),
    .Q_N(_07145_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 _14965_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net1090),
    .D(net2802),
    .Q_N(_07146_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 _14966_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net1091),
    .D(net2614),
    .Q_N(_07147_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 _14967_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net1092),
    .D(net2525),
    .Q_N(_07148_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 _14968_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net1093),
    .D(net2714),
    .Q_N(_07149_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 _14969_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net1094),
    .D(net2490),
    .Q_N(_07150_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 _14970_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net1095),
    .D(net2470),
    .Q_N(_07151_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 _14971_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net1096),
    .D(net2533),
    .Q_N(_07152_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 _14972_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net1097),
    .D(net2684),
    .Q_N(_07153_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 _14973_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net1098),
    .D(net2584),
    .Q_N(_07154_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 _14974_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net1099),
    .D(_00094_),
    .Q_N(_07155_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 _14975_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net1100),
    .D(_00095_),
    .Q_N(_07156_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 _14976_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net1101),
    .D(_00096_),
    .Q_N(_07157_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 _14977_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net1102),
    .D(_00097_),
    .Q_N(_07158_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 _14978_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net1103),
    .D(net2811),
    .Q_N(_07159_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ));
 sg13g2_dfrbp_1 _14979_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net1104),
    .D(net2841),
    .Q_N(_07160_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ));
 sg13g2_dfrbp_1 _14980_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net1105),
    .D(net2842),
    .Q_N(_07161_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ));
 sg13g2_dfrbp_1 _14981_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1106),
    .D(net2826),
    .Q_N(_07162_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ));
 sg13g2_dfrbp_1 _14982_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1107),
    .D(net2830),
    .Q_N(_07163_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ));
 sg13g2_dfrbp_1 _14983_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net1108),
    .D(net2798),
    .Q_N(_07164_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ));
 sg13g2_dfrbp_1 _14984_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net1109),
    .D(net2827),
    .Q_N(_07165_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ));
 sg13g2_dfrbp_1 _14985_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net1110),
    .D(net2809),
    .Q_N(_07166_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ));
 sg13g2_dfrbp_1 _14986_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net1111),
    .D(net2817),
    .Q_N(_07167_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ));
 sg13g2_dfrbp_1 _14987_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net1112),
    .D(net2793),
    .Q_N(_07168_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ));
 sg13g2_dfrbp_1 _14988_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net1113),
    .D(net2806),
    .Q_N(_07169_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ));
 sg13g2_dfrbp_1 _14989_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net1114),
    .D(net2797),
    .Q_N(_07170_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ));
 sg13g2_dfrbp_1 _14990_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net1115),
    .D(net2799),
    .Q_N(_07171_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ));
 sg13g2_dfrbp_1 _14991_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net1116),
    .D(net2821),
    .Q_N(_07172_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ));
 sg13g2_dfrbp_1 _14992_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net1117),
    .D(net2812),
    .Q_N(_07173_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ));
 sg13g2_dfrbp_1 _14993_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net1118),
    .D(net2824),
    .Q_N(_07174_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ));
 sg13g2_dfrbp_1 _14994_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net1119),
    .D(net2816),
    .Q_N(_07175_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ));
 sg13g2_dfrbp_1 _14995_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net1120),
    .D(net2818),
    .Q_N(_07176_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ));
 sg13g2_dfrbp_1 _14996_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net1121),
    .D(net2808),
    .Q_N(_07177_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ));
 sg13g2_dfrbp_1 _14997_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net1122),
    .D(net2810),
    .Q_N(_07178_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ));
 sg13g2_dfrbp_1 _14998_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net1123),
    .D(net2839),
    .Q_N(_07179_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ));
 sg13g2_dfrbp_1 _14999_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net1124),
    .D(net2836),
    .Q_N(_07180_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ));
 sg13g2_dfrbp_1 _15000_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net1125),
    .D(net2840),
    .Q_N(_07181_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ));
 sg13g2_dfrbp_1 _15001_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net1126),
    .D(net2835),
    .Q_N(_07182_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ));
 sg13g2_dfrbp_1 _15002_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net1127),
    .D(net2673),
    .Q_N(_07183_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ));
 sg13g2_dfrbp_1 _15003_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net1128),
    .D(net2581),
    .Q_N(_07184_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_dfrbp_1 _15004_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net1129),
    .D(net2796),
    .Q_N(_07185_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ));
 sg13g2_dfrbp_1 _15005_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net1130),
    .D(net2774),
    .Q_N(_07186_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_dfrbp_1 _15006_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net1138),
    .D(\i_tinyqv.cpu.i_core.cy_out ),
    .Q_N(_00128_),
    .Q(\i_tinyqv.cpu.i_core.cy ));
 sg13g2_dfrbp_1 _15007_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net1555),
    .D(\i_tinyqv.cpu.i_core.cmp_out ),
    .Q_N(_06711_),
    .Q(\i_tinyqv.cpu.i_core.cmp ));
 sg13g2_dfrbp_1 _15008_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net1554),
    .D(net3293),
    .Q_N(_06710_),
    .Q(\i_tinyqv.cpu.i_core.load_done ));
 sg13g2_dfrbp_1 _15009_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net1553),
    .D(net3769),
    .Q_N(_00122_),
    .Q(\i_tinyqv.cpu.i_core.cycle[0] ));
 sg13g2_dfrbp_1 _15010_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net1551),
    .D(_00605_),
    .Q_N(_06709_),
    .Q(\i_tinyqv.cpu.i_core.cycle[1] ));
 sg13g2_dfrbp_1 _15011_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net1549),
    .D(net3396),
    .Q_N(_06708_),
    .Q(\i_tinyqv.cpu.i_core.is_double_fault_r ));
 sg13g2_dfrbp_1 _15012_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net1548),
    .D(net2832),
    .Q_N(_00271_),
    .Q(\i_tinyqv.cpu.i_core.time_hi[0] ));
 sg13g2_dfrbp_1 _15013_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net1546),
    .D(net3212),
    .Q_N(_06707_),
    .Q(\i_tinyqv.cpu.i_core.time_hi[1] ));
 sg13g2_dfrbp_1 _15014_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net1158),
    .D(net3424),
    .Q_N(_07187_),
    .Q(\i_tinyqv.cpu.i_core.time_hi[2] ));
 sg13g2_dfrbp_1 _15015_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net1544),
    .D(_00065_),
    .Q_N(_00264_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.add ));
 sg13g2_dfrbp_1 _15016_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net1542),
    .D(_00610_),
    .Q_N(_06706_),
    .Q(\i_tinyqv.cpu.i_core.mcause[0] ));
 sg13g2_dfrbp_1 _15017_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net1540),
    .D(net3600),
    .Q_N(_06705_),
    .Q(\i_tinyqv.cpu.i_core.mcause[1] ));
 sg13g2_dfrbp_1 _15018_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net1538),
    .D(_00612_),
    .Q_N(_06704_),
    .Q(\i_tinyqv.cpu.i_core.mcause[2] ));
 sg13g2_dfrbp_1 _15019_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net1536),
    .D(_00613_),
    .Q_N(_06703_),
    .Q(\i_tinyqv.cpu.i_core.mcause[3] ));
 sg13g2_dfrbp_1 _15020_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net1534),
    .D(_00614_),
    .Q_N(_06702_),
    .Q(\i_tinyqv.cpu.i_core.mcause[4] ));
 sg13g2_dfrbp_1 _15021_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net1532),
    .D(_00615_),
    .Q_N(_06701_),
    .Q(\i_tinyqv.cpu.i_core.mcause[5] ));
 sg13g2_dfrbp_1 _15022_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net1530),
    .D(net3302),
    .Q_N(_06700_),
    .Q(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ));
 sg13g2_dfrbp_1 _15023_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net1529),
    .D(net3276),
    .Q_N(_06699_),
    .Q(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ));
 sg13g2_dfrbp_1 _15024_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net1528),
    .D(_00618_),
    .Q_N(_06698_),
    .Q(\i_tinyqv.cpu.i_core.mepc[20] ));
 sg13g2_dfrbp_1 _15025_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net1526),
    .D(_00619_),
    .Q_N(_06697_),
    .Q(\i_tinyqv.cpu.i_core.mepc[21] ));
 sg13g2_dfrbp_1 _15026_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net1524),
    .D(_00620_),
    .Q_N(_06696_),
    .Q(\i_tinyqv.cpu.i_core.mepc[22] ));
 sg13g2_dfrbp_1 _15027_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net1522),
    .D(_00621_),
    .Q_N(_06695_),
    .Q(\i_tinyqv.cpu.i_core.mepc[23] ));
 sg13g2_dfrbp_1 _15028_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net1520),
    .D(_00622_),
    .Q_N(_06694_),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mte ));
 sg13g2_dfrbp_1 _15029_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net1518),
    .D(_00623_),
    .Q_N(_06693_),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mie ));
 sg13g2_dfrbp_1 _15030_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net1516),
    .D(net3526),
    .Q_N(_06692_),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mpie ));
 sg13g2_dfrbp_1 _15031_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net1514),
    .D(net3036),
    .Q_N(_00255_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[0] ));
 sg13g2_dfrbp_1 _15032_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net1513),
    .D(_00626_),
    .Q_N(_06691_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[1] ));
 sg13g2_dfrbp_1 _15033_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net1512),
    .D(_00627_),
    .Q_N(_06690_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[2] ));
 sg13g2_dfrbp_1 _15034_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net1159),
    .D(_00628_),
    .Q_N(_07188_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[3] ));
 sg13g2_dfrbp_1 _15035_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net1160),
    .D(_00090_),
    .Q_N(_07189_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ));
 sg13g2_dfrbp_1 _15036_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net1161),
    .D(_00091_),
    .Q_N(_07190_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ));
 sg13g2_dfrbp_1 _15037_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net1162),
    .D(_00092_),
    .Q_N(_07191_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ));
 sg13g2_dfrbp_1 _15038_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net1263),
    .D(_00093_),
    .Q_N(_07192_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ));
 sg13g2_dfrbp_1 _15039_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net1511),
    .D(net534),
    .Q_N(_00194_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.rstn ));
 sg13g2_dfrbp_1 _15040_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1510),
    .D(_00629_),
    .Q_N(_06689_),
    .Q(\i_uart_tx.data_to_send[0] ));
 sg13g2_dfrbp_1 _15041_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1508),
    .D(net3528),
    .Q_N(_06688_),
    .Q(\i_uart_tx.data_to_send[1] ));
 sg13g2_dfrbp_1 _15042_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net1506),
    .D(net3495),
    .Q_N(_06687_),
    .Q(\i_uart_tx.data_to_send[2] ));
 sg13g2_dfrbp_1 _15043_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1504),
    .D(_00632_),
    .Q_N(_06686_),
    .Q(\i_uart_tx.data_to_send[3] ));
 sg13g2_dfrbp_1 _15044_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net1502),
    .D(net3430),
    .Q_N(_06685_),
    .Q(\i_uart_tx.data_to_send[4] ));
 sg13g2_dfrbp_1 _15045_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net1500),
    .D(_00634_),
    .Q_N(_06684_),
    .Q(\i_uart_tx.data_to_send[5] ));
 sg13g2_dfrbp_1 _15046_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1498),
    .D(net3454),
    .Q_N(_06683_),
    .Q(\i_uart_tx.data_to_send[6] ));
 sg13g2_dfrbp_1 _15047_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1496),
    .D(net2999),
    .Q_N(_06682_),
    .Q(\i_uart_tx.data_to_send[7] ));
 sg13g2_dfrbp_1 _15048_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net1494),
    .D(net2834),
    .Q_N(_00270_),
    .Q(\i_uart_tx.cycle_counter[0] ));
 sg13g2_dfrbp_1 _15049_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1492),
    .D(net3140),
    .Q_N(_06681_),
    .Q(\i_uart_tx.cycle_counter[1] ));
 sg13g2_dfrbp_1 _15050_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1490),
    .D(_00639_),
    .Q_N(_06680_),
    .Q(\i_uart_tx.cycle_counter[2] ));
 sg13g2_dfrbp_1 _15051_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net1488),
    .D(_00640_),
    .Q_N(_06679_),
    .Q(\i_uart_tx.cycle_counter[3] ));
 sg13g2_dfrbp_1 _15052_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net1486),
    .D(_00641_),
    .Q_N(_06678_),
    .Q(\i_uart_tx.cycle_counter[4] ));
 sg13g2_dfrbp_1 _15053_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net1484),
    .D(_00642_),
    .Q_N(_06677_),
    .Q(\i_uart_tx.cycle_counter[5] ));
 sg13g2_dfrbp_1 _15054_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net1482),
    .D(_00643_),
    .Q_N(_06676_),
    .Q(\i_uart_tx.cycle_counter[6] ));
 sg13g2_dfrbp_1 _15055_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net1480),
    .D(net3518),
    .Q_N(_06675_),
    .Q(\i_uart_tx.cycle_counter[7] ));
 sg13g2_dfrbp_1 _15056_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1478),
    .D(_00645_),
    .Q_N(_06674_),
    .Q(\i_uart_tx.cycle_counter[8] ));
 sg13g2_dfrbp_1 _15057_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net1476),
    .D(_00646_),
    .Q_N(_06673_),
    .Q(\i_uart_tx.cycle_counter[9] ));
 sg13g2_dfrbp_1 _15058_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net1474),
    .D(_00647_),
    .Q_N(_06672_),
    .Q(\i_uart_tx.cycle_counter[10] ));
 sg13g2_dfrbp_1 _15059_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1472),
    .D(_00648_),
    .Q_N(_06671_),
    .Q(\i_uart_tx.fsm_state[0] ));
 sg13g2_dfrbp_1 _15060_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net1470),
    .D(_00649_),
    .Q_N(_06670_),
    .Q(\i_uart_tx.fsm_state[1] ));
 sg13g2_dfrbp_1 _15061_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1468),
    .D(_00650_),
    .Q_N(_06669_),
    .Q(\i_uart_tx.fsm_state[2] ));
 sg13g2_dfrbp_1 _15062_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1466),
    .D(_00651_),
    .Q_N(_06668_),
    .Q(\i_uart_tx.fsm_state[3] ));
 sg13g2_dfrbp_1 _15063_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1464),
    .D(net3421),
    .Q_N(_06667_),
    .Q(\i_uart_rx.recieved_data[0] ));
 sg13g2_dfrbp_1 _15064_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net1463),
    .D(_00653_),
    .Q_N(_06666_),
    .Q(\i_uart_rx.recieved_data[1] ));
 sg13g2_dfrbp_1 _15065_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net1462),
    .D(_00654_),
    .Q_N(_06665_),
    .Q(\i_uart_rx.recieved_data[2] ));
 sg13g2_dfrbp_1 _15066_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net1461),
    .D(net3512),
    .Q_N(_06664_),
    .Q(\i_uart_rx.recieved_data[3] ));
 sg13g2_dfrbp_1 _15067_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net1460),
    .D(net3487),
    .Q_N(_06663_),
    .Q(\i_uart_rx.recieved_data[4] ));
 sg13g2_dfrbp_1 _15068_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net1459),
    .D(_00657_),
    .Q_N(_06662_),
    .Q(\i_uart_rx.recieved_data[5] ));
 sg13g2_dfrbp_1 _15069_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net1458),
    .D(_00658_),
    .Q_N(_06661_),
    .Q(\i_uart_rx.recieved_data[6] ));
 sg13g2_dfrbp_1 _15070_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net1457),
    .D(net3339),
    .Q_N(_06660_),
    .Q(\i_uart_rx.recieved_data[7] ));
 sg13g2_dfrbp_1 _15071_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net1456),
    .D(_00660_),
    .Q_N(_06659_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[0] ));
 sg13g2_dfrbp_1 _15072_ (.CLK(clknet_leaf_139_clk_regs),
    .RESET_B(net1454),
    .D(net3389),
    .Q_N(_06658_),
    .Q(\i_tinyqv.cpu.i_core.load_top_bit ));
 sg13g2_dfrbp_1 _15073_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1452),
    .D(_00662_),
    .Q_N(_00269_),
    .Q(\i_uart_rx.cycle_counter[0] ));
 sg13g2_dfrbp_1 _15074_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1451),
    .D(net3337),
    .Q_N(_06657_),
    .Q(\i_uart_rx.cycle_counter[1] ));
 sg13g2_dfrbp_1 _15075_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net1450),
    .D(_00664_),
    .Q_N(_06656_),
    .Q(\i_uart_rx.cycle_counter[2] ));
 sg13g2_dfrbp_1 _15076_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1449),
    .D(_00665_),
    .Q_N(_06655_),
    .Q(\i_uart_rx.cycle_counter[3] ));
 sg13g2_dfrbp_1 _15077_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1448),
    .D(_00666_),
    .Q_N(_06654_),
    .Q(\i_uart_rx.cycle_counter[4] ));
 sg13g2_dfrbp_1 _15078_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1447),
    .D(_00667_),
    .Q_N(_06653_),
    .Q(\i_uart_rx.cycle_counter[5] ));
 sg13g2_dfrbp_1 _15079_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1446),
    .D(_00668_),
    .Q_N(_06652_),
    .Q(\i_uart_rx.cycle_counter[6] ));
 sg13g2_dfrbp_1 _15080_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1445),
    .D(_00669_),
    .Q_N(_06651_),
    .Q(\i_uart_rx.cycle_counter[7] ));
 sg13g2_dfrbp_1 _15081_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1444),
    .D(_00670_),
    .Q_N(_06650_),
    .Q(\i_uart_rx.cycle_counter[8] ));
 sg13g2_dfrbp_1 _15082_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1443),
    .D(_00671_),
    .Q_N(_06649_),
    .Q(\i_uart_rx.cycle_counter[9] ));
 sg13g2_dfrbp_1 _15083_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1442),
    .D(_00672_),
    .Q_N(_06648_),
    .Q(\i_uart_rx.cycle_counter[10] ));
 sg13g2_dfrbp_1 _15084_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1441),
    .D(net3318),
    .Q_N(_06647_),
    .Q(\i_uart_rx.bit_sample ));
 sg13g2_dfrbp_1 _15085_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net1439),
    .D(_00674_),
    .Q_N(_06646_),
    .Q(\i_uart_rx.uart_rts ));
 sg13g2_dfrbp_1 _15086_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1438),
    .D(net3753),
    .Q_N(_00243_),
    .Q(\i_uart_rx.fsm_state[0] ));
 sg13g2_dfrbp_1 _15087_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1436),
    .D(_00676_),
    .Q_N(_06645_),
    .Q(\i_uart_rx.fsm_state[1] ));
 sg13g2_dfrbp_1 _15088_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1434),
    .D(net3643),
    .Q_N(_06644_),
    .Q(\i_uart_rx.fsm_state[2] ));
 sg13g2_dfrbp_1 _15089_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1432),
    .D(net3904),
    .Q_N(_06643_),
    .Q(\i_uart_rx.fsm_state[3] ));
 sg13g2_dfrbp_1 _15090_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net1430),
    .D(_00679_),
    .Q_N(_00244_),
    .Q(\i_uart_rx.rxd_reg[0] ));
 sg13g2_dfrbp_1 _15091_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1429),
    .D(_00680_),
    .Q_N(_06642_),
    .Q(\i_uart_rx.rxd_reg[1] ));
 sg13g2_dfrbp_1 _15092_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net1428),
    .D(net2838),
    .Q_N(_06641_),
    .Q(\i_tinyqv.mem.q_ctrl.stop_txn_reg ));
 sg13g2_dfrbp_1 _15093_ (.CLK(clknet_leaf_140_clk_regs),
    .RESET_B(net1427),
    .D(net3387),
    .Q_N(_06640_),
    .Q(\i_tinyqv.cpu.instr_data[3][0] ));
 sg13g2_dfrbp_1 _15094_ (.CLK(clknet_leaf_141_clk_regs),
    .RESET_B(net1426),
    .D(net3200),
    .Q_N(_00140_),
    .Q(\i_tinyqv.cpu.instr_data[3][1] ));
 sg13g2_dfrbp_1 _15095_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net1425),
    .D(net3559),
    .Q_N(_06639_),
    .Q(\i_tinyqv.cpu.instr_data[2][2] ));
 sg13g2_dfrbp_1 _15096_ (.CLK(clknet_leaf_132_clk_regs),
    .RESET_B(net1424),
    .D(net3476),
    .Q_N(_06638_),
    .Q(\i_tinyqv.cpu.instr_data[2][3] ));
 sg13g2_dfrbp_1 _15097_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net1423),
    .D(net3219),
    .Q_N(_00145_),
    .Q(\i_tinyqv.cpu.instr_data[2][4] ));
 sg13g2_dfrbp_1 _15098_ (.CLK(clknet_leaf_149_clk_regs),
    .RESET_B(net1422),
    .D(net3090),
    .Q_N(_00149_),
    .Q(\i_tinyqv.cpu.instr_data[2][5] ));
 sg13g2_dfrbp_1 _15099_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net1421),
    .D(net3063),
    .Q_N(_00153_),
    .Q(\i_tinyqv.cpu.instr_data[2][6] ));
 sg13g2_dfrbp_1 _15100_ (.CLK(clknet_leaf_149_clk_regs),
    .RESET_B(net1420),
    .D(net3074),
    .Q_N(_00170_),
    .Q(\i_tinyqv.cpu.instr_data[2][7] ));
 sg13g2_dfrbp_1 _15101_ (.CLK(clknet_leaf_148_clk_regs),
    .RESET_B(net1419),
    .D(net3107),
    .Q_N(_00174_),
    .Q(\i_tinyqv.cpu.instr_data[2][8] ));
 sg13g2_dfrbp_1 _15102_ (.CLK(clknet_leaf_148_clk_regs),
    .RESET_B(net1418),
    .D(net3039),
    .Q_N(_00178_),
    .Q(\i_tinyqv.cpu.instr_data[2][9] ));
 sg13g2_dfrbp_1 _15103_ (.CLK(clknet_leaf_151_clk_regs),
    .RESET_B(net1417),
    .D(net3026),
    .Q_N(_00182_),
    .Q(\i_tinyqv.cpu.instr_data[2][10] ));
 sg13g2_dfrbp_1 _15104_ (.CLK(clknet_leaf_147_clk_regs),
    .RESET_B(net1416),
    .D(net3044),
    .Q_N(_00190_),
    .Q(\i_tinyqv.cpu.instr_data[2][11] ));
 sg13g2_dfrbp_1 _15105_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net1415),
    .D(net3181),
    .Q_N(_00186_),
    .Q(\i_tinyqv.cpu.instr_data[2][12] ));
 sg13g2_dfrbp_1 _15106_ (.CLK(clknet_leaf_145_clk_regs),
    .RESET_B(net1414),
    .D(net3032),
    .Q_N(_00157_),
    .Q(\i_tinyqv.cpu.instr_data[2][13] ));
 sg13g2_dfrbp_1 _15107_ (.CLK(clknet_leaf_151_clk_regs),
    .RESET_B(net1413),
    .D(net3024),
    .Q_N(_00161_),
    .Q(\i_tinyqv.cpu.instr_data[2][14] ));
 sg13g2_dfrbp_1 _15108_ (.CLK(clknet_leaf_150_clk_regs),
    .RESET_B(net1412),
    .D(net3124),
    .Q_N(_00165_),
    .Q(\i_tinyqv.cpu.instr_data[2][15] ));
 sg13g2_dfrbp_1 _15109_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net1411),
    .D(_00698_),
    .Q_N(_06637_),
    .Q(\i_debug_uart_tx.data_to_send[0] ));
 sg13g2_dfrbp_1 _15110_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net1409),
    .D(_00699_),
    .Q_N(_06636_),
    .Q(\i_debug_uart_tx.data_to_send[1] ));
 sg13g2_dfrbp_1 _15111_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net1407),
    .D(_00700_),
    .Q_N(_06635_),
    .Q(\i_debug_uart_tx.data_to_send[2] ));
 sg13g2_dfrbp_1 _15112_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net1405),
    .D(_00701_),
    .Q_N(_06634_),
    .Q(\i_debug_uart_tx.data_to_send[3] ));
 sg13g2_dfrbp_1 _15113_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1403),
    .D(net3433),
    .Q_N(_06633_),
    .Q(\i_debug_uart_tx.data_to_send[4] ));
 sg13g2_dfrbp_1 _15114_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1401),
    .D(net3404),
    .Q_N(_06632_),
    .Q(\i_debug_uart_tx.data_to_send[5] ));
 sg13g2_dfrbp_1 _15115_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net1399),
    .D(net3460),
    .Q_N(_06631_),
    .Q(\i_debug_uart_tx.data_to_send[6] ));
 sg13g2_dfrbp_1 _15116_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net1397),
    .D(_00705_),
    .Q_N(_06630_),
    .Q(\i_debug_uart_tx.data_to_send[7] ));
 sg13g2_dfrbp_1 _15117_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net1395),
    .D(net2845),
    .Q_N(_00268_),
    .Q(\i_debug_uart_tx.cycle_counter[0] ));
 sg13g2_dfrbp_1 _15118_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net1393),
    .D(net3436),
    .Q_N(_06629_),
    .Q(\i_debug_uart_tx.cycle_counter[1] ));
 sg13g2_dfrbp_1 _15119_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net1391),
    .D(_00708_),
    .Q_N(_06628_),
    .Q(\i_debug_uart_tx.cycle_counter[2] ));
 sg13g2_dfrbp_1 _15120_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net1389),
    .D(_00709_),
    .Q_N(_06627_),
    .Q(\i_debug_uart_tx.cycle_counter[3] ));
 sg13g2_dfrbp_1 _15121_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net1387),
    .D(net2857),
    .Q_N(_06626_),
    .Q(\i_debug_uart_tx.cycle_counter[4] ));
 sg13g2_dfrbp_1 _15122_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net1385),
    .D(_00711_),
    .Q_N(_06625_),
    .Q(\i_debug_uart_tx.fsm_state[0] ));
 sg13g2_dfrbp_1 _15123_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net1383),
    .D(_00712_),
    .Q_N(_06624_),
    .Q(\i_debug_uart_tx.fsm_state[1] ));
 sg13g2_dfrbp_1 _15124_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net1381),
    .D(net3724),
    .Q_N(_06623_),
    .Q(\i_debug_uart_tx.fsm_state[2] ));
 sg13g2_dfrbp_1 _15125_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net1379),
    .D(_00714_),
    .Q_N(_06622_),
    .Q(\i_debug_uart_tx.fsm_state[3] ));
 sg13g2_dfrbp_1 _15126_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net1377),
    .D(_00715_),
    .Q_N(_06621_),
    .Q(\i_spi.end_txn_reg ));
 sg13g2_dfrbp_1 _15127_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net1376),
    .D(_00716_),
    .Q_N(_06620_),
    .Q(\i_spi.clock_count[0] ));
 sg13g2_dfrbp_1 _15128_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net1374),
    .D(net3383),
    .Q_N(_06619_),
    .Q(\i_spi.clock_count[1] ));
 sg13g2_dfrbp_1 _15129_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net1372),
    .D(_00718_),
    .Q_N(_06618_),
    .Q(\i_spi.clock_count[2] ));
 sg13g2_dfrbp_1 _15130_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net1370),
    .D(_00719_),
    .Q_N(_06617_),
    .Q(\i_spi.clock_count[3] ));
 sg13g2_dfrbp_1 _15131_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net1368),
    .D(_00720_),
    .Q_N(_06616_),
    .Q(\i_spi.data[0] ));
 sg13g2_dfrbp_1 _15132_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net1367),
    .D(net3462),
    .Q_N(_06615_),
    .Q(\i_spi.bits_remaining[0] ));
 sg13g2_dfrbp_1 _15133_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net1365),
    .D(net3868),
    .Q_N(_06614_),
    .Q(\i_spi.bits_remaining[1] ));
 sg13g2_dfrbp_1 _15134_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net1363),
    .D(net3705),
    .Q_N(_06613_),
    .Q(\i_spi.bits_remaining[2] ));
 sg13g2_dfrbp_1 _15135_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net1361),
    .D(_00724_),
    .Q_N(_06612_),
    .Q(\i_spi.bits_remaining[3] ));
 sg13g2_dfrbp_1 _15136_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net1359),
    .D(_00725_),
    .Q_N(_00204_),
    .Q(\i_spi.busy ));
 sg13g2_dfrbp_1 _15137_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net1358),
    .D(net3162),
    .Q_N(_06611_),
    .Q(\i_spi.spi_dc ));
 sg13g2_dfrbp_1 _15138_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net1357),
    .D(_00727_),
    .Q_N(_06610_),
    .Q(\i_spi.spi_select ));
 sg13g2_dfrbp_1 _15139_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net1355),
    .D(_00728_),
    .Q_N(_06609_),
    .Q(\i_spi.spi_clk_out ));
 sg13g2_dfrbp_1 _15140_ (.CLK(net2108),
    .RESET_B(net1353),
    .D(_00729_),
    .Q_N(_06608_),
    .Q(\i_pwm.l_pwm_level.data_out[0] ));
 sg13g2_dfrbp_1 _15141_ (.CLK(net2109),
    .RESET_B(net1351),
    .D(_00730_),
    .Q_N(_06607_),
    .Q(\i_pwm.l_pwm_level.data_out[1] ));
 sg13g2_dfrbp_1 _15142_ (.CLK(net2110),
    .RESET_B(net1349),
    .D(_00731_),
    .Q_N(_06606_),
    .Q(\i_pwm.l_pwm_level.data_out[2] ));
 sg13g2_dfrbp_1 _15143_ (.CLK(net2111),
    .RESET_B(net1347),
    .D(_00732_),
    .Q_N(_06605_),
    .Q(\i_pwm.l_pwm_level.data_out[3] ));
 sg13g2_dfrbp_1 _15144_ (.CLK(net2112),
    .RESET_B(net1345),
    .D(_00733_),
    .Q_N(_06604_),
    .Q(\i_pwm.l_pwm_level.data_out[4] ));
 sg13g2_dfrbp_1 _15145_ (.CLK(net2113),
    .RESET_B(net1343),
    .D(_00734_),
    .Q_N(_06603_),
    .Q(\i_pwm.l_pwm_level.data_out[5] ));
 sg13g2_dfrbp_1 _15146_ (.CLK(net2114),
    .RESET_B(net1341),
    .D(_00735_),
    .Q_N(_06602_),
    .Q(\i_pwm.l_pwm_level.data_out[6] ));
 sg13g2_dfrbp_1 _15147_ (.CLK(net2115),
    .RESET_B(net1339),
    .D(_00736_),
    .Q_N(_06601_),
    .Q(\i_pwm.l_pwm_level.data_out[7] ));
 sg13g2_dfrbp_1 _15148_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net1337),
    .D(_00737_),
    .Q_N(_00267_),
    .Q(\i_pwm.pwm_count[0] ));
 sg13g2_dfrbp_1 _15149_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net1336),
    .D(_00738_),
    .Q_N(_06600_),
    .Q(\i_pwm.pwm_count[1] ));
 sg13g2_dfrbp_1 _15150_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net1335),
    .D(net3586),
    .Q_N(_06599_),
    .Q(\i_pwm.pwm_count[2] ));
 sg13g2_dfrbp_1 _15151_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net1334),
    .D(_00740_),
    .Q_N(_06598_),
    .Q(\i_pwm.pwm_count[3] ));
 sg13g2_dfrbp_1 _15152_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net1333),
    .D(_00741_),
    .Q_N(_06597_),
    .Q(\i_pwm.pwm_count[4] ));
 sg13g2_dfrbp_1 _15153_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net1332),
    .D(_00742_),
    .Q_N(_06596_),
    .Q(\i_pwm.pwm_count[5] ));
 sg13g2_dfrbp_1 _15154_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net1331),
    .D(_00743_),
    .Q_N(_06595_),
    .Q(\i_pwm.pwm_count[6] ));
 sg13g2_dfrbp_1 _15155_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net1330),
    .D(_00744_),
    .Q_N(_06594_),
    .Q(\i_pwm.pwm_count[7] ));
 sg13g2_dfrbp_1 _15156_ (.CLK(net2116),
    .RESET_B(net1329),
    .D(_00745_),
    .Q_N(_06593_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15157_ (.CLK(net2117),
    .RESET_B(net1327),
    .D(_00746_),
    .Q_N(_06592_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15158_ (.CLK(net2118),
    .RESET_B(net1325),
    .D(_00747_),
    .Q_N(_06591_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15159_ (.CLK(net2119),
    .RESET_B(net1323),
    .D(_00748_),
    .Q_N(_06590_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15160_ (.CLK(net2120),
    .RESET_B(net1321),
    .D(_00749_),
    .Q_N(_06589_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15161_ (.CLK(net2121),
    .RESET_B(net1319),
    .D(_00750_),
    .Q_N(_06588_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15162_ (.CLK(net2122),
    .RESET_B(net1316),
    .D(_00751_),
    .Q_N(_06587_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15163_ (.CLK(net2123),
    .RESET_B(net1317),
    .D(_00752_),
    .Q_N(_07193_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15164_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net1314),
    .D(_00018_),
    .Q_N(_06586_),
    .Q(\i_pwm.pwm ));
 sg13g2_dfrbp_1 _15165_ (.CLK(clknet_leaf_152_clk_regs),
    .RESET_B(net1312),
    .D(net3696),
    .Q_N(_06585_),
    .Q(\i_time.l_mtimecmp.data_out[16] ));
 sg13g2_dfrbp_1 _15166_ (.CLK(clknet_leaf_152_clk_regs),
    .RESET_B(net1311),
    .D(net3661),
    .Q_N(_06584_),
    .Q(\i_time.l_mtimecmp.data_out[17] ));
 sg13g2_dfrbp_1 _15167_ (.CLK(clknet_leaf_152_clk_regs),
    .RESET_B(net1310),
    .D(net3648),
    .Q_N(_06583_),
    .Q(\i_time.l_mtimecmp.data_out[18] ));
 sg13g2_dfrbp_1 _15168_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net1309),
    .D(net3537),
    .Q_N(_06582_),
    .Q(\i_time.l_mtimecmp.data_out[19] ));
 sg13g2_dfrbp_1 _15169_ (.CLK(clknet_leaf_152_clk_regs),
    .RESET_B(net1308),
    .D(net3572),
    .Q_N(_06581_),
    .Q(\i_time.l_mtimecmp.data_out[20] ));
 sg13g2_dfrbp_1 _15170_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net1307),
    .D(net3758),
    .Q_N(_06580_),
    .Q(\i_time.l_mtimecmp.data_out[21] ));
 sg13g2_dfrbp_1 _15171_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net1306),
    .D(net3637),
    .Q_N(_06579_),
    .Q(\i_time.l_mtimecmp.data_out[22] ));
 sg13g2_dfrbp_1 _15172_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net1305),
    .D(net3631),
    .Q_N(_06578_),
    .Q(\i_time.l_mtimecmp.data_out[23] ));
 sg13g2_dfrbp_1 _15173_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net1304),
    .D(net3722),
    .Q_N(_06577_),
    .Q(\i_time.l_mtimecmp.data_out[24] ));
 sg13g2_dfrbp_1 _15174_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net1303),
    .D(net3702),
    .Q_N(_06576_),
    .Q(\i_time.l_mtimecmp.data_out[25] ));
 sg13g2_dfrbp_1 _15175_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net1302),
    .D(_00763_),
    .Q_N(_06575_),
    .Q(\i_time.l_mtimecmp.data_out[26] ));
 sg13g2_dfrbp_1 _15176_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net1301),
    .D(net3798),
    .Q_N(_06574_),
    .Q(\i_time.l_mtimecmp.data_out[27] ));
 sg13g2_dfrbp_1 _15177_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net1300),
    .D(net3726),
    .Q_N(_06573_),
    .Q(\i_time.l_mtimecmp.data_out[28] ));
 sg13g2_dfrbp_1 _15178_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net1299),
    .D(net3593),
    .Q_N(_06572_),
    .Q(\i_time.l_mtimecmp.data_out[29] ));
 sg13g2_dfrbp_1 _15179_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net1298),
    .D(net3657),
    .Q_N(_06571_),
    .Q(\i_time.l_mtimecmp.data_out[30] ));
 sg13g2_dfrbp_1 _15180_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net1297),
    .D(net3776),
    .Q_N(_06570_),
    .Q(\i_time.l_mtimecmp.data_out[31] ));
 sg13g2_dfrbp_1 _15181_ (.CLK(net2124),
    .RESET_B(net1296),
    .D(_00769_),
    .Q_N(_06569_),
    .Q(\i_spi.read_latency ));
 sg13g2_dfrbp_1 _15182_ (.CLK(net2125),
    .RESET_B(net1294),
    .D(_00770_),
    .Q_N(_06568_),
    .Q(\i_spi.clock_divider[0] ));
 sg13g2_dfrbp_1 _15183_ (.CLK(net2126),
    .RESET_B(net1292),
    .D(_00771_),
    .Q_N(_06567_),
    .Q(\i_spi.clock_divider[1] ));
 sg13g2_dfrbp_1 _15184_ (.CLK(net2127),
    .RESET_B(net1290),
    .D(_00772_),
    .Q_N(_06566_),
    .Q(\i_spi.clock_divider[2] ));
 sg13g2_dfrbp_1 _15185_ (.CLK(net2128),
    .RESET_B(net1288),
    .D(_00773_),
    .Q_N(_06565_),
    .Q(\i_spi.clock_divider[3] ));
 sg13g2_dfrbp_1 _15186_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net1286),
    .D(_00774_),
    .Q_N(_00241_),
    .Q(\i_time.mtime[0] ));
 sg13g2_dfrbp_1 _15187_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net1284),
    .D(_00775_),
    .Q_N(_06564_),
    .Q(\i_time.mtime[1] ));
 sg13g2_dfrbp_1 _15188_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net1282),
    .D(_00776_),
    .Q_N(_06563_),
    .Q(\i_time.mtime[2] ));
 sg13g2_dfrbp_1 _15189_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1280),
    .D(_00777_),
    .Q_N(_06562_),
    .Q(\i_time.mtime[3] ));
 sg13g2_dfrbp_1 _15190_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1278),
    .D(_00778_),
    .Q_N(_06561_),
    .Q(\i_time.mtime[4] ));
 sg13g2_dfrbp_1 _15191_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1276),
    .D(_00779_),
    .Q_N(_06560_),
    .Q(\i_time.mtime[5] ));
 sg13g2_dfrbp_1 _15192_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1274),
    .D(_00780_),
    .Q_N(_06559_),
    .Q(\i_time.mtime[6] ));
 sg13g2_dfrbp_1 _15193_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1272),
    .D(_00781_),
    .Q_N(_06558_),
    .Q(\i_time.mtime[7] ));
 sg13g2_dfrbp_1 _15194_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net1270),
    .D(_00782_),
    .Q_N(_06557_),
    .Q(\i_time.mtime[8] ));
 sg13g2_dfrbp_1 _15195_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net1268),
    .D(net4109),
    .Q_N(_06556_),
    .Q(\i_time.mtime[9] ));
 sg13g2_dfrbp_1 _15196_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net1266),
    .D(_00784_),
    .Q_N(_06555_),
    .Q(\i_time.mtime[10] ));
 sg13g2_dfrbp_1 _15197_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net1264),
    .D(_00785_),
    .Q_N(_06554_),
    .Q(\i_time.mtime[11] ));
 sg13g2_dfrbp_1 _15198_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net1261),
    .D(_00786_),
    .Q_N(_06553_),
    .Q(\i_time.mtime[12] ));
 sg13g2_dfrbp_1 _15199_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1259),
    .D(_00787_),
    .Q_N(_06552_),
    .Q(\i_time.mtime[13] ));
 sg13g2_dfrbp_1 _15200_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1257),
    .D(_00788_),
    .Q_N(_06551_),
    .Q(\i_time.mtime[14] ));
 sg13g2_dfrbp_1 _15201_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1255),
    .D(_00789_),
    .Q_N(_06550_),
    .Q(\i_time.mtime[15] ));
 sg13g2_dfrbp_1 _15202_ (.CLK(clknet_leaf_152_clk_regs),
    .RESET_B(net1253),
    .D(_00790_),
    .Q_N(_06549_),
    .Q(\i_time.mtime[16] ));
 sg13g2_dfrbp_1 _15203_ (.CLK(clknet_leaf_152_clk_regs),
    .RESET_B(net1251),
    .D(_00791_),
    .Q_N(_06548_),
    .Q(\i_time.mtime[17] ));
 sg13g2_dfrbp_1 _15204_ (.CLK(clknet_leaf_152_clk_regs),
    .RESET_B(net1249),
    .D(_00792_),
    .Q_N(_06547_),
    .Q(\i_time.mtime[18] ));
 sg13g2_dfrbp_1 _15205_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net1247),
    .D(_00793_),
    .Q_N(_06546_),
    .Q(\i_time.mtime[19] ));
 sg13g2_dfrbp_1 _15206_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net1245),
    .D(_00794_),
    .Q_N(_06545_),
    .Q(\i_time.mtime[20] ));
 sg13g2_dfrbp_1 _15207_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net1243),
    .D(_00795_),
    .Q_N(_06544_),
    .Q(\i_time.mtime[21] ));
 sg13g2_dfrbp_1 _15208_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net1241),
    .D(net4027),
    .Q_N(_06543_),
    .Q(\i_time.mtime[22] ));
 sg13g2_dfrbp_1 _15209_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net1239),
    .D(net4025),
    .Q_N(_06542_),
    .Q(\i_time.mtime[23] ));
 sg13g2_dfrbp_1 _15210_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net1237),
    .D(_00798_),
    .Q_N(_06541_),
    .Q(\i_time.mtime[24] ));
 sg13g2_dfrbp_1 _15211_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net1235),
    .D(_00799_),
    .Q_N(_06540_),
    .Q(\i_time.mtime[25] ));
 sg13g2_dfrbp_1 _15212_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net1233),
    .D(_00800_),
    .Q_N(_06539_),
    .Q(\i_time.mtime[26] ));
 sg13g2_dfrbp_1 _15213_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net1231),
    .D(_00801_),
    .Q_N(_06538_),
    .Q(\i_time.mtime[27] ));
 sg13g2_dfrbp_1 _15214_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net1229),
    .D(_00802_),
    .Q_N(_06537_),
    .Q(\i_time.mtime[28] ));
 sg13g2_dfrbp_1 _15215_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net1227),
    .D(_00803_),
    .Q_N(_06536_),
    .Q(\i_time.mtime[29] ));
 sg13g2_dfrbp_1 _15216_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net1225),
    .D(_00804_),
    .Q_N(_06535_),
    .Q(\i_time.mtime[30] ));
 sg13g2_dfrbp_1 _15217_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net1595),
    .D(net3865),
    .Q_N(_07194_),
    .Q(\i_time.mtime[31] ));
 sg13g2_dfrbp_1 _15218_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net1223),
    .D(_00063_),
    .Q_N(_06534_),
    .Q(\i_time.timer_interrupt ));
 sg13g2_dfrbp_1 _15219_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net1221),
    .D(_00806_),
    .Q_N(_06533_),
    .Q(\i_game.game_latch_sync[0] ));
 sg13g2_dfrbp_1 _15220_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net1220),
    .D(_00807_),
    .Q_N(_06532_),
    .Q(\i_game.game_latch_sync[1] ));
 sg13g2_dfrbp_1 _15221_ (.CLK(game_clk),
    .RESET_B(net524),
    .D(_00317_),
    .Q_N(\i_game.l_data.data_in[0] ),
    .Q(_00272_));
 sg13g2_dfrbp_1 _15222_ (.CLK(game_clk),
    .RESET_B(net523),
    .D(_00318_),
    .Q_N(\i_game.l_data.data_in[1] ),
    .Q(_00273_));
 sg13g2_dfrbp_1 _15223_ (.CLK(game_clk),
    .RESET_B(net524),
    .D(_00319_),
    .Q_N(\i_game.l_data.data_in[2] ),
    .Q(_00274_));
 sg13g2_dfrbp_1 _15224_ (.CLK(game_clk),
    .RESET_B(net523),
    .D(_00320_),
    .Q_N(\i_game.l_data.data_in[3] ),
    .Q(_00275_));
 sg13g2_dfrbp_1 _15225_ (.CLK(game_clk),
    .RESET_B(net523),
    .D(_00321_),
    .Q_N(\i_game.l_data.data_in[4] ),
    .Q(_00276_));
 sg13g2_dfrbp_1 _15226_ (.CLK(game_clk),
    .RESET_B(net523),
    .D(_00322_),
    .Q_N(\i_game.l_data.data_in[5] ),
    .Q(_00277_));
 sg13g2_dfrbp_1 _15227_ (.CLK(game_clk),
    .RESET_B(net523),
    .D(_00323_),
    .Q_N(\i_game.l_data.data_in[6] ),
    .Q(_00278_));
 sg13g2_dfrbp_1 _15228_ (.CLK(game_clk),
    .RESET_B(net519),
    .D(_00324_),
    .Q_N(\i_game.l_data.data_in[7] ),
    .Q(_00279_));
 sg13g2_dfrbp_1 _15229_ (.CLK(game_clk),
    .RESET_B(net519),
    .D(_00325_),
    .Q_N(\i_game.l_data.data_in[8] ),
    .Q(_00280_));
 sg13g2_dfrbp_1 _15230_ (.CLK(game_clk),
    .RESET_B(net519),
    .D(_00326_),
    .Q_N(\i_game.l_data.data_in[9] ),
    .Q(_00281_));
 sg13g2_dfrbp_1 _15231_ (.CLK(game_clk),
    .RESET_B(net520),
    .D(_00327_),
    .Q_N(\i_game.l_data.data_in[10] ),
    .Q(_00282_));
 sg13g2_dfrbp_1 _15232_ (.CLK(game_clk),
    .RESET_B(net520),
    .D(_00328_),
    .Q_N(\i_game.l_data.data_in[11] ),
    .Q(_00283_));
 sg13g2_dfrbp_1 _15233_ (.CLK(game_clk),
    .RESET_B(net519),
    .D(_00329_),
    .Q_N(\i_game.l_data.data_in[12] ),
    .Q(_00284_));
 sg13g2_dfrbp_1 _15234_ (.CLK(game_clk),
    .RESET_B(net519),
    .D(_00330_),
    .Q_N(\i_game.l_data.data_in[13] ),
    .Q(_00285_));
 sg13g2_dfrbp_1 _15235_ (.CLK(game_clk),
    .RESET_B(net523),
    .D(_00331_),
    .Q_N(\i_game.l_data.data_in[14] ),
    .Q(_00286_));
 sg13g2_dfrbp_1 _15236_ (.CLK(game_clk),
    .RESET_B(net523),
    .D(_00332_),
    .Q_N(\i_game.l_data.data_in[15] ),
    .Q(_00287_));
 sg13g2_dfrbp_1 _15237_ (.CLK(game_clk),
    .RESET_B(net523),
    .D(_00333_),
    .Q_N(\i_game.l_data.data_in[16] ),
    .Q(_00288_));
 sg13g2_dfrbp_1 _15238_ (.CLK(game_clk),
    .RESET_B(net518),
    .D(_00334_),
    .Q_N(\i_game.l_data.data_in[17] ),
    .Q(_00289_));
 sg13g2_dfrbp_1 _15239_ (.CLK(game_clk),
    .RESET_B(net519),
    .D(_00335_),
    .Q_N(\i_game.l_data.data_in[18] ),
    .Q(_00290_));
 sg13g2_dfrbp_1 _15240_ (.CLK(game_clk),
    .RESET_B(net518),
    .D(_00336_),
    .Q_N(\i_game.l_data.data_in[19] ),
    .Q(_00291_));
 sg13g2_dfrbp_1 _15241_ (.CLK(game_clk),
    .RESET_B(net519),
    .D(_00337_),
    .Q_N(\i_game.l_data.data_in[20] ),
    .Q(_00292_));
 sg13g2_dfrbp_1 _15242_ (.CLK(game_clk),
    .RESET_B(net519),
    .D(_00338_),
    .Q_N(\i_game.l_data.data_in[21] ),
    .Q(_00293_));
 sg13g2_dfrbp_1 _15243_ (.CLK(game_clk),
    .RESET_B(net518),
    .D(_00339_),
    .Q_N(\i_game.l_data.data_in[22] ),
    .Q(_00294_));
 sg13g2_dfrbp_1 _15244_ (.CLK(game_clk),
    .RESET_B(net520),
    .D(_00340_),
    .Q_N(\i_game.l_data.data_in[23] ),
    .Q(_00295_));
 sg13g2_dfrbp_1 _15245_ (.CLK(net2129),
    .RESET_B(net1195),
    .D(_00808_),
    .Q_N(_06531_),
    .Q(\i_game.data_latch_wen ));
 sg13g2_dfrbp_1 _15246_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net1193),
    .D(net3828),
    .Q_N(_06530_),
    .Q(debug_uart_txd));
 sg13g2_dfrbp_1 _15247_ (.CLK(net2130),
    .RESET_B(net1192),
    .D(_00810_),
    .Q_N(_06529_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15248_ (.CLK(net2131),
    .RESET_B(net1190),
    .D(_00811_),
    .Q_N(_06528_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15249_ (.CLK(net2132),
    .RESET_B(net1188),
    .D(_00812_),
    .Q_N(_06527_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15250_ (.CLK(net2133),
    .RESET_B(net1186),
    .D(_00813_),
    .Q_N(_06526_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15251_ (.CLK(net2134),
    .RESET_B(net1184),
    .D(_00814_),
    .Q_N(_06525_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15252_ (.CLK(net2135),
    .RESET_B(net1182),
    .D(_00815_),
    .Q_N(_06524_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15253_ (.CLK(net2136),
    .RESET_B(net1180),
    .D(_00816_),
    .Q_N(_06523_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15254_ (.CLK(net2137),
    .RESET_B(net1178),
    .D(_00817_),
    .Q_N(_06522_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15255_ (.CLK(net2138),
    .RESET_B(net1176),
    .D(_00818_),
    .Q_N(_06521_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15256_ (.CLK(net2139),
    .RESET_B(net1174),
    .D(_00819_),
    .Q_N(_06520_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15257_ (.CLK(net2140),
    .RESET_B(net1172),
    .D(_00820_),
    .Q_N(_06519_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15258_ (.CLK(net2141),
    .RESET_B(net1170),
    .D(_00821_),
    .Q_N(_06518_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15259_ (.CLK(net2142),
    .RESET_B(net1168),
    .D(_00822_),
    .Q_N(_06517_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15260_ (.CLK(net2143),
    .RESET_B(net1166),
    .D(_00823_),
    .Q_N(_06516_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15261_ (.CLK(net2144),
    .RESET_B(net1164),
    .D(_00824_),
    .Q_N(_06515_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15262_ (.CLK(net2145),
    .RESET_B(net1157),
    .D(_00825_),
    .Q_N(_06514_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15263_ (.CLK(net2146),
    .RESET_B(net1155),
    .D(_00826_),
    .Q_N(_06513_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15264_ (.CLK(net2147),
    .RESET_B(net1153),
    .D(_00827_),
    .Q_N(_06512_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15265_ (.CLK(net2148),
    .RESET_B(net1151),
    .D(_00828_),
    .Q_N(_06511_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15266_ (.CLK(net2149),
    .RESET_B(net1149),
    .D(_00829_),
    .Q_N(_06510_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15267_ (.CLK(net2150),
    .RESET_B(net1147),
    .D(_00830_),
    .Q_N(_06509_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15268_ (.CLK(net2151),
    .RESET_B(net1145),
    .D(_00831_),
    .Q_N(_06508_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15269_ (.CLK(net2152),
    .RESET_B(net1143),
    .D(_00832_),
    .Q_N(_06507_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15270_ (.CLK(net2153),
    .RESET_B(net1141),
    .D(_00833_),
    .Q_N(_06506_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15271_ (.CLK(net2154),
    .RESET_B(net1139),
    .D(_00834_),
    .Q_N(_06505_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15272_ (.CLK(net2155),
    .RESET_B(net1136),
    .D(_00835_),
    .Q_N(_06504_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15273_ (.CLK(net2156),
    .RESET_B(net1134),
    .D(_00836_),
    .Q_N(_06503_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15274_ (.CLK(net2157),
    .RESET_B(net1132),
    .D(_00837_),
    .Q_N(_06502_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15275_ (.CLK(net2158),
    .RESET_B(net716),
    .D(_00838_),
    .Q_N(_06501_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15276_ (.CLK(net2159),
    .RESET_B(net714),
    .D(_00839_),
    .Q_N(_06500_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15277_ (.CLK(net2160),
    .RESET_B(net712),
    .D(_00840_),
    .Q_N(_06499_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15278_ (.CLK(net2161),
    .RESET_B(net682),
    .D(_00841_),
    .Q_N(_06498_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15279_ (.CLK(net2162),
    .RESET_B(net680),
    .D(_00842_),
    .Q_N(_06497_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15280_ (.CLK(net2163),
    .RESET_B(net678),
    .D(_00843_),
    .Q_N(_06496_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15281_ (.CLK(net2164),
    .RESET_B(net2094),
    .D(_00844_),
    .Q_N(_06495_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15282_ (.CLK(net2165),
    .RESET_B(net2092),
    .D(_00845_),
    .Q_N(_06494_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15283_ (.CLK(net2166),
    .RESET_B(net2090),
    .D(_00846_),
    .Q_N(_06493_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15284_ (.CLK(net2167),
    .RESET_B(net2088),
    .D(_00847_),
    .Q_N(_06492_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15285_ (.CLK(net2168),
    .RESET_B(net2086),
    .D(_00848_),
    .Q_N(_06491_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15286_ (.CLK(net2169),
    .RESET_B(net2084),
    .D(_00849_),
    .Q_N(_06490_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15287_ (.CLK(net2170),
    .RESET_B(net2082),
    .D(_00850_),
    .Q_N(_06489_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15288_ (.CLK(net2171),
    .RESET_B(net2080),
    .D(_00851_),
    .Q_N(_06488_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15289_ (.CLK(net2172),
    .RESET_B(net2078),
    .D(_00852_),
    .Q_N(_06487_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15290_ (.CLK(net2173),
    .RESET_B(net2076),
    .D(_00853_),
    .Q_N(_06486_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15291_ (.CLK(net2174),
    .RESET_B(net2074),
    .D(_00854_),
    .Q_N(_06485_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15292_ (.CLK(net2175),
    .RESET_B(net2072),
    .D(_00855_),
    .Q_N(_06484_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15293_ (.CLK(net2176),
    .RESET_B(net2070),
    .D(_00856_),
    .Q_N(_06483_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15294_ (.CLK(net2177),
    .RESET_B(net2068),
    .D(_00857_),
    .Q_N(_06482_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15295_ (.CLK(net2178),
    .RESET_B(net2066),
    .D(_00858_),
    .Q_N(_06481_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15296_ (.CLK(net2179),
    .RESET_B(net2064),
    .D(_00859_),
    .Q_N(_06480_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15297_ (.CLK(net2180),
    .RESET_B(net2062),
    .D(_00860_),
    .Q_N(_06479_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15298_ (.CLK(net2181),
    .RESET_B(net2060),
    .D(_00861_),
    .Q_N(_06478_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15299_ (.CLK(net2182),
    .RESET_B(net2058),
    .D(_00862_),
    .Q_N(_06477_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15300_ (.CLK(net2183),
    .RESET_B(net2056),
    .D(_00863_),
    .Q_N(_06476_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15301_ (.CLK(net2184),
    .RESET_B(net2054),
    .D(_00864_),
    .Q_N(_06475_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15302_ (.CLK(net2185),
    .RESET_B(net2052),
    .D(_00865_),
    .Q_N(_06474_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15303_ (.CLK(net2186),
    .RESET_B(net2050),
    .D(_00866_),
    .Q_N(_06473_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15304_ (.CLK(net2187),
    .RESET_B(net2048),
    .D(_00867_),
    .Q_N(_06472_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15305_ (.CLK(net2188),
    .RESET_B(net2046),
    .D(_00868_),
    .Q_N(_06471_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15306_ (.CLK(net2189),
    .RESET_B(net2044),
    .D(_00869_),
    .Q_N(_06470_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15307_ (.CLK(net2190),
    .RESET_B(net2042),
    .D(_00870_),
    .Q_N(_06469_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15308_ (.CLK(net2191),
    .RESET_B(net2040),
    .D(_00871_),
    .Q_N(_06468_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15309_ (.CLK(net2192),
    .RESET_B(net2038),
    .D(_00872_),
    .Q_N(_06467_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15310_ (.CLK(net2193),
    .RESET_B(net2036),
    .D(_00873_),
    .Q_N(_06466_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15311_ (.CLK(net2194),
    .RESET_B(net2034),
    .D(_00874_),
    .Q_N(_06465_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15312_ (.CLK(net2195),
    .RESET_B(net2032),
    .D(_00875_),
    .Q_N(_06464_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15313_ (.CLK(net2196),
    .RESET_B(net2030),
    .D(_00876_),
    .Q_N(_06463_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15314_ (.CLK(net2197),
    .RESET_B(net2028),
    .D(_00877_),
    .Q_N(_06462_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15315_ (.CLK(net2198),
    .RESET_B(net2026),
    .D(_00878_),
    .Q_N(_06461_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15316_ (.CLK(net2199),
    .RESET_B(net2024),
    .D(_00879_),
    .Q_N(_06460_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15317_ (.CLK(net2200),
    .RESET_B(net2022),
    .D(_00880_),
    .Q_N(_06459_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15318_ (.CLK(net2201),
    .RESET_B(net2019),
    .D(_00881_),
    .Q_N(_06458_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15319_ (.CLK(net2202),
    .RESET_B(net2017),
    .D(_00882_),
    .Q_N(_06457_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15320_ (.CLK(net2203),
    .RESET_B(net2015),
    .D(_00883_),
    .Q_N(_06456_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15321_ (.CLK(net2204),
    .RESET_B(net2013),
    .D(_00884_),
    .Q_N(_06455_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15322_ (.CLK(net2205),
    .RESET_B(net2011),
    .D(_00885_),
    .Q_N(_06454_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15323_ (.CLK(net2206),
    .RESET_B(net2009),
    .D(_00886_),
    .Q_N(_06453_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15324_ (.CLK(net2207),
    .RESET_B(net2007),
    .D(_00887_),
    .Q_N(_06452_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15325_ (.CLK(net2208),
    .RESET_B(net2005),
    .D(_00888_),
    .Q_N(_06451_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15326_ (.CLK(net2209),
    .RESET_B(net2003),
    .D(_00889_),
    .Q_N(_06450_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15327_ (.CLK(net2210),
    .RESET_B(net2001),
    .D(_00890_),
    .Q_N(_06449_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15328_ (.CLK(net2211),
    .RESET_B(net1999),
    .D(_00891_),
    .Q_N(_06448_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15329_ (.CLK(net2212),
    .RESET_B(net1997),
    .D(_00892_),
    .Q_N(_06447_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15330_ (.CLK(net2213),
    .RESET_B(net1995),
    .D(_00893_),
    .Q_N(_06446_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15331_ (.CLK(net2214),
    .RESET_B(net1993),
    .D(_00894_),
    .Q_N(_06445_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15332_ (.CLK(net2215),
    .RESET_B(net1991),
    .D(_00895_),
    .Q_N(_06444_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15333_ (.CLK(net2216),
    .RESET_B(net1989),
    .D(_00896_),
    .Q_N(_06443_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15334_ (.CLK(net2217),
    .RESET_B(net1987),
    .D(_00897_),
    .Q_N(_06442_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15335_ (.CLK(net2218),
    .RESET_B(net1985),
    .D(_00898_),
    .Q_N(_06441_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15336_ (.CLK(net2219),
    .RESET_B(net1983),
    .D(_00899_),
    .Q_N(_06440_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15337_ (.CLK(net2220),
    .RESET_B(net1981),
    .D(_00900_),
    .Q_N(_06439_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15338_ (.CLK(net2221),
    .RESET_B(net1979),
    .D(_00901_),
    .Q_N(_06438_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15339_ (.CLK(net2222),
    .RESET_B(net1977),
    .D(_00902_),
    .Q_N(_06437_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15340_ (.CLK(net2223),
    .RESET_B(net1975),
    .D(_00903_),
    .Q_N(_06436_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15341_ (.CLK(net2224),
    .RESET_B(net1973),
    .D(_00904_),
    .Q_N(_06435_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15342_ (.CLK(net2225),
    .RESET_B(net1971),
    .D(_00905_),
    .Q_N(_06434_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15343_ (.CLK(net2226),
    .RESET_B(net1969),
    .D(_00906_),
    .Q_N(_06433_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15344_ (.CLK(net2227),
    .RESET_B(net1967),
    .D(_00907_),
    .Q_N(_06432_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15345_ (.CLK(net2228),
    .RESET_B(net1965),
    .D(_00908_),
    .Q_N(_06431_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15346_ (.CLK(net2229),
    .RESET_B(net1963),
    .D(_00909_),
    .Q_N(_06430_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15347_ (.CLK(net2230),
    .RESET_B(net1961),
    .D(_00910_),
    .Q_N(_06429_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15348_ (.CLK(net2231),
    .RESET_B(net1959),
    .D(_00911_),
    .Q_N(_06428_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15349_ (.CLK(net2232),
    .RESET_B(net1957),
    .D(_00912_),
    .Q_N(_06427_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15350_ (.CLK(net2233),
    .RESET_B(net1955),
    .D(_00913_),
    .Q_N(_06426_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15351_ (.CLK(net2234),
    .RESET_B(net1953),
    .D(_00914_),
    .Q_N(_06425_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15352_ (.CLK(net2235),
    .RESET_B(net1951),
    .D(_00915_),
    .Q_N(_06424_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15353_ (.CLK(net2236),
    .RESET_B(net1949),
    .D(_00916_),
    .Q_N(_06423_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15354_ (.CLK(net2237),
    .RESET_B(net1947),
    .D(_00917_),
    .Q_N(_06422_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15355_ (.CLK(net2238),
    .RESET_B(net1945),
    .D(_00918_),
    .Q_N(_06421_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15356_ (.CLK(net2239),
    .RESET_B(net1943),
    .D(_00919_),
    .Q_N(_06420_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15357_ (.CLK(net2240),
    .RESET_B(net1941),
    .D(_00920_),
    .Q_N(_06419_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15358_ (.CLK(net2241),
    .RESET_B(net1939),
    .D(_00921_),
    .Q_N(_06418_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15359_ (.CLK(net2242),
    .RESET_B(net1937),
    .D(_00922_),
    .Q_N(_06417_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15360_ (.CLK(net2243),
    .RESET_B(net1935),
    .D(_00923_),
    .Q_N(_06416_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15361_ (.CLK(net2244),
    .RESET_B(net1933),
    .D(_00924_),
    .Q_N(_06415_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15362_ (.CLK(net2245),
    .RESET_B(net1931),
    .D(_00925_),
    .Q_N(_06414_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15363_ (.CLK(net2246),
    .RESET_B(net1929),
    .D(_00926_),
    .Q_N(_06413_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15364_ (.CLK(net2247),
    .RESET_B(net1927),
    .D(_00927_),
    .Q_N(_06412_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15365_ (.CLK(net2248),
    .RESET_B(net1925),
    .D(_00928_),
    .Q_N(_06411_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15366_ (.CLK(net2249),
    .RESET_B(net1923),
    .D(_00929_),
    .Q_N(_06410_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15367_ (.CLK(net2250),
    .RESET_B(net1921),
    .D(_00930_),
    .Q_N(_06409_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15368_ (.CLK(net2251),
    .RESET_B(net1919),
    .D(_00931_),
    .Q_N(_06408_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15369_ (.CLK(net2252),
    .RESET_B(net1917),
    .D(_00932_),
    .Q_N(_06407_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15370_ (.CLK(net2253),
    .RESET_B(net1915),
    .D(_00933_),
    .Q_N(_06406_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15371_ (.CLK(net2254),
    .RESET_B(net1913),
    .D(_00934_),
    .Q_N(_06405_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15372_ (.CLK(net2255),
    .RESET_B(net1911),
    .D(_00935_),
    .Q_N(_06404_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15373_ (.CLK(net2256),
    .RESET_B(net1909),
    .D(_00936_),
    .Q_N(_06403_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15374_ (.CLK(net2257),
    .RESET_B(net1907),
    .D(_00937_),
    .Q_N(_06402_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15375_ (.CLK(net2258),
    .RESET_B(net1905),
    .D(_00938_),
    .Q_N(_06401_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15376_ (.CLK(net2259),
    .RESET_B(net1903),
    .D(_00939_),
    .Q_N(_06400_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15377_ (.CLK(net2260),
    .RESET_B(net1901),
    .D(_00940_),
    .Q_N(_06399_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15378_ (.CLK(net2261),
    .RESET_B(net1899),
    .D(_00941_),
    .Q_N(_06398_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15379_ (.CLK(net2262),
    .RESET_B(net1897),
    .D(_00942_),
    .Q_N(_06397_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15380_ (.CLK(net2263),
    .RESET_B(net1895),
    .D(_00943_),
    .Q_N(_06396_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15381_ (.CLK(net2264),
    .RESET_B(net1893),
    .D(_00944_),
    .Q_N(_06395_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15382_ (.CLK(net2265),
    .RESET_B(net1891),
    .D(_00945_),
    .Q_N(_06394_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15383_ (.CLK(net2266),
    .RESET_B(net1889),
    .D(_00946_),
    .Q_N(_06393_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15384_ (.CLK(net2267),
    .RESET_B(net1887),
    .D(_00947_),
    .Q_N(_06392_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15385_ (.CLK(net2268),
    .RESET_B(net1885),
    .D(_00948_),
    .Q_N(_06391_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15386_ (.CLK(net2269),
    .RESET_B(net1883),
    .D(_00949_),
    .Q_N(_06390_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15387_ (.CLK(net2270),
    .RESET_B(net1881),
    .D(_00950_),
    .Q_N(_06389_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15388_ (.CLK(net2271),
    .RESET_B(net1879),
    .D(_00951_),
    .Q_N(_06388_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15389_ (.CLK(net2272),
    .RESET_B(net1877),
    .D(_00952_),
    .Q_N(_06387_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15390_ (.CLK(net2273),
    .RESET_B(net1875),
    .D(_00953_),
    .Q_N(_06386_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15391_ (.CLK(net2274),
    .RESET_B(net1873),
    .D(_00954_),
    .Q_N(_06385_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15392_ (.CLK(net2275),
    .RESET_B(net1871),
    .D(_00955_),
    .Q_N(_06384_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15393_ (.CLK(net2276),
    .RESET_B(net1869),
    .D(_00956_),
    .Q_N(_06383_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15394_ (.CLK(net2277),
    .RESET_B(net1867),
    .D(_00957_),
    .Q_N(_06382_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15395_ (.CLK(net2278),
    .RESET_B(net1865),
    .D(_00958_),
    .Q_N(_06381_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15396_ (.CLK(net2279),
    .RESET_B(net1863),
    .D(_00959_),
    .Q_N(_06380_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15397_ (.CLK(net2280),
    .RESET_B(net1861),
    .D(_00960_),
    .Q_N(_06379_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15398_ (.CLK(net2281),
    .RESET_B(net1859),
    .D(_00961_),
    .Q_N(_06378_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15399_ (.CLK(net2282),
    .RESET_B(net1857),
    .D(_00962_),
    .Q_N(_06377_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15400_ (.CLK(net2283),
    .RESET_B(net1855),
    .D(_00963_),
    .Q_N(_06376_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15401_ (.CLK(net2284),
    .RESET_B(net1853),
    .D(_00964_),
    .Q_N(_06375_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15402_ (.CLK(net2285),
    .RESET_B(net1851),
    .D(_00965_),
    .Q_N(_06374_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15403_ (.CLK(net2286),
    .RESET_B(net1849),
    .D(_00966_),
    .Q_N(_06373_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15404_ (.CLK(net2287),
    .RESET_B(net1847),
    .D(_00967_),
    .Q_N(_06372_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15405_ (.CLK(net2288),
    .RESET_B(net1845),
    .D(_00968_),
    .Q_N(_06371_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15406_ (.CLK(net2289),
    .RESET_B(net1843),
    .D(_00969_),
    .Q_N(_06370_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15407_ (.CLK(net2290),
    .RESET_B(net1841),
    .D(_00970_),
    .Q_N(_06369_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15408_ (.CLK(net2291),
    .RESET_B(net1839),
    .D(_00971_),
    .Q_N(_06368_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15409_ (.CLK(net2292),
    .RESET_B(net1837),
    .D(_00972_),
    .Q_N(_06367_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15410_ (.CLK(net2293),
    .RESET_B(net1822),
    .D(_00973_),
    .Q_N(_06366_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15411_ (.CLK(net2294),
    .RESET_B(net1820),
    .D(_00974_),
    .Q_N(_06365_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15412_ (.CLK(net2295),
    .RESET_B(net1818),
    .D(_00975_),
    .Q_N(_06364_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15413_ (.CLK(net2296),
    .RESET_B(net1816),
    .D(_00976_),
    .Q_N(_06363_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15414_ (.CLK(net2297),
    .RESET_B(net1814),
    .D(_00977_),
    .Q_N(_06362_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15415_ (.CLK(net2298),
    .RESET_B(net1812),
    .D(_00978_),
    .Q_N(_00256_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15416_ (.CLK(net2299),
    .RESET_B(net1810),
    .D(_00979_),
    .Q_N(_00257_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15417_ (.CLK(net2300),
    .RESET_B(net1808),
    .D(_00980_),
    .Q_N(_00258_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15418_ (.CLK(net2301),
    .RESET_B(net1806),
    .D(_00981_),
    .Q_N(_00259_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15419_ (.CLK(net2302),
    .RESET_B(net1804),
    .D(_00982_),
    .Q_N(_00260_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15420_ (.CLK(net2303),
    .RESET_B(net1802),
    .D(_00983_),
    .Q_N(_00261_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15421_ (.CLK(net2304),
    .RESET_B(net1800),
    .D(_00984_),
    .Q_N(_00262_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15422_ (.CLK(net2305),
    .RESET_B(net1798),
    .D(_00985_),
    .Q_N(_00263_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15423_ (.CLK(net2306),
    .RESET_B(net1796),
    .D(_00986_),
    .Q_N(_06361_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15424_ (.CLK(net2307),
    .RESET_B(net1794),
    .D(_00987_),
    .Q_N(_06360_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15425_ (.CLK(net2308),
    .RESET_B(net1792),
    .D(_00988_),
    .Q_N(_06359_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15426_ (.CLK(net2309),
    .RESET_B(net1790),
    .D(_00989_),
    .Q_N(_06358_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15427_ (.CLK(net2310),
    .RESET_B(net1788),
    .D(_00990_),
    .Q_N(_06357_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15428_ (.CLK(net2311),
    .RESET_B(net1786),
    .D(_00991_),
    .Q_N(_06356_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15429_ (.CLK(net2312),
    .RESET_B(net1784),
    .D(_00992_),
    .Q_N(_06355_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15430_ (.CLK(net2313),
    .RESET_B(net1782),
    .D(_00993_),
    .Q_N(_06354_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15431_ (.CLK(net2314),
    .RESET_B(net1780),
    .D(_00994_),
    .Q_N(_06353_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15432_ (.CLK(net2315),
    .RESET_B(net1778),
    .D(_00995_),
    .Q_N(_06352_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15433_ (.CLK(net2316),
    .RESET_B(net1776),
    .D(_00996_),
    .Q_N(_06351_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15434_ (.CLK(net2317),
    .RESET_B(net1774),
    .D(_00997_),
    .Q_N(_06350_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15435_ (.CLK(net2318),
    .RESET_B(net1772),
    .D(_00998_),
    .Q_N(_06349_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15436_ (.CLK(net2319),
    .RESET_B(net1770),
    .D(_00999_),
    .Q_N(_06348_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15437_ (.CLK(net2320),
    .RESET_B(net1768),
    .D(_01000_),
    .Q_N(_06347_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15438_ (.CLK(net2321),
    .RESET_B(net1766),
    .D(_01001_),
    .Q_N(_06346_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15439_ (.CLK(net2322),
    .RESET_B(net1764),
    .D(_01002_),
    .Q_N(_06345_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15440_ (.CLK(net2323),
    .RESET_B(net1762),
    .D(_01003_),
    .Q_N(_06344_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15441_ (.CLK(net2324),
    .RESET_B(net1760),
    .D(_01004_),
    .Q_N(_06343_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15442_ (.CLK(net2325),
    .RESET_B(net1758),
    .D(_01005_),
    .Q_N(_06342_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15443_ (.CLK(net2326),
    .RESET_B(net1756),
    .D(_01006_),
    .Q_N(_06341_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15444_ (.CLK(net2327),
    .RESET_B(net1754),
    .D(_01007_),
    .Q_N(_06340_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15445_ (.CLK(net2328),
    .RESET_B(net1752),
    .D(_01008_),
    .Q_N(_06339_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15446_ (.CLK(net2329),
    .RESET_B(net1750),
    .D(_01009_),
    .Q_N(_06338_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15447_ (.CLK(net2330),
    .RESET_B(net1748),
    .D(_01010_),
    .Q_N(_06337_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15448_ (.CLK(net2331),
    .RESET_B(net1746),
    .D(_01011_),
    .Q_N(_06336_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15449_ (.CLK(net2332),
    .RESET_B(net1744),
    .D(_01012_),
    .Q_N(_06335_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15450_ (.CLK(net2333),
    .RESET_B(net1742),
    .D(_01013_),
    .Q_N(_06334_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15451_ (.CLK(net2334),
    .RESET_B(net1740),
    .D(_01014_),
    .Q_N(_06333_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15452_ (.CLK(net2335),
    .RESET_B(net1738),
    .D(_01015_),
    .Q_N(_06332_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15453_ (.CLK(net2336),
    .RESET_B(net1736),
    .D(_01016_),
    .Q_N(_06331_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15454_ (.CLK(net2337),
    .RESET_B(net1734),
    .D(_01017_),
    .Q_N(_06330_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15455_ (.CLK(net2338),
    .RESET_B(net1732),
    .D(_01018_),
    .Q_N(_06329_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15456_ (.CLK(net2339),
    .RESET_B(net1730),
    .D(_01019_),
    .Q_N(_06328_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15457_ (.CLK(net2340),
    .RESET_B(net1728),
    .D(_01020_),
    .Q_N(_06327_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15458_ (.CLK(net2341),
    .RESET_B(net1726),
    .D(_01021_),
    .Q_N(_06326_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15459_ (.CLK(net2342),
    .RESET_B(net1724),
    .D(_01022_),
    .Q_N(_06325_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15460_ (.CLK(net2343),
    .RESET_B(net1722),
    .D(_01023_),
    .Q_N(_06324_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15461_ (.CLK(net2344),
    .RESET_B(net1720),
    .D(_01024_),
    .Q_N(_06323_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15462_ (.CLK(net2345),
    .RESET_B(net1718),
    .D(_01025_),
    .Q_N(_06322_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15463_ (.CLK(net2346),
    .RESET_B(net1716),
    .D(_01026_),
    .Q_N(_06321_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15464_ (.CLK(net2347),
    .RESET_B(net1714),
    .D(_01027_),
    .Q_N(_06320_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15465_ (.CLK(net2348),
    .RESET_B(net1712),
    .D(_01028_),
    .Q_N(_06319_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15466_ (.CLK(net2349),
    .RESET_B(net1710),
    .D(_01029_),
    .Q_N(_06318_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15467_ (.CLK(net2350),
    .RESET_B(net1708),
    .D(_01030_),
    .Q_N(_06317_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15468_ (.CLK(net2351),
    .RESET_B(net1706),
    .D(_01031_),
    .Q_N(_06316_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15469_ (.CLK(net2352),
    .RESET_B(net1704),
    .D(_01032_),
    .Q_N(_06315_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15470_ (.CLK(net2353),
    .RESET_B(net1702),
    .D(_01033_),
    .Q_N(_06314_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15471_ (.CLK(net2354),
    .RESET_B(net1700),
    .D(_01034_),
    .Q_N(_06313_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15472_ (.CLK(net2355),
    .RESET_B(net1698),
    .D(_01035_),
    .Q_N(_06312_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15473_ (.CLK(net2356),
    .RESET_B(net1696),
    .D(_01036_),
    .Q_N(_06311_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15474_ (.CLK(net2357),
    .RESET_B(net1694),
    .D(_01037_),
    .Q_N(_06310_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15475_ (.CLK(net2358),
    .RESET_B(net1692),
    .D(_01038_),
    .Q_N(_06309_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15476_ (.CLK(net2359),
    .RESET_B(net1690),
    .D(_01039_),
    .Q_N(_06308_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15477_ (.CLK(net2360),
    .RESET_B(net1688),
    .D(_01040_),
    .Q_N(_06307_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15478_ (.CLK(net2361),
    .RESET_B(net1666),
    .D(_01041_),
    .Q_N(_06306_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15479_ (.CLK(net2362),
    .RESET_B(net1664),
    .D(_01042_),
    .Q_N(_06305_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15480_ (.CLK(net2363),
    .RESET_B(net1658),
    .D(_01043_),
    .Q_N(_06304_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15481_ (.CLK(net2364),
    .RESET_B(net1656),
    .D(_01044_),
    .Q_N(_06303_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15482_ (.CLK(net2365),
    .RESET_B(net1654),
    .D(_01045_),
    .Q_N(_06302_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15483_ (.CLK(net2366),
    .RESET_B(net1652),
    .D(_01046_),
    .Q_N(_06301_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15484_ (.CLK(net2367),
    .RESET_B(net1650),
    .D(_01047_),
    .Q_N(_06300_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15485_ (.CLK(net2368),
    .RESET_B(net1648),
    .D(_01048_),
    .Q_N(_06299_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15486_ (.CLK(net2369),
    .RESET_B(net1646),
    .D(_01049_),
    .Q_N(_06298_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15487_ (.CLK(net2370),
    .RESET_B(net1644),
    .D(_01050_),
    .Q_N(_06297_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[0] ));
 sg13g2_dfrbp_1 _15488_ (.CLK(net2371),
    .RESET_B(net1642),
    .D(_01051_),
    .Q_N(_06296_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[1] ));
 sg13g2_dfrbp_1 _15489_ (.CLK(net2372),
    .RESET_B(net1640),
    .D(_01052_),
    .Q_N(_06295_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[2] ));
 sg13g2_dfrbp_1 _15490_ (.CLK(net2373),
    .RESET_B(net1638),
    .D(_01053_),
    .Q_N(_06294_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[3] ));
 sg13g2_dfrbp_1 _15491_ (.CLK(net2374),
    .RESET_B(net1636),
    .D(_01054_),
    .Q_N(_06293_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[4] ));
 sg13g2_dfrbp_1 _15492_ (.CLK(net2375),
    .RESET_B(net1634),
    .D(_01055_),
    .Q_N(_06292_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[5] ));
 sg13g2_dfrbp_1 _15493_ (.CLK(net2376),
    .RESET_B(net1632),
    .D(_01056_),
    .Q_N(_06291_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[6] ));
 sg13g2_dfrbp_1 _15494_ (.CLK(net2377),
    .RESET_B(net1630),
    .D(_01057_),
    .Q_N(_06290_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[7] ));
 sg13g2_dfrbp_1 _15495_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net1596),
    .D(net3946),
    .Q_N(_07195_),
    .Q(\i_latch_mem.data_ready ));
 sg13g2_dfrbp_1 _15496_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net1597),
    .D(_00031_),
    .Q_N(_07196_),
    .Q(\i_latch_mem.data_out[0] ));
 sg13g2_dfrbp_1 _15497_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net1598),
    .D(_00042_),
    .Q_N(_07197_),
    .Q(\i_latch_mem.data_out[1] ));
 sg13g2_dfrbp_1 _15498_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net1599),
    .D(_00053_),
    .Q_N(_07198_),
    .Q(\i_latch_mem.data_out[2] ));
 sg13g2_dfrbp_1 _15499_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net1600),
    .D(_00056_),
    .Q_N(_07199_),
    .Q(\i_latch_mem.data_out[3] ));
 sg13g2_dfrbp_1 _15500_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net1601),
    .D(_00057_),
    .Q_N(_07200_),
    .Q(\i_latch_mem.data_out[4] ));
 sg13g2_dfrbp_1 _15501_ (.CLK(clknet_leaf_143_clk_regs),
    .RESET_B(net1602),
    .D(_00058_),
    .Q_N(_07201_),
    .Q(\i_latch_mem.data_out[5] ));
 sg13g2_dfrbp_1 _15502_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net1603),
    .D(_00059_),
    .Q_N(_07202_),
    .Q(\i_latch_mem.data_out[6] ));
 sg13g2_dfrbp_1 _15503_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net1604),
    .D(_00060_),
    .Q_N(_07203_),
    .Q(\i_latch_mem.data_out[7] ));
 sg13g2_dfrbp_1 _15504_ (.CLK(clknet_leaf_144_clk_regs),
    .RESET_B(net1605),
    .D(net3427),
    .Q_N(_07204_),
    .Q(\i_latch_mem.data_out[8] ));
 sg13g2_dfrbp_1 _15505_ (.CLK(clknet_leaf_143_clk_regs),
    .RESET_B(net1606),
    .D(net3353),
    .Q_N(_07205_),
    .Q(\i_latch_mem.data_out[9] ));
 sg13g2_dfrbp_1 _15506_ (.CLK(clknet_leaf_144_clk_regs),
    .RESET_B(net1607),
    .D(net3011),
    .Q_N(_07206_),
    .Q(\i_latch_mem.data_out[10] ));
 sg13g2_dfrbp_1 _15507_ (.CLK(clknet_leaf_144_clk_regs),
    .RESET_B(net1608),
    .D(net3002),
    .Q_N(_07207_),
    .Q(\i_latch_mem.data_out[11] ));
 sg13g2_dfrbp_1 _15508_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net1609),
    .D(net3143),
    .Q_N(_07208_),
    .Q(\i_latch_mem.data_out[12] ));
 sg13g2_dfrbp_1 _15509_ (.CLK(clknet_leaf_144_clk_regs),
    .RESET_B(net1610),
    .D(net3607),
    .Q_N(_07209_),
    .Q(\i_latch_mem.data_out[13] ));
 sg13g2_dfrbp_1 _15510_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net1611),
    .D(net3230),
    .Q_N(_07210_),
    .Q(\i_latch_mem.data_out[14] ));
 sg13g2_dfrbp_1 _15511_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net1612),
    .D(net3183),
    .Q_N(_07211_),
    .Q(\i_latch_mem.data_out[15] ));
 sg13g2_dfrbp_1 _15512_ (.CLK(clknet_leaf_142_clk_regs),
    .RESET_B(net1613),
    .D(_00038_),
    .Q_N(_07212_),
    .Q(\i_latch_mem.data_out[16] ));
 sg13g2_dfrbp_1 _15513_ (.CLK(clknet_leaf_142_clk_regs),
    .RESET_B(net1614),
    .D(_00039_),
    .Q_N(_07213_),
    .Q(\i_latch_mem.data_out[17] ));
 sg13g2_dfrbp_1 _15514_ (.CLK(clknet_leaf_143_clk_regs),
    .RESET_B(net1615),
    .D(_00040_),
    .Q_N(_07214_),
    .Q(\i_latch_mem.data_out[18] ));
 sg13g2_dfrbp_1 _15515_ (.CLK(clknet_leaf_143_clk_regs),
    .RESET_B(net1616),
    .D(_00041_),
    .Q_N(_07215_),
    .Q(\i_latch_mem.data_out[19] ));
 sg13g2_dfrbp_1 _15516_ (.CLK(clknet_leaf_143_clk_regs),
    .RESET_B(net1617),
    .D(_00043_),
    .Q_N(_07216_),
    .Q(\i_latch_mem.data_out[20] ));
 sg13g2_dfrbp_1 _15517_ (.CLK(clknet_leaf_143_clk_regs),
    .RESET_B(net1618),
    .D(_00044_),
    .Q_N(_07217_),
    .Q(\i_latch_mem.data_out[21] ));
 sg13g2_dfrbp_1 _15518_ (.CLK(clknet_leaf_142_clk_regs),
    .RESET_B(net1619),
    .D(_00045_),
    .Q_N(_07218_),
    .Q(\i_latch_mem.data_out[22] ));
 sg13g2_dfrbp_1 _15519_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net1620),
    .D(_00046_),
    .Q_N(_07219_),
    .Q(\i_latch_mem.data_out[23] ));
 sg13g2_dfrbp_1 _15520_ (.CLK(clknet_leaf_144_clk_regs),
    .RESET_B(net1621),
    .D(net3221),
    .Q_N(_07220_),
    .Q(\i_latch_mem.data_out[24] ));
 sg13g2_dfrbp_1 _15521_ (.CLK(clknet_leaf_143_clk_regs),
    .RESET_B(net1622),
    .D(net3239),
    .Q_N(_07221_),
    .Q(\i_latch_mem.data_out[25] ));
 sg13g2_dfrbp_1 _15522_ (.CLK(clknet_leaf_144_clk_regs),
    .RESET_B(net1623),
    .D(net3256),
    .Q_N(_07222_),
    .Q(\i_latch_mem.data_out[26] ));
 sg13g2_dfrbp_1 _15523_ (.CLK(clknet_leaf_144_clk_regs),
    .RESET_B(net1624),
    .D(net3289),
    .Q_N(_07223_),
    .Q(\i_latch_mem.data_out[27] ));
 sg13g2_dfrbp_1 _15524_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net1625),
    .D(net3248),
    .Q_N(_07224_),
    .Q(\i_latch_mem.data_out[28] ));
 sg13g2_dfrbp_1 _15525_ (.CLK(clknet_leaf_143_clk_regs),
    .RESET_B(net1626),
    .D(net3269),
    .Q_N(_07225_),
    .Q(\i_latch_mem.data_out[29] ));
 sg13g2_dfrbp_1 _15526_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net1659),
    .D(net3258),
    .Q_N(_07226_),
    .Q(\i_latch_mem.data_out[30] ));
 sg13g2_dfrbp_1 _15527_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net1628),
    .D(net3232),
    .Q_N(_06289_),
    .Q(\i_latch_mem.data_out[31] ));
 sg13g2_dfrbp_1 _15528_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1627),
    .D(_01059_),
    .Q_N(_06288_),
    .Q(\controller1_data[0] ));
 sg13g2_dfrbp_1 _15529_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1594),
    .D(_01060_),
    .Q_N(_06287_),
    .Q(\controller1_data[1] ));
 sg13g2_dfrbp_1 _15530_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1593),
    .D(_01061_),
    .Q_N(_06286_),
    .Q(\controller1_data[2] ));
 sg13g2_dfrbp_1 _15531_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1592),
    .D(_01062_),
    .Q_N(_06285_),
    .Q(\controller1_data[3] ));
 sg13g2_dfrbp_1 _15532_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net1591),
    .D(_01063_),
    .Q_N(_06284_),
    .Q(\controller1_data[4] ));
 sg13g2_dfrbp_1 _15533_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net1590),
    .D(_01064_),
    .Q_N(_06283_),
    .Q(\controller1_data[5] ));
 sg13g2_dfrbp_1 _15534_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net1589),
    .D(_01065_),
    .Q_N(_06282_),
    .Q(\controller1_data[6] ));
 sg13g2_dfrbp_1 _15535_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net1588),
    .D(_01066_),
    .Q_N(_06281_),
    .Q(\controller1_data[7] ));
 sg13g2_dfrbp_1 _15536_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net1587),
    .D(_01067_),
    .Q_N(_06280_),
    .Q(\controller1_data[8] ));
 sg13g2_dfrbp_1 _15537_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net1586),
    .D(_01068_),
    .Q_N(_06279_),
    .Q(\controller1_data[9] ));
 sg13g2_dfrbp_1 _15538_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net1585),
    .D(_01069_),
    .Q_N(_06278_),
    .Q(\controller1_data[10] ));
 sg13g2_dfrbp_1 _15539_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net1584),
    .D(_01070_),
    .Q_N(_06277_),
    .Q(\controller1_data[11] ));
 sg13g2_dfrbp_1 _15540_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net1583),
    .D(_01071_),
    .Q_N(_06276_),
    .Q(\controller2_data[0] ));
 sg13g2_dfrbp_1 _15541_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net1582),
    .D(_01072_),
    .Q_N(_06275_),
    .Q(\controller2_data[1] ));
 sg13g2_dfrbp_1 _15542_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1581),
    .D(_01073_),
    .Q_N(_06274_),
    .Q(\controller2_data[2] ));
 sg13g2_dfrbp_1 _15543_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net1580),
    .D(_01074_),
    .Q_N(_06273_),
    .Q(\controller2_data[3] ));
 sg13g2_dfrbp_1 _15544_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net1579),
    .D(_01075_),
    .Q_N(_06272_),
    .Q(\controller2_data[4] ));
 sg13g2_dfrbp_1 _15545_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1578),
    .D(_01076_),
    .Q_N(_06271_),
    .Q(\controller2_data[5] ));
 sg13g2_dfrbp_1 _15546_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1577),
    .D(_01077_),
    .Q_N(_06270_),
    .Q(\controller2_data[6] ));
 sg13g2_dfrbp_1 _15547_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net1576),
    .D(_01078_),
    .Q_N(_06269_),
    .Q(\controller2_data[7] ));
 sg13g2_dfrbp_1 _15548_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1575),
    .D(_01079_),
    .Q_N(_06268_),
    .Q(\controller2_data[8] ));
 sg13g2_dfrbp_1 _15549_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net1574),
    .D(_01080_),
    .Q_N(_06267_),
    .Q(\controller2_data[9] ));
 sg13g2_dfrbp_1 _15550_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net1573),
    .D(_01081_),
    .Q_N(_06266_),
    .Q(\controller2_data[10] ));
 sg13g2_dfrbp_1 _15551_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net1572),
    .D(_01082_),
    .Q_N(_06265_),
    .Q(\controller2_data[11] ));
 sg13g2_dfrbp_1 _15552_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net1571),
    .D(_01083_),
    .Q_N(_06264_),
    .Q(\i_latch_mem.cycle[1] ));
 sg13g2_dfrbp_1 _15553_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net1569),
    .D(_01084_),
    .Q_N(_06263_),
    .Q(\i_tinyqv.cpu.i_core.mie[4] ));
 sg13g2_dfrbp_1 _15554_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net1567),
    .D(net3157),
    .Q_N(_00166_),
    .Q(\i_tinyqv.cpu.i_core.mie[3] ));
 sg13g2_dfrbp_1 _15555_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net1552),
    .D(_01086_),
    .Q_N(_06262_),
    .Q(\i_tinyqv.cpu.i_core.mie[2] ));
 sg13g2_dfrbp_1 _15556_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net1547),
    .D(net3688),
    .Q_N(_06261_),
    .Q(\i_tinyqv.cpu.i_core.mie[1] ));
 sg13g2_dfrbp_1 _15557_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net1543),
    .D(_01088_),
    .Q_N(_06260_),
    .Q(\i_tinyqv.cpu.i_core.mie[0] ));
 sg13g2_dfrbp_1 _15558_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net1539),
    .D(net3764),
    .Q_N(_06259_),
    .Q(\i_tinyqv.cpu.i_core.mip[1] ));
 sg13g2_dfrbp_1 _15559_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net1660),
    .D(net3774),
    .Q_N(_07227_),
    .Q(\i_tinyqv.cpu.i_core.mip[0] ));
 sg13g2_dfrbp_1 _15560_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net1661),
    .D(\debug_rd[0] ),
    .Q_N(_07228_),
    .Q(\debug_rd_r[0] ));
 sg13g2_dfrbp_1 _15561_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1662),
    .D(\debug_rd[1] ),
    .Q_N(_07229_),
    .Q(\debug_rd_r[1] ));
 sg13g2_dfrbp_1 _15562_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net1668),
    .D(\debug_rd[2] ),
    .Q_N(_07230_),
    .Q(\debug_rd_r[2] ));
 sg13g2_dfrbp_1 _15563_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1535),
    .D(\debug_rd[3] ),
    .Q_N(_06258_),
    .Q(\debug_rd_r[3] ));
 sg13g2_dfrbp_1 _15564_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net1531),
    .D(_01091_),
    .Q_N(_06257_),
    .Q(\i_uart_tx.txd_reg ));
 sg13g2_dfrbp_1 _15565_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net1527),
    .D(_01092_),
    .Q_N(_06256_),
    .Q(debug_register_data));
 sg13g2_dfrbp_1 _15566_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net1525),
    .D(_01093_),
    .Q_N(_06255_),
    .Q(\mhz_clk_sync[0] ));
 sg13g2_dfrbp_1 _15567_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net1523),
    .D(_01094_),
    .Q_N(_06254_),
    .Q(\mhz_clk_sync[1] ));
 sg13g2_dfrbp_1 _15568_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net1669),
    .D(_01095_),
    .Q_N(_07231_),
    .Q(\mhz_clk_sync[2] ));
 sg13g2_dfrbp_1 _15569_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net1670),
    .D(_00008_),
    .Q_N(_07232_),
    .Q(\gpio_out_sel[0] ));
 sg13g2_dfrbp_1 _15570_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net1671),
    .D(net3557),
    .Q_N(_07233_),
    .Q(\gpio_out_sel[1] ));
 sg13g2_dfrbp_1 _15571_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net1672),
    .D(net3699),
    .Q_N(_07234_),
    .Q(\gpio_out_sel[2] ));
 sg13g2_dfrbp_1 _15572_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net1673),
    .D(_00011_),
    .Q_N(_07235_),
    .Q(\gpio_out_sel[3] ));
 sg13g2_dfrbp_1 _15573_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net1674),
    .D(net3743),
    .Q_N(_07236_),
    .Q(\gpio_out_sel[4] ));
 sg13g2_dfrbp_1 _15574_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net1675),
    .D(net3578),
    .Q_N(_07237_),
    .Q(\gpio_out_sel[5] ));
 sg13g2_dfrbp_1 _15575_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net1676),
    .D(net3567),
    .Q_N(_07238_),
    .Q(\gpio_out_sel[6] ));
 sg13g2_dfrbp_1 _15576_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net1677),
    .D(net3878),
    .Q_N(_07239_),
    .Q(\gpio_out_sel[7] ));
 sg13g2_dfrbp_1 _15577_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net1678),
    .D(net3634),
    .Q_N(_07240_),
    .Q(\gpio_out_sel[8] ));
 sg13g2_dfrbp_1 _15578_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net1679),
    .D(net3809),
    .Q_N(_07241_),
    .Q(\gpio_out_sel[9] ));
 sg13g2_dfrbp_1 _15579_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net1680),
    .D(_00000_),
    .Q_N(_07242_),
    .Q(\gpio_out[0] ));
 sg13g2_dfrbp_1 _15580_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net1681),
    .D(_00001_),
    .Q_N(_07243_),
    .Q(\gpio_out[1] ));
 sg13g2_dfrbp_1 _15581_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net1682),
    .D(_00002_),
    .Q_N(_07244_),
    .Q(\gpio_out[2] ));
 sg13g2_dfrbp_1 _15582_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net1683),
    .D(_00003_),
    .Q_N(_07245_),
    .Q(\gpio_out[3] ));
 sg13g2_dfrbp_1 _15583_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net1684),
    .D(_00004_),
    .Q_N(_07246_),
    .Q(\gpio_out[4] ));
 sg13g2_dfrbp_1 _15584_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net1685),
    .D(_00005_),
    .Q_N(_07247_),
    .Q(\gpio_out[5] ));
 sg13g2_dfrbp_1 _15585_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net1686),
    .D(_00006_),
    .Q_N(_07248_),
    .Q(\gpio_out[6] ));
 sg13g2_dfrbp_1 _15586_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net1687),
    .D(_00007_),
    .Q_N(_07249_),
    .Q(\gpio_out[7] ));
 sg13g2_dfrbp_1 _15587_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net1823),
    .D(net2),
    .Q_N(_07250_),
    .Q(\i_tinyqv.cpu.i_core.interrupt_req[0] ));
 sg13g2_dfrbp_1 _15588_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1521),
    .D(net3),
    .Q_N(_06253_),
    .Q(\i_tinyqv.cpu.i_core.interrupt_req[1] ));
 sg13g2_dfrbp_1 _15589_ (.CLK(net2378),
    .RESET_B(net1519),
    .D(net1),
    .Q_N(_00195_),
    .Q(\i_debug_uart_tx.resetn ));
 sg13g2_dfrbp_1 _15590_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net1517),
    .D(net3489),
    .Q_N(_06252_),
    .Q(\i_tinyqv.cpu.instr_data[0][2] ));
 sg13g2_dfrbp_1 _15591_ (.CLK(clknet_leaf_132_clk_regs),
    .RESET_B(net1515),
    .D(net3449),
    .Q_N(_06251_),
    .Q(\i_tinyqv.cpu.instr_data[0][3] ));
 sg13g2_dfrbp_1 _15592_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net1509),
    .D(net3061),
    .Q_N(_00143_),
    .Q(\i_tinyqv.cpu.instr_data[0][4] ));
 sg13g2_dfrbp_1 _15593_ (.CLK(clknet_leaf_149_clk_regs),
    .RESET_B(net1507),
    .D(net3109),
    .Q_N(_00147_),
    .Q(\i_tinyqv.cpu.instr_data[0][5] ));
 sg13g2_dfrbp_1 _15594_ (.CLK(clknet_leaf_149_clk_regs),
    .RESET_B(net1505),
    .D(net3122),
    .Q_N(_00151_),
    .Q(\i_tinyqv.cpu.instr_data[0][6] ));
 sg13g2_dfrbp_1 _15595_ (.CLK(clknet_leaf_148_clk_regs),
    .RESET_B(net1503),
    .D(net3071),
    .Q_N(_00168_),
    .Q(\i_tinyqv.cpu.instr_data[0][7] ));
 sg13g2_dfrbp_1 _15596_ (.CLK(clknet_leaf_148_clk_regs),
    .RESET_B(net1501),
    .D(net3177),
    .Q_N(_00172_),
    .Q(\i_tinyqv.cpu.instr_data[0][8] ));
 sg13g2_dfrbp_1 _15597_ (.CLK(clknet_leaf_147_clk_regs),
    .RESET_B(net1499),
    .D(net3055),
    .Q_N(_00176_),
    .Q(\i_tinyqv.cpu.instr_data[0][9] ));
 sg13g2_dfrbp_1 _15598_ (.CLK(clknet_leaf_150_clk_regs),
    .RESET_B(net1497),
    .D(net3145),
    .Q_N(_00180_),
    .Q(\i_tinyqv.cpu.instr_data[0][10] ));
 sg13g2_dfrbp_1 _15599_ (.CLK(clknet_leaf_147_clk_regs),
    .RESET_B(net1495),
    .D(net3098),
    .Q_N(_00188_),
    .Q(\i_tinyqv.cpu.instr_data[0][11] ));
 sg13g2_dfrbp_1 _15600_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net1493),
    .D(net3195),
    .Q_N(_00184_),
    .Q(\i_tinyqv.cpu.instr_data[0][12] ));
 sg13g2_dfrbp_1 _15601_ (.CLK(clknet_leaf_145_clk_regs),
    .RESET_B(net1491),
    .D(net3126),
    .Q_N(_00155_),
    .Q(\i_tinyqv.cpu.instr_data[0][13] ));
 sg13g2_dfrbp_1 _15602_ (.CLK(clknet_leaf_148_clk_regs),
    .RESET_B(net1489),
    .D(net3067),
    .Q_N(_00159_),
    .Q(\i_tinyqv.cpu.instr_data[0][14] ));
 sg13g2_dfrbp_1 _15603_ (.CLK(clknet_leaf_150_clk_regs),
    .RESET_B(net1487),
    .D(net3159),
    .Q_N(_00163_),
    .Q(\i_tinyqv.cpu.instr_data[0][15] ));
 sg13g2_dfrbp_1 _15604_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net1485),
    .D(net3718),
    .Q_N(_06250_),
    .Q(\i_tinyqv.cpu.instr_data[3][2] ));
 sg13g2_dfrbp_1 _15605_ (.CLK(clknet_leaf_147_clk_regs),
    .RESET_B(net1483),
    .D(net3378),
    .Q_N(_06249_),
    .Q(\i_tinyqv.cpu.instr_data[3][3] ));
 sg13g2_dfrbp_1 _15606_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net1481),
    .D(net3357),
    .Q_N(_00144_),
    .Q(\i_tinyqv.cpu.instr_data[3][4] ));
 sg13g2_dfrbp_1 _15607_ (.CLK(clknet_leaf_149_clk_regs),
    .RESET_B(net1479),
    .D(net2900),
    .Q_N(_00148_),
    .Q(\i_tinyqv.cpu.instr_data[3][5] ));
 sg13g2_dfrbp_1 _15608_ (.CLK(clknet_leaf_149_clk_regs),
    .RESET_B(net1477),
    .D(net3341),
    .Q_N(_00152_),
    .Q(\i_tinyqv.cpu.instr_data[3][6] ));
 sg13g2_dfrbp_1 _15609_ (.CLK(clknet_leaf_149_clk_regs),
    .RESET_B(net1475),
    .D(net3304),
    .Q_N(_00169_),
    .Q(\i_tinyqv.cpu.instr_data[3][7] ));
 sg13g2_dfrbp_1 _15610_ (.CLK(clknet_leaf_146_clk_regs),
    .RESET_B(net1473),
    .D(net2881),
    .Q_N(_00173_),
    .Q(\i_tinyqv.cpu.instr_data[3][8] ));
 sg13g2_dfrbp_1 _15611_ (.CLK(clknet_leaf_145_clk_regs),
    .RESET_B(net1471),
    .D(net2911),
    .Q_N(_00177_),
    .Q(\i_tinyqv.cpu.instr_data[3][9] ));
 sg13g2_dfrbp_1 _15612_ (.CLK(clknet_leaf_150_clk_regs),
    .RESET_B(net1469),
    .D(net2975),
    .Q_N(_00181_),
    .Q(\i_tinyqv.cpu.instr_data[3][10] ));
 sg13g2_dfrbp_1 _15613_ (.CLK(clknet_leaf_146_clk_regs),
    .RESET_B(net1467),
    .D(net2854),
    .Q_N(_00189_),
    .Q(\i_tinyqv.cpu.instr_data[3][11] ));
 sg13g2_dfrbp_1 _15614_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net1465),
    .D(net2898),
    .Q_N(_00185_),
    .Q(\i_tinyqv.cpu.instr_data[3][12] ));
 sg13g2_dfrbp_1 _15615_ (.CLK(clknet_leaf_146_clk_regs),
    .RESET_B(net1455),
    .D(net2888),
    .Q_N(_00156_),
    .Q(\i_tinyqv.cpu.instr_data[3][13] ));
 sg13g2_dfrbp_1 _15616_ (.CLK(clknet_leaf_148_clk_regs),
    .RESET_B(net1453),
    .D(net2921),
    .Q_N(_00160_),
    .Q(\i_tinyqv.cpu.instr_data[3][14] ));
 sg13g2_dfrbp_1 _15617_ (.CLK(clknet_leaf_150_clk_regs),
    .RESET_B(net1440),
    .D(net2951),
    .Q_N(_00164_),
    .Q(\i_tinyqv.cpu.instr_data[3][15] ));
 sg13g2_dfrbp_1 _15618_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net1437),
    .D(net3683),
    .Q_N(_00242_),
    .Q(\i_latch_mem.cycle[0] ));
 sg13g2_dfrbp_1 _15619_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net1435),
    .D(_01125_),
    .Q_N(_06248_),
    .Q(\i_spi.data[1] ));
 sg13g2_dfrbp_1 _15620_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net1433),
    .D(net3715),
    .Q_N(_06247_),
    .Q(\i_spi.data[2] ));
 sg13g2_dfrbp_1 _15621_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net1431),
    .D(net3681),
    .Q_N(_06246_),
    .Q(\i_spi.data[3] ));
 sg13g2_dfrbp_1 _15622_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net1410),
    .D(_01128_),
    .Q_N(_06245_),
    .Q(\i_spi.data[4] ));
 sg13g2_dfrbp_1 _15623_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net1408),
    .D(net3532),
    .Q_N(_06244_),
    .Q(\i_spi.data[5] ));
 sg13g2_dfrbp_1 _15624_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net1406),
    .D(_01130_),
    .Q_N(_06243_),
    .Q(\i_spi.data[6] ));
 sg13g2_dfrbp_1 _15625_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net1404),
    .D(net3286),
    .Q_N(_06242_),
    .Q(\i_spi.data[7] ));
 sg13g2_dfrbp_1 _15626_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net1402),
    .D(_01132_),
    .Q_N(_06241_),
    .Q(\addr[24] ));
 sg13g2_dfrbp_1 _15627_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net1398),
    .D(_01133_),
    .Q_N(_06240_),
    .Q(\addr[25] ));
 sg13g2_dfrbp_1 _15628_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net1394),
    .D(_01134_),
    .Q_N(_06239_),
    .Q(\addr[26] ));
 sg13g2_dfrbp_1 _15629_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net1390),
    .D(_01135_),
    .Q_N(_00191_),
    .Q(\addr[27] ));
 sg13g2_dfrbp_1 _15630_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net1386),
    .D(_01136_),
    .Q_N(_06238_),
    .Q(\addr[0] ));
 sg13g2_dfrbp_1 _15631_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net1384),
    .D(_01137_),
    .Q_N(_06237_),
    .Q(\addr[1] ));
 sg13g2_dfrbp_1 _15632_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net1382),
    .D(_01138_),
    .Q_N(_06236_),
    .Q(\addr[2] ));
 sg13g2_dfrbp_1 _15633_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net1380),
    .D(_01139_),
    .Q_N(_00198_),
    .Q(\addr[3] ));
 sg13g2_dfrbp_1 _15634_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net1378),
    .D(_01140_),
    .Q_N(_06235_),
    .Q(\addr[4] ));
 sg13g2_dfrbp_1 _15635_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net1375),
    .D(_01141_),
    .Q_N(_06234_),
    .Q(\addr[5] ));
 sg13g2_dfrbp_1 _15636_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net1373),
    .D(_01142_),
    .Q_N(_06233_),
    .Q(\addr[6] ));
 sg13g2_dfrbp_1 _15637_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net1371),
    .D(net3330),
    .Q_N(_06232_),
    .Q(\addr[7] ));
 sg13g2_dfrbp_1 _15638_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net1369),
    .D(_01144_),
    .Q_N(_06231_),
    .Q(\addr[8] ));
 sg13g2_dfrbp_1 _15639_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net1366),
    .D(_01145_),
    .Q_N(_06230_),
    .Q(\addr[9] ));
 sg13g2_dfrbp_1 _15640_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1364),
    .D(_01146_),
    .Q_N(_06229_),
    .Q(\addr[10] ));
 sg13g2_dfrbp_1 _15641_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net1362),
    .D(net3605),
    .Q_N(_06228_),
    .Q(\addr[11] ));
 sg13g2_dfrbp_1 _15642_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1360),
    .D(_01148_),
    .Q_N(_06227_),
    .Q(\addr[12] ));
 sg13g2_dfrbp_1 _15643_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1356),
    .D(net3711),
    .Q_N(_06226_),
    .Q(\addr[13] ));
 sg13g2_dfrbp_1 _15644_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1354),
    .D(_01150_),
    .Q_N(_06225_),
    .Q(\addr[14] ));
 sg13g2_dfrbp_1 _15645_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1352),
    .D(net3617),
    .Q_N(_06224_),
    .Q(\addr[15] ));
 sg13g2_dfrbp_1 _15646_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net1350),
    .D(_01152_),
    .Q_N(_06223_),
    .Q(\addr[16] ));
 sg13g2_dfrbp_1 _15647_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net1348),
    .D(_01153_),
    .Q_N(_06222_),
    .Q(\addr[17] ));
 sg13g2_dfrbp_1 _15648_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net1346),
    .D(_01154_),
    .Q_N(_06221_),
    .Q(\addr[18] ));
 sg13g2_dfrbp_1 _15649_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net1344),
    .D(_01155_),
    .Q_N(_06220_),
    .Q(\addr[19] ));
 sg13g2_dfrbp_1 _15650_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net1342),
    .D(net3497),
    .Q_N(_06219_),
    .Q(\addr[20] ));
 sg13g2_dfrbp_1 _15651_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net1340),
    .D(_01157_),
    .Q_N(_06218_),
    .Q(\addr[21] ));
 sg13g2_dfrbp_1 _15652_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net1338),
    .D(_01158_),
    .Q_N(_06217_),
    .Q(\addr[22] ));
 sg13g2_dfrbp_1 _15653_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net1328),
    .D(_01159_),
    .Q_N(_00201_),
    .Q(\addr[23] ));
 sg13g2_dfrbp_1 _15654_ (.CLK(clknet_leaf_130_clk_regs),
    .RESET_B(net1326),
    .D(net3419),
    .Q_N(_06216_),
    .Q(\i_tinyqv.cpu.instr_data[1][2] ));
 sg13g2_dfrbp_1 _15655_ (.CLK(clknet_leaf_147_clk_regs),
    .RESET_B(net1324),
    .D(net3464),
    .Q_N(_06215_),
    .Q(\i_tinyqv.cpu.instr_data[1][3] ));
 sg13g2_dfrbp_1 _15656_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net1322),
    .D(net3057),
    .Q_N(_00142_),
    .Q(\i_tinyqv.cpu.instr_data[1][4] ));
 sg13g2_dfrbp_1 _15657_ (.CLK(clknet_leaf_149_clk_regs),
    .RESET_B(net1320),
    .D(net3198),
    .Q_N(_00146_),
    .Q(\i_tinyqv.cpu.instr_data[1][5] ));
 sg13g2_dfrbp_1 _15658_ (.CLK(clknet_leaf_131_clk_regs),
    .RESET_B(net1318),
    .D(net3059),
    .Q_N(_00150_),
    .Q(\i_tinyqv.cpu.instr_data[1][6] ));
 sg13g2_dfrbp_1 _15659_ (.CLK(clknet_leaf_148_clk_regs),
    .RESET_B(net1315),
    .D(net3069),
    .Q_N(_00167_),
    .Q(\i_tinyqv.cpu.instr_data[1][7] ));
 sg13g2_dfrbp_1 _15660_ (.CLK(clknet_leaf_145_clk_regs),
    .RESET_B(net1313),
    .D(net3080),
    .Q_N(_00171_),
    .Q(\i_tinyqv.cpu.instr_data[1][8] ));
 sg13g2_dfrbp_1 _15661_ (.CLK(clknet_leaf_145_clk_regs),
    .RESET_B(net1295),
    .D(net3018),
    .Q_N(_00175_),
    .Q(\i_tinyqv.cpu.instr_data[1][9] ));
 sg13g2_dfrbp_1 _15662_ (.CLK(clknet_leaf_150_clk_regs),
    .RESET_B(net1293),
    .D(net3129),
    .Q_N(_00179_),
    .Q(\i_tinyqv.cpu.instr_data[1][10] ));
 sg13g2_dfrbp_1 _15663_ (.CLK(clknet_leaf_147_clk_regs),
    .RESET_B(net1291),
    .D(net3148),
    .Q_N(_00187_),
    .Q(\i_tinyqv.cpu.instr_data[1][11] ));
 sg13g2_dfrbp_1 _15664_ (.CLK(clknet_leaf_148_clk_regs),
    .RESET_B(net1289),
    .D(net3119),
    .Q_N(_00183_),
    .Q(\i_tinyqv.cpu.instr_data[1][12] ));
 sg13g2_dfrbp_1 _15665_ (.CLK(clknet_leaf_145_clk_regs),
    .RESET_B(net1287),
    .D(net3034),
    .Q_N(_00154_),
    .Q(\i_tinyqv.cpu.instr_data[1][13] ));
 sg13g2_dfrbp_1 _15666_ (.CLK(clknet_leaf_150_clk_regs),
    .RESET_B(net1285),
    .D(net3151),
    .Q_N(_00158_),
    .Q(\i_tinyqv.cpu.instr_data[1][14] ));
 sg13g2_dfrbp_1 _15667_ (.CLK(clknet_leaf_150_clk_regs),
    .RESET_B(net1283),
    .D(net3190),
    .Q_N(_00162_),
    .Q(\i_tinyqv.cpu.instr_data[1][15] ));
 sg13g2_dfrbp_1 _15668_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1281),
    .D(net3738),
    .Q_N(_00206_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[0] ));
 sg13g2_dfrbp_1 _15669_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1279),
    .D(net3924),
    .Q_N(_00237_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[1] ));
 sg13g2_dfrbp_1 _15670_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net1277),
    .D(net3919),
    .Q_N(_00235_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[2] ));
 sg13g2_dfrbp_1 _15671_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1275),
    .D(net3913),
    .Q_N(_00209_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[3] ));
 sg13g2_dfrbp_1 _15672_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net1273),
    .D(net4036),
    .Q_N(_00211_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[4] ));
 sg13g2_dfrbp_1 _15673_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net1271),
    .D(net4065),
    .Q_N(_00213_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[5] ));
 sg13g2_dfrbp_1 _15674_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net1269),
    .D(_01180_),
    .Q_N(_00215_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[6] ));
 sg13g2_dfrbp_1 _15675_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net1267),
    .D(net4072),
    .Q_N(_00217_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[7] ));
 sg13g2_dfrbp_1 _15676_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net1265),
    .D(net4020),
    .Q_N(_00219_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[8] ));
 sg13g2_dfrbp_1 _15677_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net1262),
    .D(net4038),
    .Q_N(_00221_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[9] ));
 sg13g2_dfrbp_1 _15678_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net1260),
    .D(net3965),
    .Q_N(_00223_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[10] ));
 sg13g2_dfrbp_1 _15679_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net1258),
    .D(net3953),
    .Q_N(_00225_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[11] ));
 sg13g2_dfrbp_1 _15680_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net1256),
    .D(net3440),
    .Q_N(_00227_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[12] ));
 sg13g2_dfrbp_1 _15681_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net1254),
    .D(net3685),
    .Q_N(_00229_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[13] ));
 sg13g2_dfrbp_1 _15682_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net1252),
    .D(net3408),
    .Q_N(_00231_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[14] ));
 sg13g2_dfrbp_1 _15683_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net1250),
    .D(net3466),
    .Q_N(_00233_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[15] ));
 sg13g2_dfrbp_1 _15684_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net1248),
    .D(net3406),
    .Q_N(_00232_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[16] ));
 sg13g2_dfrbp_1 _15685_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net1246),
    .D(net3669),
    .Q_N(_00230_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[17] ));
 sg13g2_dfrbp_1 _15686_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net1244),
    .D(_01192_),
    .Q_N(_00228_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[18] ));
 sg13g2_dfrbp_1 _15687_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net1242),
    .D(_01193_),
    .Q_N(_00226_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[19] ));
 sg13g2_dfrbp_1 _15688_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net1240),
    .D(_01194_),
    .Q_N(_00224_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[20] ));
 sg13g2_dfrbp_1 _15689_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net1238),
    .D(_01195_),
    .Q_N(_00222_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[21] ));
 sg13g2_dfrbp_1 _15690_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net1236),
    .D(net3539),
    .Q_N(_00220_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[22] ));
 sg13g2_dfrbp_1 _15691_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net1234),
    .D(_01197_),
    .Q_N(_00218_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[23] ));
 sg13g2_dfrbp_1 _15692_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net1232),
    .D(net3481),
    .Q_N(_00216_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[24] ));
 sg13g2_dfrbp_1 _15693_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net1230),
    .D(_01199_),
    .Q_N(_00214_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[25] ));
 sg13g2_dfrbp_1 _15694_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1228),
    .D(_01200_),
    .Q_N(_00212_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[26] ));
 sg13g2_dfrbp_1 _15695_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net1226),
    .D(_01201_),
    .Q_N(_00210_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[27] ));
 sg13g2_dfrbp_1 _15696_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net1224),
    .D(_01202_),
    .Q_N(_00236_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[30] ));
 sg13g2_dfrbp_1 _15697_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1222),
    .D(_01203_),
    .Q_N(_00238_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[31] ));
 sg13g2_dfrbp_1 _15698_ (.CLK(clknet_leaf_141_clk_regs),
    .RESET_B(net1219),
    .D(net3898),
    .Q_N(_06214_),
    .Q(\i_tinyqv.cpu.instr_data[0][0] ));
 sg13g2_dfrbp_1 _15699_ (.CLK(clknet_leaf_147_clk_regs),
    .RESET_B(net1217),
    .D(_01205_),
    .Q_N(_00139_),
    .Q(\i_tinyqv.cpu.instr_data[0][1] ));
 sg13g2_dfrbp_1 _15700_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net1215),
    .D(net3509),
    .Q_N(_06213_),
    .Q(\i_tinyqv.cpu.i_core.mepc[0] ));
 sg13g2_dfrbp_1 _15701_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net1214),
    .D(_01207_),
    .Q_N(_06212_),
    .Q(\i_tinyqv.cpu.i_core.mepc[1] ));
 sg13g2_dfrbp_1 _15702_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net1213),
    .D(net3624),
    .Q_N(_06211_),
    .Q(\i_tinyqv.cpu.i_core.mepc[2] ));
 sg13g2_dfrbp_1 _15703_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net1212),
    .D(net3720),
    .Q_N(_06210_),
    .Q(\i_tinyqv.cpu.i_core.mepc[3] ));
 sg13g2_dfrbp_1 _15704_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1211),
    .D(_01210_),
    .Q_N(_06209_),
    .Q(\i_tinyqv.cpu.i_core.mepc[4] ));
 sg13g2_dfrbp_1 _15705_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net1210),
    .D(_01211_),
    .Q_N(_06208_),
    .Q(\i_tinyqv.cpu.i_core.mepc[5] ));
 sg13g2_dfrbp_1 _15706_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net1209),
    .D(_01212_),
    .Q_N(_06207_),
    .Q(\i_tinyqv.cpu.i_core.mepc[6] ));
 sg13g2_dfrbp_1 _15707_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net1208),
    .D(net3628),
    .Q_N(_06206_),
    .Q(\i_tinyqv.cpu.i_core.mepc[7] ));
 sg13g2_dfrbp_1 _15708_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1207),
    .D(net3547),
    .Q_N(_06205_),
    .Q(\i_tinyqv.cpu.i_core.mepc[8] ));
 sg13g2_dfrbp_1 _15709_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net1206),
    .D(_01215_),
    .Q_N(_06204_),
    .Q(\i_tinyqv.cpu.i_core.mepc[9] ));
 sg13g2_dfrbp_1 _15710_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net1205),
    .D(_01216_),
    .Q_N(_06203_),
    .Q(\i_tinyqv.cpu.i_core.mepc[10] ));
 sg13g2_dfrbp_1 _15711_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net1204),
    .D(_01217_),
    .Q_N(_06202_),
    .Q(\i_tinyqv.cpu.i_core.mepc[11] ));
 sg13g2_dfrbp_1 _15712_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net1203),
    .D(_01218_),
    .Q_N(_06201_),
    .Q(\i_tinyqv.cpu.i_core.mepc[12] ));
 sg13g2_dfrbp_1 _15713_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net1202),
    .D(net3499),
    .Q_N(_06200_),
    .Q(\i_tinyqv.cpu.i_core.mepc[13] ));
 sg13g2_dfrbp_1 _15714_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net1201),
    .D(net3530),
    .Q_N(_06199_),
    .Q(\i_tinyqv.cpu.i_core.mepc[14] ));
 sg13g2_dfrbp_1 _15715_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net1200),
    .D(_01221_),
    .Q_N(_06198_),
    .Q(\i_tinyqv.cpu.i_core.mepc[15] ));
 sg13g2_dfrbp_1 _15716_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1199),
    .D(net3541),
    .Q_N(_06197_),
    .Q(\i_tinyqv.cpu.i_core.mepc[16] ));
 sg13g2_dfrbp_1 _15717_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net1198),
    .D(net3580),
    .Q_N(_06196_),
    .Q(\i_tinyqv.cpu.i_core.mepc[17] ));
 sg13g2_dfrbp_1 _15718_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net1197),
    .D(_01224_),
    .Q_N(_06195_),
    .Q(\i_tinyqv.cpu.i_core.mepc[18] ));
 sg13g2_dfrbp_1 _15719_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net1196),
    .D(_01225_),
    .Q_N(_06194_),
    .Q(\i_tinyqv.cpu.i_core.mepc[19] ));
 sg13g2_dfrbp_1 _15720_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net1194),
    .D(_01226_),
    .Q_N(_06193_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ));
 sg13g2_dfrbp_1 _15721_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net1191),
    .D(_01227_),
    .Q_N(_06192_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ));
 sg13g2_dfrbp_1 _15722_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net1189),
    .D(_01228_),
    .Q_N(_06191_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[2] ));
 sg13g2_dfrbp_1 _15723_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net1824),
    .D(_01229_),
    .Q_N(_07251_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[3] ));
 sg13g2_dfrbp_1 _15724_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1825),
    .D(_00019_),
    .Q_N(_07252_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[0] ));
 sg13g2_dfrbp_1 _15725_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net1826),
    .D(_00022_),
    .Q_N(_07253_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[1] ));
 sg13g2_dfrbp_1 _15726_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net1827),
    .D(_00023_),
    .Q_N(_07254_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[2] ));
 sg13g2_dfrbp_1 _15727_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net1828),
    .D(_00024_),
    .Q_N(_07255_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[3] ));
 sg13g2_dfrbp_1 _15728_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net1829),
    .D(_00025_),
    .Q_N(_07256_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[4] ));
 sg13g2_dfrbp_1 _15729_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net1830),
    .D(_00026_),
    .Q_N(_07257_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[5] ));
 sg13g2_dfrbp_1 _15730_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net1831),
    .D(_00027_),
    .Q_N(_07258_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[6] ));
 sg13g2_dfrbp_1 _15731_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net1832),
    .D(_00028_),
    .Q_N(_07259_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[7] ));
 sg13g2_dfrbp_1 _15732_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net1833),
    .D(_00029_),
    .Q_N(_07260_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[8] ));
 sg13g2_dfrbp_1 _15733_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net1834),
    .D(_00030_),
    .Q_N(_07261_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[9] ));
 sg13g2_dfrbp_1 _15734_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net1836),
    .D(_00020_),
    .Q_N(_07262_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[10] ));
 sg13g2_dfrbp_1 _15735_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net1187),
    .D(_00021_),
    .Q_N(_06190_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[11] ));
 sg13g2_dfrbp_1 _15736_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net2020),
    .D(net3350),
    .Q_N(_07263_),
    .Q(\i_tinyqv.mem.data_stall ));
 sg13g2_dfrbp_1 _15737_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net1185),
    .D(net3855),
    .Q_N(_00192_),
    .Q(\i_tinyqv.mem.qspi_write_done ));
 sg13g2_dfrbp_1 _15738_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net1181),
    .D(_01231_),
    .Q_N(_06189_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[12] ));
 sg13g2_dfrbp_1 _15739_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net1179),
    .D(_01232_),
    .Q_N(_06188_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[13] ));
 sg13g2_dfrbp_1 _15740_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net1177),
    .D(_01233_),
    .Q_N(_06187_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[14] ));
 sg13g2_dfrbp_1 _15741_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net1175),
    .D(_01234_),
    .Q_N(_06186_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[15] ));
 sg13g2_dfrbp_1 _15742_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net1173),
    .D(_01235_),
    .Q_N(_00196_),
    .Q(\i_tinyqv.mem.qspi_data_byte_idx[0] ));
 sg13g2_dfrbp_1 _15743_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net1169),
    .D(_01236_),
    .Q_N(_06185_),
    .Q(\i_tinyqv.mem.qspi_data_byte_idx[1] ));
 sg13g2_dfrbp_1 _15744_ (.CLK(clknet_leaf_140_clk_regs),
    .RESET_B(net1165),
    .D(_01237_),
    .Q_N(_06184_),
    .Q(\i_tinyqv.cpu.instr_data_in[0] ));
 sg13g2_dfrbp_1 _15745_ (.CLK(clknet_leaf_140_clk_regs),
    .RESET_B(net1163),
    .D(_01238_),
    .Q_N(_06183_),
    .Q(\i_tinyqv.cpu.instr_data_in[1] ));
 sg13g2_dfrbp_1 _15746_ (.CLK(clknet_leaf_140_clk_regs),
    .RESET_B(net1156),
    .D(_01239_),
    .Q_N(_06182_),
    .Q(\i_tinyqv.cpu.instr_data_in[2] ));
 sg13g2_dfrbp_1 _15747_ (.CLK(clknet_leaf_146_clk_regs),
    .RESET_B(net1154),
    .D(_01240_),
    .Q_N(_06181_),
    .Q(\i_tinyqv.cpu.instr_data_in[3] ));
 sg13g2_dfrbp_1 _15748_ (.CLK(clknet_leaf_139_clk_regs),
    .RESET_B(net1152),
    .D(net3789),
    .Q_N(_06180_),
    .Q(\i_tinyqv.cpu.instr_data_in[4] ));
 sg13g2_dfrbp_1 _15749_ (.CLK(clknet_leaf_140_clk_regs),
    .RESET_B(net1150),
    .D(net3787),
    .Q_N(_06179_),
    .Q(\i_tinyqv.cpu.instr_data_in[5] ));
 sg13g2_dfrbp_1 _15750_ (.CLK(clknet_leaf_140_clk_regs),
    .RESET_B(net1148),
    .D(net3948),
    .Q_N(_06178_),
    .Q(\i_tinyqv.cpu.instr_data_in[6] ));
 sg13g2_dfrbp_1 _15751_ (.CLK(clknet_leaf_140_clk_regs),
    .RESET_B(net1146),
    .D(net3936),
    .Q_N(_06177_),
    .Q(\i_tinyqv.cpu.instr_data_in[7] ));
 sg13g2_dfrbp_1 _15752_ (.CLK(clknet_leaf_139_clk_regs),
    .RESET_B(net1144),
    .D(_01245_),
    .Q_N(_06176_),
    .Q(\i_tinyqv.mem.qspi_data_buf[8] ));
 sg13g2_dfrbp_1 _15753_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net1142),
    .D(_01246_),
    .Q_N(_06175_),
    .Q(\i_tinyqv.mem.qspi_data_buf[9] ));
 sg13g2_dfrbp_1 _15754_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net1140),
    .D(_01247_),
    .Q_N(_06174_),
    .Q(\i_tinyqv.mem.qspi_data_buf[10] ));
 sg13g2_dfrbp_1 _15755_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net1137),
    .D(net3367),
    .Q_N(_06173_),
    .Q(\i_tinyqv.mem.qspi_data_buf[11] ));
 sg13g2_dfrbp_1 _15756_ (.CLK(clknet_leaf_139_clk_regs),
    .RESET_B(net1135),
    .D(_01249_),
    .Q_N(_06172_),
    .Q(\i_tinyqv.mem.qspi_data_buf[12] ));
 sg13g2_dfrbp_1 _15757_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net1133),
    .D(net3359),
    .Q_N(_06171_),
    .Q(\i_tinyqv.mem.qspi_data_buf[13] ));
 sg13g2_dfrbp_1 _15758_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net1131),
    .D(net3413),
    .Q_N(_06170_),
    .Q(\i_tinyqv.mem.qspi_data_buf[14] ));
 sg13g2_dfrbp_1 _15759_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net715),
    .D(net3411),
    .Q_N(_06169_),
    .Q(\i_tinyqv.mem.qspi_data_buf[15] ));
 sg13g2_dfrbp_1 _15760_ (.CLK(clknet_leaf_146_clk_regs),
    .RESET_B(net713),
    .D(net3309),
    .Q_N(_06168_),
    .Q(\i_tinyqv.mem.data_from_read[16] ));
 sg13g2_dfrbp_1 _15761_ (.CLK(clknet_leaf_145_clk_regs),
    .RESET_B(net711),
    .D(net2989),
    .Q_N(_06167_),
    .Q(\i_tinyqv.mem.data_from_read[17] ));
 sg13g2_dfrbp_1 _15762_ (.CLK(clknet_leaf_144_clk_regs),
    .RESET_B(net681),
    .D(net3155),
    .Q_N(_06166_),
    .Q(\i_tinyqv.mem.data_from_read[18] ));
 sg13g2_dfrbp_1 _15763_ (.CLK(clknet_leaf_146_clk_regs),
    .RESET_B(net679),
    .D(net3361),
    .Q_N(_06165_),
    .Q(\i_tinyqv.mem.data_from_read[19] ));
 sg13g2_dfrbp_1 _15764_ (.CLK(clknet_leaf_142_clk_regs),
    .RESET_B(net2095),
    .D(net2997),
    .Q_N(_06164_),
    .Q(\i_tinyqv.mem.data_from_read[20] ));
 sg13g2_dfrbp_1 _15765_ (.CLK(clknet_leaf_142_clk_regs),
    .RESET_B(net2093),
    .D(net3093),
    .Q_N(_06163_),
    .Q(\i_tinyqv.mem.data_from_read[21] ));
 sg13g2_dfrbp_1 _15766_ (.CLK(clknet_leaf_145_clk_regs),
    .RESET_B(net2091),
    .D(net3078),
    .Q_N(_06162_),
    .Q(\i_tinyqv.mem.data_from_read[22] ));
 sg13g2_dfrbp_1 _15767_ (.CLK(clknet_leaf_141_clk_regs),
    .RESET_B(net2089),
    .D(net3332),
    .Q_N(_06161_),
    .Q(\i_tinyqv.mem.data_from_read[23] ));
 sg13g2_dfrbp_1 _15768_ (.CLK(clknet_leaf_141_clk_regs),
    .RESET_B(net2087),
    .D(_01261_),
    .Q_N(_06160_),
    .Q(\i_tinyqv.mem.qspi_data_buf[24] ));
 sg13g2_dfrbp_1 _15769_ (.CLK(clknet_leaf_141_clk_regs),
    .RESET_B(net2085),
    .D(_01262_),
    .Q_N(_06159_),
    .Q(\i_tinyqv.mem.qspi_data_buf[25] ));
 sg13g2_dfrbp_1 _15770_ (.CLK(clknet_leaf_146_clk_regs),
    .RESET_B(net2083),
    .D(_01263_),
    .Q_N(_06158_),
    .Q(\i_tinyqv.mem.qspi_data_buf[26] ));
 sg13g2_dfrbp_1 _15771_ (.CLK(clknet_leaf_141_clk_regs),
    .RESET_B(net2081),
    .D(_01264_),
    .Q_N(_06157_),
    .Q(\i_tinyqv.mem.qspi_data_buf[27] ));
 sg13g2_dfrbp_1 _15772_ (.CLK(clknet_leaf_142_clk_regs),
    .RESET_B(net2079),
    .D(_01265_),
    .Q_N(_06156_),
    .Q(\i_tinyqv.mem.qspi_data_buf[28] ));
 sg13g2_dfrbp_1 _15773_ (.CLK(clknet_leaf_141_clk_regs),
    .RESET_B(net2077),
    .D(_01266_),
    .Q_N(_06155_),
    .Q(\i_tinyqv.mem.qspi_data_buf[29] ));
 sg13g2_dfrbp_1 _15774_ (.CLK(clknet_leaf_142_clk_regs),
    .RESET_B(net2075),
    .D(_01267_),
    .Q_N(_06154_),
    .Q(\i_tinyqv.mem.qspi_data_buf[30] ));
 sg13g2_dfrbp_1 _15775_ (.CLK(clknet_leaf_146_clk_regs),
    .RESET_B(net2073),
    .D(_01268_),
    .Q_N(_06153_),
    .Q(\i_tinyqv.mem.qspi_data_buf[31] ));
 sg13g2_dfrbp_1 _15776_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net2071),
    .D(_01269_),
    .Q_N(_06152_),
    .Q(\i_tinyqv.cpu.instr_fetch_started ));
 sg13g2_dfrbp_1 _15777_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net2069),
    .D(_01270_),
    .Q_N(_00133_),
    .Q(\i_tinyqv.mem.instr_active ));
 sg13g2_dfrbp_1 _15778_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net2065),
    .D(_01271_),
    .Q_N(_06151_),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ));
 sg13g2_dfrbp_1 _15779_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net2063),
    .D(_01272_),
    .Q_N(_06150_),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ));
 sg13g2_dfrbp_1 _15780_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net2061),
    .D(net3901),
    .Q_N(_06149_),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ));
 sg13g2_dfrbp_1 _15781_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net2059),
    .D(_01274_),
    .Q_N(_06148_),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ));
 sg13g2_dfrbp_1 _15782_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net2057),
    .D(_01275_),
    .Q_N(_06147_),
    .Q(\i_tinyqv.mem.q_ctrl.data_req ));
 sg13g2_dfrbp_1 _15783_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net2055),
    .D(_01276_),
    .Q_N(_00199_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_clk_pos ));
 sg13g2_dfrbp_1 _15784_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net2051),
    .D(_01277_),
    .Q_N(_06146_),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ));
 sg13g2_dfrbp_1 _15785_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net2047),
    .D(_01278_),
    .Q_N(_06145_),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ));
 sg13g2_dfrbp_1 _15786_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net2043),
    .D(_01279_),
    .Q_N(_06144_),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ));
 sg13g2_dfrbp_1 _15787_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net2039),
    .D(_01280_),
    .Q_N(_00200_),
    .Q(\i_tinyqv.mem.q_ctrl.is_writing ));
 sg13g2_dfrbp_1 _15788_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net2035),
    .D(_01281_),
    .Q_N(_06143_),
    .Q(\i_tinyqv.mem.q_ctrl.data_ready ));
 sg13g2_dfrbp_1 _15789_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net2033),
    .D(_01282_),
    .Q_N(_00253_),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[0] ));
 sg13g2_dfrbp_1 _15790_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net2029),
    .D(_01283_),
    .Q_N(_06142_),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[1] ));
 sg13g2_dfrbp_1 _15791_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net2025),
    .D(_01284_),
    .Q_N(_00193_),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[2] ));
 sg13g2_dfrbp_1 _15792_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net2021),
    .D(_01285_),
    .Q_N(_06141_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ));
 sg13g2_dfrbp_1 _15793_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net2016),
    .D(_01286_),
    .Q_N(_06140_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _15794_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net2012),
    .D(_01287_),
    .Q_N(_06139_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _15795_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net2008),
    .D(_01288_),
    .Q_N(_06138_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ));
 sg13g2_dfrbp_1 _15796_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net2004),
    .D(_01289_),
    .Q_N(_00208_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[28] ));
 sg13g2_dfrbp_1 _15797_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net2000),
    .D(_01290_),
    .Q_N(_00234_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[29] ));
 sg13g2_dfrbp_1 _15798_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net1996),
    .D(net3271),
    .Q_N(_06137_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ));
 sg13g2_dfrbp_1 _15799_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net1994),
    .D(net3250),
    .Q_N(_06136_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ));
 sg13g2_dfrbp_1 _15800_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net1992),
    .D(net3344),
    .Q_N(_06135_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ));
 sg13g2_dfrbp_1 _15801_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net1990),
    .D(net3264),
    .Q_N(_06134_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ));
 sg13g2_dfrbp_1 _15802_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net1988),
    .D(_01295_),
    .Q_N(_00245_),
    .Q(\i_tinyqv.cpu.instr_data_in[8] ));
 sg13g2_dfrbp_1 _15803_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net1986),
    .D(_01296_),
    .Q_N(_00246_),
    .Q(\i_tinyqv.cpu.instr_data_in[9] ));
 sg13g2_dfrbp_1 _15804_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net1984),
    .D(_01297_),
    .Q_N(_00247_),
    .Q(\i_tinyqv.cpu.instr_data_in[10] ));
 sg13g2_dfrbp_1 _15805_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net1982),
    .D(_01298_),
    .Q_N(_00248_),
    .Q(\i_tinyqv.cpu.instr_data_in[11] ));
 sg13g2_dfrbp_1 _15806_ (.CLK(clknet_leaf_139_clk_regs),
    .RESET_B(net1980),
    .D(_01299_),
    .Q_N(_00249_),
    .Q(\i_tinyqv.cpu.instr_data_in[12] ));
 sg13g2_dfrbp_1 _15807_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net1978),
    .D(_01300_),
    .Q_N(_00250_),
    .Q(\i_tinyqv.cpu.instr_data_in[13] ));
 sg13g2_dfrbp_1 _15808_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net1976),
    .D(_01301_),
    .Q_N(_00251_),
    .Q(\i_tinyqv.cpu.instr_data_in[14] ));
 sg13g2_dfrbp_1 _15809_ (.CLK(clknet_leaf_142_clk_regs),
    .RESET_B(net1974),
    .D(_01302_),
    .Q_N(_00252_),
    .Q(\i_tinyqv.cpu.instr_data_in[15] ));
 sg13g2_dfrbp_1 _15810_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1972),
    .D(_01303_),
    .Q_N(_06133_),
    .Q(\i_tinyqv.mem.q_ctrl.last_ram_b_sel ));
 sg13g2_dfrbp_1 _15811_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net1970),
    .D(_01304_),
    .Q_N(_06132_),
    .Q(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ));
 sg13g2_dfrbp_1 _15812_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net1968),
    .D(_01305_),
    .Q_N(_06131_),
    .Q(\i_tinyqv.cpu.instr_fetch_stopped ));
 sg13g2_dfrbp_1 _15813_ (.CLK(net2379),
    .RESET_B(net1966),
    .D(\i_tinyqv.mem.q_ctrl.spi_clk_pos ),
    .Q_N(_06130_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_clk_neg ));
 sg13g2_dfrbp_1 _15814_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net1964),
    .D(_01306_),
    .Q_N(_06129_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_clk_use_neg ));
 sg13g2_dfrbp_1 _15815_ (.CLK(clknet_leaf_140_clk_regs),
    .RESET_B(net1962),
    .D(net3805),
    .Q_N(_06128_),
    .Q(\i_tinyqv.cpu.instr_data[2][0] ));
 sg13g2_dfrbp_1 _15816_ (.CLK(clknet_leaf_132_clk_regs),
    .RESET_B(net1958),
    .D(net3690),
    .Q_N(_00141_),
    .Q(\i_tinyqv.cpu.instr_data[2][1] ));
 sg13g2_dfrbp_1 _15817_ (.CLK(clknet_leaf_141_clk_regs),
    .RESET_B(net1954),
    .D(net3876),
    .Q_N(_06127_),
    .Q(\i_tinyqv.cpu.instr_data[1][0] ));
 sg13g2_dfrbp_1 _15818_ (.CLK(clknet_leaf_147_clk_regs),
    .RESET_B(net1950),
    .D(_01310_),
    .Q_N(_00138_),
    .Q(\i_tinyqv.cpu.instr_data[1][1] ));
 sg13g2_dfrbp_1 _15819_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net1946),
    .D(_01311_),
    .Q_N(_00131_),
    .Q(\i_tinyqv.cpu.instr_write_offset[1] ));
 sg13g2_dfrbp_1 _15820_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net1944),
    .D(_01312_),
    .Q_N(_00197_),
    .Q(\i_tinyqv.cpu.instr_write_offset[2] ));
 sg13g2_dfrbp_1 _15821_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net1942),
    .D(net3280),
    .Q_N(_06126_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[1] ));
 sg13g2_dfrbp_1 _15822_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net1938),
    .D(_01314_),
    .Q_N(_06125_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[2] ));
 sg13g2_dfrbp_1 _15823_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net1934),
    .D(_01315_),
    .Q_N(_06124_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[3] ));
 sg13g2_dfrbp_1 _15824_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net1930),
    .D(_01316_),
    .Q_N(_06123_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[4] ));
 sg13g2_dfrbp_1 _15825_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net1928),
    .D(_01317_),
    .Q_N(_06122_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[5] ));
 sg13g2_dfrbp_1 _15826_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net1926),
    .D(net3458),
    .Q_N(_06121_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[6] ));
 sg13g2_dfrbp_1 _15827_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1924),
    .D(net3551),
    .Q_N(_06120_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[7] ));
 sg13g2_dfrbp_1 _15828_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net1922),
    .D(net3471),
    .Q_N(_06119_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[8] ));
 sg13g2_dfrbp_1 _15829_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net1920),
    .D(net3347),
    .Q_N(_06118_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[9] ));
 sg13g2_dfrbp_1 _15830_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1918),
    .D(net3713),
    .Q_N(_06117_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[10] ));
 sg13g2_dfrbp_1 _15831_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net1916),
    .D(net3020),
    .Q_N(_06116_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[11] ));
 sg13g2_dfrbp_1 _15832_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1914),
    .D(net3442),
    .Q_N(_06115_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[12] ));
 sg13g2_dfrbp_1 _15833_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net1912),
    .D(net3380),
    .Q_N(_06114_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[13] ));
 sg13g2_dfrbp_1 _15834_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net1910),
    .D(net3254),
    .Q_N(_06113_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[14] ));
 sg13g2_dfrbp_1 _15835_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net1908),
    .D(net3355),
    .Q_N(_06112_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[15] ));
 sg13g2_dfrbp_1 _15836_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net1906),
    .D(net3501),
    .Q_N(_06111_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[16] ));
 sg13g2_dfrbp_1 _15837_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net1904),
    .D(net3469),
    .Q_N(_06110_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[17] ));
 sg13g2_dfrbp_1 _15838_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net1902),
    .D(net3320),
    .Q_N(_06109_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[18] ));
 sg13g2_dfrbp_1 _15839_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net1900),
    .D(net3322),
    .Q_N(_06108_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[19] ));
 sg13g2_dfrbp_1 _15840_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net1898),
    .D(_01332_),
    .Q_N(_06107_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[20] ));
 sg13g2_dfrbp_1 _15841_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net1896),
    .D(net3394),
    .Q_N(_06106_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[21] ));
 sg13g2_dfrbp_1 _15842_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net1894),
    .D(_01334_),
    .Q_N(_06105_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[22] ));
 sg13g2_dfrbp_1 _15843_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net1892),
    .D(net3708),
    .Q_N(_06104_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[23] ));
 sg13g2_dfrbp_1 _15844_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net1890),
    .D(_01336_),
    .Q_N(_00136_),
    .Q(\i_tinyqv.cpu.pc[1] ));
 sg13g2_dfrbp_1 _15845_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net1886),
    .D(_01337_),
    .Q_N(_00137_),
    .Q(\i_tinyqv.cpu.pc[2] ));
 sg13g2_dfrbp_1 _15846_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net1882),
    .D(_01338_),
    .Q_N(_06103_),
    .Q(\i_time.l_mtimecmp.data_out[0] ));
 sg13g2_dfrbp_1 _15847_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net1880),
    .D(net3474),
    .Q_N(_06102_),
    .Q(\i_time.l_mtimecmp.data_out[1] ));
 sg13g2_dfrbp_1 _15848_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net1878),
    .D(net3619),
    .Q_N(_06101_),
    .Q(\i_time.l_mtimecmp.data_out[2] ));
 sg13g2_dfrbp_1 _15849_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net1876),
    .D(_01341_),
    .Q_N(_06100_),
    .Q(\i_time.l_mtimecmp.data_out[3] ));
 sg13g2_dfrbp_1 _15850_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net1874),
    .D(_01342_),
    .Q_N(_06099_),
    .Q(\i_time.l_mtimecmp.data_out[4] ));
 sg13g2_dfrbp_1 _15851_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net1872),
    .D(_01343_),
    .Q_N(_06098_),
    .Q(\i_time.l_mtimecmp.data_out[5] ));
 sg13g2_dfrbp_1 _15852_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net1870),
    .D(net3484),
    .Q_N(_06097_),
    .Q(\i_time.l_mtimecmp.data_out[6] ));
 sg13g2_dfrbp_1 _15853_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1868),
    .D(net3675),
    .Q_N(_06096_),
    .Q(\i_time.l_mtimecmp.data_out[7] ));
 sg13g2_dfrbp_1 _15854_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net1866),
    .D(net3663),
    .Q_N(_06095_),
    .Q(\i_time.l_mtimecmp.data_out[8] ));
 sg13g2_dfrbp_1 _15855_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net1864),
    .D(net3831),
    .Q_N(_06094_),
    .Q(\i_time.l_mtimecmp.data_out[9] ));
 sg13g2_dfrbp_1 _15856_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net1862),
    .D(net3779),
    .Q_N(_06093_),
    .Q(\i_time.l_mtimecmp.data_out[10] ));
 sg13g2_dfrbp_1 _15857_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net1860),
    .D(net3748),
    .Q_N(_06092_),
    .Q(\i_time.l_mtimecmp.data_out[11] ));
 sg13g2_dfrbp_1 _15858_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1858),
    .D(_01350_),
    .Q_N(_06091_),
    .Q(\i_time.l_mtimecmp.data_out[12] ));
 sg13g2_dfrbp_1 _15859_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1856),
    .D(net3729),
    .Q_N(_06090_),
    .Q(\i_time.l_mtimecmp.data_out[13] ));
 sg13g2_dfrbp_1 _15860_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1854),
    .D(net3815),
    .Q_N(_06089_),
    .Q(\i_time.l_mtimecmp.data_out[14] ));
 sg13g2_dfrbp_1 _15861_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1852),
    .D(net3545),
    .Q_N(_06088_),
    .Q(\i_time.l_mtimecmp.data_out[15] ));
 sg13g2_dfrbp_1 _15862_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net1850),
    .D(_01354_),
    .Q_N(_06087_),
    .Q(\i_tinyqv.cpu.instr_data_start[3] ));
 sg13g2_dfrbp_1 _15863_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net1846),
    .D(_01355_),
    .Q_N(_00203_),
    .Q(\i_tinyqv.cpu.instr_data_start[4] ));
 sg13g2_dfrbp_1 _15864_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net1842),
    .D(_01356_),
    .Q_N(_06086_),
    .Q(\i_tinyqv.cpu.instr_data_start[5] ));
 sg13g2_dfrbp_1 _15865_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net1838),
    .D(_01357_),
    .Q_N(_06085_),
    .Q(\i_tinyqv.cpu.instr_data_start[6] ));
 sg13g2_dfrbp_1 _15866_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net1821),
    .D(_01358_),
    .Q_N(_06084_),
    .Q(\i_tinyqv.cpu.instr_data_start[7] ));
 sg13g2_dfrbp_1 _15867_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net1817),
    .D(_01359_),
    .Q_N(_06083_),
    .Q(\i_tinyqv.cpu.instr_data_start[8] ));
 sg13g2_dfrbp_1 _15868_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net1813),
    .D(_01360_),
    .Q_N(_06082_),
    .Q(\i_tinyqv.cpu.instr_data_start[9] ));
 sg13g2_dfrbp_1 _15869_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1809),
    .D(_01361_),
    .Q_N(_06081_),
    .Q(\i_tinyqv.cpu.instr_data_start[10] ));
 sg13g2_dfrbp_1 _15870_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net1805),
    .D(_01362_),
    .Q_N(_00239_),
    .Q(\i_tinyqv.cpu.instr_data_start[11] ));
 sg13g2_dfrbp_1 _15871_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net1801),
    .D(_01363_),
    .Q_N(_06080_),
    .Q(\i_tinyqv.cpu.instr_data_start[12] ));
 sg13g2_dfrbp_1 _15872_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net1797),
    .D(_01364_),
    .Q_N(_06079_),
    .Q(\i_tinyqv.cpu.instr_data_start[13] ));
 sg13g2_dfrbp_1 _15873_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net1793),
    .D(_01365_),
    .Q_N(_06078_),
    .Q(\i_tinyqv.cpu.instr_data_start[14] ));
 sg13g2_dfrbp_1 _15874_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net1789),
    .D(_01366_),
    .Q_N(_06077_),
    .Q(\i_tinyqv.cpu.instr_data_start[15] ));
 sg13g2_dfrbp_1 _15875_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net1785),
    .D(_01367_),
    .Q_N(_06076_),
    .Q(\i_tinyqv.cpu.instr_data_start[16] ));
 sg13g2_dfrbp_1 _15876_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net1781),
    .D(_01368_),
    .Q_N(_06075_),
    .Q(\i_tinyqv.cpu.instr_data_start[17] ));
 sg13g2_dfrbp_1 _15877_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net1777),
    .D(_01369_),
    .Q_N(_06074_),
    .Q(\i_tinyqv.cpu.instr_data_start[18] ));
 sg13g2_dfrbp_1 _15878_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net1773),
    .D(_01370_),
    .Q_N(_00207_),
    .Q(\i_tinyqv.cpu.instr_data_start[19] ));
 sg13g2_dfrbp_1 _15879_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net1769),
    .D(_01371_),
    .Q_N(_06073_),
    .Q(\i_tinyqv.cpu.instr_data_start[20] ));
 sg13g2_dfrbp_1 _15880_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net1765),
    .D(_01372_),
    .Q_N(_06072_),
    .Q(\i_tinyqv.cpu.instr_data_start[21] ));
 sg13g2_dfrbp_1 _15881_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net1761),
    .D(_01373_),
    .Q_N(_06071_),
    .Q(\i_tinyqv.cpu.instr_data_start[22] ));
 sg13g2_dfrbp_1 _15882_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net1757),
    .D(_01374_),
    .Q_N(_00202_),
    .Q(\i_tinyqv.cpu.instr_data_start[23] ));
 sg13g2_dfrbp_1 _15883_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net1753),
    .D(net3839),
    .Q_N(_00132_),
    .Q(\i_tinyqv.cpu.instr_fetch_running ));
 sg13g2_dfrbp_1 _15884_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net1749),
    .D(_01376_),
    .Q_N(_00134_),
    .Q(\i_tinyqv.cpu.was_early_branch ));
 sg13g2_dfrbp_1 _15885_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1745),
    .D(_01377_),
    .Q_N(_06070_),
    .Q(\data_to_write[0] ));
 sg13g2_dfrbp_1 _15886_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1741),
    .D(_01378_),
    .Q_N(_06069_),
    .Q(\data_to_write[1] ));
 sg13g2_dfrbp_1 _15887_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1737),
    .D(_01379_),
    .Q_N(_06068_),
    .Q(\data_to_write[2] ));
 sg13g2_dfrbp_1 _15888_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1733),
    .D(_01380_),
    .Q_N(_06067_),
    .Q(\data_to_write[3] ));
 sg13g2_dfrbp_1 _15889_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1729),
    .D(_01381_),
    .Q_N(_06066_),
    .Q(\data_to_write[4] ));
 sg13g2_dfrbp_1 _15890_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1725),
    .D(_01382_),
    .Q_N(_06065_),
    .Q(\data_to_write[5] ));
 sg13g2_dfrbp_1 _15891_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1721),
    .D(_01383_),
    .Q_N(_06064_),
    .Q(\data_to_write[6] ));
 sg13g2_dfrbp_1 _15892_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net1717),
    .D(_01384_),
    .Q_N(_00240_),
    .Q(\data_to_write[7] ));
 sg13g2_dfrbp_1 _15893_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1713),
    .D(_01385_),
    .Q_N(_06063_),
    .Q(\data_to_write[8] ));
 sg13g2_dfrbp_1 _15894_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1709),
    .D(_01386_),
    .Q_N(_06062_),
    .Q(\data_to_write[9] ));
 sg13g2_dfrbp_1 _15895_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net1705),
    .D(_01387_),
    .Q_N(_06061_),
    .Q(\data_to_write[10] ));
 sg13g2_dfrbp_1 _15896_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1701),
    .D(_01388_),
    .Q_N(_06060_),
    .Q(\data_to_write[11] ));
 sg13g2_dfrbp_1 _15897_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net1697),
    .D(_01389_),
    .Q_N(_06059_),
    .Q(\data_to_write[12] ));
 sg13g2_dfrbp_1 _15898_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net1693),
    .D(_01390_),
    .Q_N(_06058_),
    .Q(\data_to_write[13] ));
 sg13g2_dfrbp_1 _15899_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net1689),
    .D(_01391_),
    .Q_N(_06057_),
    .Q(\data_to_write[14] ));
 sg13g2_dfrbp_1 _15900_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net1665),
    .D(_01392_),
    .Q_N(_06056_),
    .Q(\data_to_write[15] ));
 sg13g2_dfrbp_1 _15901_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net1657),
    .D(_01393_),
    .Q_N(_06055_),
    .Q(\data_to_write[16] ));
 sg13g2_dfrbp_1 _15902_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1653),
    .D(_01394_),
    .Q_N(_06054_),
    .Q(\data_to_write[17] ));
 sg13g2_dfrbp_1 _15903_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net1649),
    .D(_01395_),
    .Q_N(_06053_),
    .Q(\data_to_write[18] ));
 sg13g2_dfrbp_1 _15904_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net1645),
    .D(_01396_),
    .Q_N(_06052_),
    .Q(\data_to_write[19] ));
 sg13g2_dfrbp_1 _15905_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net1641),
    .D(_01397_),
    .Q_N(_06051_),
    .Q(\data_to_write[20] ));
 sg13g2_dfrbp_1 _15906_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net1637),
    .D(_01398_),
    .Q_N(_06050_),
    .Q(\data_to_write[21] ));
 sg13g2_dfrbp_1 _15907_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1633),
    .D(_01399_),
    .Q_N(_06049_),
    .Q(\data_to_write[22] ));
 sg13g2_dfrbp_1 _15908_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net1629),
    .D(_01400_),
    .Q_N(_06048_),
    .Q(\data_to_write[23] ));
 sg13g2_dfrbp_1 _15909_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1568),
    .D(_01401_),
    .Q_N(_06047_),
    .Q(\data_to_write[24] ));
 sg13g2_dfrbp_1 _15910_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1550),
    .D(_01402_),
    .Q_N(_06046_),
    .Q(\data_to_write[25] ));
 sg13g2_dfrbp_1 _15911_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net1541),
    .D(_01403_),
    .Q_N(_06045_),
    .Q(\data_to_write[26] ));
 sg13g2_dfrbp_1 _15912_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1533),
    .D(_01404_),
    .Q_N(_06044_),
    .Q(\data_to_write[27] ));
 sg13g2_dfrbp_1 _15913_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net1396),
    .D(_01405_),
    .Q_N(_06043_),
    .Q(\data_to_write[28] ));
 sg13g2_dfrbp_1 _15914_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net1388),
    .D(_01406_),
    .Q_N(_06042_),
    .Q(\data_to_write[29] ));
 sg13g2_dfrbp_1 _15915_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net1216),
    .D(_01407_),
    .Q_N(_06041_),
    .Q(\data_to_write[30] ));
 sg13g2_dfrbp_1 _15916_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1171),
    .D(_01408_),
    .Q_N(_06040_),
    .Q(\data_to_write[31] ));
 sg13g2_dfrbp_1 _15917_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net2067),
    .D(_01409_),
    .Q_N(_06039_),
    .Q(\i_tinyqv.cpu.data_write_n[0] ));
 sg13g2_dfrbp_1 _15918_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net2049),
    .D(_01410_),
    .Q_N(_06038_),
    .Q(\i_tinyqv.cpu.data_write_n[1] ));
 sg13g2_dfrbp_1 _15919_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net2041),
    .D(_01411_),
    .Q_N(_06037_),
    .Q(\i_tinyqv.cpu.data_read_n[0] ));
 sg13g2_dfrbp_1 _15920_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net1791),
    .D(net3860),
    .Q_N(_07264_),
    .Q(\i_tinyqv.cpu.data_read_n[1] ));
 sg13g2_dfrbp_1 _15921_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net2031),
    .D(_00064_),
    .Q_N(_06036_),
    .Q(debug_data_continue));
 sg13g2_dfrbp_1 _15922_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net2023),
    .D(net3791),
    .Q_N(_00119_),
    .Q(\i_tinyqv.cpu.no_write_in_progress ));
 sg13g2_dfrbp_1 _15923_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net2014),
    .D(net3179),
    .Q_N(_06035_),
    .Q(\i_tinyqv.cpu.load_started ));
 sg13g2_dfrbp_1 _15924_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net2006),
    .D(net3857),
    .Q_N(_00266_),
    .Q(\i_tinyqv.cpu.counter[2] ));
 sg13g2_dfrbp_1 _15925_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net2002),
    .D(_01416_),
    .Q_N(_00124_),
    .Q(\i_tinyqv.cpu.counter[3] ));
 sg13g2_dfrbp_1 _15926_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net1998),
    .D(_01417_),
    .Q_N(_00120_),
    .Q(\i_tinyqv.cpu.counter[4] ));
 sg13g2_dfrbp_1 _15927_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net1960),
    .D(net3050),
    .Q_N(_00205_),
    .Q(\i_tinyqv.cpu.data_ready_sync ));
 sg13g2_dfrbp_1 _15928_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net1952),
    .D(net3824),
    .Q_N(_06034_),
    .Q(\i_tinyqv.cpu.data_ready_latch ));
 sg13g2_dfrbp_1 _15929_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net1948),
    .D(_01420_),
    .Q_N(_06033_),
    .Q(\i_tinyqv.cpu.is_load ));
 sg13g2_dfrbp_1 _15930_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net1936),
    .D(_01421_),
    .Q_N(_06032_),
    .Q(\i_tinyqv.cpu.is_alu_imm ));
 sg13g2_dfrbp_1 _15931_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net1888),
    .D(_01422_),
    .Q_N(_06031_),
    .Q(\i_tinyqv.cpu.is_auipc ));
 sg13g2_dfrbp_1 _15932_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net1848),
    .D(_01423_),
    .Q_N(_06030_),
    .Q(\i_tinyqv.cpu.is_store ));
 sg13g2_dfrbp_1 _15933_ (.CLK(clknet_leaf_129_clk_regs),
    .RESET_B(net1840),
    .D(_01424_),
    .Q_N(_06029_),
    .Q(\i_tinyqv.cpu.is_alu_reg ));
 sg13g2_dfrbp_1 _15934_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net1819),
    .D(_01425_),
    .Q_N(_06028_),
    .Q(\i_tinyqv.cpu.is_lui ));
 sg13g2_dfrbp_1 _15935_ (.CLK(clknet_leaf_125_clk_regs),
    .RESET_B(net1811),
    .D(_01426_),
    .Q_N(_06027_),
    .Q(\i_tinyqv.cpu.is_branch ));
 sg13g2_dfrbp_1 _15936_ (.CLK(clknet_leaf_128_clk_regs),
    .RESET_B(net1803),
    .D(_01427_),
    .Q_N(_06026_),
    .Q(\i_tinyqv.cpu.is_jalr ));
 sg13g2_dfrbp_1 _15937_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net1795),
    .D(net3679),
    .Q_N(_06025_),
    .Q(\i_tinyqv.cpu.is_jal ));
 sg13g2_dfrbp_1 _15938_ (.CLK(clknet_leaf_124_clk_regs),
    .RESET_B(net1787),
    .D(_01429_),
    .Q_N(_06024_),
    .Q(\i_tinyqv.cpu.is_system ));
 sg13g2_dfrbp_1 _15939_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net1779),
    .D(_01430_),
    .Q_N(_06023_),
    .Q(\i_tinyqv.cpu.instr_len[1] ));
 sg13g2_dfrbp_1 _15940_ (.CLK(clknet_leaf_139_clk_regs),
    .RESET_B(net1771),
    .D(_01431_),
    .Q_N(_06022_),
    .Q(\i_tinyqv.cpu.instr_len[2] ));
 sg13g2_dfrbp_1 _15941_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net1763),
    .D(_01432_),
    .Q_N(_06021_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[0] ));
 sg13g2_dfrbp_1 _15942_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net1759),
    .D(_01433_),
    .Q_N(_06020_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[1] ));
 sg13g2_dfrbp_1 _15943_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net1755),
    .D(_01434_),
    .Q_N(_06019_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[2] ));
 sg13g2_dfrbp_1 _15944_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net1751),
    .D(_01435_),
    .Q_N(_06018_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[3] ));
 sg13g2_dfrbp_1 _15945_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net1747),
    .D(_01436_),
    .Q_N(_06017_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[4] ));
 sg13g2_dfrbp_1 _15946_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net1743),
    .D(_01437_),
    .Q_N(_06016_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[5] ));
 sg13g2_dfrbp_1 _15947_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net1739),
    .D(_01438_),
    .Q_N(_06015_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[6] ));
 sg13g2_dfrbp_1 _15948_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net1735),
    .D(_01439_),
    .Q_N(_06014_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[7] ));
 sg13g2_dfrbp_1 _15949_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net1731),
    .D(_01440_),
    .Q_N(_06013_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[8] ));
 sg13g2_dfrbp_1 _15950_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net1727),
    .D(_01441_),
    .Q_N(_06012_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[9] ));
 sg13g2_dfrbp_1 _15951_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net1723),
    .D(_01442_),
    .Q_N(_06011_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[10] ));
 sg13g2_dfrbp_1 _15952_ (.CLK(clknet_leaf_134_clk_regs),
    .RESET_B(net1719),
    .D(_01443_),
    .Q_N(_06010_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[11] ));
 sg13g2_dfrbp_1 _15953_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net1715),
    .D(_01444_),
    .Q_N(_06009_),
    .Q(\i_tinyqv.cpu.imm[12] ));
 sg13g2_dfrbp_1 _15954_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net1711),
    .D(_01445_),
    .Q_N(_06008_),
    .Q(\i_tinyqv.cpu.imm[13] ));
 sg13g2_dfrbp_1 _15955_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net1707),
    .D(_01446_),
    .Q_N(_06007_),
    .Q(\i_tinyqv.cpu.imm[14] ));
 sg13g2_dfrbp_1 _15956_ (.CLK(clknet_leaf_135_clk_regs),
    .RESET_B(net1703),
    .D(_01447_),
    .Q_N(_06006_),
    .Q(\i_tinyqv.cpu.imm[15] ));
 sg13g2_dfrbp_1 _15957_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net1699),
    .D(_01448_),
    .Q_N(_06005_),
    .Q(\i_tinyqv.cpu.imm[16] ));
 sg13g2_dfrbp_1 _15958_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net1695),
    .D(_01449_),
    .Q_N(_06004_),
    .Q(\i_tinyqv.cpu.imm[17] ));
 sg13g2_dfrbp_1 _15959_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net1691),
    .D(_01450_),
    .Q_N(_06003_),
    .Q(\i_tinyqv.cpu.imm[18] ));
 sg13g2_dfrbp_1 _15960_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net1667),
    .D(net3993),
    .Q_N(_06002_),
    .Q(\i_tinyqv.cpu.imm[19] ));
 sg13g2_dfrbp_1 _15961_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net1663),
    .D(_01452_),
    .Q_N(_06001_),
    .Q(\i_tinyqv.cpu.imm[20] ));
 sg13g2_dfrbp_1 _15962_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net1655),
    .D(_01453_),
    .Q_N(_06000_),
    .Q(\i_tinyqv.cpu.imm[21] ));
 sg13g2_dfrbp_1 _15963_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net1651),
    .D(_01454_),
    .Q_N(_05999_),
    .Q(\i_tinyqv.cpu.imm[22] ));
 sg13g2_dfrbp_1 _15964_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net1647),
    .D(_01455_),
    .Q_N(_05998_),
    .Q(\i_tinyqv.cpu.imm[23] ));
 sg13g2_dfrbp_1 _15965_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net1643),
    .D(_01456_),
    .Q_N(_05997_),
    .Q(\i_tinyqv.cpu.imm[24] ));
 sg13g2_dfrbp_1 _15966_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net1639),
    .D(_01457_),
    .Q_N(_05996_),
    .Q(\i_tinyqv.cpu.imm[25] ));
 sg13g2_dfrbp_1 _15967_ (.CLK(clknet_leaf_132_clk_regs),
    .RESET_B(net1635),
    .D(_01458_),
    .Q_N(_05995_),
    .Q(\i_tinyqv.cpu.imm[26] ));
 sg13g2_dfrbp_1 _15968_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net1631),
    .D(_01459_),
    .Q_N(_05994_),
    .Q(\i_tinyqv.cpu.imm[27] ));
 sg13g2_dfrbp_1 _15969_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net1570),
    .D(_01460_),
    .Q_N(_05993_),
    .Q(\i_tinyqv.cpu.imm[28] ));
 sg13g2_dfrbp_1 _15970_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net1566),
    .D(_01461_),
    .Q_N(_05992_),
    .Q(\i_tinyqv.cpu.imm[29] ));
 sg13g2_dfrbp_1 _15971_ (.CLK(clknet_leaf_136_clk_regs),
    .RESET_B(net1545),
    .D(_01462_),
    .Q_N(_05991_),
    .Q(\i_tinyqv.cpu.imm[30] ));
 sg13g2_dfrbp_1 _15972_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net1537),
    .D(_01463_),
    .Q_N(_05990_),
    .Q(\i_tinyqv.cpu.imm[31] ));
 sg13g2_dfrbp_1 _15973_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net1400),
    .D(_01464_),
    .Q_N(_05989_),
    .Q(\i_tinyqv.cpu.alu_op[0] ));
 sg13g2_dfrbp_1 _15974_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net1392),
    .D(_01465_),
    .Q_N(_00125_),
    .Q(\i_tinyqv.cpu.alu_op[1] ));
 sg13g2_dfrbp_1 _15975_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net1218),
    .D(_01466_),
    .Q_N(_00130_),
    .Q(\i_tinyqv.cpu.alu_op[2] ));
 sg13g2_dfrbp_1 _15976_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net1183),
    .D(_01467_),
    .Q_N(_00121_),
    .Q(\i_tinyqv.cpu.alu_op[3] ));
 sg13g2_dfrbp_1 _15977_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net1167),
    .D(_01468_),
    .Q_N(_05988_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[0] ));
 sg13g2_dfrbp_1 _15978_ (.CLK(clknet_leaf_138_clk_regs),
    .RESET_B(net2053),
    .D(_01469_),
    .Q_N(_05987_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[1] ));
 sg13g2_dfrbp_1 _15979_ (.CLK(clknet_leaf_137_clk_regs),
    .RESET_B(net2045),
    .D(_01470_),
    .Q_N(_05986_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[2] ));
 sg13g2_dfrbp_1 _15980_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net2037),
    .D(_01471_),
    .Q_N(_05985_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ));
 sg13g2_dfrbp_1 _15981_ (.CLK(clknet_leaf_123_clk_regs),
    .RESET_B(net2027),
    .D(_01472_),
    .Q_N(_05984_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ));
 sg13g2_dfrbp_1 _15982_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net2018),
    .D(_01473_),
    .Q_N(_05983_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ));
 sg13g2_dfrbp_1 _15983_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net2010),
    .D(_01474_),
    .Q_N(_05982_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ));
 sg13g2_dfrbp_1 _15984_ (.CLK(clknet_leaf_123_clk_regs),
    .RESET_B(net1956),
    .D(_01475_),
    .Q_N(_05981_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ));
 sg13g2_dfrbp_1 _15985_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net1940),
    .D(_01476_),
    .Q_N(_05980_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ));
 sg13g2_dfrbp_1 _15986_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net1932),
    .D(_01477_),
    .Q_N(_05979_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ));
 sg13g2_dfrbp_1 _15987_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net1884),
    .D(_01478_),
    .Q_N(_05978_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ));
 sg13g2_dfrbp_1 _15988_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net1844),
    .D(net3445),
    .Q_N(_00254_),
    .Q(\i_tinyqv.cpu.additional_mem_ops[0] ));
 sg13g2_dfrbp_1 _15989_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net1815),
    .D(_01480_),
    .Q_N(_05977_),
    .Q(\i_tinyqv.cpu.additional_mem_ops[1] ));
 sg13g2_dfrbp_1 _15990_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net1799),
    .D(_01481_),
    .Q_N(_05976_),
    .Q(\i_tinyqv.cpu.additional_mem_ops[2] ));
 sg13g2_dfrbp_1 _15991_ (.CLK(clknet_leaf_133_clk_regs),
    .RESET_B(net1783),
    .D(net3894),
    .Q_N(_05975_),
    .Q(\i_tinyqv.cpu.mem_op_increment_reg ));
 sg13g2_dfrbp_1 _15992_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net1767),
    .D(_01483_),
    .Q_N(_00129_),
    .Q(\i_tinyqv.cpu.i_core.is_interrupt ));
 sg13g2_dfrbp_1 _15993_ (.CLK(clknet_leaf_139_clk_regs),
    .RESET_B(net1807),
    .D(net4102),
    .Q_N(_00135_),
    .Q(debug_instr_valid));
 sg13g2_dfrbp_1 _15994_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net1775),
    .D(net2829),
    .Q_N(_05974_),
    .Q(\i_time.time_pulse ));
 sg13g2_dfrbp_1 _15995_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net1835),
    .D(_01486_),
    .Q_N(_05973_),
    .Q(\i_tinyqv.cpu.instr_write_offset[3] ));
 sg13g2_tiehi _14539__664 (.L_HI(net664));
 sg13g2_tiehi _14540__665 (.L_HI(net665));
 sg13g2_tiehi _14541__666 (.L_HI(net666));
 sg13g2_tiehi _14542__667 (.L_HI(net667));
 sg13g2_tiehi _14543__668 (.L_HI(net668));
 sg13g2_tiehi _14544__669 (.L_HI(net669));
 sg13g2_tiehi _14545__670 (.L_HI(net670));
 sg13g2_tiehi _14546__671 (.L_HI(net671));
 sg13g2_tiehi _14547__672 (.L_HI(net672));
 sg13g2_tiehi _14548__673 (.L_HI(net673));
 sg13g2_tiehi _14549__674 (.L_HI(net674));
 sg13g2_tiehi _14550__675 (.L_HI(net675));
 sg13g2_tiehi _14551__676 (.L_HI(net676));
 sg13g2_tiehi _14552__677 (.L_HI(net677));
 sg13g2_tiehi _15280__678 (.L_HI(net678));
 sg13g2_tiehi _15763__679 (.L_HI(net679));
 sg13g2_tiehi _15279__680 (.L_HI(net680));
 sg13g2_tiehi _15762__681 (.L_HI(net681));
 sg13g2_tiehi _15278__682 (.L_HI(net682));
 sg13g2_tiehi _14553__683 (.L_HI(net683));
 sg13g2_tiehi _14559__684 (.L_HI(net684));
 sg13g2_tiehi _14560__685 (.L_HI(net685));
 sg13g2_tiehi _14561__686 (.L_HI(net686));
 sg13g2_tiehi _14562__687 (.L_HI(net687));
 sg13g2_tiehi _14563__688 (.L_HI(net688));
 sg13g2_tiehi _14564__689 (.L_HI(net689));
 sg13g2_tiehi _14565__690 (.L_HI(net690));
 sg13g2_tiehi _14566__691 (.L_HI(net691));
 sg13g2_tiehi _14567__692 (.L_HI(net692));
 sg13g2_tiehi _14568__693 (.L_HI(net693));
 sg13g2_tiehi _14569__694 (.L_HI(net694));
 sg13g2_tiehi _14570__695 (.L_HI(net695));
 sg13g2_tiehi _14571__696 (.L_HI(net696));
 sg13g2_tiehi _14572__697 (.L_HI(net697));
 sg13g2_tiehi _14573__698 (.L_HI(net698));
 sg13g2_tiehi _14574__699 (.L_HI(net699));
 sg13g2_tiehi _14575__700 (.L_HI(net700));
 sg13g2_tiehi _14576__701 (.L_HI(net701));
 sg13g2_tiehi _14577__702 (.L_HI(net702));
 sg13g2_tiehi _14578__703 (.L_HI(net703));
 sg13g2_tiehi _14579__704 (.L_HI(net704));
 sg13g2_tiehi _14580__705 (.L_HI(net705));
 sg13g2_tiehi _14581__706 (.L_HI(net706));
 sg13g2_tiehi _14582__707 (.L_HI(net707));
 sg13g2_tiehi _14583__708 (.L_HI(net708));
 sg13g2_tiehi _14584__709 (.L_HI(net709));
 sg13g2_tiehi _14585__710 (.L_HI(net710));
 sg13g2_tiehi _15761__711 (.L_HI(net711));
 sg13g2_tiehi _15277__712 (.L_HI(net712));
 sg13g2_tiehi _15760__713 (.L_HI(net713));
 sg13g2_tiehi _15276__714 (.L_HI(net714));
 sg13g2_tiehi _15759__715 (.L_HI(net715));
 sg13g2_tiehi _15275__716 (.L_HI(net716));
 sg13g2_tiehi _14586__717 (.L_HI(net717));
 sg13g2_tiehi _14593__718 (.L_HI(net718));
 sg13g2_tiehi _14594__719 (.L_HI(net719));
 sg13g2_tiehi _14595__720 (.L_HI(net720));
 sg13g2_tiehi _14596__721 (.L_HI(net721));
 sg13g2_tiehi _14597__722 (.L_HI(net722));
 sg13g2_tiehi _14598__723 (.L_HI(net723));
 sg13g2_tiehi _14599__724 (.L_HI(net724));
 sg13g2_tiehi _14600__725 (.L_HI(net725));
 sg13g2_tiehi _14601__726 (.L_HI(net726));
 sg13g2_tiehi _14602__727 (.L_HI(net727));
 sg13g2_tiehi _14603__728 (.L_HI(net728));
 sg13g2_tiehi _14604__729 (.L_HI(net729));
 sg13g2_tiehi _14605__730 (.L_HI(net730));
 sg13g2_tiehi _14606__731 (.L_HI(net731));
 sg13g2_tiehi _14607__732 (.L_HI(net732));
 sg13g2_tiehi _14608__733 (.L_HI(net733));
 sg13g2_tiehi _14609__734 (.L_HI(net734));
 sg13g2_tiehi _14610__735 (.L_HI(net735));
 sg13g2_tiehi _14611__736 (.L_HI(net736));
 sg13g2_tiehi _14612__737 (.L_HI(net737));
 sg13g2_tiehi _14613__738 (.L_HI(net738));
 sg13g2_tiehi _14614__739 (.L_HI(net739));
 sg13g2_tiehi _14615__740 (.L_HI(net740));
 sg13g2_tiehi _14616__741 (.L_HI(net741));
 sg13g2_tiehi _14617__742 (.L_HI(net742));
 sg13g2_tiehi _14618__743 (.L_HI(net743));
 sg13g2_tiehi _14619__744 (.L_HI(net744));
 sg13g2_tiehi _14620__745 (.L_HI(net745));
 sg13g2_tiehi _14621__746 (.L_HI(net746));
 sg13g2_tiehi _14622__747 (.L_HI(net747));
 sg13g2_tiehi _14623__748 (.L_HI(net748));
 sg13g2_tiehi _14624__749 (.L_HI(net749));
 sg13g2_tiehi _14625__750 (.L_HI(net750));
 sg13g2_tiehi _14626__751 (.L_HI(net751));
 sg13g2_tiehi _14627__752 (.L_HI(net752));
 sg13g2_tiehi _14628__753 (.L_HI(net753));
 sg13g2_tiehi _14629__754 (.L_HI(net754));
 sg13g2_tiehi _14630__755 (.L_HI(net755));
 sg13g2_tiehi _14631__756 (.L_HI(net756));
 sg13g2_tiehi _14632__757 (.L_HI(net757));
 sg13g2_tiehi _14633__758 (.L_HI(net758));
 sg13g2_tiehi _14634__759 (.L_HI(net759));
 sg13g2_tiehi _14635__760 (.L_HI(net760));
 sg13g2_tiehi _14636__761 (.L_HI(net761));
 sg13g2_tiehi _14637__762 (.L_HI(net762));
 sg13g2_tiehi _14638__763 (.L_HI(net763));
 sg13g2_tiehi _14639__764 (.L_HI(net764));
 sg13g2_tiehi _14640__765 (.L_HI(net765));
 sg13g2_tiehi _14641__766 (.L_HI(net766));
 sg13g2_tiehi _14642__767 (.L_HI(net767));
 sg13g2_tiehi _14643__768 (.L_HI(net768));
 sg13g2_tiehi _14644__769 (.L_HI(net769));
 sg13g2_tiehi _14645__770 (.L_HI(net770));
 sg13g2_tiehi _14646__771 (.L_HI(net771));
 sg13g2_tiehi _14647__772 (.L_HI(net772));
 sg13g2_tiehi _14648__773 (.L_HI(net773));
 sg13g2_tiehi _14649__774 (.L_HI(net774));
 sg13g2_tiehi _14650__775 (.L_HI(net775));
 sg13g2_tiehi _14651__776 (.L_HI(net776));
 sg13g2_tiehi _14652__777 (.L_HI(net777));
 sg13g2_tiehi _14653__778 (.L_HI(net778));
 sg13g2_tiehi _14654__779 (.L_HI(net779));
 sg13g2_tiehi _14655__780 (.L_HI(net780));
 sg13g2_tiehi _14656__781 (.L_HI(net781));
 sg13g2_tiehi _14657__782 (.L_HI(net782));
 sg13g2_tiehi _14658__783 (.L_HI(net783));
 sg13g2_tiehi _14659__784 (.L_HI(net784));
 sg13g2_tiehi _14660__785 (.L_HI(net785));
 sg13g2_tiehi _14661__786 (.L_HI(net786));
 sg13g2_tiehi _14662__787 (.L_HI(net787));
 sg13g2_tiehi _14663__788 (.L_HI(net788));
 sg13g2_tiehi _14664__789 (.L_HI(net789));
 sg13g2_tiehi _14665__790 (.L_HI(net790));
 sg13g2_tiehi _14666__791 (.L_HI(net791));
 sg13g2_tiehi _14667__792 (.L_HI(net792));
 sg13g2_tiehi _14668__793 (.L_HI(net793));
 sg13g2_tiehi _14669__794 (.L_HI(net794));
 sg13g2_tiehi _14670__795 (.L_HI(net795));
 sg13g2_tiehi _14671__796 (.L_HI(net796));
 sg13g2_tiehi _14672__797 (.L_HI(net797));
 sg13g2_tiehi _14673__798 (.L_HI(net798));
 sg13g2_tiehi _14674__799 (.L_HI(net799));
 sg13g2_tiehi _14675__800 (.L_HI(net800));
 sg13g2_tiehi _14676__801 (.L_HI(net801));
 sg13g2_tiehi _14677__802 (.L_HI(net802));
 sg13g2_tiehi _14678__803 (.L_HI(net803));
 sg13g2_tiehi _14679__804 (.L_HI(net804));
 sg13g2_tiehi _14680__805 (.L_HI(net805));
 sg13g2_tiehi _14681__806 (.L_HI(net806));
 sg13g2_tiehi _14682__807 (.L_HI(net807));
 sg13g2_tiehi _14683__808 (.L_HI(net808));
 sg13g2_tiehi _14684__809 (.L_HI(net809));
 sg13g2_tiehi _14685__810 (.L_HI(net810));
 sg13g2_tiehi _14686__811 (.L_HI(net811));
 sg13g2_tiehi _14687__812 (.L_HI(net812));
 sg13g2_tiehi _14688__813 (.L_HI(net813));
 sg13g2_tiehi _14689__814 (.L_HI(net814));
 sg13g2_tiehi _14690__815 (.L_HI(net815));
 sg13g2_tiehi _14691__816 (.L_HI(net816));
 sg13g2_tiehi _14692__817 (.L_HI(net817));
 sg13g2_tiehi _14693__818 (.L_HI(net818));
 sg13g2_tiehi _14694__819 (.L_HI(net819));
 sg13g2_tiehi _14695__820 (.L_HI(net820));
 sg13g2_tiehi _14696__821 (.L_HI(net821));
 sg13g2_tiehi _14697__822 (.L_HI(net822));
 sg13g2_tiehi _14698__823 (.L_HI(net823));
 sg13g2_tiehi _14699__824 (.L_HI(net824));
 sg13g2_tiehi _14700__825 (.L_HI(net825));
 sg13g2_tiehi _14701__826 (.L_HI(net826));
 sg13g2_tiehi _14702__827 (.L_HI(net827));
 sg13g2_tiehi _14703__828 (.L_HI(net828));
 sg13g2_tiehi _14704__829 (.L_HI(net829));
 sg13g2_tiehi _14705__830 (.L_HI(net830));
 sg13g2_tiehi _14706__831 (.L_HI(net831));
 sg13g2_tiehi _14707__832 (.L_HI(net832));
 sg13g2_tiehi _14708__833 (.L_HI(net833));
 sg13g2_tiehi _14709__834 (.L_HI(net834));
 sg13g2_tiehi _14710__835 (.L_HI(net835));
 sg13g2_tiehi _14711__836 (.L_HI(net836));
 sg13g2_tiehi _14712__837 (.L_HI(net837));
 sg13g2_tiehi _14713__838 (.L_HI(net838));
 sg13g2_tiehi _14714__839 (.L_HI(net839));
 sg13g2_tiehi _14715__840 (.L_HI(net840));
 sg13g2_tiehi _14716__841 (.L_HI(net841));
 sg13g2_tiehi _14717__842 (.L_HI(net842));
 sg13g2_tiehi _14718__843 (.L_HI(net843));
 sg13g2_tiehi _14719__844 (.L_HI(net844));
 sg13g2_tiehi _14720__845 (.L_HI(net845));
 sg13g2_tiehi _14721__846 (.L_HI(net846));
 sg13g2_tiehi _14722__847 (.L_HI(net847));
 sg13g2_tiehi _14723__848 (.L_HI(net848));
 sg13g2_tiehi _14724__849 (.L_HI(net849));
 sg13g2_tiehi _14725__850 (.L_HI(net850));
 sg13g2_tiehi _14726__851 (.L_HI(net851));
 sg13g2_tiehi _14727__852 (.L_HI(net852));
 sg13g2_tiehi _14728__853 (.L_HI(net853));
 sg13g2_tiehi _14729__854 (.L_HI(net854));
 sg13g2_tiehi _14730__855 (.L_HI(net855));
 sg13g2_tiehi _14731__856 (.L_HI(net856));
 sg13g2_tiehi _14732__857 (.L_HI(net857));
 sg13g2_tiehi _14733__858 (.L_HI(net858));
 sg13g2_tiehi _14734__859 (.L_HI(net859));
 sg13g2_tiehi _14735__860 (.L_HI(net860));
 sg13g2_tiehi _14736__861 (.L_HI(net861));
 sg13g2_tiehi _14737__862 (.L_HI(net862));
 sg13g2_tiehi _14738__863 (.L_HI(net863));
 sg13g2_tiehi _14739__864 (.L_HI(net864));
 sg13g2_tiehi _14740__865 (.L_HI(net865));
 sg13g2_tiehi _14741__866 (.L_HI(net866));
 sg13g2_tiehi _14742__867 (.L_HI(net867));
 sg13g2_tiehi _14743__868 (.L_HI(net868));
 sg13g2_tiehi _14744__869 (.L_HI(net869));
 sg13g2_tiehi _14745__870 (.L_HI(net870));
 sg13g2_tiehi _14746__871 (.L_HI(net871));
 sg13g2_tiehi _14747__872 (.L_HI(net872));
 sg13g2_tiehi _14748__873 (.L_HI(net873));
 sg13g2_tiehi _14749__874 (.L_HI(net874));
 sg13g2_tiehi _14750__875 (.L_HI(net875));
 sg13g2_tiehi _14751__876 (.L_HI(net876));
 sg13g2_tiehi _14752__877 (.L_HI(net877));
 sg13g2_tiehi _14753__878 (.L_HI(net878));
 sg13g2_tiehi _14754__879 (.L_HI(net879));
 sg13g2_tiehi _14755__880 (.L_HI(net880));
 sg13g2_tiehi _14756__881 (.L_HI(net881));
 sg13g2_tiehi _14757__882 (.L_HI(net882));
 sg13g2_tiehi _14758__883 (.L_HI(net883));
 sg13g2_tiehi _14759__884 (.L_HI(net884));
 sg13g2_tiehi _14760__885 (.L_HI(net885));
 sg13g2_tiehi _14761__886 (.L_HI(net886));
 sg13g2_tiehi _14762__887 (.L_HI(net887));
 sg13g2_tiehi _14763__888 (.L_HI(net888));
 sg13g2_tiehi _14764__889 (.L_HI(net889));
 sg13g2_tiehi _14765__890 (.L_HI(net890));
 sg13g2_tiehi _14766__891 (.L_HI(net891));
 sg13g2_tiehi _14767__892 (.L_HI(net892));
 sg13g2_tiehi _14768__893 (.L_HI(net893));
 sg13g2_tiehi _14769__894 (.L_HI(net894));
 sg13g2_tiehi _14770__895 (.L_HI(net895));
 sg13g2_tiehi _14771__896 (.L_HI(net896));
 sg13g2_tiehi _14772__897 (.L_HI(net897));
 sg13g2_tiehi _14773__898 (.L_HI(net898));
 sg13g2_tiehi _14774__899 (.L_HI(net899));
 sg13g2_tiehi _14775__900 (.L_HI(net900));
 sg13g2_tiehi _14776__901 (.L_HI(net901));
 sg13g2_tiehi _14777__902 (.L_HI(net902));
 sg13g2_tiehi _14778__903 (.L_HI(net903));
 sg13g2_tiehi _14779__904 (.L_HI(net904));
 sg13g2_tiehi _14780__905 (.L_HI(net905));
 sg13g2_tiehi _14781__906 (.L_HI(net906));
 sg13g2_tiehi _14782__907 (.L_HI(net907));
 sg13g2_tiehi _14783__908 (.L_HI(net908));
 sg13g2_tiehi _14784__909 (.L_HI(net909));
 sg13g2_tiehi _14785__910 (.L_HI(net910));
 sg13g2_tiehi _14786__911 (.L_HI(net911));
 sg13g2_tiehi _14787__912 (.L_HI(net912));
 sg13g2_tiehi _14788__913 (.L_HI(net913));
 sg13g2_tiehi _14789__914 (.L_HI(net914));
 sg13g2_tiehi _14790__915 (.L_HI(net915));
 sg13g2_tiehi _14791__916 (.L_HI(net916));
 sg13g2_tiehi _14792__917 (.L_HI(net917));
 sg13g2_tiehi _14793__918 (.L_HI(net918));
 sg13g2_tiehi _14794__919 (.L_HI(net919));
 sg13g2_tiehi _14795__920 (.L_HI(net920));
 sg13g2_tiehi _14796__921 (.L_HI(net921));
 sg13g2_tiehi _14797__922 (.L_HI(net922));
 sg13g2_tiehi _14798__923 (.L_HI(net923));
 sg13g2_tiehi _14799__924 (.L_HI(net924));
 sg13g2_tiehi _14800__925 (.L_HI(net925));
 sg13g2_tiehi _14801__926 (.L_HI(net926));
 sg13g2_tiehi _14802__927 (.L_HI(net927));
 sg13g2_tiehi _14803__928 (.L_HI(net928));
 sg13g2_tiehi _14804__929 (.L_HI(net929));
 sg13g2_tiehi _14805__930 (.L_HI(net930));
 sg13g2_tiehi _14806__931 (.L_HI(net931));
 sg13g2_tiehi _14807__932 (.L_HI(net932));
 sg13g2_tiehi _14808__933 (.L_HI(net933));
 sg13g2_tiehi _14809__934 (.L_HI(net934));
 sg13g2_tiehi _14810__935 (.L_HI(net935));
 sg13g2_tiehi _14811__936 (.L_HI(net936));
 sg13g2_tiehi _14812__937 (.L_HI(net937));
 sg13g2_tiehi _14813__938 (.L_HI(net938));
 sg13g2_tiehi _14814__939 (.L_HI(net939));
 sg13g2_tiehi _14815__940 (.L_HI(net940));
 sg13g2_tiehi _14816__941 (.L_HI(net941));
 sg13g2_tiehi _14817__942 (.L_HI(net942));
 sg13g2_tiehi _14818__943 (.L_HI(net943));
 sg13g2_tiehi _14819__944 (.L_HI(net944));
 sg13g2_tiehi _14820__945 (.L_HI(net945));
 sg13g2_tiehi _14821__946 (.L_HI(net946));
 sg13g2_tiehi _14822__947 (.L_HI(net947));
 sg13g2_tiehi _14823__948 (.L_HI(net948));
 sg13g2_tiehi _14824__949 (.L_HI(net949));
 sg13g2_tiehi _14825__950 (.L_HI(net950));
 sg13g2_tiehi _14826__951 (.L_HI(net951));
 sg13g2_tiehi _14827__952 (.L_HI(net952));
 sg13g2_tiehi _14828__953 (.L_HI(net953));
 sg13g2_tiehi _14829__954 (.L_HI(net954));
 sg13g2_tiehi _14830__955 (.L_HI(net955));
 sg13g2_tiehi _14831__956 (.L_HI(net956));
 sg13g2_tiehi _14832__957 (.L_HI(net957));
 sg13g2_tiehi _14833__958 (.L_HI(net958));
 sg13g2_tiehi _14834__959 (.L_HI(net959));
 sg13g2_tiehi _14835__960 (.L_HI(net960));
 sg13g2_tiehi _14836__961 (.L_HI(net961));
 sg13g2_tiehi _14837__962 (.L_HI(net962));
 sg13g2_tiehi _14838__963 (.L_HI(net963));
 sg13g2_tiehi _14839__964 (.L_HI(net964));
 sg13g2_tiehi _14840__965 (.L_HI(net965));
 sg13g2_tiehi _14841__966 (.L_HI(net966));
 sg13g2_tiehi _14842__967 (.L_HI(net967));
 sg13g2_tiehi _14843__968 (.L_HI(net968));
 sg13g2_tiehi _14844__969 (.L_HI(net969));
 sg13g2_tiehi _14845__970 (.L_HI(net970));
 sg13g2_tiehi _14846__971 (.L_HI(net971));
 sg13g2_tiehi _14847__972 (.L_HI(net972));
 sg13g2_tiehi _14848__973 (.L_HI(net973));
 sg13g2_tiehi _14849__974 (.L_HI(net974));
 sg13g2_tiehi _14850__975 (.L_HI(net975));
 sg13g2_tiehi _14851__976 (.L_HI(net976));
 sg13g2_tiehi _14852__977 (.L_HI(net977));
 sg13g2_tiehi _14853__978 (.L_HI(net978));
 sg13g2_tiehi _14854__979 (.L_HI(net979));
 sg13g2_tiehi _14855__980 (.L_HI(net980));
 sg13g2_tiehi _14856__981 (.L_HI(net981));
 sg13g2_tiehi _14857__982 (.L_HI(net982));
 sg13g2_tiehi _14858__983 (.L_HI(net983));
 sg13g2_tiehi _14859__984 (.L_HI(net984));
 sg13g2_tiehi _14860__985 (.L_HI(net985));
 sg13g2_tiehi _14861__986 (.L_HI(net986));
 sg13g2_tiehi _14862__987 (.L_HI(net987));
 sg13g2_tiehi _14863__988 (.L_HI(net988));
 sg13g2_tiehi _14864__989 (.L_HI(net989));
 sg13g2_tiehi _14865__990 (.L_HI(net990));
 sg13g2_tiehi _14866__991 (.L_HI(net991));
 sg13g2_tiehi _14867__992 (.L_HI(net992));
 sg13g2_tiehi _14868__993 (.L_HI(net993));
 sg13g2_tiehi _14869__994 (.L_HI(net994));
 sg13g2_tiehi _14870__995 (.L_HI(net995));
 sg13g2_tiehi _14871__996 (.L_HI(net996));
 sg13g2_tiehi _14872__997 (.L_HI(net997));
 sg13g2_tiehi _14873__998 (.L_HI(net998));
 sg13g2_tiehi _14874__999 (.L_HI(net999));
 sg13g2_tiehi _14875__1000 (.L_HI(net1000));
 sg13g2_tiehi _14876__1001 (.L_HI(net1001));
 sg13g2_tiehi _14877__1002 (.L_HI(net1002));
 sg13g2_tiehi _14878__1003 (.L_HI(net1003));
 sg13g2_tiehi _14879__1004 (.L_HI(net1004));
 sg13g2_tiehi _14880__1005 (.L_HI(net1005));
 sg13g2_tiehi _14881__1006 (.L_HI(net1006));
 sg13g2_tiehi _14882__1007 (.L_HI(net1007));
 sg13g2_tiehi _14883__1008 (.L_HI(net1008));
 sg13g2_tiehi _14884__1009 (.L_HI(net1009));
 sg13g2_tiehi _14885__1010 (.L_HI(net1010));
 sg13g2_tiehi _14886__1011 (.L_HI(net1011));
 sg13g2_tiehi _14887__1012 (.L_HI(net1012));
 sg13g2_tiehi _14888__1013 (.L_HI(net1013));
 sg13g2_tiehi _14889__1014 (.L_HI(net1014));
 sg13g2_tiehi _14890__1015 (.L_HI(net1015));
 sg13g2_tiehi _14891__1016 (.L_HI(net1016));
 sg13g2_tiehi _14892__1017 (.L_HI(net1017));
 sg13g2_tiehi _14893__1018 (.L_HI(net1018));
 sg13g2_tiehi _14894__1019 (.L_HI(net1019));
 sg13g2_tiehi _14895__1020 (.L_HI(net1020));
 sg13g2_tiehi _14896__1021 (.L_HI(net1021));
 sg13g2_tiehi _14897__1022 (.L_HI(net1022));
 sg13g2_tiehi _14898__1023 (.L_HI(net1023));
 sg13g2_tiehi _14899__1024 (.L_HI(net1024));
 sg13g2_tiehi _14900__1025 (.L_HI(net1025));
 sg13g2_tiehi _14901__1026 (.L_HI(net1026));
 sg13g2_tiehi _14902__1027 (.L_HI(net1027));
 sg13g2_tiehi _14903__1028 (.L_HI(net1028));
 sg13g2_tiehi _14904__1029 (.L_HI(net1029));
 sg13g2_tiehi _14905__1030 (.L_HI(net1030));
 sg13g2_tiehi _14906__1031 (.L_HI(net1031));
 sg13g2_tiehi _14907__1032 (.L_HI(net1032));
 sg13g2_tiehi _14908__1033 (.L_HI(net1033));
 sg13g2_tiehi _14909__1034 (.L_HI(net1034));
 sg13g2_tiehi _14910__1035 (.L_HI(net1035));
 sg13g2_tiehi _14911__1036 (.L_HI(net1036));
 sg13g2_tiehi _14912__1037 (.L_HI(net1037));
 sg13g2_tiehi _14913__1038 (.L_HI(net1038));
 sg13g2_tiehi _14914__1039 (.L_HI(net1039));
 sg13g2_tiehi _14915__1040 (.L_HI(net1040));
 sg13g2_tiehi _14916__1041 (.L_HI(net1041));
 sg13g2_tiehi _14917__1042 (.L_HI(net1042));
 sg13g2_tiehi _14918__1043 (.L_HI(net1043));
 sg13g2_tiehi _14919__1044 (.L_HI(net1044));
 sg13g2_tiehi _14920__1045 (.L_HI(net1045));
 sg13g2_tiehi _14921__1046 (.L_HI(net1046));
 sg13g2_tiehi _14922__1047 (.L_HI(net1047));
 sg13g2_tiehi _14923__1048 (.L_HI(net1048));
 sg13g2_tiehi _14924__1049 (.L_HI(net1049));
 sg13g2_tiehi _14925__1050 (.L_HI(net1050));
 sg13g2_tiehi _14926__1051 (.L_HI(net1051));
 sg13g2_tiehi _14927__1052 (.L_HI(net1052));
 sg13g2_tiehi _14928__1053 (.L_HI(net1053));
 sg13g2_tiehi _14929__1054 (.L_HI(net1054));
 sg13g2_tiehi _14930__1055 (.L_HI(net1055));
 sg13g2_tiehi _14931__1056 (.L_HI(net1056));
 sg13g2_tiehi _14932__1057 (.L_HI(net1057));
 sg13g2_tiehi _14933__1058 (.L_HI(net1058));
 sg13g2_tiehi _14934__1059 (.L_HI(net1059));
 sg13g2_tiehi _14935__1060 (.L_HI(net1060));
 sg13g2_tiehi _14936__1061 (.L_HI(net1061));
 sg13g2_tiehi _14937__1062 (.L_HI(net1062));
 sg13g2_tiehi _14938__1063 (.L_HI(net1063));
 sg13g2_tiehi _14939__1064 (.L_HI(net1064));
 sg13g2_tiehi _14940__1065 (.L_HI(net1065));
 sg13g2_tiehi _14941__1066 (.L_HI(net1066));
 sg13g2_tiehi _14942__1067 (.L_HI(net1067));
 sg13g2_tiehi _14943__1068 (.L_HI(net1068));
 sg13g2_tiehi _14944__1069 (.L_HI(net1069));
 sg13g2_tiehi _14945__1070 (.L_HI(net1070));
 sg13g2_tiehi _14946__1071 (.L_HI(net1071));
 sg13g2_tiehi _14947__1072 (.L_HI(net1072));
 sg13g2_tiehi _14948__1073 (.L_HI(net1073));
 sg13g2_tiehi _14949__1074 (.L_HI(net1074));
 sg13g2_tiehi _14950__1075 (.L_HI(net1075));
 sg13g2_tiehi _14951__1076 (.L_HI(net1076));
 sg13g2_tiehi _14952__1077 (.L_HI(net1077));
 sg13g2_tiehi _14953__1078 (.L_HI(net1078));
 sg13g2_tiehi _14954__1079 (.L_HI(net1079));
 sg13g2_tiehi _14955__1080 (.L_HI(net1080));
 sg13g2_tiehi _14956__1081 (.L_HI(net1081));
 sg13g2_tiehi _14957__1082 (.L_HI(net1082));
 sg13g2_tiehi _14958__1083 (.L_HI(net1083));
 sg13g2_tiehi _14959__1084 (.L_HI(net1084));
 sg13g2_tiehi _14960__1085 (.L_HI(net1085));
 sg13g2_tiehi _14961__1086 (.L_HI(net1086));
 sg13g2_tiehi _14962__1087 (.L_HI(net1087));
 sg13g2_tiehi _14963__1088 (.L_HI(net1088));
 sg13g2_tiehi _14964__1089 (.L_HI(net1089));
 sg13g2_tiehi _14965__1090 (.L_HI(net1090));
 sg13g2_tiehi _14966__1091 (.L_HI(net1091));
 sg13g2_tiehi _14967__1092 (.L_HI(net1092));
 sg13g2_tiehi _14968__1093 (.L_HI(net1093));
 sg13g2_tiehi _14969__1094 (.L_HI(net1094));
 sg13g2_tiehi _14970__1095 (.L_HI(net1095));
 sg13g2_tiehi _14971__1096 (.L_HI(net1096));
 sg13g2_tiehi _14972__1097 (.L_HI(net1097));
 sg13g2_tiehi _14973__1098 (.L_HI(net1098));
 sg13g2_tiehi _14974__1099 (.L_HI(net1099));
 sg13g2_tiehi _14975__1100 (.L_HI(net1100));
 sg13g2_tiehi _14976__1101 (.L_HI(net1101));
 sg13g2_tiehi _14977__1102 (.L_HI(net1102));
 sg13g2_tiehi _14978__1103 (.L_HI(net1103));
 sg13g2_tiehi _14979__1104 (.L_HI(net1104));
 sg13g2_tiehi _14980__1105 (.L_HI(net1105));
 sg13g2_tiehi _14981__1106 (.L_HI(net1106));
 sg13g2_tiehi _14982__1107 (.L_HI(net1107));
 sg13g2_tiehi _14983__1108 (.L_HI(net1108));
 sg13g2_tiehi _14984__1109 (.L_HI(net1109));
 sg13g2_tiehi _14985__1110 (.L_HI(net1110));
 sg13g2_tiehi _14986__1111 (.L_HI(net1111));
 sg13g2_tiehi _14987__1112 (.L_HI(net1112));
 sg13g2_tiehi _14988__1113 (.L_HI(net1113));
 sg13g2_tiehi _14989__1114 (.L_HI(net1114));
 sg13g2_tiehi _14990__1115 (.L_HI(net1115));
 sg13g2_tiehi _14991__1116 (.L_HI(net1116));
 sg13g2_tiehi _14992__1117 (.L_HI(net1117));
 sg13g2_tiehi _14993__1118 (.L_HI(net1118));
 sg13g2_tiehi _14994__1119 (.L_HI(net1119));
 sg13g2_tiehi _14995__1120 (.L_HI(net1120));
 sg13g2_tiehi _14996__1121 (.L_HI(net1121));
 sg13g2_tiehi _14997__1122 (.L_HI(net1122));
 sg13g2_tiehi _14998__1123 (.L_HI(net1123));
 sg13g2_tiehi _14999__1124 (.L_HI(net1124));
 sg13g2_tiehi _15000__1125 (.L_HI(net1125));
 sg13g2_tiehi _15001__1126 (.L_HI(net1126));
 sg13g2_tiehi _15002__1127 (.L_HI(net1127));
 sg13g2_tiehi _15003__1128 (.L_HI(net1128));
 sg13g2_tiehi _15004__1129 (.L_HI(net1129));
 sg13g2_tiehi _15005__1130 (.L_HI(net1130));
 sg13g2_tiehi _15758__1131 (.L_HI(net1131));
 sg13g2_tiehi _15274__1132 (.L_HI(net1132));
 sg13g2_tiehi _15757__1133 (.L_HI(net1133));
 sg13g2_tiehi _15273__1134 (.L_HI(net1134));
 sg13g2_tiehi _15756__1135 (.L_HI(net1135));
 sg13g2_tiehi _15272__1136 (.L_HI(net1136));
 sg13g2_tiehi _15755__1137 (.L_HI(net1137));
 sg13g2_tiehi _15006__1138 (.L_HI(net1138));
 sg13g2_tiehi _15271__1139 (.L_HI(net1139));
 sg13g2_tiehi _15754__1140 (.L_HI(net1140));
 sg13g2_tiehi _15270__1141 (.L_HI(net1141));
 sg13g2_tiehi _15753__1142 (.L_HI(net1142));
 sg13g2_tiehi _15269__1143 (.L_HI(net1143));
 sg13g2_tiehi _15752__1144 (.L_HI(net1144));
 sg13g2_tiehi _15268__1145 (.L_HI(net1145));
 sg13g2_tiehi _15751__1146 (.L_HI(net1146));
 sg13g2_tiehi _15267__1147 (.L_HI(net1147));
 sg13g2_tiehi _15750__1148 (.L_HI(net1148));
 sg13g2_tiehi _15266__1149 (.L_HI(net1149));
 sg13g2_tiehi _15749__1150 (.L_HI(net1150));
 sg13g2_tiehi _15265__1151 (.L_HI(net1151));
 sg13g2_tiehi _15748__1152 (.L_HI(net1152));
 sg13g2_tiehi _15264__1153 (.L_HI(net1153));
 sg13g2_tiehi _15747__1154 (.L_HI(net1154));
 sg13g2_tiehi _15263__1155 (.L_HI(net1155));
 sg13g2_tiehi _15746__1156 (.L_HI(net1156));
 sg13g2_tiehi _15262__1157 (.L_HI(net1157));
 sg13g2_tiehi _15014__1158 (.L_HI(net1158));
 sg13g2_tiehi _15034__1159 (.L_HI(net1159));
 sg13g2_tiehi _15035__1160 (.L_HI(net1160));
 sg13g2_tiehi _15036__1161 (.L_HI(net1161));
 sg13g2_tiehi _15037__1162 (.L_HI(net1162));
 sg13g2_tiehi _15745__1163 (.L_HI(net1163));
 sg13g2_tiehi _15261__1164 (.L_HI(net1164));
 sg13g2_tiehi _15744__1165 (.L_HI(net1165));
 sg13g2_tiehi _15260__1166 (.L_HI(net1166));
 sg13g2_tiehi _15977__1167 (.L_HI(net1167));
 sg13g2_tiehi _15259__1168 (.L_HI(net1168));
 sg13g2_tiehi _15743__1169 (.L_HI(net1169));
 sg13g2_tiehi _15258__1170 (.L_HI(net1170));
 sg13g2_tiehi _15916__1171 (.L_HI(net1171));
 sg13g2_tiehi _15257__1172 (.L_HI(net1172));
 sg13g2_tiehi _15742__1173 (.L_HI(net1173));
 sg13g2_tiehi _15256__1174 (.L_HI(net1174));
 sg13g2_tiehi _15741__1175 (.L_HI(net1175));
 sg13g2_tiehi _15255__1176 (.L_HI(net1176));
 sg13g2_tiehi _15740__1177 (.L_HI(net1177));
 sg13g2_tiehi _15254__1178 (.L_HI(net1178));
 sg13g2_tiehi _15739__1179 (.L_HI(net1179));
 sg13g2_tiehi _15253__1180 (.L_HI(net1180));
 sg13g2_tiehi _15738__1181 (.L_HI(net1181));
 sg13g2_tiehi _15252__1182 (.L_HI(net1182));
 sg13g2_tiehi _15976__1183 (.L_HI(net1183));
 sg13g2_tiehi _15251__1184 (.L_HI(net1184));
 sg13g2_tiehi _15737__1185 (.L_HI(net1185));
 sg13g2_tiehi _15250__1186 (.L_HI(net1186));
 sg13g2_tiehi _15735__1187 (.L_HI(net1187));
 sg13g2_tiehi _15249__1188 (.L_HI(net1188));
 sg13g2_tiehi _15722__1189 (.L_HI(net1189));
 sg13g2_tiehi _15248__1190 (.L_HI(net1190));
 sg13g2_tiehi _15721__1191 (.L_HI(net1191));
 sg13g2_tiehi _15247__1192 (.L_HI(net1192));
 sg13g2_tiehi _15246__1193 (.L_HI(net1193));
 sg13g2_tiehi _15720__1194 (.L_HI(net1194));
 sg13g2_tiehi _15245__1195 (.L_HI(net1195));
 sg13g2_tiehi _15719__1196 (.L_HI(net1196));
 sg13g2_tiehi _15718__1197 (.L_HI(net1197));
 sg13g2_tiehi _15717__1198 (.L_HI(net1198));
 sg13g2_tiehi _15716__1199 (.L_HI(net1199));
 sg13g2_tiehi _15715__1200 (.L_HI(net1200));
 sg13g2_tiehi _15714__1201 (.L_HI(net1201));
 sg13g2_tiehi _15713__1202 (.L_HI(net1202));
 sg13g2_tiehi _15712__1203 (.L_HI(net1203));
 sg13g2_tiehi _15711__1204 (.L_HI(net1204));
 sg13g2_tiehi _15710__1205 (.L_HI(net1205));
 sg13g2_tiehi _15709__1206 (.L_HI(net1206));
 sg13g2_tiehi _15708__1207 (.L_HI(net1207));
 sg13g2_tiehi _15707__1208 (.L_HI(net1208));
 sg13g2_tiehi _15706__1209 (.L_HI(net1209));
 sg13g2_tiehi _15705__1210 (.L_HI(net1210));
 sg13g2_tiehi _15704__1211 (.L_HI(net1211));
 sg13g2_tiehi _15703__1212 (.L_HI(net1212));
 sg13g2_tiehi _15702__1213 (.L_HI(net1213));
 sg13g2_tiehi _15701__1214 (.L_HI(net1214));
 sg13g2_tiehi _15700__1215 (.L_HI(net1215));
 sg13g2_tiehi _15915__1216 (.L_HI(net1216));
 sg13g2_tiehi _15699__1217 (.L_HI(net1217));
 sg13g2_tiehi _15975__1218 (.L_HI(net1218));
 sg13g2_tiehi _15698__1219 (.L_HI(net1219));
 sg13g2_tiehi _15220__1220 (.L_HI(net1220));
 sg13g2_tiehi _15219__1221 (.L_HI(net1221));
 sg13g2_tiehi _15697__1222 (.L_HI(net1222));
 sg13g2_tiehi _15218__1223 (.L_HI(net1223));
 sg13g2_tiehi _15696__1224 (.L_HI(net1224));
 sg13g2_tiehi _15216__1225 (.L_HI(net1225));
 sg13g2_tiehi _15695__1226 (.L_HI(net1226));
 sg13g2_tiehi _15215__1227 (.L_HI(net1227));
 sg13g2_tiehi _15694__1228 (.L_HI(net1228));
 sg13g2_tiehi _15214__1229 (.L_HI(net1229));
 sg13g2_tiehi _15693__1230 (.L_HI(net1230));
 sg13g2_tiehi _15213__1231 (.L_HI(net1231));
 sg13g2_tiehi _15692__1232 (.L_HI(net1232));
 sg13g2_tiehi _15212__1233 (.L_HI(net1233));
 sg13g2_tiehi _15691__1234 (.L_HI(net1234));
 sg13g2_tiehi _15211__1235 (.L_HI(net1235));
 sg13g2_tiehi _15690__1236 (.L_HI(net1236));
 sg13g2_tiehi _15210__1237 (.L_HI(net1237));
 sg13g2_tiehi _15689__1238 (.L_HI(net1238));
 sg13g2_tiehi _15209__1239 (.L_HI(net1239));
 sg13g2_tiehi _15688__1240 (.L_HI(net1240));
 sg13g2_tiehi _15208__1241 (.L_HI(net1241));
 sg13g2_tiehi _15687__1242 (.L_HI(net1242));
 sg13g2_tiehi _15207__1243 (.L_HI(net1243));
 sg13g2_tiehi _15686__1244 (.L_HI(net1244));
 sg13g2_tiehi _15206__1245 (.L_HI(net1245));
 sg13g2_tiehi _15685__1246 (.L_HI(net1246));
 sg13g2_tiehi _15205__1247 (.L_HI(net1247));
 sg13g2_tiehi _15684__1248 (.L_HI(net1248));
 sg13g2_tiehi _15204__1249 (.L_HI(net1249));
 sg13g2_tiehi _15683__1250 (.L_HI(net1250));
 sg13g2_tiehi _15203__1251 (.L_HI(net1251));
 sg13g2_tiehi _15682__1252 (.L_HI(net1252));
 sg13g2_tiehi _15202__1253 (.L_HI(net1253));
 sg13g2_tiehi _15681__1254 (.L_HI(net1254));
 sg13g2_tiehi _15201__1255 (.L_HI(net1255));
 sg13g2_tiehi _15680__1256 (.L_HI(net1256));
 sg13g2_tiehi _15200__1257 (.L_HI(net1257));
 sg13g2_tiehi _15679__1258 (.L_HI(net1258));
 sg13g2_tiehi _15199__1259 (.L_HI(net1259));
 sg13g2_tiehi _15678__1260 (.L_HI(net1260));
 sg13g2_tiehi _15198__1261 (.L_HI(net1261));
 sg13g2_tiehi _15677__1262 (.L_HI(net1262));
 sg13g2_tiehi _15038__1263 (.L_HI(net1263));
 sg13g2_tiehi _15197__1264 (.L_HI(net1264));
 sg13g2_tiehi _15676__1265 (.L_HI(net1265));
 sg13g2_tiehi _15196__1266 (.L_HI(net1266));
 sg13g2_tiehi _15675__1267 (.L_HI(net1267));
 sg13g2_tiehi _15195__1268 (.L_HI(net1268));
 sg13g2_tiehi _15674__1269 (.L_HI(net1269));
 sg13g2_tiehi _15194__1270 (.L_HI(net1270));
 sg13g2_tiehi _15673__1271 (.L_HI(net1271));
 sg13g2_tiehi _15193__1272 (.L_HI(net1272));
 sg13g2_tiehi _15672__1273 (.L_HI(net1273));
 sg13g2_tiehi _15192__1274 (.L_HI(net1274));
 sg13g2_tiehi _15671__1275 (.L_HI(net1275));
 sg13g2_tiehi _15191__1276 (.L_HI(net1276));
 sg13g2_tiehi _15670__1277 (.L_HI(net1277));
 sg13g2_tiehi _15190__1278 (.L_HI(net1278));
 sg13g2_tiehi _15669__1279 (.L_HI(net1279));
 sg13g2_tiehi _15189__1280 (.L_HI(net1280));
 sg13g2_tiehi _15668__1281 (.L_HI(net1281));
 sg13g2_tiehi _15188__1282 (.L_HI(net1282));
 sg13g2_tiehi _15667__1283 (.L_HI(net1283));
 sg13g2_tiehi _15187__1284 (.L_HI(net1284));
 sg13g2_tiehi _15666__1285 (.L_HI(net1285));
 sg13g2_tiehi _15186__1286 (.L_HI(net1286));
 sg13g2_tiehi _15665__1287 (.L_HI(net1287));
 sg13g2_tiehi _15185__1288 (.L_HI(net1288));
 sg13g2_tiehi _15664__1289 (.L_HI(net1289));
 sg13g2_tiehi _15184__1290 (.L_HI(net1290));
 sg13g2_tiehi _15663__1291 (.L_HI(net1291));
 sg13g2_tiehi _15183__1292 (.L_HI(net1292));
 sg13g2_tiehi _15662__1293 (.L_HI(net1293));
 sg13g2_tiehi _15182__1294 (.L_HI(net1294));
 sg13g2_tiehi _15661__1295 (.L_HI(net1295));
 sg13g2_tiehi _15181__1296 (.L_HI(net1296));
 sg13g2_tiehi _15180__1297 (.L_HI(net1297));
 sg13g2_tiehi _15179__1298 (.L_HI(net1298));
 sg13g2_tiehi _15178__1299 (.L_HI(net1299));
 sg13g2_tiehi _15177__1300 (.L_HI(net1300));
 sg13g2_tiehi _15176__1301 (.L_HI(net1301));
 sg13g2_tiehi _15175__1302 (.L_HI(net1302));
 sg13g2_tiehi _15174__1303 (.L_HI(net1303));
 sg13g2_tiehi _15173__1304 (.L_HI(net1304));
 sg13g2_tiehi _15172__1305 (.L_HI(net1305));
 sg13g2_tiehi _15171__1306 (.L_HI(net1306));
 sg13g2_tiehi _15170__1307 (.L_HI(net1307));
 sg13g2_tiehi _15169__1308 (.L_HI(net1308));
 sg13g2_tiehi _15168__1309 (.L_HI(net1309));
 sg13g2_tiehi _15167__1310 (.L_HI(net1310));
 sg13g2_tiehi _15166__1311 (.L_HI(net1311));
 sg13g2_tiehi _15165__1312 (.L_HI(net1312));
 sg13g2_tiehi _15660__1313 (.L_HI(net1313));
 sg13g2_tiehi _15164__1314 (.L_HI(net1314));
 sg13g2_tiehi _15659__1315 (.L_HI(net1315));
 sg13g2_tiehi _15162__1316 (.L_HI(net1316));
 sg13g2_tiehi _15163__1317 (.L_HI(net1317));
 sg13g2_tiehi _15658__1318 (.L_HI(net1318));
 sg13g2_tiehi _15161__1319 (.L_HI(net1319));
 sg13g2_tiehi _15657__1320 (.L_HI(net1320));
 sg13g2_tiehi _15160__1321 (.L_HI(net1321));
 sg13g2_tiehi _15656__1322 (.L_HI(net1322));
 sg13g2_tiehi _15159__1323 (.L_HI(net1323));
 sg13g2_tiehi _15655__1324 (.L_HI(net1324));
 sg13g2_tiehi _15158__1325 (.L_HI(net1325));
 sg13g2_tiehi _15654__1326 (.L_HI(net1326));
 sg13g2_tiehi _15157__1327 (.L_HI(net1327));
 sg13g2_tiehi _15653__1328 (.L_HI(net1328));
 sg13g2_tiehi _15156__1329 (.L_HI(net1329));
 sg13g2_tiehi _15155__1330 (.L_HI(net1330));
 sg13g2_tiehi _15154__1331 (.L_HI(net1331));
 sg13g2_tiehi _15153__1332 (.L_HI(net1332));
 sg13g2_tiehi _15152__1333 (.L_HI(net1333));
 sg13g2_tiehi _15151__1334 (.L_HI(net1334));
 sg13g2_tiehi _15150__1335 (.L_HI(net1335));
 sg13g2_tiehi _15149__1336 (.L_HI(net1336));
 sg13g2_tiehi _15148__1337 (.L_HI(net1337));
 sg13g2_tiehi _15652__1338 (.L_HI(net1338));
 sg13g2_tiehi _15147__1339 (.L_HI(net1339));
 sg13g2_tiehi _15651__1340 (.L_HI(net1340));
 sg13g2_tiehi _15146__1341 (.L_HI(net1341));
 sg13g2_tiehi _15650__1342 (.L_HI(net1342));
 sg13g2_tiehi _15145__1343 (.L_HI(net1343));
 sg13g2_tiehi _15649__1344 (.L_HI(net1344));
 sg13g2_tiehi _15144__1345 (.L_HI(net1345));
 sg13g2_tiehi _15648__1346 (.L_HI(net1346));
 sg13g2_tiehi _15143__1347 (.L_HI(net1347));
 sg13g2_tiehi _15647__1348 (.L_HI(net1348));
 sg13g2_tiehi _15142__1349 (.L_HI(net1349));
 sg13g2_tiehi _15646__1350 (.L_HI(net1350));
 sg13g2_tiehi _15141__1351 (.L_HI(net1351));
 sg13g2_tiehi _15645__1352 (.L_HI(net1352));
 sg13g2_tiehi _15140__1353 (.L_HI(net1353));
 sg13g2_tiehi _15644__1354 (.L_HI(net1354));
 sg13g2_tiehi _15139__1355 (.L_HI(net1355));
 sg13g2_tiehi _15643__1356 (.L_HI(net1356));
 sg13g2_tiehi _15138__1357 (.L_HI(net1357));
 sg13g2_tiehi _15137__1358 (.L_HI(net1358));
 sg13g2_tiehi _15136__1359 (.L_HI(net1359));
 sg13g2_tiehi _15642__1360 (.L_HI(net1360));
 sg13g2_tiehi _15135__1361 (.L_HI(net1361));
 sg13g2_tiehi _15641__1362 (.L_HI(net1362));
 sg13g2_tiehi _15134__1363 (.L_HI(net1363));
 sg13g2_tiehi _15640__1364 (.L_HI(net1364));
 sg13g2_tiehi _15133__1365 (.L_HI(net1365));
 sg13g2_tiehi _15639__1366 (.L_HI(net1366));
 sg13g2_tiehi _15132__1367 (.L_HI(net1367));
 sg13g2_tiehi _15131__1368 (.L_HI(net1368));
 sg13g2_tiehi _15638__1369 (.L_HI(net1369));
 sg13g2_tiehi _15130__1370 (.L_HI(net1370));
 sg13g2_tiehi _15637__1371 (.L_HI(net1371));
 sg13g2_tiehi _15129__1372 (.L_HI(net1372));
 sg13g2_tiehi _15636__1373 (.L_HI(net1373));
 sg13g2_tiehi _15128__1374 (.L_HI(net1374));
 sg13g2_tiehi _15635__1375 (.L_HI(net1375));
 sg13g2_tiehi _15127__1376 (.L_HI(net1376));
 sg13g2_tiehi _15126__1377 (.L_HI(net1377));
 sg13g2_tiehi _15634__1378 (.L_HI(net1378));
 sg13g2_tiehi _15125__1379 (.L_HI(net1379));
 sg13g2_tiehi _15633__1380 (.L_HI(net1380));
 sg13g2_tiehi _15124__1381 (.L_HI(net1381));
 sg13g2_tiehi _15632__1382 (.L_HI(net1382));
 sg13g2_tiehi _15123__1383 (.L_HI(net1383));
 sg13g2_tiehi _15631__1384 (.L_HI(net1384));
 sg13g2_tiehi _15122__1385 (.L_HI(net1385));
 sg13g2_tiehi _15630__1386 (.L_HI(net1386));
 sg13g2_tiehi _15121__1387 (.L_HI(net1387));
 sg13g2_tiehi _15914__1388 (.L_HI(net1388));
 sg13g2_tiehi _15120__1389 (.L_HI(net1389));
 sg13g2_tiehi _15629__1390 (.L_HI(net1390));
 sg13g2_tiehi _15119__1391 (.L_HI(net1391));
 sg13g2_tiehi _15974__1392 (.L_HI(net1392));
 sg13g2_tiehi _15118__1393 (.L_HI(net1393));
 sg13g2_tiehi _15628__1394 (.L_HI(net1394));
 sg13g2_tiehi _15117__1395 (.L_HI(net1395));
 sg13g2_tiehi _15913__1396 (.L_HI(net1396));
 sg13g2_tiehi _15116__1397 (.L_HI(net1397));
 sg13g2_tiehi _15627__1398 (.L_HI(net1398));
 sg13g2_tiehi _15115__1399 (.L_HI(net1399));
 sg13g2_tiehi _15973__1400 (.L_HI(net1400));
 sg13g2_tiehi _15114__1401 (.L_HI(net1401));
 sg13g2_tiehi _15626__1402 (.L_HI(net1402));
 sg13g2_tiehi _15113__1403 (.L_HI(net1403));
 sg13g2_tiehi _15625__1404 (.L_HI(net1404));
 sg13g2_tiehi _15112__1405 (.L_HI(net1405));
 sg13g2_tiehi _15624__1406 (.L_HI(net1406));
 sg13g2_tiehi _15111__1407 (.L_HI(net1407));
 sg13g2_tiehi _15623__1408 (.L_HI(net1408));
 sg13g2_tiehi _15110__1409 (.L_HI(net1409));
 sg13g2_tiehi _15622__1410 (.L_HI(net1410));
 sg13g2_tiehi _15109__1411 (.L_HI(net1411));
 sg13g2_tiehi _15108__1412 (.L_HI(net1412));
 sg13g2_tiehi _15107__1413 (.L_HI(net1413));
 sg13g2_tiehi _15106__1414 (.L_HI(net1414));
 sg13g2_tiehi _15105__1415 (.L_HI(net1415));
 sg13g2_tiehi _15104__1416 (.L_HI(net1416));
 sg13g2_tiehi _15103__1417 (.L_HI(net1417));
 sg13g2_tiehi _15102__1418 (.L_HI(net1418));
 sg13g2_tiehi _15101__1419 (.L_HI(net1419));
 sg13g2_tiehi _15100__1420 (.L_HI(net1420));
 sg13g2_tiehi _15099__1421 (.L_HI(net1421));
 sg13g2_tiehi _15098__1422 (.L_HI(net1422));
 sg13g2_tiehi _15097__1423 (.L_HI(net1423));
 sg13g2_tiehi _15096__1424 (.L_HI(net1424));
 sg13g2_tiehi _15095__1425 (.L_HI(net1425));
 sg13g2_tiehi _15094__1426 (.L_HI(net1426));
 sg13g2_tiehi _15093__1427 (.L_HI(net1427));
 sg13g2_tiehi _15092__1428 (.L_HI(net1428));
 sg13g2_tiehi _15091__1429 (.L_HI(net1429));
 sg13g2_tiehi _15090__1430 (.L_HI(net1430));
 sg13g2_tiehi _15621__1431 (.L_HI(net1431));
 sg13g2_tiehi _15089__1432 (.L_HI(net1432));
 sg13g2_tiehi _15620__1433 (.L_HI(net1433));
 sg13g2_tiehi _15088__1434 (.L_HI(net1434));
 sg13g2_tiehi _15619__1435 (.L_HI(net1435));
 sg13g2_tiehi _15087__1436 (.L_HI(net1436));
 sg13g2_tiehi _15618__1437 (.L_HI(net1437));
 sg13g2_tiehi _15086__1438 (.L_HI(net1438));
 sg13g2_tiehi _15085__1439 (.L_HI(net1439));
 sg13g2_tiehi _15617__1440 (.L_HI(net1440));
 sg13g2_tiehi _15084__1441 (.L_HI(net1441));
 sg13g2_tiehi _15083__1442 (.L_HI(net1442));
 sg13g2_tiehi _15082__1443 (.L_HI(net1443));
 sg13g2_tiehi _15081__1444 (.L_HI(net1444));
 sg13g2_tiehi _15080__1445 (.L_HI(net1445));
 sg13g2_tiehi _15079__1446 (.L_HI(net1446));
 sg13g2_tiehi _15078__1447 (.L_HI(net1447));
 sg13g2_tiehi _15077__1448 (.L_HI(net1448));
 sg13g2_tiehi _15076__1449 (.L_HI(net1449));
 sg13g2_tiehi _15075__1450 (.L_HI(net1450));
 sg13g2_tiehi _15074__1451 (.L_HI(net1451));
 sg13g2_tiehi _15073__1452 (.L_HI(net1452));
 sg13g2_tiehi _15616__1453 (.L_HI(net1453));
 sg13g2_tiehi _15072__1454 (.L_HI(net1454));
 sg13g2_tiehi _15615__1455 (.L_HI(net1455));
 sg13g2_tiehi _15071__1456 (.L_HI(net1456));
 sg13g2_tiehi _15070__1457 (.L_HI(net1457));
 sg13g2_tiehi _15069__1458 (.L_HI(net1458));
 sg13g2_tiehi _15068__1459 (.L_HI(net1459));
 sg13g2_tiehi _15067__1460 (.L_HI(net1460));
 sg13g2_tiehi _15066__1461 (.L_HI(net1461));
 sg13g2_tiehi _15065__1462 (.L_HI(net1462));
 sg13g2_tiehi _15064__1463 (.L_HI(net1463));
 sg13g2_tiehi _15063__1464 (.L_HI(net1464));
 sg13g2_tiehi _15614__1465 (.L_HI(net1465));
 sg13g2_tiehi _15062__1466 (.L_HI(net1466));
 sg13g2_tiehi _15613__1467 (.L_HI(net1467));
 sg13g2_tiehi _15061__1468 (.L_HI(net1468));
 sg13g2_tiehi _15612__1469 (.L_HI(net1469));
 sg13g2_tiehi _15060__1470 (.L_HI(net1470));
 sg13g2_tiehi _15611__1471 (.L_HI(net1471));
 sg13g2_tiehi _15059__1472 (.L_HI(net1472));
 sg13g2_tiehi _15610__1473 (.L_HI(net1473));
 sg13g2_tiehi _15058__1474 (.L_HI(net1474));
 sg13g2_tiehi _15609__1475 (.L_HI(net1475));
 sg13g2_tiehi _15057__1476 (.L_HI(net1476));
 sg13g2_tiehi _15608__1477 (.L_HI(net1477));
 sg13g2_tiehi _15056__1478 (.L_HI(net1478));
 sg13g2_tiehi _15607__1479 (.L_HI(net1479));
 sg13g2_tiehi _15055__1480 (.L_HI(net1480));
 sg13g2_tiehi _15606__1481 (.L_HI(net1481));
 sg13g2_tiehi _15054__1482 (.L_HI(net1482));
 sg13g2_tiehi _15605__1483 (.L_HI(net1483));
 sg13g2_tiehi _15053__1484 (.L_HI(net1484));
 sg13g2_tiehi _15604__1485 (.L_HI(net1485));
 sg13g2_tiehi _15052__1486 (.L_HI(net1486));
 sg13g2_tiehi _15603__1487 (.L_HI(net1487));
 sg13g2_tiehi _15051__1488 (.L_HI(net1488));
 sg13g2_tiehi _15602__1489 (.L_HI(net1489));
 sg13g2_tiehi _15050__1490 (.L_HI(net1490));
 sg13g2_tiehi _15601__1491 (.L_HI(net1491));
 sg13g2_tiehi _15049__1492 (.L_HI(net1492));
 sg13g2_tiehi _15600__1493 (.L_HI(net1493));
 sg13g2_tiehi _15048__1494 (.L_HI(net1494));
 sg13g2_tiehi _15599__1495 (.L_HI(net1495));
 sg13g2_tiehi _15047__1496 (.L_HI(net1496));
 sg13g2_tiehi _15598__1497 (.L_HI(net1497));
 sg13g2_tiehi _15046__1498 (.L_HI(net1498));
 sg13g2_tiehi _15597__1499 (.L_HI(net1499));
 sg13g2_tiehi _15045__1500 (.L_HI(net1500));
 sg13g2_tiehi _15596__1501 (.L_HI(net1501));
 sg13g2_tiehi _15044__1502 (.L_HI(net1502));
 sg13g2_tiehi _15595__1503 (.L_HI(net1503));
 sg13g2_tiehi _15043__1504 (.L_HI(net1504));
 sg13g2_tiehi _15594__1505 (.L_HI(net1505));
 sg13g2_tiehi _15042__1506 (.L_HI(net1506));
 sg13g2_tiehi _15593__1507 (.L_HI(net1507));
 sg13g2_tiehi _15041__1508 (.L_HI(net1508));
 sg13g2_tiehi _15592__1509 (.L_HI(net1509));
 sg13g2_tiehi _15040__1510 (.L_HI(net1510));
 sg13g2_tiehi _15039__1511 (.L_HI(net1511));
 sg13g2_tiehi _15033__1512 (.L_HI(net1512));
 sg13g2_tiehi _15032__1513 (.L_HI(net1513));
 sg13g2_tiehi _15031__1514 (.L_HI(net1514));
 sg13g2_tiehi _15591__1515 (.L_HI(net1515));
 sg13g2_tiehi _15030__1516 (.L_HI(net1516));
 sg13g2_tiehi _15590__1517 (.L_HI(net1517));
 sg13g2_tiehi _15029__1518 (.L_HI(net1518));
 sg13g2_tiehi _15589__1519 (.L_HI(net1519));
 sg13g2_tiehi _15028__1520 (.L_HI(net1520));
 sg13g2_tiehi _15588__1521 (.L_HI(net1521));
 sg13g2_tiehi _15027__1522 (.L_HI(net1522));
 sg13g2_tiehi _15567__1523 (.L_HI(net1523));
 sg13g2_tiehi _15026__1524 (.L_HI(net1524));
 sg13g2_tiehi _15566__1525 (.L_HI(net1525));
 sg13g2_tiehi _15025__1526 (.L_HI(net1526));
 sg13g2_tiehi _15565__1527 (.L_HI(net1527));
 sg13g2_tiehi _15024__1528 (.L_HI(net1528));
 sg13g2_tiehi _15023__1529 (.L_HI(net1529));
 sg13g2_tiehi _15022__1530 (.L_HI(net1530));
 sg13g2_tiehi _15564__1531 (.L_HI(net1531));
 sg13g2_tiehi _15021__1532 (.L_HI(net1532));
 sg13g2_tiehi _15912__1533 (.L_HI(net1533));
 sg13g2_tiehi _15020__1534 (.L_HI(net1534));
 sg13g2_tiehi _15563__1535 (.L_HI(net1535));
 sg13g2_tiehi _15019__1536 (.L_HI(net1536));
 sg13g2_tiehi _15972__1537 (.L_HI(net1537));
 sg13g2_tiehi _15018__1538 (.L_HI(net1538));
 sg13g2_tiehi _15558__1539 (.L_HI(net1539));
 sg13g2_tiehi _15017__1540 (.L_HI(net1540));
 sg13g2_tiehi _15911__1541 (.L_HI(net1541));
 sg13g2_tiehi _15016__1542 (.L_HI(net1542));
 sg13g2_tiehi _15557__1543 (.L_HI(net1543));
 sg13g2_tiehi _15015__1544 (.L_HI(net1544));
 sg13g2_tiehi _15971__1545 (.L_HI(net1545));
 sg13g2_tiehi _15013__1546 (.L_HI(net1546));
 sg13g2_tiehi _15556__1547 (.L_HI(net1547));
 sg13g2_tiehi _15012__1548 (.L_HI(net1548));
 sg13g2_tiehi _15011__1549 (.L_HI(net1549));
 sg13g2_tiehi _15910__1550 (.L_HI(net1550));
 sg13g2_tiehi _15010__1551 (.L_HI(net1551));
 sg13g2_tiehi _15555__1552 (.L_HI(net1552));
 sg13g2_tiehi _15009__1553 (.L_HI(net1553));
 sg13g2_tiehi _15008__1554 (.L_HI(net1554));
 sg13g2_tiehi _15007__1555 (.L_HI(net1555));
 sg13g2_tiehi _14592__1556 (.L_HI(net1556));
 sg13g2_tiehi _14591__1557 (.L_HI(net1557));
 sg13g2_tiehi _14590__1558 (.L_HI(net1558));
 sg13g2_tiehi _14589__1559 (.L_HI(net1559));
 sg13g2_tiehi _14588__1560 (.L_HI(net1560));
 sg13g2_tiehi _14587__1561 (.L_HI(net1561));
 sg13g2_tiehi _14558__1562 (.L_HI(net1562));
 sg13g2_tiehi _14557__1563 (.L_HI(net1563));
 sg13g2_tiehi _14556__1564 (.L_HI(net1564));
 sg13g2_tiehi _14555__1565 (.L_HI(net1565));
 sg13g2_tiehi _15970__1566 (.L_HI(net1566));
 sg13g2_tiehi _15554__1567 (.L_HI(net1567));
 sg13g2_tiehi _15909__1568 (.L_HI(net1568));
 sg13g2_tiehi _15553__1569 (.L_HI(net1569));
 sg13g2_tiehi _15969__1570 (.L_HI(net1570));
 sg13g2_tiehi _15552__1571 (.L_HI(net1571));
 sg13g2_tiehi _15551__1572 (.L_HI(net1572));
 sg13g2_tiehi _15550__1573 (.L_HI(net1573));
 sg13g2_tiehi _15549__1574 (.L_HI(net1574));
 sg13g2_tiehi _15548__1575 (.L_HI(net1575));
 sg13g2_tiehi _15547__1576 (.L_HI(net1576));
 sg13g2_tiehi _15546__1577 (.L_HI(net1577));
 sg13g2_tiehi _15545__1578 (.L_HI(net1578));
 sg13g2_tiehi _15544__1579 (.L_HI(net1579));
 sg13g2_tiehi _15543__1580 (.L_HI(net1580));
 sg13g2_tiehi _15542__1581 (.L_HI(net1581));
 sg13g2_tiehi _15541__1582 (.L_HI(net1582));
 sg13g2_tiehi _15540__1583 (.L_HI(net1583));
 sg13g2_tiehi _15539__1584 (.L_HI(net1584));
 sg13g2_tiehi _15538__1585 (.L_HI(net1585));
 sg13g2_tiehi _15537__1586 (.L_HI(net1586));
 sg13g2_tiehi _15536__1587 (.L_HI(net1587));
 sg13g2_tiehi _15535__1588 (.L_HI(net1588));
 sg13g2_tiehi _15534__1589 (.L_HI(net1589));
 sg13g2_tiehi _15533__1590 (.L_HI(net1590));
 sg13g2_tiehi _15532__1591 (.L_HI(net1591));
 sg13g2_tiehi _15531__1592 (.L_HI(net1592));
 sg13g2_tiehi _15530__1593 (.L_HI(net1593));
 sg13g2_tiehi _15529__1594 (.L_HI(net1594));
 sg13g2_tiehi _15217__1595 (.L_HI(net1595));
 sg13g2_tiehi _15495__1596 (.L_HI(net1596));
 sg13g2_tiehi _15496__1597 (.L_HI(net1597));
 sg13g2_tiehi _15497__1598 (.L_HI(net1598));
 sg13g2_tiehi _15498__1599 (.L_HI(net1599));
 sg13g2_tiehi _15499__1600 (.L_HI(net1600));
 sg13g2_tiehi _15500__1601 (.L_HI(net1601));
 sg13g2_tiehi _15501__1602 (.L_HI(net1602));
 sg13g2_tiehi _15502__1603 (.L_HI(net1603));
 sg13g2_tiehi _15503__1604 (.L_HI(net1604));
 sg13g2_tiehi _15504__1605 (.L_HI(net1605));
 sg13g2_tiehi _15505__1606 (.L_HI(net1606));
 sg13g2_tiehi _15506__1607 (.L_HI(net1607));
 sg13g2_tiehi _15507__1608 (.L_HI(net1608));
 sg13g2_tiehi _15508__1609 (.L_HI(net1609));
 sg13g2_tiehi _15509__1610 (.L_HI(net1610));
 sg13g2_tiehi _15510__1611 (.L_HI(net1611));
 sg13g2_tiehi _15511__1612 (.L_HI(net1612));
 sg13g2_tiehi _15512__1613 (.L_HI(net1613));
 sg13g2_tiehi _15513__1614 (.L_HI(net1614));
 sg13g2_tiehi _15514__1615 (.L_HI(net1615));
 sg13g2_tiehi _15515__1616 (.L_HI(net1616));
 sg13g2_tiehi _15516__1617 (.L_HI(net1617));
 sg13g2_tiehi _15517__1618 (.L_HI(net1618));
 sg13g2_tiehi _15518__1619 (.L_HI(net1619));
 sg13g2_tiehi _15519__1620 (.L_HI(net1620));
 sg13g2_tiehi _15520__1621 (.L_HI(net1621));
 sg13g2_tiehi _15521__1622 (.L_HI(net1622));
 sg13g2_tiehi _15522__1623 (.L_HI(net1623));
 sg13g2_tiehi _15523__1624 (.L_HI(net1624));
 sg13g2_tiehi _15524__1625 (.L_HI(net1625));
 sg13g2_tiehi _15525__1626 (.L_HI(net1626));
 sg13g2_tiehi _15528__1627 (.L_HI(net1627));
 sg13g2_tiehi _15527__1628 (.L_HI(net1628));
 sg13g2_tiehi _15908__1629 (.L_HI(net1629));
 sg13g2_tiehi _15494__1630 (.L_HI(net1630));
 sg13g2_tiehi _15968__1631 (.L_HI(net1631));
 sg13g2_tiehi _15493__1632 (.L_HI(net1632));
 sg13g2_tiehi _15907__1633 (.L_HI(net1633));
 sg13g2_tiehi _15492__1634 (.L_HI(net1634));
 sg13g2_tiehi _15967__1635 (.L_HI(net1635));
 sg13g2_tiehi _15491__1636 (.L_HI(net1636));
 sg13g2_tiehi _15906__1637 (.L_HI(net1637));
 sg13g2_tiehi _15490__1638 (.L_HI(net1638));
 sg13g2_tiehi _15966__1639 (.L_HI(net1639));
 sg13g2_tiehi _15489__1640 (.L_HI(net1640));
 sg13g2_tiehi _15905__1641 (.L_HI(net1641));
 sg13g2_tiehi _15488__1642 (.L_HI(net1642));
 sg13g2_tiehi _15965__1643 (.L_HI(net1643));
 sg13g2_tiehi _15487__1644 (.L_HI(net1644));
 sg13g2_tiehi _15904__1645 (.L_HI(net1645));
 sg13g2_tiehi _15486__1646 (.L_HI(net1646));
 sg13g2_tiehi _15964__1647 (.L_HI(net1647));
 sg13g2_tiehi _15485__1648 (.L_HI(net1648));
 sg13g2_tiehi _15903__1649 (.L_HI(net1649));
 sg13g2_tiehi _15484__1650 (.L_HI(net1650));
 sg13g2_tiehi _15963__1651 (.L_HI(net1651));
 sg13g2_tiehi _15483__1652 (.L_HI(net1652));
 sg13g2_tiehi _15902__1653 (.L_HI(net1653));
 sg13g2_tiehi _15482__1654 (.L_HI(net1654));
 sg13g2_tiehi _15962__1655 (.L_HI(net1655));
 sg13g2_tiehi _15481__1656 (.L_HI(net1656));
 sg13g2_tiehi _15901__1657 (.L_HI(net1657));
 sg13g2_tiehi _15480__1658 (.L_HI(net1658));
 sg13g2_tiehi _15526__1659 (.L_HI(net1659));
 sg13g2_tiehi _15559__1660 (.L_HI(net1660));
 sg13g2_tiehi _15560__1661 (.L_HI(net1661));
 sg13g2_tiehi _15561__1662 (.L_HI(net1662));
 sg13g2_tiehi _15961__1663 (.L_HI(net1663));
 sg13g2_tiehi _15479__1664 (.L_HI(net1664));
 sg13g2_tiehi _15900__1665 (.L_HI(net1665));
 sg13g2_tiehi _15478__1666 (.L_HI(net1666));
 sg13g2_tiehi _15960__1667 (.L_HI(net1667));
 sg13g2_tiehi _15562__1668 (.L_HI(net1668));
 sg13g2_tiehi _15568__1669 (.L_HI(net1669));
 sg13g2_tiehi _15569__1670 (.L_HI(net1670));
 sg13g2_tiehi _15570__1671 (.L_HI(net1671));
 sg13g2_tiehi _15571__1672 (.L_HI(net1672));
 sg13g2_tiehi _15572__1673 (.L_HI(net1673));
 sg13g2_tiehi _15573__1674 (.L_HI(net1674));
 sg13g2_tiehi _15574__1675 (.L_HI(net1675));
 sg13g2_tiehi _15575__1676 (.L_HI(net1676));
 sg13g2_tiehi _15576__1677 (.L_HI(net1677));
 sg13g2_tiehi _15577__1678 (.L_HI(net1678));
 sg13g2_tiehi _15578__1679 (.L_HI(net1679));
 sg13g2_tiehi _15579__1680 (.L_HI(net1680));
 sg13g2_tiehi _15580__1681 (.L_HI(net1681));
 sg13g2_tiehi _15581__1682 (.L_HI(net1682));
 sg13g2_tiehi _15582__1683 (.L_HI(net1683));
 sg13g2_tiehi _15583__1684 (.L_HI(net1684));
 sg13g2_tiehi _15584__1685 (.L_HI(net1685));
 sg13g2_tiehi _15585__1686 (.L_HI(net1686));
 sg13g2_tiehi _15586__1687 (.L_HI(net1687));
 sg13g2_tiehi _15477__1688 (.L_HI(net1688));
 sg13g2_tiehi _15899__1689 (.L_HI(net1689));
 sg13g2_tiehi _15476__1690 (.L_HI(net1690));
 sg13g2_tiehi _15959__1691 (.L_HI(net1691));
 sg13g2_tiehi _15475__1692 (.L_HI(net1692));
 sg13g2_tiehi _15898__1693 (.L_HI(net1693));
 sg13g2_tiehi _15474__1694 (.L_HI(net1694));
 sg13g2_tiehi _15958__1695 (.L_HI(net1695));
 sg13g2_tiehi _15473__1696 (.L_HI(net1696));
 sg13g2_tiehi _15897__1697 (.L_HI(net1697));
 sg13g2_tiehi _15472__1698 (.L_HI(net1698));
 sg13g2_tiehi _15957__1699 (.L_HI(net1699));
 sg13g2_tiehi _15471__1700 (.L_HI(net1700));
 sg13g2_tiehi _15896__1701 (.L_HI(net1701));
 sg13g2_tiehi _15470__1702 (.L_HI(net1702));
 sg13g2_tiehi _15956__1703 (.L_HI(net1703));
 sg13g2_tiehi _15469__1704 (.L_HI(net1704));
 sg13g2_tiehi _15895__1705 (.L_HI(net1705));
 sg13g2_tiehi _15468__1706 (.L_HI(net1706));
 sg13g2_tiehi _15955__1707 (.L_HI(net1707));
 sg13g2_tiehi _15467__1708 (.L_HI(net1708));
 sg13g2_tiehi _15894__1709 (.L_HI(net1709));
 sg13g2_tiehi _15466__1710 (.L_HI(net1710));
 sg13g2_tiehi _15954__1711 (.L_HI(net1711));
 sg13g2_tiehi _15465__1712 (.L_HI(net1712));
 sg13g2_tiehi _15893__1713 (.L_HI(net1713));
 sg13g2_tiehi _15464__1714 (.L_HI(net1714));
 sg13g2_tiehi _15953__1715 (.L_HI(net1715));
 sg13g2_tiehi _15463__1716 (.L_HI(net1716));
 sg13g2_tiehi _15892__1717 (.L_HI(net1717));
 sg13g2_tiehi _15462__1718 (.L_HI(net1718));
 sg13g2_tiehi _15952__1719 (.L_HI(net1719));
 sg13g2_tiehi _15461__1720 (.L_HI(net1720));
 sg13g2_tiehi _15891__1721 (.L_HI(net1721));
 sg13g2_tiehi _15460__1722 (.L_HI(net1722));
 sg13g2_tiehi _15951__1723 (.L_HI(net1723));
 sg13g2_tiehi _15459__1724 (.L_HI(net1724));
 sg13g2_tiehi _15890__1725 (.L_HI(net1725));
 sg13g2_tiehi _15458__1726 (.L_HI(net1726));
 sg13g2_tiehi _15950__1727 (.L_HI(net1727));
 sg13g2_tiehi _15457__1728 (.L_HI(net1728));
 sg13g2_tiehi _15889__1729 (.L_HI(net1729));
 sg13g2_tiehi _15456__1730 (.L_HI(net1730));
 sg13g2_tiehi _15949__1731 (.L_HI(net1731));
 sg13g2_tiehi _15455__1732 (.L_HI(net1732));
 sg13g2_tiehi _15888__1733 (.L_HI(net1733));
 sg13g2_tiehi _15454__1734 (.L_HI(net1734));
 sg13g2_tiehi _15948__1735 (.L_HI(net1735));
 sg13g2_tiehi _15453__1736 (.L_HI(net1736));
 sg13g2_tiehi _15887__1737 (.L_HI(net1737));
 sg13g2_tiehi _15452__1738 (.L_HI(net1738));
 sg13g2_tiehi _15947__1739 (.L_HI(net1739));
 sg13g2_tiehi _15451__1740 (.L_HI(net1740));
 sg13g2_tiehi _15886__1741 (.L_HI(net1741));
 sg13g2_tiehi _15450__1742 (.L_HI(net1742));
 sg13g2_tiehi _15946__1743 (.L_HI(net1743));
 sg13g2_tiehi _15449__1744 (.L_HI(net1744));
 sg13g2_tiehi _15885__1745 (.L_HI(net1745));
 sg13g2_tiehi _15448__1746 (.L_HI(net1746));
 sg13g2_tiehi _15945__1747 (.L_HI(net1747));
 sg13g2_tiehi _15447__1748 (.L_HI(net1748));
 sg13g2_tiehi _15884__1749 (.L_HI(net1749));
 sg13g2_tiehi _15446__1750 (.L_HI(net1750));
 sg13g2_tiehi _15944__1751 (.L_HI(net1751));
 sg13g2_tiehi _15445__1752 (.L_HI(net1752));
 sg13g2_tiehi _15883__1753 (.L_HI(net1753));
 sg13g2_tiehi _15444__1754 (.L_HI(net1754));
 sg13g2_tiehi _15943__1755 (.L_HI(net1755));
 sg13g2_tiehi _15443__1756 (.L_HI(net1756));
 sg13g2_tiehi _15882__1757 (.L_HI(net1757));
 sg13g2_tiehi _15442__1758 (.L_HI(net1758));
 sg13g2_tiehi _15942__1759 (.L_HI(net1759));
 sg13g2_tiehi _15441__1760 (.L_HI(net1760));
 sg13g2_tiehi _15881__1761 (.L_HI(net1761));
 sg13g2_tiehi _15440__1762 (.L_HI(net1762));
 sg13g2_tiehi _15941__1763 (.L_HI(net1763));
 sg13g2_tiehi _15439__1764 (.L_HI(net1764));
 sg13g2_tiehi _15880__1765 (.L_HI(net1765));
 sg13g2_tiehi _15438__1766 (.L_HI(net1766));
 sg13g2_tiehi _15992__1767 (.L_HI(net1767));
 sg13g2_tiehi _15437__1768 (.L_HI(net1768));
 sg13g2_tiehi _15879__1769 (.L_HI(net1769));
 sg13g2_tiehi _15436__1770 (.L_HI(net1770));
 sg13g2_tiehi _15940__1771 (.L_HI(net1771));
 sg13g2_tiehi _15435__1772 (.L_HI(net1772));
 sg13g2_tiehi _15878__1773 (.L_HI(net1773));
 sg13g2_tiehi _15434__1774 (.L_HI(net1774));
 sg13g2_tiehi _15994__1775 (.L_HI(net1775));
 sg13g2_tiehi _15433__1776 (.L_HI(net1776));
 sg13g2_tiehi _15877__1777 (.L_HI(net1777));
 sg13g2_tiehi _15432__1778 (.L_HI(net1778));
 sg13g2_tiehi _15939__1779 (.L_HI(net1779));
 sg13g2_tiehi _15431__1780 (.L_HI(net1780));
 sg13g2_tiehi _15876__1781 (.L_HI(net1781));
 sg13g2_tiehi _15430__1782 (.L_HI(net1782));
 sg13g2_tiehi _15991__1783 (.L_HI(net1783));
 sg13g2_tiehi _15429__1784 (.L_HI(net1784));
 sg13g2_tiehi _15875__1785 (.L_HI(net1785));
 sg13g2_tiehi _15428__1786 (.L_HI(net1786));
 sg13g2_tiehi _15938__1787 (.L_HI(net1787));
 sg13g2_tiehi _15427__1788 (.L_HI(net1788));
 sg13g2_tiehi _15874__1789 (.L_HI(net1789));
 sg13g2_tiehi _15426__1790 (.L_HI(net1790));
 sg13g2_tiehi _15920__1791 (.L_HI(net1791));
 sg13g2_tiehi _15425__1792 (.L_HI(net1792));
 sg13g2_tiehi _15873__1793 (.L_HI(net1793));
 sg13g2_tiehi _15424__1794 (.L_HI(net1794));
 sg13g2_tiehi _15937__1795 (.L_HI(net1795));
 sg13g2_tiehi _15423__1796 (.L_HI(net1796));
 sg13g2_tiehi _15872__1797 (.L_HI(net1797));
 sg13g2_tiehi _15422__1798 (.L_HI(net1798));
 sg13g2_tiehi _15990__1799 (.L_HI(net1799));
 sg13g2_tiehi _15421__1800 (.L_HI(net1800));
 sg13g2_tiehi _15871__1801 (.L_HI(net1801));
 sg13g2_tiehi _15420__1802 (.L_HI(net1802));
 sg13g2_tiehi _15936__1803 (.L_HI(net1803));
 sg13g2_tiehi _15419__1804 (.L_HI(net1804));
 sg13g2_tiehi _15870__1805 (.L_HI(net1805));
 sg13g2_tiehi _15418__1806 (.L_HI(net1806));
 sg13g2_tiehi _15993__1807 (.L_HI(net1807));
 sg13g2_tiehi _15417__1808 (.L_HI(net1808));
 sg13g2_tiehi _15869__1809 (.L_HI(net1809));
 sg13g2_tiehi _15416__1810 (.L_HI(net1810));
 sg13g2_tiehi _15935__1811 (.L_HI(net1811));
 sg13g2_tiehi _15415__1812 (.L_HI(net1812));
 sg13g2_tiehi _15868__1813 (.L_HI(net1813));
 sg13g2_tiehi _15414__1814 (.L_HI(net1814));
 sg13g2_tiehi _15989__1815 (.L_HI(net1815));
 sg13g2_tiehi _15413__1816 (.L_HI(net1816));
 sg13g2_tiehi _15867__1817 (.L_HI(net1817));
 sg13g2_tiehi _15412__1818 (.L_HI(net1818));
 sg13g2_tiehi _15934__1819 (.L_HI(net1819));
 sg13g2_tiehi _15411__1820 (.L_HI(net1820));
 sg13g2_tiehi _15866__1821 (.L_HI(net1821));
 sg13g2_tiehi _15410__1822 (.L_HI(net1822));
 sg13g2_tiehi _15587__1823 (.L_HI(net1823));
 sg13g2_tiehi _15723__1824 (.L_HI(net1824));
 sg13g2_tiehi _15724__1825 (.L_HI(net1825));
 sg13g2_tiehi _15725__1826 (.L_HI(net1826));
 sg13g2_tiehi _15726__1827 (.L_HI(net1827));
 sg13g2_tiehi _15727__1828 (.L_HI(net1828));
 sg13g2_tiehi _15728__1829 (.L_HI(net1829));
 sg13g2_tiehi _15729__1830 (.L_HI(net1830));
 sg13g2_tiehi _15730__1831 (.L_HI(net1831));
 sg13g2_tiehi _15731__1832 (.L_HI(net1832));
 sg13g2_tiehi _15732__1833 (.L_HI(net1833));
 sg13g2_tiehi _15733__1834 (.L_HI(net1834));
 sg13g2_tiehi _15995__1835 (.L_HI(net1835));
 sg13g2_tiehi _15734__1836 (.L_HI(net1836));
 sg13g2_tiehi _15409__1837 (.L_HI(net1837));
 sg13g2_tiehi _15865__1838 (.L_HI(net1838));
 sg13g2_tiehi _15408__1839 (.L_HI(net1839));
 sg13g2_tiehi _15933__1840 (.L_HI(net1840));
 sg13g2_tiehi _15407__1841 (.L_HI(net1841));
 sg13g2_tiehi _15864__1842 (.L_HI(net1842));
 sg13g2_tiehi _15406__1843 (.L_HI(net1843));
 sg13g2_tiehi _15988__1844 (.L_HI(net1844));
 sg13g2_tiehi _15405__1845 (.L_HI(net1845));
 sg13g2_tiehi _15863__1846 (.L_HI(net1846));
 sg13g2_tiehi _15404__1847 (.L_HI(net1847));
 sg13g2_tiehi _15932__1848 (.L_HI(net1848));
 sg13g2_tiehi _15403__1849 (.L_HI(net1849));
 sg13g2_tiehi _15862__1850 (.L_HI(net1850));
 sg13g2_tiehi _15402__1851 (.L_HI(net1851));
 sg13g2_tiehi _15861__1852 (.L_HI(net1852));
 sg13g2_tiehi _15401__1853 (.L_HI(net1853));
 sg13g2_tiehi _15860__1854 (.L_HI(net1854));
 sg13g2_tiehi _15400__1855 (.L_HI(net1855));
 sg13g2_tiehi _15859__1856 (.L_HI(net1856));
 sg13g2_tiehi _15399__1857 (.L_HI(net1857));
 sg13g2_tiehi _15858__1858 (.L_HI(net1858));
 sg13g2_tiehi _15398__1859 (.L_HI(net1859));
 sg13g2_tiehi _15857__1860 (.L_HI(net1860));
 sg13g2_tiehi _15397__1861 (.L_HI(net1861));
 sg13g2_tiehi _15856__1862 (.L_HI(net1862));
 sg13g2_tiehi _15396__1863 (.L_HI(net1863));
 sg13g2_tiehi _15855__1864 (.L_HI(net1864));
 sg13g2_tiehi _15395__1865 (.L_HI(net1865));
 sg13g2_tiehi _15854__1866 (.L_HI(net1866));
 sg13g2_tiehi _15394__1867 (.L_HI(net1867));
 sg13g2_tiehi _15853__1868 (.L_HI(net1868));
 sg13g2_tiehi _15393__1869 (.L_HI(net1869));
 sg13g2_tiehi _15852__1870 (.L_HI(net1870));
 sg13g2_tiehi _15392__1871 (.L_HI(net1871));
 sg13g2_tiehi _15851__1872 (.L_HI(net1872));
 sg13g2_tiehi _15391__1873 (.L_HI(net1873));
 sg13g2_tiehi _15850__1874 (.L_HI(net1874));
 sg13g2_tiehi _15390__1875 (.L_HI(net1875));
 sg13g2_tiehi _15849__1876 (.L_HI(net1876));
 sg13g2_tiehi _15389__1877 (.L_HI(net1877));
 sg13g2_tiehi _15848__1878 (.L_HI(net1878));
 sg13g2_tiehi _15388__1879 (.L_HI(net1879));
 sg13g2_tiehi _15847__1880 (.L_HI(net1880));
 sg13g2_tiehi _15387__1881 (.L_HI(net1881));
 sg13g2_tiehi _15846__1882 (.L_HI(net1882));
 sg13g2_tiehi _15386__1883 (.L_HI(net1883));
 sg13g2_tiehi _15987__1884 (.L_HI(net1884));
 sg13g2_tiehi _15385__1885 (.L_HI(net1885));
 sg13g2_tiehi _15845__1886 (.L_HI(net1886));
 sg13g2_tiehi _15384__1887 (.L_HI(net1887));
 sg13g2_tiehi _15931__1888 (.L_HI(net1888));
 sg13g2_tiehi _15383__1889 (.L_HI(net1889));
 sg13g2_tiehi _15844__1890 (.L_HI(net1890));
 sg13g2_tiehi _15382__1891 (.L_HI(net1891));
 sg13g2_tiehi _15843__1892 (.L_HI(net1892));
 sg13g2_tiehi _15381__1893 (.L_HI(net1893));
 sg13g2_tiehi _15842__1894 (.L_HI(net1894));
 sg13g2_tiehi _15380__1895 (.L_HI(net1895));
 sg13g2_tiehi _15841__1896 (.L_HI(net1896));
 sg13g2_tiehi _15379__1897 (.L_HI(net1897));
 sg13g2_tiehi _15840__1898 (.L_HI(net1898));
 sg13g2_tiehi _15378__1899 (.L_HI(net1899));
 sg13g2_tiehi _15839__1900 (.L_HI(net1900));
 sg13g2_tiehi _15377__1901 (.L_HI(net1901));
 sg13g2_tiehi _15838__1902 (.L_HI(net1902));
 sg13g2_tiehi _15376__1903 (.L_HI(net1903));
 sg13g2_tiehi _15837__1904 (.L_HI(net1904));
 sg13g2_tiehi _15375__1905 (.L_HI(net1905));
 sg13g2_tiehi _15836__1906 (.L_HI(net1906));
 sg13g2_tiehi _15374__1907 (.L_HI(net1907));
 sg13g2_tiehi _15835__1908 (.L_HI(net1908));
 sg13g2_tiehi _15373__1909 (.L_HI(net1909));
 sg13g2_tiehi _15834__1910 (.L_HI(net1910));
 sg13g2_tiehi _15372__1911 (.L_HI(net1911));
 sg13g2_tiehi _15833__1912 (.L_HI(net1912));
 sg13g2_tiehi _15371__1913 (.L_HI(net1913));
 sg13g2_tiehi _15832__1914 (.L_HI(net1914));
 sg13g2_tiehi _15370__1915 (.L_HI(net1915));
 sg13g2_tiehi _15831__1916 (.L_HI(net1916));
 sg13g2_tiehi _15369__1917 (.L_HI(net1917));
 sg13g2_tiehi _15830__1918 (.L_HI(net1918));
 sg13g2_tiehi _15368__1919 (.L_HI(net1919));
 sg13g2_tiehi _15829__1920 (.L_HI(net1920));
 sg13g2_tiehi _15367__1921 (.L_HI(net1921));
 sg13g2_tiehi _15828__1922 (.L_HI(net1922));
 sg13g2_tiehi _15366__1923 (.L_HI(net1923));
 sg13g2_tiehi _15827__1924 (.L_HI(net1924));
 sg13g2_tiehi _15365__1925 (.L_HI(net1925));
 sg13g2_tiehi _15826__1926 (.L_HI(net1926));
 sg13g2_tiehi _15364__1927 (.L_HI(net1927));
 sg13g2_tiehi _15825__1928 (.L_HI(net1928));
 sg13g2_tiehi _15363__1929 (.L_HI(net1929));
 sg13g2_tiehi _15824__1930 (.L_HI(net1930));
 sg13g2_tiehi _15362__1931 (.L_HI(net1931));
 sg13g2_tiehi _15986__1932 (.L_HI(net1932));
 sg13g2_tiehi _15361__1933 (.L_HI(net1933));
 sg13g2_tiehi _15823__1934 (.L_HI(net1934));
 sg13g2_tiehi _15360__1935 (.L_HI(net1935));
 sg13g2_tiehi _15930__1936 (.L_HI(net1936));
 sg13g2_tiehi _15359__1937 (.L_HI(net1937));
 sg13g2_tiehi _15822__1938 (.L_HI(net1938));
 sg13g2_tiehi _15358__1939 (.L_HI(net1939));
 sg13g2_tiehi _15985__1940 (.L_HI(net1940));
 sg13g2_tiehi _15357__1941 (.L_HI(net1941));
 sg13g2_tiehi _15821__1942 (.L_HI(net1942));
 sg13g2_tiehi _15356__1943 (.L_HI(net1943));
 sg13g2_tiehi _15820__1944 (.L_HI(net1944));
 sg13g2_tiehi _15355__1945 (.L_HI(net1945));
 sg13g2_tiehi _15819__1946 (.L_HI(net1946));
 sg13g2_tiehi _15354__1947 (.L_HI(net1947));
 sg13g2_tiehi _15929__1948 (.L_HI(net1948));
 sg13g2_tiehi _15353__1949 (.L_HI(net1949));
 sg13g2_tiehi _15818__1950 (.L_HI(net1950));
 sg13g2_tiehi _15352__1951 (.L_HI(net1951));
 sg13g2_tiehi _15928__1952 (.L_HI(net1952));
 sg13g2_tiehi _15351__1953 (.L_HI(net1953));
 sg13g2_tiehi _15817__1954 (.L_HI(net1954));
 sg13g2_tiehi _15350__1955 (.L_HI(net1955));
 sg13g2_tiehi _15984__1956 (.L_HI(net1956));
 sg13g2_tiehi _15349__1957 (.L_HI(net1957));
 sg13g2_tiehi _15816__1958 (.L_HI(net1958));
 sg13g2_tiehi _15348__1959 (.L_HI(net1959));
 sg13g2_tiehi _15927__1960 (.L_HI(net1960));
 sg13g2_tiehi _15347__1961 (.L_HI(net1961));
 sg13g2_tiehi _15815__1962 (.L_HI(net1962));
 sg13g2_tiehi _15346__1963 (.L_HI(net1963));
 sg13g2_tiehi _15814__1964 (.L_HI(net1964));
 sg13g2_tiehi _15345__1965 (.L_HI(net1965));
 sg13g2_tiehi _15813__1966 (.L_HI(net1966));
 sg13g2_tiehi _15344__1967 (.L_HI(net1967));
 sg13g2_tiehi _15812__1968 (.L_HI(net1968));
 sg13g2_tiehi _15343__1969 (.L_HI(net1969));
 sg13g2_tiehi _15811__1970 (.L_HI(net1970));
 sg13g2_tiehi _15342__1971 (.L_HI(net1971));
 sg13g2_tiehi _15810__1972 (.L_HI(net1972));
 sg13g2_tiehi _15341__1973 (.L_HI(net1973));
 sg13g2_tiehi _15809__1974 (.L_HI(net1974));
 sg13g2_tiehi _15340__1975 (.L_HI(net1975));
 sg13g2_tiehi _15808__1976 (.L_HI(net1976));
 sg13g2_tiehi _15339__1977 (.L_HI(net1977));
 sg13g2_tiehi _15807__1978 (.L_HI(net1978));
 sg13g2_tiehi _15338__1979 (.L_HI(net1979));
 sg13g2_tiehi _15806__1980 (.L_HI(net1980));
 sg13g2_tiehi _15337__1981 (.L_HI(net1981));
 sg13g2_tiehi _15805__1982 (.L_HI(net1982));
 sg13g2_tiehi _15336__1983 (.L_HI(net1983));
 sg13g2_tiehi _15804__1984 (.L_HI(net1984));
 sg13g2_tiehi _15335__1985 (.L_HI(net1985));
 sg13g2_tiehi _15803__1986 (.L_HI(net1986));
 sg13g2_tiehi _15334__1987 (.L_HI(net1987));
 sg13g2_tiehi _15802__1988 (.L_HI(net1988));
 sg13g2_tiehi _15333__1989 (.L_HI(net1989));
 sg13g2_tiehi _15801__1990 (.L_HI(net1990));
 sg13g2_tiehi _15332__1991 (.L_HI(net1991));
 sg13g2_tiehi _15800__1992 (.L_HI(net1992));
 sg13g2_tiehi _15331__1993 (.L_HI(net1993));
 sg13g2_tiehi _15799__1994 (.L_HI(net1994));
 sg13g2_tiehi _15330__1995 (.L_HI(net1995));
 sg13g2_tiehi _15798__1996 (.L_HI(net1996));
 sg13g2_tiehi _15329__1997 (.L_HI(net1997));
 sg13g2_tiehi _15926__1998 (.L_HI(net1998));
 sg13g2_tiehi _15328__1999 (.L_HI(net1999));
 sg13g2_tiehi _15797__2000 (.L_HI(net2000));
 sg13g2_tiehi _15327__2001 (.L_HI(net2001));
 sg13g2_tiehi _15925__2002 (.L_HI(net2002));
 sg13g2_tiehi _15326__2003 (.L_HI(net2003));
 sg13g2_tiehi _15796__2004 (.L_HI(net2004));
 sg13g2_tiehi _15325__2005 (.L_HI(net2005));
 sg13g2_tiehi _15924__2006 (.L_HI(net2006));
 sg13g2_tiehi _15324__2007 (.L_HI(net2007));
 sg13g2_tiehi _15795__2008 (.L_HI(net2008));
 sg13g2_tiehi _15323__2009 (.L_HI(net2009));
 sg13g2_tiehi _15983__2010 (.L_HI(net2010));
 sg13g2_tiehi _15322__2011 (.L_HI(net2011));
 sg13g2_tiehi _15794__2012 (.L_HI(net2012));
 sg13g2_tiehi _15321__2013 (.L_HI(net2013));
 sg13g2_tiehi _15923__2014 (.L_HI(net2014));
 sg13g2_tiehi _15320__2015 (.L_HI(net2015));
 sg13g2_tiehi _15793__2016 (.L_HI(net2016));
 sg13g2_tiehi _15319__2017 (.L_HI(net2017));
 sg13g2_tiehi _15982__2018 (.L_HI(net2018));
 sg13g2_tiehi _15318__2019 (.L_HI(net2019));
 sg13g2_tiehi _15736__2020 (.L_HI(net2020));
 sg13g2_tiehi _15792__2021 (.L_HI(net2021));
 sg13g2_tiehi _15317__2022 (.L_HI(net2022));
 sg13g2_tiehi _15922__2023 (.L_HI(net2023));
 sg13g2_tiehi _15316__2024 (.L_HI(net2024));
 sg13g2_tiehi _15791__2025 (.L_HI(net2025));
 sg13g2_tiehi _15315__2026 (.L_HI(net2026));
 sg13g2_tiehi _15981__2027 (.L_HI(net2027));
 sg13g2_tiehi _15314__2028 (.L_HI(net2028));
 sg13g2_tiehi _15790__2029 (.L_HI(net2029));
 sg13g2_tiehi _15313__2030 (.L_HI(net2030));
 sg13g2_tiehi _15921__2031 (.L_HI(net2031));
 sg13g2_tiehi _15312__2032 (.L_HI(net2032));
 sg13g2_tiehi _15789__2033 (.L_HI(net2033));
 sg13g2_tiehi _15311__2034 (.L_HI(net2034));
 sg13g2_tiehi _15788__2035 (.L_HI(net2035));
 sg13g2_tiehi _15310__2036 (.L_HI(net2036));
 sg13g2_tiehi _15980__2037 (.L_HI(net2037));
 sg13g2_tiehi _15309__2038 (.L_HI(net2038));
 sg13g2_tiehi _15787__2039 (.L_HI(net2039));
 sg13g2_tiehi _15308__2040 (.L_HI(net2040));
 sg13g2_tiehi _15919__2041 (.L_HI(net2041));
 sg13g2_tiehi _15307__2042 (.L_HI(net2042));
 sg13g2_tiehi _15786__2043 (.L_HI(net2043));
 sg13g2_tiehi _15306__2044 (.L_HI(net2044));
 sg13g2_tiehi _15979__2045 (.L_HI(net2045));
 sg13g2_tiehi _15305__2046 (.L_HI(net2046));
 sg13g2_tiehi _15785__2047 (.L_HI(net2047));
 sg13g2_tiehi _15304__2048 (.L_HI(net2048));
 sg13g2_tiehi _15918__2049 (.L_HI(net2049));
 sg13g2_tiehi _15303__2050 (.L_HI(net2050));
 sg13g2_tiehi _15784__2051 (.L_HI(net2051));
 sg13g2_tiehi _15302__2052 (.L_HI(net2052));
 sg13g2_tiehi _15978__2053 (.L_HI(net2053));
 sg13g2_tiehi _15301__2054 (.L_HI(net2054));
 sg13g2_tiehi _15783__2055 (.L_HI(net2055));
 sg13g2_tiehi _15300__2056 (.L_HI(net2056));
 sg13g2_tiehi _15782__2057 (.L_HI(net2057));
 sg13g2_tiehi _15299__2058 (.L_HI(net2058));
 sg13g2_tiehi _15781__2059 (.L_HI(net2059));
 sg13g2_tiehi _15298__2060 (.L_HI(net2060));
 sg13g2_tiehi _15780__2061 (.L_HI(net2061));
 sg13g2_tiehi _15297__2062 (.L_HI(net2062));
 sg13g2_tiehi _15779__2063 (.L_HI(net2063));
 sg13g2_tiehi _15296__2064 (.L_HI(net2064));
 sg13g2_tiehi _15778__2065 (.L_HI(net2065));
 sg13g2_tiehi _15295__2066 (.L_HI(net2066));
 sg13g2_tiehi _15917__2067 (.L_HI(net2067));
 sg13g2_tiehi _15294__2068 (.L_HI(net2068));
 sg13g2_tiehi _15777__2069 (.L_HI(net2069));
 sg13g2_tiehi _15293__2070 (.L_HI(net2070));
 sg13g2_tiehi _15776__2071 (.L_HI(net2071));
 sg13g2_tiehi _15292__2072 (.L_HI(net2072));
 sg13g2_tiehi _15775__2073 (.L_HI(net2073));
 sg13g2_tiehi _15291__2074 (.L_HI(net2074));
 sg13g2_tiehi _15774__2075 (.L_HI(net2075));
 sg13g2_tiehi _15290__2076 (.L_HI(net2076));
 sg13g2_tiehi _15773__2077 (.L_HI(net2077));
 sg13g2_tiehi _15289__2078 (.L_HI(net2078));
 sg13g2_tiehi _15772__2079 (.L_HI(net2079));
 sg13g2_tiehi _15288__2080 (.L_HI(net2080));
 sg13g2_tiehi _15771__2081 (.L_HI(net2081));
 sg13g2_tiehi _15287__2082 (.L_HI(net2082));
 sg13g2_tiehi _15770__2083 (.L_HI(net2083));
 sg13g2_tiehi _15286__2084 (.L_HI(net2084));
 sg13g2_tiehi _15769__2085 (.L_HI(net2085));
 sg13g2_tiehi _15285__2086 (.L_HI(net2086));
 sg13g2_tiehi _15768__2087 (.L_HI(net2087));
 sg13g2_tiehi _15284__2088 (.L_HI(net2088));
 sg13g2_tiehi _15767__2089 (.L_HI(net2089));
 sg13g2_tiehi _15283__2090 (.L_HI(net2090));
 sg13g2_tiehi _15766__2091 (.L_HI(net2091));
 sg13g2_tiehi _15282__2092 (.L_HI(net2092));
 sg13g2_tiehi _15765__2093 (.L_HI(net2093));
 sg13g2_tiehi _15281__2094 (.L_HI(net2094));
 sg13g2_tiehi _15764__2095 (.L_HI(net2095));
 sg13g2_tiehi _14554__2096 (.L_HI(net2096));
 sg13g2_tiehi _14527__2097 (.L_HI(net2097));
 sg13g2_tiehi _14528__2098 (.L_HI(net2098));
 sg13g2_tiehi _14529__2099 (.L_HI(net2099));
 sg13g2_tiehi _14530__2100 (.L_HI(net2100));
 sg13g2_tiehi _14531__2101 (.L_HI(net2101));
 sg13g2_tiehi _14532__2102 (.L_HI(net2102));
 sg13g2_tiehi _14533__2103 (.L_HI(net2103));
 sg13g2_tiehi _14534__2104 (.L_HI(net2104));
 sg13g2_tiehi _14535__2105 (.L_HI(net2105));
 sg13g2_tiehi _14536__2106 (.L_HI(net2106));
 sg13g2_tiehi _14537__2107 (.L_HI(net2107));
 sg13g2_inv_1 _08955__1 (.Y(net2108),
    .A(clknet_leaf_17_clk));
 sg13g2_buf_4 fanout656 (.X(net656),
    .A(net658));
 sg13g2_buf_2 _17442_ (.A(net1),
    .X(uio_oe[0]));
 sg13g2_buf_2 _17443_ (.A(uio_oe[5]),
    .X(uio_oe[1]));
 sg13g2_buf_2 _17444_ (.A(uio_oe[5]),
    .X(uio_oe[2]));
 sg13g2_buf_2 _17445_ (.A(net1),
    .X(uio_oe[3]));
 sg13g2_buf_2 _17446_ (.A(uio_oe[5]),
    .X(uio_oe[4]));
 sg13g2_buf_2 _17447_ (.A(net1),
    .X(uio_oe[6]));
 sg13g2_buf_2 _17448_ (.A(net1),
    .X(uio_oe[7]));
 sg13g2_buf_2 fanout655 (.A(net3907),
    .X(net655));
 sg13g2_buf_1 fanout654 (.A(net655),
    .X(net654));
 sg13g2_buf_2 fanout653 (.A(net654),
    .X(net653));
 sg13g2_buf_2 fanout652 (.A(net3907),
    .X(net652));
 sg13g2_buf_8 game_clk_buf (.A(net7),
    .X(game_clk));
 sg13g2_buf_2 fanout651 (.A(net652),
    .X(net651));
 sg13g2_buf_2 fanout650 (.A(net651),
    .X(net650));
 sg13g2_buf_2 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(net3917));
 sg13g2_buf_4 fanout647 (.X(net647),
    .A(net648));
 sg13g2_buf_1 fanout646 (.A(\i_spi.busy ),
    .X(net646));
 sg13g2_buf_1 fanout645 (.A(net646),
    .X(net645));
 sg13g2_buf_1 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_1 fanout643 (.A(net644),
    .X(net643));
 sg13g2_buf_2 fanout642 (.A(net644),
    .X(net642));
 sg13g2_buf_2 fanout641 (.A(net646),
    .X(net641));
 sg13g2_buf_4 fanout640 (.X(net640),
    .A(\i_latch_mem.cycle[1] ));
 sg13g2_buf_4 fanout639 (.X(net639),
    .A(\i_latch_mem.cycle[0] ));
 sg13g2_buf_4 fanout638 (.X(net638),
    .A(\addr[26] ));
 sg13g2_buf_4 fanout637 (.X(net637),
    .A(net638));
 sg13g2_buf_2 fanout636 (.A(net638),
    .X(net636));
 sg13g2_buf_1 fanout635 (.A(net636),
    .X(net635));
 sg13g2_buf_2 fanout634 (.A(net635),
    .X(net634));
 sg13g2_buf_4 fanout633 (.X(net633),
    .A(\addr[2] ));
 sg13g2_buf_4 fanout632 (.X(net632),
    .A(net633));
 sg13g2_buf_2 fanout631 (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .X(net631));
 sg13g2_buf_2 fanout630 (.A(net631),
    .X(net630));
 sg13g2_buf_2 fanout629 (.A(net630),
    .X(net629));
 sg13g2_buf_2 fanout628 (.A(net629),
    .X(net628));
 sg13g2_buf_2 fanout627 (.A(net4125),
    .X(net627));
 sg13g2_buf_2 fanout626 (.A(net627),
    .X(net626));
 sg13g2_buf_2 fanout625 (.A(net626),
    .X(net625));
 sg13g2_buf_2 fanout624 (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .X(net624));
 sg13g2_buf_2 fanout623 (.A(net624),
    .X(net623));
 sg13g2_buf_2 fanout622 (.A(net623),
    .X(net622));
 sg13g2_buf_2 fanout621 (.A(net624),
    .X(net621));
 sg13g2_buf_2 fanout620 (.A(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .X(net620));
 sg13g2_buf_4 fanout619 (.X(net619),
    .A(net4118));
 sg13g2_buf_1 fanout618 (.A(net3933),
    .X(net618));
 sg13g2_buf_2 fanout617 (.A(net3933),
    .X(net617));
 sg13g2_buf_4 fanout616 (.X(net616),
    .A(\i_tinyqv.mem.q_ctrl.fsm_state[0] ));
 sg13g2_buf_2 fanout615 (.A(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .X(net615));
 sg13g2_buf_4 fanout614 (.X(net614),
    .A(\i_tinyqv.cpu.instr_data_start[13] ));
 sg13g2_buf_2 fanout613 (.A(\i_tinyqv.cpu.instr_data_start[14] ),
    .X(net613));
 sg13g2_buf_2 fanout612 (.A(\i_tinyqv.cpu.instr_data_start[16] ),
    .X(net612));
 sg13g2_buf_2 fanout611 (.A(\i_tinyqv.cpu.instr_data_start[17] ),
    .X(net611));
 sg13g2_buf_4 fanout610 (.X(net610),
    .A(net4123));
 sg13g2_buf_2 fanout609 (.A(\i_tinyqv.cpu.instr_data_start[21] ),
    .X(net609));
 sg13g2_buf_2 fanout608 (.A(\i_tinyqv.cpu.was_early_branch ),
    .X(net608));
 sg13g2_buf_1 fanout607 (.A(net608),
    .X(net607));
 sg13g2_buf_1 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_2 fanout605 (.A(net606),
    .X(net605));
 sg13g2_buf_4 fanout604 (.X(net604),
    .A(net4098));
 sg13g2_buf_1 fanout603 (.A(net604),
    .X(net603));
 sg13g2_buf_2 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_4 fanout601 (.X(net601),
    .A(net4124));
 sg13g2_buf_4 fanout600 (.X(net600),
    .A(net4126));
 sg13g2_buf_4 fanout599 (.X(net599),
    .A(\data_to_write[4] ));
 sg13g2_buf_8 fanout598 (.A(\data_to_write[5] ),
    .X(net598));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(\data_to_write[6] ));
 sg13g2_buf_4 fanout596 (.X(net596),
    .A(\i_tinyqv.cpu.counter[2] ));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(net596));
 sg13g2_buf_1 fanout594 (.A(net595),
    .X(net594));
 sg13g2_buf_2 fanout593 (.A(net594),
    .X(net593));
 sg13g2_buf_4 fanout592 (.X(net592),
    .A(\i_tinyqv.cpu.counter[2] ));
 sg13g2_buf_4 fanout591 (.X(net591),
    .A(\i_tinyqv.cpu.counter[2] ));
 sg13g2_buf_2 fanout590 (.A(net592),
    .X(net590));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(\i_tinyqv.cpu.counter[3] ));
 sg13g2_buf_4 fanout588 (.X(net588),
    .A(net589));
 sg13g2_buf_2 fanout587 (.A(\i_tinyqv.cpu.counter[4] ),
    .X(net587));
 sg13g2_buf_2 fanout586 (.A(net587),
    .X(net586));
 sg13g2_buf_2 fanout585 (.A(net587),
    .X(net585));
 sg13g2_buf_2 fanout584 (.A(net587),
    .X(net584));
 sg13g2_buf_4 fanout583 (.X(net583),
    .A(net587));
 sg13g2_buf_4 fanout582 (.X(net582),
    .A(\i_tinyqv.cpu.i_core.imm_lo[2] ));
 sg13g2_buf_4 fanout581 (.X(net581),
    .A(\i_tinyqv.cpu.alu_op[0] ));
 sg13g2_buf_2 fanout580 (.A(\i_tinyqv.cpu.alu_op[2] ),
    .X(net580));
 sg13g2_buf_2 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_2 fanout578 (.A(net579),
    .X(net578));
 sg13g2_buf_8 fanout577 (.A(net579),
    .X(net577));
 sg13g2_buf_4 fanout576 (.X(net576),
    .A(net580));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(net580));
 sg13g2_buf_2 fanout574 (.A(net4127),
    .X(net574));
 sg13g2_buf_2 fanout573 (.A(net574),
    .X(net573));
 sg13g2_buf_2 fanout572 (.A(net574),
    .X(net572));
 sg13g2_buf_2 fanout571 (.A(net4101),
    .X(net571));
 sg13g2_buf_2 fanout570 (.A(net571),
    .X(net570));
 sg13g2_buf_2 fanout569 (.A(net570),
    .X(net569));
 sg13g2_buf_4 fanout568 (.X(net568),
    .A(net571));
 sg13g2_buf_2 fanout567 (.A(_02128_),
    .X(net567));
 sg13g2_buf_2 fanout566 (.A(net567),
    .X(net566));
 sg13g2_buf_2 fanout565 (.A(_02129_),
    .X(net565));
 sg13g2_buf_2 fanout564 (.A(_02132_),
    .X(net564));
 sg13g2_buf_2 fanout563 (.A(_02132_),
    .X(net563));
 sg13g2_buf_2 fanout562 (.A(_02135_),
    .X(net562));
 sg13g2_buf_2 fanout561 (.A(_02135_),
    .X(net561));
 sg13g2_buf_2 fanout560 (.A(_02137_),
    .X(net560));
 sg13g2_buf_2 fanout559 (.A(_02140_),
    .X(net559));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_2 fanout557 (.A(_02185_),
    .X(net557));
 sg13g2_buf_2 fanout556 (.A(net557),
    .X(net556));
 sg13g2_buf_1 fanout555 (.A(_02186_),
    .X(net555));
 sg13g2_buf_2 fanout554 (.A(_02186_),
    .X(net554));
 sg13g2_buf_1 fanout553 (.A(_02189_),
    .X(net553));
 sg13g2_buf_2 fanout552 (.A(_02189_),
    .X(net552));
 sg13g2_buf_2 fanout551 (.A(_02192_),
    .X(net551));
 sg13g2_buf_1 fanout550 (.A(_02193_),
    .X(net550));
 sg13g2_buf_2 fanout549 (.A(_02193_),
    .X(net549));
 sg13g2_buf_2 fanout548 (.A(_02196_),
    .X(net548));
 sg13g2_buf_2 fanout547 (.A(_04925_),
    .X(net547));
 sg13g2_buf_1 fanout546 (.A(\i_game.data_latch_wen ),
    .X(net546));
 sg13g2_buf_2 fanout545 (.A(net546),
    .X(net545));
 sg13g2_buf_2 fanout544 (.A(net546),
    .X(net544));
 sg13g2_buf_1 fanout543 (.A(net546),
    .X(net543));
 sg13g2_buf_2 fanout542 (.A(net546),
    .X(net542));
 sg13g2_buf_2 fanout541 (.A(\i_game.data_latch_wen ),
    .X(net541));
 sg13g2_buf_2 fanout540 (.A(net541),
    .X(net540));
 sg13g2_buf_2 fanout539 (.A(net541),
    .X(net539));
 sg13g2_buf_1 fanout538 (.A(\i_debug_uart_tx.resetn ),
    .X(net538));
 sg13g2_buf_4 fanout537 (.X(net537),
    .A(net538));
 sg13g2_buf_2 fanout536 (.A(net538),
    .X(net536));
 sg13g2_buf_2 fanout535 (.A(net538),
    .X(net535));
 sg13g2_buf_2 fanout534 (.A(\i_debug_uart_tx.resetn ),
    .X(net534));
 sg13g2_buf_1 fanout533 (.A(net534),
    .X(net533));
 sg13g2_buf_2 fanout532 (.A(net534),
    .X(net532));
 sg13g2_buf_4 fanout531 (.X(net531),
    .A(\i_debug_uart_tx.resetn ));
 sg13g2_buf_2 fanout530 (.A(net531),
    .X(net530));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(net530));
 sg13g2_buf_2 fanout528 (.A(net529),
    .X(net528));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527));
 sg13g2_buf_2 fanout526 (.A(net530),
    .X(net526));
 sg13g2_buf_2 fanout525 (.A(net526),
    .X(net525));
 sg13g2_buf_2 fanout524 (.A(net530),
    .X(net524));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(net524));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(net531));
 sg13g2_buf_2 fanout521 (.A(net522),
    .X(net521));
 sg13g2_buf_4 fanout520 (.X(net520),
    .A(net531));
 sg13g2_buf_4 fanout519 (.X(net519),
    .A(net520));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(net520));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(_00195_));
 sg13g2_buf_4 fanout516 (.X(net516),
    .A(net4131));
 sg13g2_buf_2 fanout515 (.A(_01522_),
    .X(net515));
 sg13g2_buf_2 fanout514 (.A(_01577_),
    .X(net514));
 sg13g2_buf_2 fanout513 (.A(net514),
    .X(net513));
 sg13g2_buf_4 fanout512 (.X(net512),
    .A(net513));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(net512));
 sg13g2_buf_4 fanout510 (.X(net510),
    .A(net513));
 sg13g2_buf_2 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_4 fanout508 (.X(net508),
    .A(net514));
 sg13g2_buf_1 fanout507 (.A(net508),
    .X(net507));
 sg13g2_buf_2 fanout506 (.A(net508),
    .X(net506));
 sg13g2_buf_1 fanout505 (.A(_01667_),
    .X(net505));
 sg13g2_buf_2 fanout504 (.A(net505),
    .X(net504));
 sg13g2_buf_2 fanout503 (.A(net504),
    .X(net503));
 sg13g2_buf_2 fanout502 (.A(net503),
    .X(net502));
 sg13g2_buf_2 fanout501 (.A(net505),
    .X(net501));
 sg13g2_buf_2 fanout500 (.A(_01727_),
    .X(net500));
 sg13g2_buf_2 fanout499 (.A(net500),
    .X(net499));
 sg13g2_buf_1 fanout498 (.A(net499),
    .X(net498));
 sg13g2_buf_2 fanout497 (.A(net499),
    .X(net497));
 sg13g2_buf_4 fanout496 (.X(net496),
    .A(_01729_));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(_01731_));
 sg13g2_buf_2 fanout494 (.A(net495),
    .X(net494));
 sg13g2_buf_1 fanout493 (.A(net495),
    .X(net493));
 sg13g2_buf_2 fanout492 (.A(net493),
    .X(net492));
 sg13g2_buf_2 fanout491 (.A(net492),
    .X(net491));
 sg13g2_buf_4 fanout490 (.X(net490),
    .A(_01733_));
 sg13g2_buf_2 fanout489 (.A(net490),
    .X(net489));
 sg13g2_buf_1 fanout488 (.A(net489),
    .X(net488));
 sg13g2_buf_2 fanout487 (.A(net489),
    .X(net487));
 sg13g2_buf_4 fanout486 (.X(net486),
    .A(_03624_));
 sg13g2_buf_2 fanout485 (.A(_04892_),
    .X(net485));
 sg13g2_buf_2 fanout484 (.A(net485),
    .X(net484));
 sg13g2_buf_2 fanout483 (.A(_04901_),
    .X(net483));
 sg13g2_buf_1 fanout482 (.A(_05027_),
    .X(net482));
 sg13g2_buf_2 fanout481 (.A(_05027_),
    .X(net481));
 sg13g2_buf_2 fanout480 (.A(_05028_),
    .X(net480));
 sg13g2_buf_2 fanout479 (.A(net480),
    .X(net479));
 sg13g2_buf_2 fanout478 (.A(_01512_),
    .X(net478));
 sg13g2_buf_2 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_2 fanout476 (.A(_01580_),
    .X(net476));
 sg13g2_buf_2 fanout475 (.A(net476),
    .X(net475));
 sg13g2_buf_4 fanout474 (.X(net474),
    .A(net475));
 sg13g2_buf_8 fanout473 (.A(_01582_),
    .X(net473));
 sg13g2_buf_4 fanout472 (.X(net472),
    .A(net473));
 sg13g2_buf_4 fanout471 (.X(net471),
    .A(_02163_));
 sg13g2_buf_2 fanout470 (.A(net471),
    .X(net470));
 sg13g2_buf_1 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_2 fanout468 (.A(net470),
    .X(net468));
 sg13g2_buf_4 fanout467 (.X(net467),
    .A(_02165_));
 sg13g2_buf_2 fanout466 (.A(net467),
    .X(net466));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(net466));
 sg13g2_buf_4 fanout464 (.X(net464),
    .A(_02166_));
 sg13g2_buf_4 fanout463 (.X(net463),
    .A(_02168_));
 sg13g2_buf_4 fanout462 (.X(net462),
    .A(net463));
 sg13g2_buf_4 fanout461 (.X(net461),
    .A(net462));
 sg13g2_buf_2 fanout460 (.A(_02170_),
    .X(net460));
 sg13g2_buf_2 fanout459 (.A(net460),
    .X(net459));
 sg13g2_buf_2 fanout458 (.A(net459),
    .X(net458));
 sg13g2_buf_4 fanout457 (.X(net457),
    .A(net459));
 sg13g2_buf_4 fanout456 (.X(net456),
    .A(_02231_));
 sg13g2_buf_2 fanout455 (.A(_02232_),
    .X(net455));
 sg13g2_buf_2 fanout454 (.A(net455),
    .X(net454));
 sg13g2_buf_2 fanout453 (.A(net454),
    .X(net453));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(net453));
 sg13g2_buf_2 fanout451 (.A(_03477_),
    .X(net451));
 sg13g2_buf_2 fanout450 (.A(_03477_),
    .X(net450));
 sg13g2_buf_4 fanout449 (.X(net449),
    .A(_03478_));
 sg13g2_buf_1 fanout448 (.A(net449),
    .X(net448));
 sg13g2_buf_2 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_2 fanout446 (.A(net447),
    .X(net446));
 sg13g2_buf_2 fanout445 (.A(net449),
    .X(net445));
 sg13g2_buf_2 fanout444 (.A(net445),
    .X(net444));
 sg13g2_buf_1 fanout443 (.A(net449),
    .X(net443));
 sg13g2_buf_1 fanout442 (.A(net443),
    .X(net442));
 sg13g2_buf_2 fanout441 (.A(net443),
    .X(net441));
 sg13g2_buf_1 fanout440 (.A(net443),
    .X(net440));
 sg13g2_buf_2 fanout439 (.A(net443),
    .X(net439));
 sg13g2_buf_4 fanout438 (.X(net438),
    .A(_03480_));
 sg13g2_buf_1 fanout437 (.A(_03481_),
    .X(net437));
 sg13g2_buf_4 fanout436 (.X(net436),
    .A(net437));
 sg13g2_buf_1 fanout435 (.A(net437),
    .X(net435));
 sg13g2_buf_2 fanout434 (.A(net435),
    .X(net434));
 sg13g2_buf_2 fanout433 (.A(_03602_),
    .X(net433));
 sg13g2_buf_2 fanout432 (.A(_04866_),
    .X(net432));
 sg13g2_buf_2 fanout431 (.A(net432),
    .X(net431));
 sg13g2_buf_2 fanout430 (.A(_04874_),
    .X(net430));
 sg13g2_buf_2 fanout429 (.A(_04874_),
    .X(net429));
 sg13g2_buf_2 fanout428 (.A(_04986_),
    .X(net428));
 sg13g2_buf_2 fanout427 (.A(_01525_),
    .X(net427));
 sg13g2_buf_2 fanout426 (.A(_01710_),
    .X(net426));
 sg13g2_buf_4 fanout425 (.X(net425),
    .A(net426));
 sg13g2_buf_4 fanout424 (.X(net424),
    .A(_01710_));
 sg13g2_buf_2 fanout423 (.A(net424),
    .X(net423));
 sg13g2_buf_2 fanout422 (.A(_01710_),
    .X(net422));
 sg13g2_buf_4 fanout421 (.X(net421),
    .A(_02074_));
 sg13g2_buf_4 fanout420 (.X(net420),
    .A(net421));
 sg13g2_buf_2 fanout419 (.A(net420),
    .X(net419));
 sg13g2_buf_2 fanout418 (.A(net420),
    .X(net418));
 sg13g2_buf_2 fanout417 (.A(_02075_),
    .X(net417));
 sg13g2_buf_1 fanout416 (.A(net417),
    .X(net416));
 sg13g2_buf_2 fanout415 (.A(net417),
    .X(net415));
 sg13g2_buf_4 fanout414 (.X(net414),
    .A(_02182_));
 sg13g2_buf_2 fanout413 (.A(net414),
    .X(net413));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(net413));
 sg13g2_buf_2 fanout411 (.A(net413),
    .X(net411));
 sg13g2_buf_2 fanout410 (.A(_02183_),
    .X(net410));
 sg13g2_buf_1 fanout409 (.A(net410),
    .X(net409));
 sg13g2_buf_2 fanout408 (.A(net410),
    .X(net408));
 sg13g2_buf_4 fanout407 (.X(net407),
    .A(_02482_));
 sg13g2_buf_2 fanout406 (.A(_02831_),
    .X(net406));
 sg13g2_buf_2 fanout405 (.A(_04225_),
    .X(net405));
 sg13g2_buf_2 fanout404 (.A(net405),
    .X(net404));
 sg13g2_buf_2 fanout403 (.A(_04251_),
    .X(net403));
 sg13g2_buf_2 fanout402 (.A(_04298_),
    .X(net402));
 sg13g2_buf_2 fanout401 (.A(_04298_),
    .X(net401));
 sg13g2_buf_2 fanout400 (.A(_04387_),
    .X(net400));
 sg13g2_buf_2 fanout399 (.A(net400),
    .X(net399));
 sg13g2_buf_2 fanout398 (.A(_01527_),
    .X(net398));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(_01527_));
 sg13g2_buf_2 fanout396 (.A(_01735_),
    .X(net396));
 sg13g2_buf_2 fanout395 (.A(net396),
    .X(net395));
 sg13g2_buf_4 fanout394 (.X(net394),
    .A(net395));
 sg13g2_buf_4 fanout393 (.X(net393),
    .A(net396));
 sg13g2_buf_4 fanout392 (.X(net392),
    .A(net393));
 sg13g2_buf_4 fanout391 (.X(net391),
    .A(net392));
 sg13g2_buf_4 fanout390 (.X(net390),
    .A(_01739_));
 sg13g2_buf_2 fanout389 (.A(net390),
    .X(net389));
 sg13g2_buf_4 fanout388 (.X(net388),
    .A(net389));
 sg13g2_buf_4 fanout387 (.X(net387),
    .A(net390));
 sg13g2_buf_2 fanout386 (.A(net390),
    .X(net386));
 sg13g2_buf_4 fanout385 (.X(net385),
    .A(net390));
 sg13g2_buf_4 fanout384 (.X(net384),
    .A(_01743_));
 sg13g2_buf_4 fanout383 (.X(net383),
    .A(net384));
 sg13g2_buf_4 fanout382 (.X(net382),
    .A(net384));
 sg13g2_buf_2 fanout381 (.A(net384),
    .X(net381));
 sg13g2_buf_4 fanout380 (.X(net380),
    .A(net381));
 sg13g2_buf_4 fanout379 (.X(net379),
    .A(_01747_));
 sg13g2_buf_2 fanout378 (.A(net379),
    .X(net378));
 sg13g2_buf_4 fanout377 (.X(net377),
    .A(net378));
 sg13g2_buf_4 fanout376 (.X(net376),
    .A(net379));
 sg13g2_buf_2 fanout375 (.A(net379),
    .X(net375));
 sg13g2_buf_4 fanout374 (.X(net374),
    .A(net379));
 sg13g2_buf_4 fanout373 (.X(net373),
    .A(_01751_));
 sg13g2_buf_4 fanout372 (.X(net372),
    .A(net373));
 sg13g2_buf_4 fanout371 (.X(net371),
    .A(net372));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(net371));
 sg13g2_buf_2 fanout369 (.A(_01755_),
    .X(net369));
 sg13g2_buf_4 fanout368 (.X(net368),
    .A(net369));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(_01755_));
 sg13g2_buf_2 fanout366 (.A(net367),
    .X(net366));
 sg13g2_buf_4 fanout365 (.X(net365),
    .A(net366));
 sg13g2_buf_2 fanout364 (.A(_01759_),
    .X(net364));
 sg13g2_buf_4 fanout363 (.X(net363),
    .A(net364));
 sg13g2_buf_2 fanout362 (.A(net364),
    .X(net362));
 sg13g2_buf_2 fanout361 (.A(net362),
    .X(net361));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(net362));
 sg13g2_buf_4 fanout359 (.X(net359),
    .A(net362));
 sg13g2_buf_4 fanout358 (.X(net358),
    .A(_01763_));
 sg13g2_buf_4 fanout357 (.X(net357),
    .A(_01763_));
 sg13g2_buf_4 fanout356 (.X(net356),
    .A(net357));
 sg13g2_buf_2 fanout355 (.A(net357),
    .X(net355));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(net357));
 sg13g2_buf_4 fanout353 (.X(net353),
    .A(_02250_));
 sg13g2_buf_1 fanout352 (.A(_02864_),
    .X(net352));
 sg13g2_buf_2 fanout351 (.A(_02864_),
    .X(net351));
 sg13g2_buf_2 fanout350 (.A(_02865_),
    .X(net350));
 sg13g2_buf_2 fanout349 (.A(net350),
    .X(net349));
 sg13g2_buf_2 fanout348 (.A(_03461_),
    .X(net348));
 sg13g2_buf_2 fanout347 (.A(net348),
    .X(net347));
 sg13g2_buf_2 fanout346 (.A(net347),
    .X(net346));
 sg13g2_buf_4 fanout345 (.X(net345),
    .A(net347));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(_03462_));
 sg13g2_buf_4 fanout343 (.X(net343),
    .A(net344));
 sg13g2_buf_2 fanout342 (.A(net343),
    .X(net342));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(net344));
 sg13g2_buf_2 fanout340 (.A(_04130_),
    .X(net340));
 sg13g2_buf_2 fanout339 (.A(_04313_),
    .X(net339));
 sg13g2_buf_4 fanout338 (.X(net338),
    .A(_05657_));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(net338));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(_02290_));
 sg13g2_buf_2 fanout335 (.A(_02290_),
    .X(net335));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(net336));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(_03485_));
 sg13g2_buf_2 fanout332 (.A(_03522_),
    .X(net332));
 sg13g2_buf_2 fanout331 (.A(_03838_),
    .X(net331));
 sg13g2_buf_2 fanout330 (.A(_04787_),
    .X(net330));
 sg13g2_buf_2 fanout329 (.A(net330),
    .X(net329));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(net329));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(net329));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(_04787_));
 sg13g2_buf_2 fanout325 (.A(net326),
    .X(net325));
 sg13g2_buf_2 fanout324 (.A(_05040_),
    .X(net324));
 sg13g2_buf_2 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(_05656_));
 sg13g2_buf_2 fanout321 (.A(net322),
    .X(net321));
 sg13g2_buf_8 fanout320 (.A(_01723_),
    .X(net320));
 sg13g2_buf_4 fanout319 (.X(net319),
    .A(_01723_));
 sg13g2_buf_4 fanout318 (.X(net318),
    .A(_01724_));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(_01724_));
 sg13g2_buf_4 fanout316 (.X(net316),
    .A(_02289_));
 sg13g2_buf_4 fanout315 (.X(net315),
    .A(net316));
 sg13g2_buf_2 fanout314 (.A(_02483_),
    .X(net314));
 sg13g2_buf_4 fanout313 (.X(net313),
    .A(net314));
 sg13g2_buf_2 fanout312 (.A(_02543_),
    .X(net312));
 sg13g2_buf_2 fanout311 (.A(_02543_),
    .X(net311));
 sg13g2_buf_2 fanout310 (.A(_02567_),
    .X(net310));
 sg13g2_buf_2 fanout309 (.A(net310),
    .X(net309));
 sg13g2_buf_2 fanout308 (.A(net310),
    .X(net308));
 sg13g2_buf_4 fanout307 (.X(net307),
    .A(_03082_));
 sg13g2_buf_2 fanout306 (.A(_02541_),
    .X(net306));
 sg13g2_buf_2 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_4 fanout304 (.X(net304),
    .A(_02545_));
 sg13g2_buf_2 fanout303 (.A(net304),
    .X(net303));
 sg13g2_buf_2 fanout302 (.A(net303),
    .X(net302));
 sg13g2_buf_4 fanout301 (.X(net301),
    .A(_03068_));
 sg13g2_buf_2 fanout300 (.A(net301),
    .X(net300));
 sg13g2_buf_2 fanout299 (.A(net300),
    .X(net299));
 sg13g2_buf_4 fanout298 (.X(net298),
    .A(net299));
 sg13g2_buf_4 fanout297 (.X(net297),
    .A(net300));
 sg13g2_buf_4 fanout296 (.X(net296),
    .A(_03069_));
 sg13g2_buf_2 fanout295 (.A(net296),
    .X(net295));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(_03070_));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(_03075_));
 sg13g2_buf_2 fanout292 (.A(_03078_),
    .X(net292));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(_03078_));
 sg13g2_buf_4 fanout290 (.X(net290),
    .A(_03080_));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(net290));
 sg13g2_buf_2 fanout288 (.A(_03083_),
    .X(net288));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(_03083_));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(_03486_));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(_03487_));
 sg13g2_buf_1 fanout284 (.A(_03537_),
    .X(net284));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(_03537_));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(_03588_));
 sg13g2_buf_2 fanout281 (.A(_03813_),
    .X(net281));
 sg13g2_buf_1 fanout280 (.A(_03813_),
    .X(net280));
 sg13g2_buf_2 fanout279 (.A(_03813_),
    .X(net279));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(_04303_));
 sg13g2_buf_2 fanout277 (.A(net278),
    .X(net277));
 sg13g2_buf_2 fanout276 (.A(net278),
    .X(net276));
 sg13g2_buf_2 fanout275 (.A(_04388_),
    .X(net275));
 sg13g2_buf_2 fanout274 (.A(net275),
    .X(net274));
 sg13g2_buf_2 fanout273 (.A(_04514_),
    .X(net273));
 sg13g2_buf_2 fanout272 (.A(net273),
    .X(net272));
 sg13g2_buf_2 fanout271 (.A(_04514_),
    .X(net271));
 sg13g2_buf_1 fanout270 (.A(net271),
    .X(net270));
 sg13g2_buf_2 fanout269 (.A(net270),
    .X(net269));
 sg13g2_buf_1 fanout268 (.A(net270),
    .X(net268));
 sg13g2_buf_2 fanout267 (.A(net270),
    .X(net267));
 sg13g2_buf_2 fanout266 (.A(_04723_),
    .X(net266));
 sg13g2_buf_2 fanout265 (.A(net266),
    .X(net265));
 sg13g2_buf_2 fanout264 (.A(net265),
    .X(net264));
 sg13g2_buf_2 fanout263 (.A(net266),
    .X(net263));
 sg13g2_buf_2 fanout262 (.A(net266),
    .X(net262));
 sg13g2_buf_2 fanout261 (.A(_04723_),
    .X(net261));
 sg13g2_buf_4 fanout260 (.X(net260),
    .A(_01725_));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(_01767_));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(_01777_));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(_01787_));
 sg13g2_buf_4 fanout256 (.X(net256),
    .A(_01800_));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(_01810_));
 sg13g2_buf_4 fanout254 (.X(net254),
    .A(_01821_));
 sg13g2_buf_2 fanout253 (.A(_01831_),
    .X(net253));
 sg13g2_buf_4 fanout252 (.X(net252),
    .A(_01842_));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(_01853_));
 sg13g2_buf_2 fanout250 (.A(net251),
    .X(net250));
 sg13g2_buf_2 fanout249 (.A(_01854_),
    .X(net249));
 sg13g2_buf_2 fanout248 (.A(net249),
    .X(net248));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(_01863_));
 sg13g2_buf_4 fanout246 (.X(net246),
    .A(_01873_));
 sg13g2_buf_4 fanout245 (.X(net245),
    .A(_01883_));
 sg13g2_buf_4 fanout244 (.X(net244),
    .A(_01893_));
 sg13g2_buf_4 fanout243 (.X(net243),
    .A(_01903_));
 sg13g2_buf_4 fanout242 (.X(net242),
    .A(_01913_));
 sg13g2_buf_2 fanout241 (.A(_01924_),
    .X(net241));
 sg13g2_buf_2 fanout240 (.A(_01924_),
    .X(net240));
 sg13g2_buf_4 fanout239 (.X(net239),
    .A(_01933_));
 sg13g2_buf_4 fanout238 (.X(net238),
    .A(_01943_));
 sg13g2_buf_4 fanout237 (.X(net237),
    .A(_01953_));
 sg13g2_buf_8 fanout236 (.A(_01963_),
    .X(net236));
 sg13g2_buf_4 fanout235 (.X(net235),
    .A(_01973_));
 sg13g2_buf_2 fanout234 (.A(_01983_),
    .X(net234));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(_01993_));
 sg13g2_buf_4 fanout232 (.X(net232),
    .A(_02003_));
 sg13g2_buf_8 fanout231 (.A(_02013_),
    .X(net231));
 sg13g2_buf_4 fanout230 (.X(net230),
    .A(_02023_));
 sg13g2_buf_8 fanout229 (.A(_02033_),
    .X(net229));
 sg13g2_buf_4 fanout228 (.X(net228),
    .A(_02043_));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(_02053_));
 sg13g2_buf_4 fanout226 (.X(net226),
    .A(_02063_));
 sg13g2_buf_4 fanout225 (.X(net225),
    .A(_02102_));
 sg13g2_buf_2 fanout224 (.A(_02115_),
    .X(net224));
 sg13g2_buf_2 fanout223 (.A(net224),
    .X(net223));
 sg13g2_buf_4 fanout222 (.X(net222),
    .A(_03087_));
 sg13g2_buf_4 fanout221 (.X(net221),
    .A(net222));
 sg13g2_buf_4 fanout220 (.X(net220),
    .A(net222));
 sg13g2_buf_2 fanout219 (.A(_03488_),
    .X(net219));
 sg13g2_buf_2 fanout218 (.A(net219),
    .X(net218));
 sg13g2_buf_2 fanout217 (.A(net218),
    .X(net217));
 sg13g2_buf_2 fanout216 (.A(net217),
    .X(net216));
 sg13g2_buf_2 fanout215 (.A(net219),
    .X(net215));
 sg13g2_buf_1 fanout214 (.A(net215),
    .X(net214));
 sg13g2_buf_2 fanout213 (.A(net219),
    .X(net213));
 sg13g2_buf_2 fanout212 (.A(_03512_),
    .X(net212));
 sg13g2_buf_4 fanout211 (.X(net211),
    .A(_03512_));
 sg13g2_buf_4 fanout210 (.X(net210),
    .A(_03517_));
 sg13g2_buf_1 fanout209 (.A(_03527_),
    .X(net209));
 sg13g2_buf_2 fanout208 (.A(net209),
    .X(net208));
 sg13g2_buf_4 fanout207 (.X(net207),
    .A(_03554_));
 sg13g2_buf_2 fanout206 (.A(_03582_),
    .X(net206));
 sg13g2_buf_4 fanout205 (.X(net205),
    .A(_03583_));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(_03593_));
 sg13g2_buf_4 fanout203 (.X(net203),
    .A(_05658_));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(net203));
 sg13g2_buf_2 fanout201 (.A(_01768_),
    .X(net201));
 sg13g2_buf_2 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_2 fanout199 (.A(_01778_),
    .X(net199));
 sg13g2_buf_2 fanout198 (.A(net199),
    .X(net198));
 sg13g2_buf_2 fanout197 (.A(_01904_),
    .X(net197));
 sg13g2_buf_2 fanout196 (.A(_01904_),
    .X(net196));
 sg13g2_buf_2 fanout195 (.A(_01914_),
    .X(net195));
 sg13g2_buf_1 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_2 fanout193 (.A(net195),
    .X(net193));
 sg13g2_buf_2 fanout192 (.A(_01954_),
    .X(net192));
 sg13g2_buf_2 fanout191 (.A(net192),
    .X(net191));
 sg13g2_buf_2 fanout190 (.A(_01974_),
    .X(net190));
 sg13g2_buf_2 fanout189 (.A(_01974_),
    .X(net189));
 sg13g2_buf_2 fanout188 (.A(_02044_),
    .X(net188));
 sg13g2_buf_2 fanout187 (.A(_02044_),
    .X(net187));
 sg13g2_buf_2 fanout186 (.A(_02064_),
    .X(net186));
 sg13g2_buf_2 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_2 fanout184 (.A(_02097_),
    .X(net184));
 sg13g2_buf_4 fanout183 (.X(net183),
    .A(_03105_));
 sg13g2_buf_2 fanout182 (.A(_03803_),
    .X(net182));
 sg13g2_buf_2 fanout181 (.A(_03803_),
    .X(net181));
 sg13g2_buf_2 fanout180 (.A(_04107_),
    .X(net180));
 sg13g2_buf_2 fanout179 (.A(_04124_),
    .X(net179));
 sg13g2_buf_2 fanout178 (.A(_04227_),
    .X(net178));
 sg13g2_buf_2 fanout177 (.A(net178),
    .X(net177));
 sg13g2_buf_2 fanout176 (.A(_04500_),
    .X(net176));
 sg13g2_buf_2 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_2 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_2 fanout173 (.A(net175),
    .X(net173));
 sg13g2_buf_2 fanout172 (.A(net175),
    .X(net172));
 sg13g2_buf_2 fanout171 (.A(net176),
    .X(net171));
 sg13g2_buf_2 fanout170 (.A(net171),
    .X(net170));
 sg13g2_buf_2 fanout169 (.A(net170),
    .X(net169));
 sg13g2_buf_2 fanout168 (.A(net176),
    .X(net168));
 sg13g2_buf_2 fanout167 (.A(net168),
    .X(net167));
 sg13g2_buf_2 fanout166 (.A(_01726_),
    .X(net166));
 sg13g2_buf_2 fanout165 (.A(_01726_),
    .X(net165));
 sg13g2_buf_2 fanout164 (.A(_01788_),
    .X(net164));
 sg13g2_buf_2 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_2 fanout162 (.A(_01801_),
    .X(net162));
 sg13g2_buf_2 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_2 fanout160 (.A(_01811_),
    .X(net160));
 sg13g2_buf_1 fanout159 (.A(net160),
    .X(net159));
 sg13g2_buf_2 fanout158 (.A(net159),
    .X(net158));
 sg13g2_buf_2 fanout157 (.A(_01822_),
    .X(net157));
 sg13g2_buf_1 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_2 fanout155 (.A(net157),
    .X(net155));
 sg13g2_buf_2 fanout154 (.A(_01832_),
    .X(net154));
 sg13g2_buf_2 fanout153 (.A(_01832_),
    .X(net153));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(_01843_));
 sg13g2_buf_2 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_2 fanout150 (.A(_01864_),
    .X(net150));
 sg13g2_buf_2 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_2 fanout148 (.A(_01874_),
    .X(net148));
 sg13g2_buf_2 fanout147 (.A(_01874_),
    .X(net147));
 sg13g2_buf_2 fanout146 (.A(_01884_),
    .X(net146));
 sg13g2_buf_2 fanout145 (.A(_01884_),
    .X(net145));
 sg13g2_buf_2 fanout144 (.A(_01894_),
    .X(net144));
 sg13g2_buf_2 fanout143 (.A(_01894_),
    .X(net143));
 sg13g2_buf_2 fanout142 (.A(_01934_),
    .X(net142));
 sg13g2_buf_2 fanout141 (.A(net142),
    .X(net141));
 sg13g2_buf_2 fanout140 (.A(_01944_),
    .X(net140));
 sg13g2_buf_2 fanout139 (.A(_01944_),
    .X(net139));
 sg13g2_buf_2 fanout138 (.A(_01964_),
    .X(net138));
 sg13g2_buf_2 fanout137 (.A(net138),
    .X(net137));
 sg13g2_buf_2 fanout136 (.A(_01984_),
    .X(net136));
 sg13g2_buf_2 fanout135 (.A(_01984_),
    .X(net135));
 sg13g2_buf_2 fanout134 (.A(_01994_),
    .X(net134));
 sg13g2_buf_2 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(_02004_));
 sg13g2_buf_2 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_2 fanout130 (.A(_02014_),
    .X(net130));
 sg13g2_buf_2 fanout129 (.A(net130),
    .X(net129));
 sg13g2_buf_2 fanout128 (.A(_02024_),
    .X(net128));
 sg13g2_buf_2 fanout127 (.A(net128),
    .X(net127));
 sg13g2_buf_2 fanout126 (.A(_02034_),
    .X(net126));
 sg13g2_buf_2 fanout125 (.A(net126),
    .X(net125));
 sg13g2_buf_2 fanout124 (.A(_02054_),
    .X(net124));
 sg13g2_buf_2 fanout123 (.A(_02054_),
    .X(net123));
 sg13g2_buf_2 fanout122 (.A(_02103_),
    .X(net122));
 sg13g2_buf_2 fanout121 (.A(net122),
    .X(net121));
 sg13g2_buf_2 fanout120 (.A(_03542_),
    .X(net120));
 sg13g2_buf_2 fanout119 (.A(_03542_),
    .X(net119));
 sg13g2_buf_2 fanout118 (.A(_03549_),
    .X(net118));
 sg13g2_buf_4 fanout117 (.X(net117),
    .A(_02982_));
 sg13g2_buf_2 fanout116 (.A(_03116_),
    .X(net116));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(_03117_));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(net115));
 sg13g2_buf_1 fanout113 (.A(_04517_),
    .X(net113));
 sg13g2_buf_2 fanout112 (.A(net113),
    .X(net112));
 sg13g2_buf_2 fanout111 (.A(net112),
    .X(net111));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(net113));
 sg13g2_buf_2 fanout109 (.A(_05628_),
    .X(net109));
 sg13g2_buf_2 fanout108 (.A(_03123_),
    .X(net108));
 sg13g2_buf_2 fanout107 (.A(_04169_),
    .X(net107));
 sg13g2_buf_2 fanout106 (.A(_03131_),
    .X(net106));
 sg13g2_buf_2 fanout105 (.A(net106),
    .X(net105));
 sg13g2_buf_2 fanout104 (.A(_05607_),
    .X(net104));
 sg13g2_buf_2 fanout103 (.A(_05608_),
    .X(net103));
 sg13g2_buf_2 fanout102 (.A(net103),
    .X(net102));
 sg13g2_buf_2 fanout101 (.A(_05615_),
    .X(net101));
 sg13g2_buf_2 fanout100 (.A(_05627_),
    .X(net100));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(_03465_));
 sg13g2_buf_1 fanout98 (.A(net99),
    .X(net98));
 sg13g2_buf_1 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_2 fanout96 (.A(net98),
    .X(net96));
 sg13g2_buf_2 fanout95 (.A(net98),
    .X(net95));
 sg13g2_buf_2 fanout94 (.A(_03466_),
    .X(net94));
 sg13g2_buf_1 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_2 fanout92 (.A(net94),
    .X(net92));
 sg13g2_buf_2 fanout91 (.A(net94),
    .X(net91));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(_04161_));
 sg13g2_buf_1 fanout89 (.A(_04162_),
    .X(net89));
 sg13g2_buf_4 fanout88 (.X(net88),
    .A(_04162_));
 sg13g2_buf_2 fanout87 (.A(_05836_),
    .X(net87));
 sg13g2_buf_2 fanout86 (.A(_03596_),
    .X(net86));
 sg13g2_buf_2 fanout85 (.A(net86),
    .X(net85));
 sg13g2_buf_2 fanout84 (.A(\debug_rd[0] ),
    .X(net84));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(\debug_rd[0] ));
 sg13g2_buf_2 fanout82 (.A(\debug_rd[2] ),
    .X(net82));
 sg13g2_buf_4 fanout81 (.X(net81),
    .A(\debug_rd[2] ));
 sg13g2_buf_4 fanout80 (.X(net80),
    .A(_03597_));
 sg13g2_buf_2 fanout79 (.A(net80),
    .X(net79));
 sg13g2_buf_2 fanout78 (.A(net80),
    .X(net78));
 sg13g2_buf_1 fanout77 (.A(_03598_),
    .X(net77));
 sg13g2_buf_2 fanout76 (.A(_03598_),
    .X(net76));
 sg13g2_buf_2 fanout75 (.A(\debug_rd[1] ),
    .X(net75));
 sg13g2_buf_4 fanout74 (.X(net74),
    .A(\debug_rd[1] ));
 sg13g2_buf_4 fanout73 (.X(net73),
    .A(_04296_));
 sg13g2_buf_2 fanout72 (.A(net73),
    .X(net72));
 sg13g2_buf_2 fanout71 (.A(_04297_),
    .X(net71));
 sg13g2_buf_4 fanout70 (.X(net70),
    .A(_04297_));
 sg13g2_buf_2 fanout69 (.A(_04363_),
    .X(net69));
 sg13g2_buf_2 fanout68 (.A(_05580_),
    .X(net68));
 sg13g2_buf_4 fanout67 (.X(net67),
    .A(_05581_));
 sg13g2_buf_2 fanout66 (.A(_05581_),
    .X(net66));
 sg13g2_buf_1 fanout65 (.A(_04166_),
    .X(net65));
 sg13g2_buf_2 fanout64 (.A(_04166_),
    .X(net64));
 sg13g2_buf_1 fanout63 (.A(_04299_),
    .X(net63));
 sg13g2_buf_2 fanout62 (.A(net63),
    .X(net62));
 sg13g2_buf_2 fanout61 (.A(net63),
    .X(net61));
 sg13g2_buf_1 fanout60 (.A(net63),
    .X(net60));
 sg13g2_buf_2 fanout59 (.A(net63),
    .X(net59));
 sg13g2_buf_4 fanout58 (.X(net58),
    .A(_05125_));
 sg13g2_buf_2 fanout57 (.A(net58),
    .X(net57));
 sg13g2_buf_2 fanout56 (.A(net57),
    .X(net56));
 sg13g2_buf_2 fanout55 (.A(_05349_),
    .X(net55));
 sg13g2_buf_2 fanout54 (.A(net55),
    .X(net54));
 sg13g2_buf_2 fanout53 (.A(net54),
    .X(net53));
 sg13g2_buf_2 fanout52 (.A(net55),
    .X(net52));
 sg13g2_buf_2 fanout51 (.A(net55),
    .X(net51));
 sg13g2_buf_4 fanout50 (.X(net50),
    .A(_05350_));
 sg13g2_buf_2 fanout49 (.A(net50),
    .X(net49));
 sg13g2_buf_2 fanout48 (.A(_05653_),
    .X(net48));
 sg13g2_buf_2 fanout47 (.A(net48),
    .X(net47));
 sg13g2_buf_2 fanout46 (.A(net47),
    .X(net46));
 sg13g2_buf_2 fanout45 (.A(net47),
    .X(net45));
 sg13g2_buf_2 fanout44 (.A(_04371_),
    .X(net44));
 sg13g2_buf_4 fanout43 (.X(net43),
    .A(net44));
 sg13g2_buf_2 fanout42 (.A(net44),
    .X(net42));
 sg13g2_buf_2 fanout41 (.A(net42),
    .X(net41));
 sg13g2_buf_2 fanout40 (.A(_04682_),
    .X(net40));
 sg13g2_buf_4 fanout39 (.X(net39),
    .A(net40));
 sg13g2_buf_2 fanout38 (.A(net40),
    .X(net38));
 sg13g2_buf_2 fanout37 (.A(net40),
    .X(net37));
 sg13g2_buf_2 fanout36 (.A(net37),
    .X(net36));
 sg13g2_buf_4 fanout35 (.X(net35),
    .A(_04776_));
 sg13g2_buf_2 fanout34 (.A(net35),
    .X(net34));
 sg13g2_buf_1 fanout33 (.A(net34),
    .X(net33));
 sg13g2_buf_2 fanout32 (.A(net34),
    .X(net32));
 sg13g2_buf_2 fanout31 (.A(net34),
    .X(net31));
 sg13g2_buf_2 fanout30 (.A(_04913_),
    .X(net30));
 sg13g2_buf_4 fanout29 (.X(net29),
    .A(_05652_));
 sg13g2_buf_1 fanout28 (.A(_05652_),
    .X(net28));
 sg13g2_buf_2 fanout27 (.A(net28),
    .X(net27));
 sg13g2_buf_1 fanout26 (.A(net28),
    .X(net26));
 sg13g2_buf_1 fanout25 (.A(net26),
    .X(net25));
 sg13g2_buf_2 fanout24 (.A(net26),
    .X(net24));
 sg13g2_buf_2 fanout23 (.A(net26),
    .X(net23));
 sg13g2_buf_2 fanout22 (.A(net23),
    .X(net22));
 sg13g2_buf_4 fanout21 (.X(net21),
    .A(net28));
 sg13g2_buf_2 fanout20 (.A(net21),
    .X(net20));
 sg13g2_buf_2 fanout19 (.A(_04366_),
    .X(net19));
 sg13g2_buf_4 fanout18 (.X(net18),
    .A(net19));
 sg13g2_buf_4 fanout17 (.X(net17),
    .A(net19));
 sg13g2_buf_2 fanout16 (.A(net17),
    .X(net16));
 sg13g2_buf_4 fanout15 (.X(net15),
    .A(\debug_rd[3] ));
 sg13g2_buf_4 fanout14 (.X(net14),
    .A(\debug_rd[3] ));
 sg13g2_buf_2 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_buf_2 input12 (.A(uio_in[4]),
    .X(net12));
 sg13g2_buf_2 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_2 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_4 input8 (.X(net8),
    .A(ui_in[6]));
 sg13g2_buf_4 input7 (.X(net7),
    .A(ui_in[5]));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[4]));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[3]));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[1]));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[0]));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 fanout657 (.A(net658),
    .X(net657));
 sg13g2_buf_4 fanout658 (.X(net658),
    .A(net659));
 sg13g2_buf_4 fanout659 (.X(net659),
    .A(net3907));
 sg13g2_buf_2 fanout660 (.A(net4122),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(net4078),
    .X(net661));
 sg13g2_buf_4 fanout662 (.X(net662),
    .A(net6));
 sg13g2_tiehi _14538__663 (.L_HI(net663));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_35_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_37_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_42_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_3_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_10_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_31_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_32_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_21_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_24_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_25_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_23_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_29_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_38_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_39_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_40_clk));
 sg13g2_inv_2 clkload21 (.A(clknet_leaf_41_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_4_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_5_clk));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_9_clk));
 sg13g2_inv_4 clkload25 (.A(clknet_leaf_12_clk));
 sg13g2_inv_2 clkload26 (.A(clknet_leaf_7_clk));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_8_clk));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_0_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_0_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_1_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_1_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_2_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_2_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_3_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_3_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_4_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_4_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_5_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_5_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_6_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_6_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_7_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_7_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_8_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_8_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_9_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_9_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_10_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_10_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_11_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_11_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_12_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_12_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_13_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_13_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_14_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_14_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_15_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_15_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_16_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_16_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_17_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_17_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_18_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_18_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_19_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_19_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_20_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_20_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_21_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_21_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_22_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_22_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_23_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_23_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_24_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_24_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_25_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_25_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_26_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_26_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_27_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_27_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_28_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_28_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_29_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_29_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_30_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_30_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_31_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_31_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_32_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_32_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_33_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_33_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_34_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_34_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_35_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_35_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_36_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_36_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_37_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_37_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_38_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_38_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_39_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_39_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_40_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_40_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_41_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_41_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_42_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_42_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_43_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_43_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_44_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_44_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_45_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_45_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_46_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_46_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_47_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_47_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_48_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_48_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_49_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_49_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_50_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_50_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_51_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_51_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_52_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_52_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_53_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_53_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_54_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_54_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_55_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_55_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_56_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_56_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_58_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_58_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_59_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_59_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_60_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_60_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_61_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_61_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_62_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_62_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_63_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_63_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_64_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_64_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_65_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_65_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_66_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_66_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_67_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_67_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_68_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_68_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_69_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_69_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_70_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_70_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_71_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_71_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_72_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_72_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_73_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_73_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_74_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_74_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_75_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_75_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_76_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_76_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_77_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_77_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_78_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_78_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_79_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_79_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_80_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_80_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_81_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_81_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_82_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_82_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_83_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_83_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_84_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_84_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_85_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_85_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_86_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_86_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_87_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_87_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_88_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_88_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_89_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_89_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_90_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_90_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_91_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_91_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_92_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_92_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_93_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_93_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_94_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_94_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_95_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_95_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_96_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_96_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_97_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_97_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_98_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_98_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_99_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_99_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_100_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_100_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_101_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_101_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_102_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_102_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_103_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_103_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_104_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_104_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_105_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_105_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_106_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_106_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_107_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_107_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_108_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_108_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_109_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_109_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_110_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_110_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_111_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_111_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_112_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_112_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_113_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_113_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_114_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_114_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_115_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_115_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_116_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_116_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_117_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_117_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_118_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_118_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_119_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_119_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_120_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_120_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_121_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_121_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_122_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_122_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_123_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_123_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_124_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_124_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_125_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_125_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_126_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_126_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_127_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_127_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_128_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_128_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_129_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_129_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_130_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_130_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_131_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_131_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_132_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_132_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_133_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_133_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_134_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_134_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_135_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_135_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_136_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_136_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_137_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_137_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_138_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_138_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_139_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_139_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_140_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_140_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_141_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_141_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_142_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_142_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_143_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_143_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_144_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_144_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_145_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_145_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_146_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_146_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_147_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_147_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_148_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_148_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_149_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_149_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_150_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_150_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_151_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_151_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_152_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_152_clk_regs));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_8 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_2 clkload30 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkload31 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkload32 (.A(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkload33 (.A(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkload34 (.A(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_1 clkload35 (.A(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_2 clkload36 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkload37 (.A(clknet_5_31__leaf_clk_regs));
 sg13g2_inv_8 clkload38 (.A(clknet_leaf_151_clk_regs));
 sg13g2_inv_1 clkload39 (.A(clknet_leaf_152_clk_regs));
 sg13g2_inv_4 clkload40 (.A(clknet_leaf_132_clk_regs));
 sg13g2_inv_2 clkload41 (.A(clknet_leaf_42_clk_regs));
 sg13g2_inv_1 clkload42 (.A(clknet_leaf_139_clk_regs));
 sg13g2_inv_4 clkload43 (.A(clknet_leaf_40_clk_regs));
 sg13g2_inv_1 clkload44 (.A(clknet_leaf_44_clk_regs));
 sg13g2_inv_2 clkload45 (.A(clknet_leaf_85_clk_regs));
 sg13g2_inv_4 clkload46 (.A(clknet_leaf_11_clk_regs));
 sg13g2_inv_1 clkload47 (.A(clknet_leaf_17_clk_regs));
 sg13g2_inv_4 clkload48 (.A(clknet_leaf_18_clk_regs));
 sg13g2_inv_1 clkload49 (.A(clknet_leaf_19_clk_regs));
 sg13g2_inv_1 clkload50 (.A(clknet_leaf_21_clk_regs));
 sg13g2_inv_1 clkload51 (.A(clknet_leaf_34_clk_regs));
 sg13g2_inv_1 clkload52 (.A(clknet_leaf_103_clk_regs));
 sg13g2_inv_1 clkload53 (.A(clknet_leaf_88_clk_regs));
 sg13g2_inv_4 clkload54 (.A(clknet_leaf_89_clk_regs));
 sg13g2_inv_4 clkload55 (.A(clknet_leaf_69_clk_regs));
 sg13g2_inv_4 clkload56 (.A(clknet_leaf_56_clk_regs));
 sg13g2_buf_8 rebuffer1 (.A(\addr[1] ),
    .X(net2380));
 sg13g2_buf_4 rebuffer2 (.X(net2381),
    .A(_02086_));
 sg13g2_dlygate4sd1_1 rebuffer3 (.A(net2381),
    .X(net2382));
 sg13g2_dlygate4sd1_1 rebuffer5 (.A(_01714_),
    .X(net2384));
 sg13g2_buf_1 rebuffer6 (.A(net2384),
    .X(net2385));
 sg13g2_dlygate4sd1_1 rebuffer7 (.A(\i_latch_mem.cycle[0] ),
    .X(net2386));
 sg13g2_dlygate4sd1_1 rebuffer8 (.A(\addr[0] ),
    .X(net2387));
 sg13g2_dlygate4sd1_1 rebuffer9 (.A(net2387),
    .X(net2388));
 sg13g2_dlygate4sd1_1 rebuffer10 (.A(\addr[0] ),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold11 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold12 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold13 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold15 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold16 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold17 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold18 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold19 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold21 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold22 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold23 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold24 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold25 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold26 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold27 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold28 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold29 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold31 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold33 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold34 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold35 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold36 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold37 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold38 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold39 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold40 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold41 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold42 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold43 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold44 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold45 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold46 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold47 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold48 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold49 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold50 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold51 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold52 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold53 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold54 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold55 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold56 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold57 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold58 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold59 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold60 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold61 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold62 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold63 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold64 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold65 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold66 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold67 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold68 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold69 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold71 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold72 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold73 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold74 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold75 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold76 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold77 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold78 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold79 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold80 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold81 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold83 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold84 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold85 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold86 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold87 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold88 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold89 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold90 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold91 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold92 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold93 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold94 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold95 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold96 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold97 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold98 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold100 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold101 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold102 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold103 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold104 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold105 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold106 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold107 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold108 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold109 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold110 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold111 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold112 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold113 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold114 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold115 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold116 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold117 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold119 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold120 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold121 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold122 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold123 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold124 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold125 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold126 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold127 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold128 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold129 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold130 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold131 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold132 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold133 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold134 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold135 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold136 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold137 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold138 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold139 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold140 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold141 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold142 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold143 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold144 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold145 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold146 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold147 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold148 (.A(\i_game.l_data.data_in[15] ),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold149 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold150 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold152 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold153 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold154 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold155 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold156 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold157 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold158 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold159 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold160 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold161 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold162 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold163 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold164 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold165 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold166 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold167 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold168 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold169 (.A(\i_game.l_data.data_in[0] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold170 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold171 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold172 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold173 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold174 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold175 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold176 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold177 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold178 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold179 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold180 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold181 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold182 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold183 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold184 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold185 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold186 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold187 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold188 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold189 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold190 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold191 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold192 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold193 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold194 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold195 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold196 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold197 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold198 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold199 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold200 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold201 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold202 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold203 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold204 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold205 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold206 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold207 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold208 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold209 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold210 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold211 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold212 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold213 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold214 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold215 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold216 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold217 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold218 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold219 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold220 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold221 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold222 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold223 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold224 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold225 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold226 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold227 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold228 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold229 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold230 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold231 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold232 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold233 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold234 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold235 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold236 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold237 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold238 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold239 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold240 (.A(\i_game.l_data.data_in[2] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold241 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold242 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold243 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold244 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold245 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold246 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold247 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold248 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold249 (.A(\i_game.l_data.data_in[14] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold250 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold251 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold252 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold253 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold254 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold255 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold256 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold257 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold258 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold259 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold260 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold261 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold262 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold263 (.A(\i_game.l_data.data_in[4] ),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold264 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold265 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold266 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold267 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold268 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold269 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold270 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold271 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold272 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold273 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold274 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold275 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold276 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold277 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold278 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold279 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold280 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold281 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold282 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold283 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold284 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold285 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold286 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold287 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold288 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold289 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold290 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold291 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold292 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold293 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold294 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold295 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold296 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold297 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold298 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold299 (.A(\i_game.l_data.data_in[21] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold300 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold301 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold302 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold303 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold304 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold305 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold306 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold307 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold308 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold309 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold310 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold311 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold312 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold313 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold314 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold315 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold316 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold317 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold318 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold319 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold320 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold321 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold322 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold323 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold324 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold325 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold326 (.A(\i_game.l_data.data_in[8] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold327 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold328 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold329 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold330 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold331 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold332 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold333 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold334 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold335 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold336 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold337 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold338 (.A(\i_game.l_data.data_in[16] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold339 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold340 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold341 (.A(\i_game.l_data.data_in[13] ),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold342 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold343 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold344 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold345 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold346 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold347 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold348 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold349 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold350 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold351 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold352 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold353 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold354 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold355 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold356 (.A(\i_game.l_data.data_in[7] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold357 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold358 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold359 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold360 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold361 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold362 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold363 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold364 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold365 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold366 (.A(\i_game.l_data.data_in[22] ),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold367 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold368 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold369 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold370 (.A(\i_game.l_data.data_in[10] ),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold371 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold372 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold373 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold374 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold375 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold376 (.A(\i_game.l_data.data_in[1] ),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold377 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold378 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold379 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold380 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold381 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold382 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold383 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold384 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold385 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold386 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold387 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold388 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold389 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold390 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold391 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold392 (.A(\i_game.l_data.data_in[20] ),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold393 (.A(\i_game.l_data.data_in[9] ),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold394 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold395 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold396 (.A(\i_game.l_data.data_in[17] ),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold397 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold398 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold399 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold400 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold401 (.A(\i_game.l_data.data_in[19] ),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold402 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold403 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold404 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold405 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold406 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold407 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold408 (.A(\i_game.l_data.data_in[3] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold409 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold410 (.A(\i_game.l_data.data_in[12] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold411 (.A(\i_game.l_data.data_in[5] ),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold412 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold413 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold414 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold415 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold416 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold417 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold418 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold419 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold420 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold421 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold422 (.A(\i_game.l_data.data_in[11] ),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold423 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold424 (.A(\i_game.l_data.data_in[18] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold425 (.A(\i_game.l_data.data_in[6] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold426 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold427 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold428 (.A(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold429 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold430 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold431 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold432 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold433 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold434 (.A(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold435 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold436 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold437 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold438 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold439 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold440 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold441 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold442 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold443 (.A(_00269_),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold444 (.A(_00267_),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold445 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold446 (.A(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold447 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold448 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold449 (.A(\mhz_clk_sync[2] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold450 (.A(_01485_),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold451 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold452 (.A(_00271_),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold453 (.A(_00607_),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold454 (.A(_00270_),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold455 (.A(_00637_),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold456 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold457 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold458 (.A(\i_tinyqv.mem.q_ctrl.stop_txn_reg ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold459 (.A(_00681_),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold460 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold461 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold462 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold463 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold464 (.A(_00268_),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold465 (.A(_04413_),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold466 (.A(_00706_),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold467 (.A(\i_game.game_latch_sync[0] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold468 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[7] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold469 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[7] ),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold470 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[0] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold471 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[1] ),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold472 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[5] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold473 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[2] ),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold474 (.A(\i_tinyqv.cpu.instr_data[3][11] ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold475 (.A(_01119_),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold476 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[0] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold477 (.A(\i_debug_uart_tx.cycle_counter[4] ),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold478 (.A(_00710_),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold479 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[4] ),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold480 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[3] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold481 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[3] ),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold482 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[0] ),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold483 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[1] ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold484 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[1] ),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold485 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[0] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold486 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[4] ),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold487 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[0] ),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold488 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[6] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold489 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[4] ),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold490 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[7] ),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold491 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[1] ),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold492 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[5] ),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold493 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[6] ),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold494 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[2] ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold495 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[0] ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold496 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[0] ),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold497 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[4] ),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold498 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[0] ),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold499 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[2] ),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold500 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[1] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold501 (.A(\i_tinyqv.cpu.instr_data[3][8] ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold502 (.A(_01116_),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold503 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[0] ),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold504 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[3] ),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold505 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[6] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold506 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[1] ),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold507 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[6] ),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold508 (.A(\i_tinyqv.cpu.instr_data[3][13] ),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold509 (.A(_01121_),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold510 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[3] ),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold511 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[0] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold512 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[2] ),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold513 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[5] ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold514 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[7] ),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold515 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[0] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold516 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[6] ),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold517 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[3] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold518 (.A(\i_tinyqv.cpu.instr_data[3][12] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold519 (.A(_01120_),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold520 (.A(\i_tinyqv.cpu.instr_data[3][5] ),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold521 (.A(_01113_),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold522 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[0] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold523 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[2] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold524 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[6] ),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold525 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[3] ),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold526 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[3] ),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold527 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[1] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold528 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[2] ),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold529 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[2] ),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold530 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[5] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold531 (.A(\i_tinyqv.cpu.instr_data[3][9] ),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold532 (.A(_01117_),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold533 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[0] ),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold534 (.A(\mhz_clk_sync[1] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold535 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[1] ),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold536 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[5] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold537 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[5] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold538 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[4] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold539 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[6] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold540 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[2] ),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold541 (.A(\i_tinyqv.cpu.instr_data[3][14] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold542 (.A(_01122_),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold543 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[6] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold544 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[1] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold545 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[1] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold546 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[7] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold547 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[7] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold548 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[6] ),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold549 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[0] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold550 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[3] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold551 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[2] ),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold552 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[3] ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold553 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[7] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold554 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[0] ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold555 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[5] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold556 (.A(\i_uart_rx.rxd_reg[1] ),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold557 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[3] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold558 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[0] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold559 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[6] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold560 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[6] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold561 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[4] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold562 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[2] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold563 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[1] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold564 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[2] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold565 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[4] ),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold566 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[3] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold567 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[3] ),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold568 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[1] ),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold569 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[5] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold570 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[7] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold571 (.A(\i_tinyqv.cpu.instr_data[3][15] ),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold572 (.A(_01123_),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold573 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[5] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold574 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[7] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold575 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[5] ),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold576 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[6] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold577 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[3] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold578 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[5] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold579 (.A(\i_pwm.l_pwm_level.data_out[0] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold580 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[4] ),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold581 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[3] ),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold582 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[4] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold583 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[4] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold584 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[5] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold585 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[2] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold586 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[7] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold587 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[7] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold588 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[7] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold589 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[3] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold590 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[5] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold591 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[7] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold592 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[2] ),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold593 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[7] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold594 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[5] ),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold595 (.A(\i_tinyqv.cpu.instr_data[3][10] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold596 (.A(_01118_),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold597 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[2] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold598 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[5] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold599 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[4] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold600 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[2] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold601 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[6] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold602 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[7] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold603 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[4] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold604 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[5] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold605 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[4] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold606 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[1] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold607 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[1] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold608 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[6] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold609 (.A(\i_tinyqv.mem.data_from_read[17] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold610 (.A(_01254_),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold611 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[7] ),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold612 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[7] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold613 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[4] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold614 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[0] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold615 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[4] ),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold616 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[4] ),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold617 (.A(\i_tinyqv.mem.data_from_read[20] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold618 (.A(_01257_),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold619 (.A(_00240_),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold620 (.A(_00636_),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold621 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[6] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold622 (.A(\i_latch_mem.data_out[11] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold623 (.A(_00033_),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold624 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[4] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold625 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[4] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold626 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[0] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold627 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[7] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold628 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[0] ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold629 (.A(\i_spi.clock_divider[0] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold630 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[6] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold631 (.A(\i_latch_mem.data_out[10] ),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold632 (.A(_00032_),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold633 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[7] ),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold634 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[7] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold635 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[6] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold636 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[5] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold637 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[7] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold638 (.A(\i_tinyqv.cpu.instr_data[1][9] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold639 (.A(_01167_),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold640 (.A(\i_tinyqv.mem.q_ctrl.addr[11] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold641 (.A(_01323_),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold642 (.A(\i_pwm.l_pwm_level.data_out[2] ),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold643 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[5] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold644 (.A(\i_tinyqv.cpu.instr_data[2][14] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold645 (.A(_00696_),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold646 (.A(\i_tinyqv.cpu.instr_data[2][10] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold647 (.A(_00692_),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold648 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[2] ),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold649 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[6] ),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold650 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[1] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold651 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[7] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold652 (.A(\i_tinyqv.cpu.instr_data[2][13] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold653 (.A(_00695_),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold654 (.A(\i_tinyqv.cpu.instr_data[1][13] ),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold655 (.A(_01171_),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold656 (.A(_00255_),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold657 (.A(_00625_),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold658 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[3] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold659 (.A(\i_tinyqv.cpu.instr_data[2][9] ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold660 (.A(_00691_),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold661 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[5] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold662 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[3] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold663 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[3] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold664 (.A(\i_tinyqv.cpu.instr_data[2][11] ),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold665 (.A(_00693_),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold666 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[2] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold667 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[6] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold668 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[2] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold669 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[0] ),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold670 (.A(\i_tinyqv.cpu.data_ready_sync ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold671 (.A(_01418_),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold672 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[0] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold673 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[4] ),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold674 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[7] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold675 (.A(\i_tinyqv.cpu.instr_data[0][9] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold676 (.A(_01103_),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold677 (.A(\i_tinyqv.cpu.instr_data[1][4] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold678 (.A(_01162_),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold679 (.A(\i_tinyqv.cpu.instr_data[1][6] ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold680 (.A(_01164_),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold681 (.A(\i_tinyqv.cpu.instr_data[0][4] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold682 (.A(_01098_),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold683 (.A(\i_tinyqv.cpu.instr_data[2][6] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold684 (.A(_00688_),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold685 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[3] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold686 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[3] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold687 (.A(\i_tinyqv.cpu.instr_data[0][14] ),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold688 (.A(_01108_),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold689 (.A(\i_tinyqv.cpu.instr_data[1][7] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold690 (.A(_01165_),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold691 (.A(\i_tinyqv.cpu.instr_data[0][7] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold692 (.A(_01101_),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold693 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[5] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold694 (.A(\i_tinyqv.cpu.instr_data[2][7] ),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold695 (.A(_00689_),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold696 (.A(\i_spi.clock_divider[2] ),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold697 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[1] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold698 (.A(\i_tinyqv.mem.data_from_read[22] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold699 (.A(_01259_),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold700 (.A(\i_tinyqv.cpu.instr_data[1][8] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold701 (.A(_01166_),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold702 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[3] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold703 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[7] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold704 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[4] ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold705 (.A(\i_pwm.l_pwm_level.data_out[1] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold707 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[4] ),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold708 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[0] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold709 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[5] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold710 (.A(\i_tinyqv.cpu.instr_data[2][5] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold711 (.A(_00687_),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold712 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[3] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold713 (.A(\i_tinyqv.mem.data_from_read[21] ),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold714 (.A(_01258_),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold715 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[6] ),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold716 (.A(\i_spi.clock_divider[1] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold717 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[0] ),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold718 (.A(\i_tinyqv.cpu.instr_data[0][11] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold719 (.A(_01105_),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold720 (.A(\mhz_clk_sync[0] ),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold721 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[7] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold722 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[6] ),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold723 (.A(\i_spi.spi_select ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold724 (.A(_04479_),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold725 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[4] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold726 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[7] ),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold727 (.A(\i_tinyqv.cpu.instr_data[2][8] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold728 (.A(_00690_),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold729 (.A(\i_tinyqv.cpu.instr_data[0][5] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold730 (.A(_01099_),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold731 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[2] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold732 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[5] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold733 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[4] ),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold734 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[1] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold735 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[1] ),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold736 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[6] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold737 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[1] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold738 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[0] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold739 (.A(\i_tinyqv.cpu.instr_data[1][12] ),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold740 (.A(_01170_),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold741 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[3] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold742 (.A(\i_tinyqv.cpu.instr_data[0][6] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold743 (.A(_01100_),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold744 (.A(\i_tinyqv.cpu.instr_data[2][15] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold745 (.A(_00697_),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold746 (.A(\i_tinyqv.cpu.instr_data[0][13] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold747 (.A(_01107_),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold748 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[3] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold749 (.A(\i_tinyqv.cpu.instr_data[1][10] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold750 (.A(_01168_),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold751 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[1] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold752 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[1] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold753 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[0] ),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold754 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[2] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold755 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[0] ),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold756 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[7] ),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold757 (.A(\gpio_out[7] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold758 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[1] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold759 (.A(\i_uart_tx.cycle_counter[1] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold760 (.A(_04254_),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold761 (.A(_00638_),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold762 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[1] ),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold763 (.A(\i_latch_mem.data_out[12] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold764 (.A(_00034_),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold765 (.A(\i_tinyqv.cpu.instr_data[0][10] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold766 (.A(_01104_),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold767 (.A(\i_spi.clock_divider[3] ),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold768 (.A(\i_tinyqv.cpu.instr_data[1][11] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold769 (.A(_01169_),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold770 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[6] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold771 (.A(\i_tinyqv.cpu.instr_data[1][14] ),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold772 (.A(_01172_),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold773 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[2] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold774 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[4] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold775 (.A(\i_tinyqv.mem.data_from_read[18] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold776 (.A(_01255_),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold777 (.A(\i_tinyqv.cpu.i_core.mie[3] ),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold778 (.A(_01085_),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold779 (.A(\i_tinyqv.cpu.instr_data[0][15] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold780 (.A(_01109_),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold781 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[6] ),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold782 (.A(\i_spi.spi_dc ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold783 (.A(_00726_),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold784 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[3] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold785 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[5] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold786 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[5] ),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold787 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[6] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold788 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[2] ),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold789 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[2] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold790 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[1] ),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold791 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[3] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold792 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[1] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold793 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[5] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold794 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[3] ),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold795 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[4] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold796 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[0] ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold797 (.A(\i_tinyqv.cpu.instr_data[0][8] ),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold798 (.A(_01102_),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold799 (.A(\i_tinyqv.cpu.load_started ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold800 (.A(_01414_),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold801 (.A(\i_tinyqv.cpu.instr_data[2][12] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold802 (.A(_00694_),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold803 (.A(\i_latch_mem.data_out[15] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold804 (.A(_00037_),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold805 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[3] ),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold806 (.A(\i_tinyqv.cpu.imm[24] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold807 (.A(\i_pwm.l_pwm_level.data_out[3] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold808 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[3] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold809 (.A(\i_pwm.l_pwm_level.data_out[7] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold810 (.A(\i_tinyqv.cpu.instr_data[1][15] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold811 (.A(_01173_),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold812 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[5] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold813 (.A(\i_tinyqv.cpu.imm[28] ),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold814 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[5] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold815 (.A(\i_tinyqv.cpu.instr_data[0][12] ),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold816 (.A(_01106_),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold817 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[4] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold818 (.A(\i_tinyqv.cpu.instr_data[1][5] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold819 (.A(_01163_),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold820 (.A(\i_tinyqv.cpu.instr_data[3][1] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold821 (.A(_00683_),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold822 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[1] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold823 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[2] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold824 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[6] ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold825 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[2] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold826 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[6] ),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold827 (.A(\addr[27] ),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold828 (.A(_04722_),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold829 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[1] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold830 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[3] ),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold831 (.A(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold832 (.A(_04103_),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold833 (.A(_00608_),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold834 (.A(\gpio_out[4] ),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold835 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[5] ),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold836 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[5] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold837 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[1] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold838 (.A(\i_tinyqv.cpu.additional_mem_ops[2] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold839 (.A(\i_tinyqv.cpu.instr_data[2][4] ),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold840 (.A(_00686_),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold841 (.A(\i_latch_mem.data_out[24] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold842 (.A(_00047_),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold843 (.A(\i_latch_mem.data_out[17] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold844 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[0] ),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold845 (.A(\i_latch_mem.data_out[3] ),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold846 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[2] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold847 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[0] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold848 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[4] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold849 (.A(\i_latch_mem.data_out[22] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold850 (.A(\i_latch_mem.data_out[14] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold851 (.A(_00036_),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold852 (.A(\i_latch_mem.data_out[31] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold853 (.A(_00055_),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold854 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[2] ),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold855 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[4] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold856 (.A(\gpio_out[3] ),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold857 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[1] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold858 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[2] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold859 (.A(\i_latch_mem.data_out[25] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold860 (.A(_00048_),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold861 (.A(\gpio_out[2] ),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold862 (.A(\gpio_out[0] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold863 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[2] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold864 (.A(\controller1_data[3] ),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold865 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[0] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold866 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[7] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold867 (.A(\i_pwm.l_pwm_level.data_out[5] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold868 (.A(\i_latch_mem.data_out[28] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold869 (.A(_00051_),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold870 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold871 (.A(_01292_),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold872 (.A(\i_time.l_mtimecmp.data_out[0] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold873 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[6] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold874 (.A(\i_tinyqv.mem.q_ctrl.addr[14] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold875 (.A(_01326_),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold876 (.A(\i_latch_mem.data_out[26] ),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold877 (.A(_00049_),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold878 (.A(\i_latch_mem.data_out[30] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold879 (.A(_00054_),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold880 (.A(\i_spi.end_txn_reg ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold881 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[6] ),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold882 (.A(\controller2_data[5] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold883 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[3] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold884 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold885 (.A(_01294_),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold886 (.A(\i_pwm.l_pwm_level.data_out[6] ),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold887 (.A(\controller2_data[9] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold888 (.A(\i_tinyqv.mem.q_ctrl.addr[0] ),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold889 (.A(\i_latch_mem.data_out[29] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold890 (.A(_00052_),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold891 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold892 (.A(_01291_),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold893 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[1] ),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold894 (.A(\controller1_data[8] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold895 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[6] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold896 (.A(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold897 (.A(_00617_),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold898 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[4] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold899 (.A(\i_latch_mem.data_out[16] ),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold900 (.A(\i_tinyqv.mem.q_ctrl.addr[1] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold901 (.A(_01313_),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold902 (.A(\controller1_data[10] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold903 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[2] ),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold904 (.A(\controller2_data[10] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold905 (.A(\i_latch_mem.data_out[7] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold906 (.A(\i_spi.data[7] ),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold907 (.A(_01131_),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold908 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[5] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold909 (.A(\i_latch_mem.data_out[27] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold910 (.A(_00050_),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold911 (.A(\gpio_out[6] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold912 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[5] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold913 (.A(\i_tinyqv.cpu.i_core.load_done ),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold914 (.A(_00603_),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold915 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[6] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold916 (.A(\addr[23] ),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold917 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[1] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold918 (.A(\i_tinyqv.cpu.i_core.mcause[3] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold919 (.A(_04121_),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold920 (.A(\i_tinyqv.cpu.i_core.mcause[4] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold921 (.A(_04122_),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold922 (.A(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold923 (.A(_00616_),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold924 (.A(\i_tinyqv.cpu.instr_data[3][7] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold925 (.A(_01115_),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold926 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[4] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold927 (.A(\i_tinyqv.mem.qspi_data_buf[28] ),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold928 (.A(\gpio_out[5] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold929 (.A(\i_tinyqv.mem.data_from_read[16] ),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold930 (.A(_01253_),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold931 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold932 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[3] ),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold933 (.A(\controller1_data[2] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold934 (.A(\i_tinyqv.cpu.imm[31] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold935 (.A(\i_tinyqv.cpu.imm[27] ),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold936 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[0] ),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold937 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[2] ),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold938 (.A(\i_uart_rx.rxd_reg[0] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold939 (.A(_00673_),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold940 (.A(\addr[18] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold941 (.A(_01330_),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold942 (.A(\addr[19] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold943 (.A(_01331_),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold944 (.A(\controller2_data[6] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold945 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[7] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold946 (.A(\gpio_out[1] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold947 (.A(\i_latch_mem.data_out[6] ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold948 (.A(\i_pwm.l_pwm_level.data_out[4] ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold949 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[7] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold950 (.A(\addr[7] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold951 (.A(_01143_),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold952 (.A(\i_tinyqv.mem.data_from_read[23] ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold953 (.A(_01260_),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold954 (.A(\i_spi.spi_clk_out ),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold955 (.A(_04481_),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold956 (.A(\i_uart_rx.cycle_counter[0] ),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold957 (.A(_04314_),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold958 (.A(_00663_),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold959 (.A(\i_uart_rx.bit_sample ),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold960 (.A(_00659_),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold961 (.A(\i_tinyqv.cpu.instr_data[3][6] ),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold962 (.A(_01114_),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold963 (.A(\i_latch_mem.data_out[4] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold964 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold965 (.A(_01293_),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold966 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[0] ),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold967 (.A(\i_tinyqv.mem.q_ctrl.addr[9] ),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold968 (.A(_01321_),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold969 (.A(\controller2_data[2] ),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold970 (.A(debug_data_continue),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold971 (.A(_01230_),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold972 (.A(\i_tinyqv.mem.qspi_data_buf[12] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold973 (.A(\i_latch_mem.data_out[9] ),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold974 (.A(_00062_),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold975 (.A(\i_tinyqv.mem.q_ctrl.addr[15] ),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold976 (.A(_01327_),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold977 (.A(\i_tinyqv.cpu.instr_data[3][4] ),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold978 (.A(_01112_),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold979 (.A(\i_tinyqv.mem.qspi_data_buf[13] ),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold980 (.A(_01250_),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold981 (.A(\i_tinyqv.mem.data_from_read[19] ),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold982 (.A(_01256_),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold983 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[4] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold984 (.A(\i_tinyqv.mem.qspi_data_buf[31] ),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold985 (.A(_04910_),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold986 (.A(\i_debug_uart_tx.data_to_send[7] ),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold987 (.A(\i_tinyqv.mem.qspi_data_buf[11] ),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold988 (.A(_01248_),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold989 (.A(\i_latch_mem.data_out[2] ),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold990 (.A(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold991 (.A(\i_tinyqv.cpu.imm[29] ),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold992 (.A(\i_latch_mem.data_out[1] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold993 (.A(\i_tinyqv.mem.q_ctrl.addr[4] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold994 (.A(\controller1_data[9] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold995 (.A(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold996 (.A(\i_latch_mem.data_out[23] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold997 (.A(\i_time.l_mtimecmp.data_out[5] ),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold998 (.A(\i_tinyqv.cpu.instr_data[3][3] ),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold999 (.A(_01111_),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\i_tinyqv.mem.q_ctrl.addr[13] ),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold1001 (.A(_01325_),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\i_spi.clock_count[1] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold1003 (.A(_04448_),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold1004 (.A(_00717_),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\i_tinyqv.cpu.i_core.mcause[5] ),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold1006 (.A(_04123_),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\i_tinyqv.cpu.instr_data[3][0] ),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold1008 (.A(_00682_),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\i_tinyqv.cpu.i_core.load_top_bit ),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold1010 (.A(_00661_),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\i_tinyqv.mem.qspi_data_buf[29] ),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold1012 (.A(_04908_),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\i_latch_mem.data_out[5] ),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold1015 (.A(_01333_),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\i_tinyqv.cpu.i_core.is_double_fault_r ),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold1017 (.A(_00606_),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\controller2_data[3] ),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\i_latch_mem.data_out[0] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\i_tinyqv.mem.qspi_data_buf[10] ),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[7] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\i_spi.read_latency ),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\i_debug_uart_tx.data_to_send[5] ),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold1024 (.A(_04406_),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold1025 (.A(_00703_),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold1027 (.A(_01190_),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold1029 (.A(_01188_),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\i_tinyqv.mem.qspi_data_buf[30] ),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\i_tinyqv.mem.qspi_data_buf[15] ),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold1032 (.A(_01252_),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\i_tinyqv.mem.qspi_data_buf[14] ),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold1034 (.A(_01251_),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[2] ),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\i_tinyqv.mem.qspi_data_buf[9] ),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\i_tinyqv.mem.qspi_data_buf[8] ),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\controller1_data[1] ),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\i_tinyqv.cpu.instr_data[1][2] ),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold1040 (.A(_01160_),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\i_uart_rx.recieved_data[1] ),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold1042 (.A(_00652_),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[6] ),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\i_tinyqv.cpu.i_core.time_hi[2] ),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold1045 (.A(_00609_),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\i_tinyqv.cpu.i_core.mepc[19] ),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\i_latch_mem.data_out[8] ),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold1048 (.A(_00061_),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\i_uart_tx.data_to_send[4] ),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold1050 (.A(_04241_),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold1051 (.A(_00633_),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\i_debug_uart_tx.data_to_send[4] ),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold1054 (.A(_00702_),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\i_debug_uart_tx.cycle_counter[1] ),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold1056 (.A(_04416_),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold1057 (.A(_00707_),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\i_tinyqv.mem.qspi_data_buf[27] ),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold1059 (.A(_04906_),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold1061 (.A(_01186_),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\i_tinyqv.mem.q_ctrl.addr[12] ),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold1063 (.A(_01324_),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\i_tinyqv.cpu.imm[30] ),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\i_tinyqv.cpu.additional_mem_ops[0] ),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold1066 (.A(_01479_),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\i_debug_uart_tx.data_to_send[2] ),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold1068 (.A(_04397_),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\i_tinyqv.cpu.instr_data[0][3] ),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold1070 (.A(_01097_),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\i_latch_mem.data_out[20] ),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\i_tinyqv.mem.q_ctrl.addr[5] ),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\i_uart_tx.data_to_send[6] ),
    .X(net3452));
 sg13g2_dlygate4sd3_1 hold1074 (.A(_04247_),
    .X(net3453));
 sg13g2_dlygate4sd3_1 hold1075 (.A(_00635_),
    .X(net3454));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\i_tinyqv.mem.qspi_data_buf[25] ),
    .X(net3455));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[5] ),
    .X(net3456));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\i_tinyqv.mem.q_ctrl.addr[6] ),
    .X(net3457));
 sg13g2_dlygate4sd3_1 hold1079 (.A(_01318_),
    .X(net3458));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\i_debug_uart_tx.data_to_send[6] ),
    .X(net3459));
 sg13g2_dlygate4sd3_1 hold1081 (.A(_00704_),
    .X(net3460));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\i_spi.bits_remaining[0] ),
    .X(net3461));
 sg13g2_dlygate4sd3_1 hold1083 (.A(_00721_),
    .X(net3462));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\i_tinyqv.cpu.instr_data[1][3] ),
    .X(net3463));
 sg13g2_dlygate4sd3_1 hold1085 (.A(_01161_),
    .X(net3464));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .X(net3465));
 sg13g2_dlygate4sd3_1 hold1087 (.A(_01189_),
    .X(net3466));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[4] ),
    .X(net3467));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\i_tinyqv.mem.q_ctrl.addr[17] ),
    .X(net3468));
 sg13g2_dlygate4sd3_1 hold1090 (.A(_01329_),
    .X(net3469));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\i_tinyqv.mem.q_ctrl.addr[8] ),
    .X(net3470));
 sg13g2_dlygate4sd3_1 hold1092 (.A(_01320_),
    .X(net3471));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\i_uart_tx.data_to_send[3] ),
    .X(net3472));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\i_time.l_mtimecmp.data_out[1] ),
    .X(net3473));
 sg13g2_dlygate4sd3_1 hold1095 (.A(_01339_),
    .X(net3474));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\i_tinyqv.cpu.instr_data[2][3] ),
    .X(net3475));
 sg13g2_dlygate4sd3_1 hold1097 (.A(_00685_),
    .X(net3476));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\controller2_data[4] ),
    .X(net3477));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\i_debug_uart_tx.data_to_send[0] ),
    .X(net3478));
 sg13g2_dlygate4sd3_1 hold1100 (.A(_04391_),
    .X(net3479));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .X(net3480));
 sg13g2_dlygate4sd3_1 hold1102 (.A(_01198_),
    .X(net3481));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\i_latch_mem.data_out[18] ),
    .X(net3482));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\i_time.l_mtimecmp.data_out[6] ),
    .X(net3483));
 sg13g2_dlygate4sd3_1 hold1105 (.A(_01344_),
    .X(net3484));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\controller2_data[1] ),
    .X(net3485));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\i_uart_rx.recieved_data[5] ),
    .X(net3486));
 sg13g2_dlygate4sd3_1 hold1108 (.A(_00656_),
    .X(net3487));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\i_tinyqv.cpu.instr_data[0][2] ),
    .X(net3488));
 sg13g2_dlygate4sd3_1 hold1110 (.A(_01096_),
    .X(net3489));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\i_uart_rx.cycle_counter[6] ),
    .X(net3490));
 sg13g2_dlygate4sd3_1 hold1112 (.A(_04323_),
    .X(net3491));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\i_tinyqv.cpu.imm[25] ),
    .X(net3492));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\controller2_data[11] ),
    .X(net3493));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\i_uart_tx.data_to_send[2] ),
    .X(net3494));
 sg13g2_dlygate4sd3_1 hold1116 (.A(_00631_),
    .X(net3495));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\addr[20] ),
    .X(net3496));
 sg13g2_dlygate4sd3_1 hold1118 (.A(_01156_),
    .X(net3497));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\i_tinyqv.cpu.i_core.mepc[13] ),
    .X(net3498));
 sg13g2_dlygate4sd3_1 hold1120 (.A(_01219_),
    .X(net3499));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\i_tinyqv.mem.q_ctrl.addr[16] ),
    .X(net3500));
 sg13g2_dlygate4sd3_1 hold1122 (.A(_01328_),
    .X(net3501));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\i_uart_tx.data_to_send[0] ),
    .X(net3502));
 sg13g2_dlygate4sd3_1 hold1124 (.A(_04229_),
    .X(net3503));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\controller1_data[4] ),
    .X(net3504));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\i_uart_rx.recieved_data[6] ),
    .X(net3505));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\i_time.l_mtimecmp.data_out[3] ),
    .X(net3506));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\addr[8] ),
    .X(net3507));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\i_tinyqv.cpu.i_core.mepc[4] ),
    .X(net3508));
 sg13g2_dlygate4sd3_1 hold1130 (.A(_01206_),
    .X(net3509));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\controller1_data[0] ),
    .X(net3510));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\i_uart_rx.recieved_data[4] ),
    .X(net3511));
 sg13g2_dlygate4sd3_1 hold1133 (.A(_00655_),
    .X(net3512));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\i_tinyqv.cpu.i_core.mem_op[2] ),
    .X(net3513));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\i_uart_tx.data_to_send[5] ),
    .X(net3514));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .X(net3515));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\i_uart_tx.cycle_counter[7] ),
    .X(net3516));
 sg13g2_dlygate4sd3_1 hold1138 (.A(_04266_),
    .X(net3517));
 sg13g2_dlygate4sd3_1 hold1139 (.A(_00644_),
    .X(net3518));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\i_tinyqv.mem.qspi_data_buf[24] ),
    .X(net3519));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\i_tinyqv.cpu.i_core.mcause[2] ),
    .X(net3520));
 sg13g2_dlygate4sd3_1 hold1142 (.A(_04120_),
    .X(net3521));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\i_latch_mem.data_out[21] ),
    .X(net3522));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\i_debug_uart_tx.data_to_send[1] ),
    .X(net3523));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\i_tinyqv.cpu.additional_mem_ops[1] ),
    .X(net3524));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .X(net3525));
 sg13g2_dlygate4sd3_1 hold1147 (.A(_00624_),
    .X(net3526));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\i_uart_tx.data_to_send[1] ),
    .X(net3527));
 sg13g2_dlygate4sd3_1 hold1149 (.A(_00630_),
    .X(net3528));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\i_tinyqv.cpu.i_core.mepc[14] ),
    .X(net3529));
 sg13g2_dlygate4sd3_1 hold1151 (.A(_01220_),
    .X(net3530));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\i_spi.data[5] ),
    .X(net3531));
 sg13g2_dlygate4sd3_1 hold1153 (.A(_01129_),
    .X(net3532));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\i_uart_tx.cycle_counter[9] ),
    .X(net3533));
 sg13g2_dlygate4sd3_1 hold1155 (.A(_04270_),
    .X(net3534));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\i_uart_rx.recieved_data[2] ),
    .X(net3535));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\i_time.l_mtimecmp.data_out[19] ),
    .X(net3536));
 sg13g2_dlygate4sd3_1 hold1158 (.A(_00756_),
    .X(net3537));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .X(net3538));
 sg13g2_dlygate4sd3_1 hold1160 (.A(_01196_),
    .X(net3539));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\i_tinyqv.cpu.i_core.mepc[16] ),
    .X(net3540));
 sg13g2_dlygate4sd3_1 hold1162 (.A(_01222_),
    .X(net3541));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\i_latch_mem.data_out[19] ),
    .X(net3542));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\i_tinyqv.cpu.i_core.mepc[9] ),
    .X(net3543));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\i_time.l_mtimecmp.data_out[15] ),
    .X(net3544));
 sg13g2_dlygate4sd3_1 hold1166 (.A(_01353_),
    .X(net3545));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\i_tinyqv.cpu.i_core.mepc[8] ),
    .X(net3546));
 sg13g2_dlygate4sd3_1 hold1168 (.A(_01214_),
    .X(net3547));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\addr[22] ),
    .X(net3548));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\gpio_out_sel[3] ),
    .X(net3549));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\i_tinyqv.mem.q_ctrl.addr[7] ),
    .X(net3550));
 sg13g2_dlygate4sd3_1 hold1172 (.A(_01319_),
    .X(net3551));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[1] ),
    .X(net3552));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\addr[25] ),
    .X(net3553));
 sg13g2_dlygate4sd3_1 hold1175 (.A(_04720_),
    .X(net3554));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\i_debug_uart_tx.data_to_send[3] ),
    .X(net3555));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\gpio_out_sel[1] ),
    .X(net3556));
 sg13g2_dlygate4sd3_1 hold1178 (.A(_00009_),
    .X(net3557));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\i_tinyqv.cpu.instr_data[2][2] ),
    .X(net3558));
 sg13g2_dlygate4sd3_1 hold1180 (.A(_00684_),
    .X(net3559));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\i_tinyqv.cpu.i_core.mepc[10] ),
    .X(net3560));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\i_tinyqv.cpu.i_core.mepc[8] ),
    .X(net3561));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\i_tinyqv.mem.qspi_data_buf[26] ),
    .X(net3562));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\controller1_data[6] ),
    .X(net3563));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\i_tinyqv.cpu.i_core.mepc[18] ),
    .X(net3564));
 sg13g2_dlygate4sd3_1 hold1186 (.A(_04768_),
    .X(net3565));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\gpio_out_sel[6] ),
    .X(net3566));
 sg13g2_dlygate4sd3_1 hold1188 (.A(_00014_),
    .X(net3567));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\i_time.l_mtimecmp.data_out[4] ),
    .X(net3568));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\controller1_data[5] ),
    .X(net3569));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\addr[16] ),
    .X(net3570));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\i_time.l_mtimecmp.data_out[20] ),
    .X(net3571));
 sg13g2_dlygate4sd3_1 hold1193 (.A(_00757_),
    .X(net3572));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\addr[17] ),
    .X(net3573));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\i_tinyqv.cpu.i_core.mepc[12] ),
    .X(net3574));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\controller1_data[11] ),
    .X(net3575));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .X(net3576));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\gpio_out_sel[5] ),
    .X(net3577));
 sg13g2_dlygate4sd3_1 hold1199 (.A(_00013_),
    .X(net3578));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\i_tinyqv.cpu.i_core.mepc[17] ),
    .X(net3579));
 sg13g2_dlygate4sd3_1 hold1201 (.A(_01223_),
    .X(net3580));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\i_uart_tx.cycle_counter[8] ),
    .X(net3581));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\i_pwm.pwm_count[3] ),
    .X(net3582));
 sg13g2_dlygate4sd3_1 hold1204 (.A(_04490_),
    .X(net3583));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\i_pwm.pwm_count[2] ),
    .X(net3584));
 sg13g2_dlygate4sd3_1 hold1206 (.A(_04488_),
    .X(net3585));
 sg13g2_dlygate4sd3_1 hold1207 (.A(_00739_),
    .X(net3586));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\i_uart_rx.recieved_data[3] ),
    .X(net3587));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .X(net3588));
 sg13g2_dlygate4sd3_1 hold1210 (.A(_00086_),
    .X(net3589));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\i_tinyqv.cpu.instr_len[1] ),
    .X(net3590));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .X(net3591));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\i_time.l_mtimecmp.data_out[29] ),
    .X(net3592));
 sg13g2_dlygate4sd3_1 hold1214 (.A(_00766_),
    .X(net3593));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\i_uart_tx.cycle_counter[3] ),
    .X(net3594));
 sg13g2_dlygate4sd3_1 hold1216 (.A(_04258_),
    .X(net3595));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\i_uart_rx.cycle_counter[7] ),
    .X(net3596));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[7] ),
    .X(net3597));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\i_tinyqv.cpu.i_core.mcause[1] ),
    .X(net3598));
 sg13g2_dlygate4sd3_1 hold1220 (.A(_04118_),
    .X(net3599));
 sg13g2_dlygate4sd3_1 hold1221 (.A(_00611_),
    .X(net3600));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\i_uart_tx.cycle_counter[6] ),
    .X(net3601));
 sg13g2_dlygate4sd3_1 hold1223 (.A(_04264_),
    .X(net3602));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .X(net3603));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\addr[11] ),
    .X(net3604));
 sg13g2_dlygate4sd3_1 hold1226 (.A(_01147_),
    .X(net3605));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\i_latch_mem.data_out[13] ),
    .X(net3606));
 sg13g2_dlygate4sd3_1 hold1228 (.A(_00035_),
    .X(net3607));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\i_uart_tx.cycle_counter[5] ),
    .X(net3608));
 sg13g2_dlygate4sd3_1 hold1230 (.A(_04262_),
    .X(net3609));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\i_uart_rx.cycle_counter[3] ),
    .X(net3610));
 sg13g2_dlygate4sd3_1 hold1232 (.A(_04318_),
    .X(net3611));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\i_uart_tx.cycle_counter[4] ),
    .X(net3612));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\i_tinyqv.cpu.i_core.cycle[1] ),
    .X(net3613));
 sg13g2_dlygate4sd3_1 hold1235 (.A(_04098_),
    .X(net3614));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\i_tinyqv.cpu.i_core.mepc[22] ),
    .X(net3615));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\addr[15] ),
    .X(net3616));
 sg13g2_dlygate4sd3_1 hold1238 (.A(_01151_),
    .X(net3617));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\i_time.l_mtimecmp.data_out[2] ),
    .X(net3618));
 sg13g2_dlygate4sd3_1 hold1240 (.A(_01340_),
    .X(net3619));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\i_tinyqv.cpu.imm[26] ),
    .X(net3620));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\i_uart_tx.cycle_counter[2] ),
    .X(net3621));
 sg13g2_dlygate4sd3_1 hold1243 (.A(_04256_),
    .X(net3622));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\i_tinyqv.cpu.i_core.mepc[6] ),
    .X(net3623));
 sg13g2_dlygate4sd3_1 hold1245 (.A(_01208_),
    .X(net3624));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\i_tinyqv.cpu.i_core.mepc[23] ),
    .X(net3625));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\addr[12] ),
    .X(net3626));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\i_tinyqv.cpu.i_core.mepc[11] ),
    .X(net3627));
 sg13g2_dlygate4sd3_1 hold1249 (.A(_01213_),
    .X(net3628));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .X(net3629));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\i_time.l_mtimecmp.data_out[23] ),
    .X(net3630));
 sg13g2_dlygate4sd3_1 hold1252 (.A(_00760_),
    .X(net3631));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\i_tinyqv.mem.q_ctrl.addr[20] ),
    .X(net3632));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\gpio_out_sel[8] ),
    .X(net3633));
 sg13g2_dlygate4sd3_1 hold1255 (.A(_00016_),
    .X(net3634));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\addr[9] ),
    .X(net3635));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\i_time.l_mtimecmp.data_out[22] ),
    .X(net3636));
 sg13g2_dlygate4sd3_1 hold1258 (.A(_00759_),
    .X(net3637));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .X(net3638));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\controller2_data[8] ),
    .X(net3639));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\i_tinyqv.cpu.i_core.mepc[15] ),
    .X(net3640));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ),
    .X(net3641));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\i_uart_rx.fsm_state[2] ),
    .X(net3642));
 sg13g2_dlygate4sd3_1 hold1264 (.A(_00677_),
    .X(net3643));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[0] ),
    .X(net3644));
 sg13g2_dlygate4sd3_1 hold1266 (.A(_04090_),
    .X(net3645));
 sg13g2_dlygate4sd3_1 hold1267 (.A(_00599_),
    .X(net3646));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\i_time.l_mtimecmp.data_out[18] ),
    .X(net3647));
 sg13g2_dlygate4sd3_1 hold1269 (.A(_00755_),
    .X(net3648));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .X(net3649));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ),
    .X(net3650));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\i_debug_uart_tx.cycle_counter[3] ),
    .X(net3651));
 sg13g2_dlygate4sd3_1 hold1273 (.A(_04420_),
    .X(net3652));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\i_spi.data[0] ),
    .X(net3653));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\i_tinyqv.mem.q_ctrl.addr[2] ),
    .X(net3654));
 sg13g2_dlygate4sd3_1 hold1276 (.A(_05130_),
    .X(net3655));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\i_time.l_mtimecmp.data_out[30] ),
    .X(net3656));
 sg13g2_dlygate4sd3_1 hold1278 (.A(_00767_),
    .X(net3657));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\i_spi.clock_count[0] ),
    .X(net3658));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\i_tinyqv.cpu.i_core.mie[0] ),
    .X(net3659));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\i_time.l_mtimecmp.data_out[17] ),
    .X(net3660));
 sg13g2_dlygate4sd3_1 hold1282 (.A(_00754_),
    .X(net3661));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\i_time.l_mtimecmp.data_out[8] ),
    .X(net3662));
 sg13g2_dlygate4sd3_1 hold1284 (.A(_01346_),
    .X(net3663));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\addr[21] ),
    .X(net3664));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .X(net3665));
 sg13g2_dlygate4sd3_1 hold1287 (.A(_00201_),
    .X(net3666));
 sg13g2_dlygate4sd3_1 hold1288 (.A(_04954_),
    .X(net3667));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .X(net3668));
 sg13g2_dlygate4sd3_1 hold1290 (.A(_01191_),
    .X(net3669));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\i_spi.bits_remaining[3] ),
    .X(net3670));
 sg13g2_dlygate4sd3_1 hold1292 (.A(_04472_),
    .X(net3671));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .X(net3672));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .X(net3673));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\i_time.l_mtimecmp.data_out[7] ),
    .X(net3674));
 sg13g2_dlygate4sd3_1 hold1296 (.A(_01345_),
    .X(net3675));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\i_tinyqv.mem.q_ctrl.addr[3] ),
    .X(net3676));
 sg13g2_dlygate4sd3_1 hold1298 (.A(_05139_),
    .X(net3677));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\i_tinyqv.cpu.is_jal ),
    .X(net3678));
 sg13g2_dlygate4sd3_1 hold1300 (.A(_01428_),
    .X(net3679));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\i_spi.data[3] ),
    .X(net3680));
 sg13g2_dlygate4sd3_1 hold1302 (.A(_01127_),
    .X(net3681));
 sg13g2_dlygate4sd3_1 hold1303 (.A(_00242_),
    .X(net3682));
 sg13g2_dlygate4sd3_1 hold1304 (.A(_01124_),
    .X(net3683));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .X(net3684));
 sg13g2_dlygate4sd3_1 hold1306 (.A(_01187_),
    .X(net3685));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\i_tinyqv.mem.q_ctrl.fsm_state[0] ),
    .X(net3686));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\i_tinyqv.cpu.i_core.mie[1] ),
    .X(net3687));
 sg13g2_dlygate4sd3_1 hold1309 (.A(_01087_),
    .X(net3688));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\i_tinyqv.cpu.instr_data_in[1] ),
    .X(net3689));
 sg13g2_dlygate4sd3_1 hold1311 (.A(_01308_),
    .X(net3690));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\i_spi.data[4] ),
    .X(net3691));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .X(net3692));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\i_debug_uart_tx.cycle_counter[2] ),
    .X(net3693));
 sg13g2_dlygate4sd3_1 hold1315 (.A(_04418_),
    .X(net3694));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\i_time.l_mtimecmp.data_out[16] ),
    .X(net3695));
 sg13g2_dlygate4sd3_1 hold1317 (.A(_00753_),
    .X(net3696));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\controller2_data[0] ),
    .X(net3697));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\gpio_out_sel[2] ),
    .X(net3698));
 sg13g2_dlygate4sd3_1 hold1320 (.A(_00010_),
    .X(net3699));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\i_tinyqv.cpu.i_core.mepc[5] ),
    .X(net3700));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\i_time.l_mtimecmp.data_out[25] ),
    .X(net3701));
 sg13g2_dlygate4sd3_1 hold1323 (.A(_00762_),
    .X(net3702));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\i_spi.bits_remaining[2] ),
    .X(net3703));
 sg13g2_dlygate4sd3_1 hold1325 (.A(_04469_),
    .X(net3704));
 sg13g2_dlygate4sd3_1 hold1326 (.A(_00723_),
    .X(net3705));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\i_tinyqv.mem.q_ctrl.addr[23] ),
    .X(net3706));
 sg13g2_dlygate4sd3_1 hold1328 (.A(_05348_),
    .X(net3707));
 sg13g2_dlygate4sd3_1 hold1329 (.A(_01335_),
    .X(net3708));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\i_uart_rx.cycle_counter[8] ),
    .X(net3709));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\addr[13] ),
    .X(net3710));
 sg13g2_dlygate4sd3_1 hold1332 (.A(_01149_),
    .X(net3711));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\addr[10] ),
    .X(net3712));
 sg13g2_dlygate4sd3_1 hold1334 (.A(_01322_),
    .X(net3713));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\i_spi.data[2] ),
    .X(net3714));
 sg13g2_dlygate4sd3_1 hold1336 (.A(_01126_),
    .X(net3715));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\i_tinyqv.cpu.i_core.mepc[10] ),
    .X(net3716));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\i_tinyqv.cpu.instr_data[3][2] ),
    .X(net3717));
 sg13g2_dlygate4sd3_1 hold1339 (.A(_01110_),
    .X(net3718));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\i_tinyqv.cpu.i_core.mepc[7] ),
    .X(net3719));
 sg13g2_dlygate4sd3_1 hold1341 (.A(_01209_),
    .X(net3720));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\i_time.l_mtimecmp.data_out[24] ),
    .X(net3721));
 sg13g2_dlygate4sd3_1 hold1343 (.A(_00761_),
    .X(net3722));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\i_debug_uart_tx.fsm_state[2] ),
    .X(net3723));
 sg13g2_dlygate4sd3_1 hold1345 (.A(_00713_),
    .X(net3724));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\i_time.l_mtimecmp.data_out[28] ),
    .X(net3725));
 sg13g2_dlygate4sd3_1 hold1347 (.A(_00765_),
    .X(net3726));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\gpio_out_sel[0] ),
    .X(net3727));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\i_time.l_mtimecmp.data_out[13] ),
    .X(net3728));
 sg13g2_dlygate4sd3_1 hold1350 (.A(_01351_),
    .X(net3729));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\i_tinyqv.cpu.instr_data[1][1] ),
    .X(net3730));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\i_tinyqv.cpu.instr_data[0][1] ),
    .X(net3731));
 sg13g2_dlygate4sd3_1 hold1353 (.A(\i_spi.data[1] ),
    .X(net3732));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\controller1_data[7] ),
    .X(net3733));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\i_tinyqv.cpu.instr_data_start[13] ),
    .X(net3734));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\i_tinyqv.mem.q_ctrl.addr[18] ),
    .X(net3735));
 sg13g2_dlygate4sd3_1 hold1357 (.A(_05340_),
    .X(net3736));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .X(net3737));
 sg13g2_dlygate4sd3_1 hold1359 (.A(_01174_),
    .X(net3738));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\i_uart_rx.cycle_counter[5] ),
    .X(net3739));
 sg13g2_dlygate4sd3_1 hold1361 (.A(_04322_),
    .X(net3740));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\controller2_data[7] ),
    .X(net3741));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\gpio_out_sel[4] ),
    .X(net3742));
 sg13g2_dlygate4sd3_1 hold1364 (.A(_00012_),
    .X(net3743));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\i_uart_rx.cycle_counter[4] ),
    .X(net3744));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\i_uart_rx.cycle_counter[2] ),
    .X(net3745));
 sg13g2_dlygate4sd3_1 hold1367 (.A(_04316_),
    .X(net3746));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\i_time.l_mtimecmp.data_out[11] ),
    .X(net3747));
 sg13g2_dlygate4sd3_1 hold1369 (.A(_01349_),
    .X(net3748));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\i_uart_tx.fsm_state[3] ),
    .X(net3749));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .X(net3750));
 sg13g2_dlygate4sd3_1 hold1372 (.A(_00243_),
    .X(net3751));
 sg13g2_dlygate4sd3_1 hold1373 (.A(_04347_),
    .X(net3752));
 sg13g2_dlygate4sd3_1 hold1374 (.A(_00675_),
    .X(net3753));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .X(net3754));
 sg13g2_dlygate4sd3_1 hold1376 (.A(_04863_),
    .X(net3755));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\i_tinyqv.cpu.i_core.mepc[20] ),
    .X(net3756));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\i_time.l_mtimecmp.data_out[21] ),
    .X(net3757));
 sg13g2_dlygate4sd3_1 hold1379 (.A(_00758_),
    .X(net3758));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\i_tinyqv.cpu.i_core.mie[4] ),
    .X(net3759));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\i_pwm.pwm_count[1] ),
    .X(net3760));
 sg13g2_dlygate4sd3_1 hold1382 (.A(_04486_),
    .X(net3761));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\i_uart_rx.cycle_counter[9] ),
    .X(net3762));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\i_tinyqv.cpu.i_core.mip[1] ),
    .X(net3763));
 sg13g2_dlygate4sd3_1 hold1385 (.A(_01089_),
    .X(net3764));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\i_spi.clock_count[3] ),
    .X(net3765));
 sg13g2_dlygate4sd3_1 hold1387 (.A(_04451_),
    .X(net3766));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .X(net3767));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\i_tinyqv.cpu.i_core.cycle[0] ),
    .X(net3768));
 sg13g2_dlygate4sd3_1 hold1390 (.A(_00604_),
    .X(net3769));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .X(net3770));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\data_to_write[19] ),
    .X(net3771));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .X(net3772));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\i_tinyqv.cpu.i_core.mip[0] ),
    .X(net3773));
 sg13g2_dlygate4sd3_1 hold1395 (.A(_01090_),
    .X(net3774));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\i_time.l_mtimecmp.data_out[31] ),
    .X(net3775));
 sg13g2_dlygate4sd3_1 hold1397 (.A(_00768_),
    .X(net3776));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .X(net3777));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\i_time.l_mtimecmp.data_out[10] ),
    .X(net3778));
 sg13g2_dlygate4sd3_1 hold1400 (.A(_01348_),
    .X(net3779));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\i_uart_rx.recieved_data[7] ),
    .X(net3780));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\i_pwm.pwm_count[5] ),
    .X(net3781));
 sg13g2_dlygate4sd3_1 hold1403 (.A(_04493_),
    .X(net3782));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\i_tinyqv.cpu.instr_len[2] ),
    .X(net3783));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .X(net3784));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\i_pwm.pwm_count[4] ),
    .X(net3785));
 sg13g2_dlygate4sd3_1 hold1407 (.A(\i_tinyqv.cpu.instr_data_in[5] ),
    .X(net3786));
 sg13g2_dlygate4sd3_1 hold1408 (.A(_01242_),
    .X(net3787));
 sg13g2_dlygate4sd3_1 hold1409 (.A(\i_tinyqv.cpu.instr_data_in[12] ),
    .X(net3788));
 sg13g2_dlygate4sd3_1 hold1410 (.A(_01241_),
    .X(net3789));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\i_tinyqv.cpu.no_write_in_progress ),
    .X(net3790));
 sg13g2_dlygate4sd3_1 hold1412 (.A(_01413_),
    .X(net3791));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\data_to_write[26] ),
    .X(net3792));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\i_spi.clock_count[2] ),
    .X(net3793));
 sg13g2_dlygate4sd3_1 hold1415 (.A(\i_debug_uart_tx.fsm_state[3] ),
    .X(net3794));
 sg13g2_dlygate4sd3_1 hold1416 (.A(_04434_),
    .X(net3795));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .X(net3796));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\i_time.l_mtimecmp.data_out[27] ),
    .X(net3797));
 sg13g2_dlygate4sd3_1 hold1419 (.A(_00764_),
    .X(net3798));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\i_tinyqv.mem.q_ctrl.spi_clk_pos ),
    .X(net3799));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\data_to_write[12] ),
    .X(net3800));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\i_tinyqv.mem.q_ctrl.spi_clk_use_neg ),
    .X(net3801));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .X(net3802));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\addr[14] ),
    .X(net3803));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\i_tinyqv.cpu.instr_data[2][0] ),
    .X(net3804));
 sg13g2_dlygate4sd3_1 hold1426 (.A(_01307_),
    .X(net3805));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\i_uart_tx.cycle_counter[10] ),
    .X(net3806));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\i_pwm.pwm_count[6] ),
    .X(net3807));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\gpio_out_sel[9] ),
    .X(net3808));
 sg13g2_dlygate4sd3_1 hold1430 (.A(_00017_),
    .X(net3809));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\i_tinyqv.cpu.i_core.mepc[1] ),
    .X(net3810));
 sg13g2_dlygate4sd3_1 hold1432 (.A(_00241_),
    .X(net3811));
 sg13g2_dlygate4sd3_1 hold1433 (.A(_04515_),
    .X(net3812));
 sg13g2_dlygate4sd3_1 hold1434 (.A(_04516_),
    .X(net3813));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\i_time.l_mtimecmp.data_out[14] ),
    .X(net3814));
 sg13g2_dlygate4sd3_1 hold1436 (.A(_01352_),
    .X(net3815));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\i_spi.data[6] ),
    .X(net3816));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\data_to_write[27] ),
    .X(net3817));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .X(net3818));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\i_tinyqv.cpu.instr_data_in[9] ),
    .X(net3819));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .X(net3820));
 sg13g2_dlygate4sd3_1 hold1442 (.A(_04973_),
    .X(net3821));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .X(net3822));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\i_tinyqv.cpu.data_ready_latch ),
    .X(net3823));
 sg13g2_dlygate4sd3_1 hold1445 (.A(_01419_),
    .X(net3824));
 sg13g2_dlygate4sd3_1 hold1446 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .X(net3825));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\i_tinyqv.cpu.instr_data_start[17] ),
    .X(net3826));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\i_debug_uart_tx.fsm_state[1] ),
    .X(net3827));
 sg13g2_dlygate4sd3_1 hold1449 (.A(_00809_),
    .X(net3828));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .X(net3829));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\i_time.l_mtimecmp.data_out[9] ),
    .X(net3830));
 sg13g2_dlygate4sd3_1 hold1452 (.A(_01347_),
    .X(net3831));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .X(net3832));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .X(net3833));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\i_time.l_mtimecmp.data_out[12] ),
    .X(net3834));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\data_to_write[13] ),
    .X(net3835));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\i_tinyqv.cpu.instr_fetch_stopped ),
    .X(net3836));
 sg13g2_dlygate4sd3_1 hold1458 (.A(_05496_),
    .X(net3837));
 sg13g2_dlygate4sd3_1 hold1459 (.A(_05497_),
    .X(net3838));
 sg13g2_dlygate4sd3_1 hold1460 (.A(_01375_),
    .X(net3839));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .X(net3840));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\i_tinyqv.cpu.imm[23] ),
    .X(net3841));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\data_to_write[16] ),
    .X(net3842));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\i_tinyqv.cpu.i_core.i_cycles.cy ),
    .X(net3843));
 sg13g2_dlygate4sd3_1 hold1465 (.A(_04073_),
    .X(net3844));
 sg13g2_dlygate4sd3_1 hold1466 (.A(_00592_),
    .X(net3845));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\i_tinyqv.cpu.data_read_n[0] ),
    .X(net3846));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\i_tinyqv.cpu.i_core.mcause[0] ),
    .X(net3847));
 sg13g2_dlygate4sd3_1 hold1469 (.A(_04115_),
    .X(net3848));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .X(net3849));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .X(net3850));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\i_tinyqv.cpu.instr_data_start[23] ),
    .X(net3851));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\i_debug_uart_tx.fsm_state[0] ),
    .X(net3852));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\i_time.mtime[19] ),
    .X(net3853));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\i_tinyqv.mem.q_ctrl.data_req ),
    .X(net3854));
 sg13g2_dlygate4sd3_1 hold1476 (.A(_00118_),
    .X(net3855));
 sg13g2_dlygate4sd3_1 hold1477 (.A(_00266_),
    .X(net3856));
 sg13g2_dlygate4sd3_1 hold1478 (.A(_01415_),
    .X(net3857));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .X(net3858));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\i_tinyqv.cpu.data_read_n[1] ),
    .X(net3859));
 sg13g2_dlygate4sd3_1 hold1481 (.A(_01412_),
    .X(net3860));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\i_tinyqv.cpu.instr_data_in[10] ),
    .X(net3861));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\i_time.l_mtimecmp.data_out[26] ),
    .X(net3862));
 sg13g2_dlygate4sd3_1 hold1484 (.A(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .X(net3863));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\data_to_write[31] ),
    .X(net3864));
 sg13g2_dlygate4sd3_1 hold1486 (.A(_00805_),
    .X(net3865));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .X(net3866));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\i_spi.bits_remaining[1] ),
    .X(net3867));
 sg13g2_dlygate4sd3_1 hold1489 (.A(_00722_),
    .X(net3868));
 sg13g2_dlygate4sd3_1 hold1490 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .X(net3869));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .X(net3870));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\i_tinyqv.cpu.i_core.mepc[21] ),
    .X(net3871));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\i_uart_rx.cycle_counter[10] ),
    .X(net3872));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\data_to_write[15] ),
    .X(net3873));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .X(net3874));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\i_tinyqv.cpu.instr_data[1][0] ),
    .X(net3875));
 sg13g2_dlygate4sd3_1 hold1497 (.A(_01309_),
    .X(net3876));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\gpio_out_sel[7] ),
    .X(net3877));
 sg13g2_dlygate4sd3_1 hold1499 (.A(_00015_),
    .X(net3878));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .X(net3879));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\i_time.mtime[3] ),
    .X(net3880));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .X(net3881));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\data_to_write[14] ),
    .X(net3882));
 sg13g2_dlygate4sd3_1 hold1504 (.A(_00200_),
    .X(net3883));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[3] ),
    .X(net3884));
 sg13g2_dlygate4sd3_1 hold1506 (.A(_00596_),
    .X(net3885));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\i_tinyqv.cpu.instr_data_in[8] ),
    .X(net3886));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\addr[24] ),
    .X(net3887));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .X(net3888));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\data_to_write[10] ),
    .X(net3889));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\i_tinyqv.cpu.imm[22] ),
    .X(net3890));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\i_tinyqv.cpu.alu_op[0] ),
    .X(net3891));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\i_pwm.pwm_count[7] ),
    .X(net3892));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\i_tinyqv.cpu.mem_op_increment_reg ),
    .X(net3893));
 sg13g2_dlygate4sd3_1 hold1515 (.A(_01482_),
    .X(net3894));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\i_tinyqv.cpu.instr_data_start[4] ),
    .X(net3895));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .X(net3896));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\i_tinyqv.cpu.instr_data[0][0] ),
    .X(net3897));
 sg13g2_dlygate4sd3_1 hold1519 (.A(_01204_),
    .X(net3898));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .X(net3899));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .X(net3900));
 sg13g2_dlygate4sd3_1 hold1522 (.A(_01273_),
    .X(net3901));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .X(net3902));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\i_uart_rx.fsm_state[3] ),
    .X(net3903));
 sg13g2_dlygate4sd3_1 hold1525 (.A(_00678_),
    .X(net3904));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .X(net3905));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .X(net3906));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\i_tinyqv.cpu.i_core.i_cycles.rstn ),
    .X(net3907));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .X(net3908));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\data_to_write[17] ),
    .X(net3909));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .X(net3910));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\data_to_write[11] ),
    .X(net3911));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .X(net3912));
 sg13g2_dlygate4sd3_1 hold1534 (.A(_01177_),
    .X(net3913));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\i_tinyqv.cpu.instr_data_in[0] ),
    .X(net3914));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .X(net3915));
 sg13g2_dlygate4sd3_1 hold1537 (.A(_04079_),
    .X(net3916));
 sg13g2_dlygate4sd3_1 hold1538 (.A(_00194_),
    .X(net3917));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .X(net3918));
 sg13g2_dlygate4sd3_1 hold1540 (.A(_01176_),
    .X(net3919));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\data_to_write[18] ),
    .X(net3920));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\data_to_write[30] ),
    .X(net3921));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .X(net3922));
 sg13g2_dlygate4sd3_1 hold1544 (.A(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .X(net3923));
 sg13g2_dlygate4sd3_1 hold1545 (.A(_01175_),
    .X(net3924));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\i_tinyqv.cpu.i_core.multiplier.accum[8] ),
    .X(net3925));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\data_to_write[24] ),
    .X(net3926));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\i_tinyqv.cpu.instr_data_start[15] ),
    .X(net3927));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\i_time.mtime[30] ),
    .X(net3928));
 sg13g2_dlygate4sd3_1 hold1550 (.A(_04608_),
    .X(net3929));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .X(net3930));
 sg13g2_dlygate4sd3_1 hold1552 (.A(\i_tinyqv.cpu.instr_data_start[18] ),
    .X(net3931));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\i_tinyqv.cpu.is_alu_reg ),
    .X(net3932));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\i_tinyqv.mem.q_ctrl.is_writing ),
    .X(net3933));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .X(net3934));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\i_tinyqv.cpu.instr_data_in[7] ),
    .X(net3935));
 sg13g2_dlygate4sd3_1 hold1557 (.A(_01244_),
    .X(net3936));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\i_tinyqv.cpu.instr_data_in[11] ),
    .X(net3937));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\i_tinyqv.cpu.instr_data_start[12] ),
    .X(net3938));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\i_tinyqv.cpu.imm[20] ),
    .X(net3939));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\i_tinyqv.cpu.instr_data_in[3] ),
    .X(net3940));
 sg13g2_dlygate4sd3_1 hold1562 (.A(\i_tinyqv.cpu.imm[18] ),
    .X(net3941));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .X(net3942));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\i_time.mtime[12] ),
    .X(net3943));
 sg13g2_dlygate4sd3_1 hold1565 (.A(_04554_),
    .X(net3944));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\i_tinyqv.cpu.data_write_n[1] ),
    .X(net3945));
 sg13g2_dlygate4sd3_1 hold1567 (.A(_01058_),
    .X(net3946));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\i_tinyqv.cpu.instr_data_in[6] ),
    .X(net3947));
 sg13g2_dlygate4sd3_1 hold1569 (.A(_01243_),
    .X(net3948));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\i_tinyqv.cpu.is_auipc ),
    .X(net3949));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .X(net3950));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\data_to_write[28] ),
    .X(net3951));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\i_tinyqv.cpu.i_core.i_shift.a[15] ),
    .X(net3952));
 sg13g2_dlygate4sd3_1 hold1574 (.A(_01185_),
    .X(net3953));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\i_time.mtime[13] ),
    .X(net3954));
 sg13g2_dlygate4sd3_1 hold1576 (.A(\i_tinyqv.cpu.imm[12] ),
    .X(net3955));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .X(net3956));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .X(net3957));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .X(net3958));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\i_time.mtime[27] ),
    .X(net3959));
 sg13g2_dlygate4sd3_1 hold1581 (.A(_04599_),
    .X(net3960));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\i_time.mtime[26] ),
    .X(net3961));
 sg13g2_dlygate4sd3_1 hold1583 (.A(_04595_),
    .X(net3962));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\i_tinyqv.cpu.imm[13] ),
    .X(net3963));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .X(net3964));
 sg13g2_dlygate4sd3_1 hold1586 (.A(_01184_),
    .X(net3965));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .X(net3966));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\i_tinyqv.cpu.instr_data_start[6] ),
    .X(net3967));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\i_tinyqv.cpu.i_core.cycle_count[2] ),
    .X(net3968));
 sg13g2_dlygate4sd3_1 hold1590 (.A(_04080_),
    .X(net3969));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .X(net3970));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\data_to_write[25] ),
    .X(net3971));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\i_tinyqv.cpu.is_system ),
    .X(net3972));
 sg13g2_dlygate4sd3_1 hold1594 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[1] ),
    .X(net3973));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\data_to_write[29] ),
    .X(net3974));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\i_tinyqv.cpu.imm[17] ),
    .X(net3975));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\i_time.mtime[11] ),
    .X(net3976));
 sg13g2_dlygate4sd3_1 hold1598 (.A(_04550_),
    .X(net3977));
 sg13g2_dlygate4sd3_1 hold1599 (.A(_00197_),
    .X(net3978));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\i_tinyqv.cpu.instr_data_start[11] ),
    .X(net3979));
 sg13g2_dlygate4sd3_1 hold1601 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .X(net3980));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .X(net3981));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .X(net3982));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\i_uart_tx.fsm_state[1] ),
    .X(net3983));
 sg13g2_dlygate4sd3_1 hold1605 (.A(\i_time.mtime[16] ),
    .X(net3984));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .X(net3985));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\i_tinyqv.cpu.instr_data_start[8] ),
    .X(net3986));
 sg13g2_dlygate4sd3_1 hold1608 (.A(\addr[5] ),
    .X(net3987));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\i_tinyqv.cpu.imm[21] ),
    .X(net3988));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .X(net3989));
 sg13g2_dlygate4sd3_1 hold1611 (.A(uio_out[6]),
    .X(net3990));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\i_tinyqv.cpu.is_lui ),
    .X(net3991));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\i_tinyqv.cpu.imm[19] ),
    .X(net3992));
 sg13g2_dlygate4sd3_1 hold1614 (.A(_01451_),
    .X(net3993));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .X(net3994));
 sg13g2_dlygate4sd3_1 hold1616 (.A(\i_time.mtime[10] ),
    .X(net3995));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .X(net3996));
 sg13g2_dlygate4sd3_1 hold1618 (.A(\i_time.mtime[29] ),
    .X(net3997));
 sg13g2_dlygate4sd3_1 hold1619 (.A(_04604_),
    .X(net3998));
 sg13g2_dlygate4sd3_1 hold1620 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .X(net3999));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\i_uart_tx.fsm_state[2] ),
    .X(net4000));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\i_time.mtime[28] ),
    .X(net4001));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\i_tinyqv.cpu.imm[15] ),
    .X(net4002));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .X(net4003));
 sg13g2_dlygate4sd3_1 hold1625 (.A(\i_tinyqv.cpu.is_alu_imm ),
    .X(net4004));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .X(net4005));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .X(net4006));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .X(net4007));
 sg13g2_dlygate4sd3_1 hold1629 (.A(\i_time.mtime[25] ),
    .X(net4008));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\i_tinyqv.cpu.i_core.mie[2] ),
    .X(net4009));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .X(net4010));
 sg13g2_dlygate4sd3_1 hold1632 (.A(net2380),
    .X(net4011));
 sg13g2_dlygate4sd3_1 hold1633 (.A(\i_time.mtime[15] ),
    .X(net4012));
 sg13g2_dlygate4sd3_1 hold1634 (.A(_04563_),
    .X(net4013));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\i_tinyqv.cpu.instr_data_start[14] ),
    .X(net4014));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\i_time.mtime[7] ),
    .X(net4015));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .X(net4016));
 sg13g2_dlygate4sd3_1 hold1638 (.A(net633),
    .X(net4017));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\i_time.mtime[14] ),
    .X(net4018));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .X(net4019));
 sg13g2_dlygate4sd3_1 hold1641 (.A(_01182_),
    .X(net4020));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .X(net4021));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .X(net4022));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .X(net4023));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\data_to_write[23] ),
    .X(net4024));
 sg13g2_dlygate4sd3_1 hold1646 (.A(_00797_),
    .X(net4025));
 sg13g2_dlygate4sd3_1 hold1647 (.A(\data_to_write[22] ),
    .X(net4026));
 sg13g2_dlygate4sd3_1 hold1648 (.A(_00796_),
    .X(net4027));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[2] ),
    .X(net4028));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\i_time.mtime[24] ),
    .X(net4029));
 sg13g2_dlygate4sd3_1 hold1651 (.A(_04590_),
    .X(net4030));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\i_tinyqv.mem.instr_active ),
    .X(net4031));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .X(net4032));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .X(net4033));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .X(net4034));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .X(net4035));
 sg13g2_dlygate4sd3_1 hold1657 (.A(_01178_),
    .X(net4036));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .X(net4037));
 sg13g2_dlygate4sd3_1 hold1659 (.A(_01183_),
    .X(net4038));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .X(net4039));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\i_tinyqv.cpu.instr_data_in[13] ),
    .X(net4040));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .X(net4041));
 sg13g2_dlygate4sd3_1 hold1663 (.A(_00129_),
    .X(net4042));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\i_tinyqv.cpu.instr_data_start[19] ),
    .X(net4043));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\i_time.mtime[17] ),
    .X(net4044));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\i_tinyqv.cpu.imm[16] ),
    .X(net4045));
 sg13g2_dlygate4sd3_1 hold1667 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .X(net4046));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .X(net4047));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\i_tinyqv.cpu.data_write_n[0] ),
    .X(net4048));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\i_time.mtime[18] ),
    .X(net4049));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\data_to_write[21] ),
    .X(net4050));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\i_uart_rx.fsm_state[1] ),
    .X(net4051));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\i_tinyqv.cpu.pc[1] ),
    .X(net4052));
 sg13g2_dlygate4sd3_1 hold1674 (.A(_00244_),
    .X(net4053));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .X(net4054));
 sg13g2_dlygate4sd3_1 hold1676 (.A(debug_register_data),
    .X(net4055));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .X(net4056));
 sg13g2_dlygate4sd3_1 hold1678 (.A(_00192_),
    .X(net4057));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\i_tinyqv.cpu.instr_data_start[7] ),
    .X(net4058));
 sg13g2_dlygate4sd3_1 hold1680 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .X(net4059));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\i_tinyqv.mem.q_ctrl.last_ram_b_sel ),
    .X(net4060));
 sg13g2_dlygate4sd3_1 hold1682 (.A(\data_to_write[20] ),
    .X(net4061));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\i_uart_tx.fsm_state[0] ),
    .X(net4062));
 sg13g2_dlygate4sd3_1 hold1684 (.A(\i_tinyqv.cpu.imm[14] ),
    .X(net4063));
 sg13g2_dlygate4sd3_1 hold1685 (.A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .X(net4064));
 sg13g2_dlygate4sd3_1 hold1686 (.A(_01179_),
    .X(net4065));
 sg13g2_dlygate4sd3_1 hold1687 (.A(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .X(net4066));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\i_time.mtime[21] ),
    .X(net4067));
 sg13g2_dlygate4sd3_1 hold1689 (.A(_04581_),
    .X(net4068));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .X(net4069));
 sg13g2_dlygate4sd3_1 hold1691 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .X(net4070));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .X(net4071));
 sg13g2_dlygate4sd3_1 hold1693 (.A(_01181_),
    .X(net4072));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .X(net4073));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .X(net4074));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\i_time.mtime[20] ),
    .X(net4075));
 sg13g2_dlygate4sd3_1 hold1697 (.A(_04578_),
    .X(net4076));
 sg13g2_dlygate4sd3_1 hold1698 (.A(\i_tinyqv.cpu.pc[2] ),
    .X(net4077));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .X(net4078));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\i_tinyqv.cpu.instr_data_in[14] ),
    .X(net4079));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\i_time.mtime[8] ),
    .X(net4080));
 sg13g2_dlygate4sd3_1 hold1702 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .X(net4081));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\i_time.mtime[4] ),
    .X(net4082));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\i_time.mtime[0] ),
    .X(net4083));
 sg13g2_dlygate4sd3_1 hold1705 (.A(_04520_),
    .X(net4084));
 sg13g2_dlygate4sd3_1 hold1706 (.A(\i_tinyqv.cpu.instr_data_in[2] ),
    .X(net4085));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .X(net4086));
 sg13g2_dlygate4sd3_1 hold1708 (.A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .X(net4087));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\addr[6] ),
    .X(net4088));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .X(net4089));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .X(net4090));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .X(net4091));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .X(net4092));
 sg13g2_dlygate4sd3_1 hold1714 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .X(net4093));
 sg13g2_dlygate4sd3_1 hold1715 (.A(_00131_),
    .X(net4094));
 sg13g2_dlygate4sd3_1 hold1716 (.A(net640),
    .X(net4095));
 sg13g2_dlygate4sd3_1 hold1717 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .X(net4096));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\i_tinyqv.cpu.is_jalr ),
    .X(net4097));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\i_tinyqv.cpu.was_early_branch ),
    .X(net4098));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\i_pwm.pwm_count[7] ),
    .X(net4099));
 sg13g2_dlygate4sd3_1 hold1721 (.A(\i_tinyqv.cpu.instr_data_in[15] ),
    .X(net4100));
 sg13g2_dlygate4sd3_1 hold1722 (.A(debug_instr_valid),
    .X(net4101));
 sg13g2_dlygate4sd3_1 hold1723 (.A(_01484_),
    .X(net4102));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\i_tinyqv.cpu.alu_op[1] ),
    .X(net4103));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .X(net4104));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\i_tinyqv.cpu.is_branch ),
    .X(net4105));
 sg13g2_dlygate4sd3_1 hold1727 (.A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .X(net4106));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\i_time.mtime[9] ),
    .X(net4107));
 sg13g2_dlygate4sd3_1 hold1729 (.A(_04545_),
    .X(net4108));
 sg13g2_dlygate4sd3_1 hold1730 (.A(_00783_),
    .X(net4109));
 sg13g2_dlygate4sd3_1 hold1731 (.A(\i_tinyqv.cpu.instr_data_start[9] ),
    .X(net4110));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\i_tinyqv.cpu.instr_data_start[3] ),
    .X(net4111));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\addr[3] ),
    .X(net4112));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .X(net4113));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\i_time.mtime[6] ),
    .X(net4114));
 sg13g2_dlygate4sd3_1 hold1736 (.A(\i_time.mtime[5] ),
    .X(net4115));
 sg13g2_dlygate4sd3_1 hold1737 (.A(uio_out[0]),
    .X(net4116));
 sg13g2_dlygate4sd3_1 hold1738 (.A(\i_tinyqv.cpu.alu_op[3] ),
    .X(net4117));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .X(net4118));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\i_time.mtime[2] ),
    .X(net4119));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\data_to_write[9] ),
    .X(net4120));
 sg13g2_dlygate4sd3_1 hold1742 (.A(\i_tinyqv.cpu.instr_data_start[10] ),
    .X(net4121));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .X(net4122));
 sg13g2_dlygate4sd3_1 hold1744 (.A(\i_tinyqv.cpu.instr_data_start[20] ),
    .X(net4123));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\data_to_write[1] ),
    .X(net4124));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .X(net4125));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\data_to_write[2] ),
    .X(net4126));
 sg13g2_dlygate4sd3_1 hold1748 (.A(\i_tinyqv.cpu.alu_op[2] ),
    .X(net4127));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .X(net4128));
 sg13g2_dlygate4sd3_1 hold1750 (.A(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .X(net4129));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\i_tinyqv.cpu.i_core.multiplier.accum[15] ),
    .X(net4130));
 sg13g2_dlygate4sd3_1 hold1752 (.A(_00195_),
    .X(net4131));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\i_uart_tx.fsm_state[0] ),
    .X(net4132));
 sg13g2_dlygate4sd3_1 hold1754 (.A(_00129_),
    .X(net4133));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .X(net4134));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\i_uart_tx.fsm_state[0] ),
    .X(net4135));
 sg13g2_antennanp ANTENNA_1 (.A(_00063_));
 sg13g2_antennanp ANTENNA_2 (.A(\debug_rd[1] ));
 sg13g2_antennanp ANTENNA_3 (.A(\debug_rd[1] ));
 sg13g2_antennanp ANTENNA_4 (.A(\debug_rd[1] ));
 sg13g2_antennanp ANTENNA_5 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_antennanp ANTENNA_6 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ));
 sg13g2_antennanp ANTENNA_7 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_antennanp ANTENNA_8 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ));
 sg13g2_antennanp ANTENNA_9 (.A(uio_out[6]));
 sg13g2_antennanp ANTENNA_10 (.A(uio_out[6]));
 sg13g2_antennanp ANTENNA_11 (.A(_00063_));
 sg13g2_antennanp ANTENNA_12 (.A(\debug_rd[0] ));
 sg13g2_antennanp ANTENNA_13 (.A(\debug_rd[0] ));
 sg13g2_antennanp ANTENNA_14 (.A(\debug_rd[0] ));
 sg13g2_antennanp ANTENNA_15 (.A(uio_out[6]));
 sg13g2_antennanp ANTENNA_16 (.A(uio_out[6]));
 sg13g2_antennanp ANTENNA_17 (.A(\debug_rd[0] ));
 sg13g2_antennanp ANTENNA_18 (.A(\debug_rd[0] ));
 sg13g2_antennanp ANTENNA_19 (.A(\debug_rd[0] ));
 sg13g2_antennanp ANTENNA_20 (.A(uio_out[6]));
 sg13g2_antennanp ANTENNA_21 (.A(uio_out[6]));
 sg13g2_antennanp ANTENNA_22 (.A(net2836));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_fill_2 FILLER_0_14 ();
 sg13g2_fill_2 FILLER_0_45 ();
 sg13g2_fill_2 FILLER_0_51 ();
 sg13g2_decap_8 FILLER_0_58 ();
 sg13g2_fill_1 FILLER_0_65 ();
 sg13g2_decap_4 FILLER_0_95 ();
 sg13g2_decap_8 FILLER_0_102 ();
 sg13g2_decap_4 FILLER_0_114 ();
 sg13g2_fill_2 FILLER_0_118 ();
 sg13g2_fill_1 FILLER_0_128 ();
 sg13g2_fill_2 FILLER_0_134 ();
 sg13g2_fill_1 FILLER_0_136 ();
 sg13g2_decap_8 FILLER_0_149 ();
 sg13g2_decap_8 FILLER_0_160 ();
 sg13g2_decap_4 FILLER_0_167 ();
 sg13g2_fill_1 FILLER_0_171 ();
 sg13g2_fill_2 FILLER_0_205 ();
 sg13g2_fill_1 FILLER_0_245 ();
 sg13g2_fill_1 FILLER_0_268 ();
 sg13g2_fill_1 FILLER_0_273 ();
 sg13g2_fill_1 FILLER_0_381 ();
 sg13g2_fill_1 FILLER_0_414 ();
 sg13g2_fill_1 FILLER_0_452 ();
 sg13g2_fill_1 FILLER_0_529 ();
 sg13g2_fill_1 FILLER_0_571 ();
 sg13g2_fill_1 FILLER_0_638 ();
 sg13g2_fill_1 FILLER_0_665 ();
 sg13g2_fill_2 FILLER_0_733 ();
 sg13g2_fill_1 FILLER_0_735 ();
 sg13g2_fill_2 FILLER_0_766 ();
 sg13g2_fill_1 FILLER_0_768 ();
 sg13g2_fill_1 FILLER_0_808 ();
 sg13g2_fill_1 FILLER_0_826 ();
 sg13g2_fill_2 FILLER_0_866 ();
 sg13g2_fill_1 FILLER_0_868 ();
 sg13g2_fill_1 FILLER_0_925 ();
 sg13g2_fill_2 FILLER_0_961 ();
 sg13g2_fill_1 FILLER_0_963 ();
 sg13g2_fill_2 FILLER_0_1046 ();
 sg13g2_fill_1 FILLER_0_1048 ();
 sg13g2_fill_2 FILLER_0_1163 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_1 FILLER_1_36 ();
 sg13g2_fill_2 FILLER_1_67 ();
 sg13g2_fill_2 FILLER_1_78 ();
 sg13g2_fill_1 FILLER_1_84 ();
 sg13g2_fill_1 FILLER_1_159 ();
 sg13g2_fill_1 FILLER_1_217 ();
 sg13g2_fill_2 FILLER_1_371 ();
 sg13g2_fill_1 FILLER_1_544 ();
 sg13g2_fill_1 FILLER_1_610 ();
 sg13g2_fill_2 FILLER_1_709 ();
 sg13g2_fill_2 FILLER_1_747 ();
 sg13g2_fill_2 FILLER_1_784 ();
 sg13g2_fill_1 FILLER_1_786 ();
 sg13g2_fill_2 FILLER_1_887 ();
 sg13g2_fill_2 FILLER_1_937 ();
 sg13g2_fill_1 FILLER_1_939 ();
 sg13g2_fill_2 FILLER_1_984 ();
 sg13g2_fill_2 FILLER_1_1073 ();
 sg13g2_fill_2 FILLER_1_1180 ();
 sg13g2_fill_1 FILLER_1_1182 ();
 sg13g2_fill_2 FILLER_1_1265 ();
 sg13g2_fill_2 FILLER_1_1300 ();
 sg13g2_fill_1 FILLER_1_1314 ();
 sg13g2_fill_2 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_28 ();
 sg13g2_fill_2 FILLER_2_38 ();
 sg13g2_fill_1 FILLER_2_48 ();
 sg13g2_decap_8 FILLER_2_75 ();
 sg13g2_fill_1 FILLER_2_82 ();
 sg13g2_fill_1 FILLER_2_120 ();
 sg13g2_fill_2 FILLER_2_134 ();
 sg13g2_fill_2 FILLER_2_188 ();
 sg13g2_fill_2 FILLER_2_213 ();
 sg13g2_fill_1 FILLER_2_224 ();
 sg13g2_fill_2 FILLER_2_229 ();
 sg13g2_fill_2 FILLER_2_250 ();
 sg13g2_fill_1 FILLER_2_282 ();
 sg13g2_fill_1 FILLER_2_288 ();
 sg13g2_fill_1 FILLER_2_308 ();
 sg13g2_fill_2 FILLER_2_349 ();
 sg13g2_fill_1 FILLER_2_382 ();
 sg13g2_fill_2 FILLER_2_391 ();
 sg13g2_fill_2 FILLER_2_412 ();
 sg13g2_fill_2 FILLER_2_478 ();
 sg13g2_fill_2 FILLER_2_682 ();
 sg13g2_fill_2 FILLER_2_787 ();
 sg13g2_fill_1 FILLER_2_789 ();
 sg13g2_fill_2 FILLER_2_825 ();
 sg13g2_fill_1 FILLER_2_827 ();
 sg13g2_fill_2 FILLER_2_1008 ();
 sg13g2_fill_1 FILLER_2_1010 ();
 sg13g2_fill_2 FILLER_2_1094 ();
 sg13g2_fill_1 FILLER_2_1096 ();
 sg13g2_fill_2 FILLER_2_1127 ();
 sg13g2_fill_1 FILLER_2_1182 ();
 sg13g2_fill_1 FILLER_2_1196 ();
 sg13g2_fill_2 FILLER_2_1227 ();
 sg13g2_fill_2 FILLER_2_1297 ();
 sg13g2_fill_1 FILLER_2_1299 ();
 sg13g2_fill_1 FILLER_2_1308 ();
 sg13g2_fill_2 FILLER_2_1313 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_10 ();
 sg13g2_fill_1 FILLER_3_12 ();
 sg13g2_fill_2 FILLER_3_21 ();
 sg13g2_fill_1 FILLER_3_86 ();
 sg13g2_fill_1 FILLER_3_94 ();
 sg13g2_fill_1 FILLER_3_150 ();
 sg13g2_fill_1 FILLER_3_214 ();
 sg13g2_fill_1 FILLER_3_294 ();
 sg13g2_fill_1 FILLER_3_372 ();
 sg13g2_fill_1 FILLER_3_436 ();
 sg13g2_fill_2 FILLER_3_497 ();
 sg13g2_fill_2 FILLER_3_555 ();
 sg13g2_fill_1 FILLER_3_572 ();
 sg13g2_fill_1 FILLER_3_578 ();
 sg13g2_fill_2 FILLER_3_633 ();
 sg13g2_fill_2 FILLER_3_680 ();
 sg13g2_fill_1 FILLER_3_718 ();
 sg13g2_fill_1 FILLER_3_755 ();
 sg13g2_fill_1 FILLER_3_847 ();
 sg13g2_fill_1 FILLER_3_874 ();
 sg13g2_fill_2 FILLER_3_883 ();
 sg13g2_fill_2 FILLER_3_911 ();
 sg13g2_fill_2 FILLER_3_949 ();
 sg13g2_fill_1 FILLER_3_951 ();
 sg13g2_fill_1 FILLER_3_965 ();
 sg13g2_fill_2 FILLER_3_992 ();
 sg13g2_fill_1 FILLER_3_994 ();
 sg13g2_fill_1 FILLER_3_1004 ();
 sg13g2_fill_2 FILLER_3_1075 ();
 sg13g2_fill_1 FILLER_3_1086 ();
 sg13g2_fill_2 FILLER_3_1100 ();
 sg13g2_fill_1 FILLER_3_1102 ();
 sg13g2_fill_2 FILLER_3_1155 ();
 sg13g2_fill_1 FILLER_3_1214 ();
 sg13g2_fill_2 FILLER_3_1237 ();
 sg13g2_fill_1 FILLER_3_1239 ();
 sg13g2_fill_2 FILLER_3_1297 ();
 sg13g2_fill_2 FILLER_3_1312 ();
 sg13g2_fill_1 FILLER_3_1314 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_45 ();
 sg13g2_decap_4 FILLER_4_183 ();
 sg13g2_fill_2 FILLER_4_187 ();
 sg13g2_fill_2 FILLER_4_224 ();
 sg13g2_fill_2 FILLER_4_229 ();
 sg13g2_fill_2 FILLER_4_235 ();
 sg13g2_fill_1 FILLER_4_312 ();
 sg13g2_fill_1 FILLER_4_367 ();
 sg13g2_fill_2 FILLER_4_421 ();
 sg13g2_fill_1 FILLER_4_437 ();
 sg13g2_fill_1 FILLER_4_500 ();
 sg13g2_fill_2 FILLER_4_546 ();
 sg13g2_fill_2 FILLER_4_663 ();
 sg13g2_fill_2 FILLER_4_734 ();
 sg13g2_fill_1 FILLER_4_783 ();
 sg13g2_decap_8 FILLER_4_788 ();
 sg13g2_decap_4 FILLER_4_795 ();
 sg13g2_fill_1 FILLER_4_812 ();
 sg13g2_fill_1 FILLER_4_905 ();
 sg13g2_fill_1 FILLER_4_925 ();
 sg13g2_fill_1 FILLER_4_987 ();
 sg13g2_fill_1 FILLER_4_997 ();
 sg13g2_fill_2 FILLER_4_1020 ();
 sg13g2_fill_1 FILLER_4_1022 ();
 sg13g2_fill_2 FILLER_4_1058 ();
 sg13g2_fill_1 FILLER_4_1060 ();
 sg13g2_fill_1 FILLER_4_1122 ();
 sg13g2_fill_2 FILLER_4_1171 ();
 sg13g2_fill_1 FILLER_4_1173 ();
 sg13g2_fill_1 FILLER_4_1200 ();
 sg13g2_fill_2 FILLER_4_1266 ();
 sg13g2_fill_2 FILLER_4_1303 ();
 sg13g2_fill_1 FILLER_4_1305 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_2 ();
 sg13g2_fill_1 FILLER_5_19 ();
 sg13g2_fill_2 FILLER_5_97 ();
 sg13g2_fill_2 FILLER_5_131 ();
 sg13g2_fill_2 FILLER_5_149 ();
 sg13g2_fill_2 FILLER_5_162 ();
 sg13g2_fill_1 FILLER_5_182 ();
 sg13g2_decap_4 FILLER_5_191 ();
 sg13g2_fill_1 FILLER_5_225 ();
 sg13g2_fill_1 FILLER_5_261 ();
 sg13g2_fill_1 FILLER_5_286 ();
 sg13g2_fill_1 FILLER_5_296 ();
 sg13g2_fill_1 FILLER_5_305 ();
 sg13g2_fill_1 FILLER_5_310 ();
 sg13g2_fill_2 FILLER_5_349 ();
 sg13g2_fill_2 FILLER_5_412 ();
 sg13g2_fill_2 FILLER_5_449 ();
 sg13g2_fill_1 FILLER_5_472 ();
 sg13g2_fill_1 FILLER_5_526 ();
 sg13g2_fill_2 FILLER_5_596 ();
 sg13g2_fill_2 FILLER_5_616 ();
 sg13g2_fill_1 FILLER_5_618 ();
 sg13g2_fill_1 FILLER_5_650 ();
 sg13g2_fill_2 FILLER_5_677 ();
 sg13g2_fill_2 FILLER_5_689 ();
 sg13g2_fill_1 FILLER_5_691 ();
 sg13g2_fill_2 FILLER_5_773 ();
 sg13g2_fill_1 FILLER_5_775 ();
 sg13g2_fill_2 FILLER_5_796 ();
 sg13g2_fill_2 FILLER_5_808 ();
 sg13g2_fill_1 FILLER_5_810 ();
 sg13g2_decap_4 FILLER_5_815 ();
 sg13g2_fill_1 FILLER_5_819 ();
 sg13g2_fill_1 FILLER_5_841 ();
 sg13g2_fill_2 FILLER_5_848 ();
 sg13g2_fill_1 FILLER_5_850 ();
 sg13g2_fill_2 FILLER_5_899 ();
 sg13g2_fill_2 FILLER_5_942 ();
 sg13g2_fill_1 FILLER_5_944 ();
 sg13g2_fill_2 FILLER_5_959 ();
 sg13g2_fill_1 FILLER_5_961 ();
 sg13g2_fill_2 FILLER_5_1040 ();
 sg13g2_fill_1 FILLER_5_1042 ();
 sg13g2_fill_2 FILLER_5_1099 ();
 sg13g2_fill_1 FILLER_5_1101 ();
 sg13g2_fill_1 FILLER_5_1132 ();
 sg13g2_fill_1 FILLER_5_1247 ();
 sg13g2_fill_2 FILLER_5_1287 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_27 ();
 sg13g2_fill_1 FILLER_6_82 ();
 sg13g2_fill_2 FILLER_6_170 ();
 sg13g2_fill_1 FILLER_6_237 ();
 sg13g2_fill_2 FILLER_6_246 ();
 sg13g2_fill_1 FILLER_6_248 ();
 sg13g2_fill_2 FILLER_6_368 ();
 sg13g2_fill_2 FILLER_6_391 ();
 sg13g2_fill_2 FILLER_6_424 ();
 sg13g2_fill_1 FILLER_6_472 ();
 sg13g2_fill_2 FILLER_6_499 ();
 sg13g2_fill_1 FILLER_6_525 ();
 sg13g2_fill_2 FILLER_6_562 ();
 sg13g2_fill_2 FILLER_6_585 ();
 sg13g2_fill_1 FILLER_6_597 ();
 sg13g2_fill_2 FILLER_6_628 ();
 sg13g2_fill_1 FILLER_6_650 ();
 sg13g2_fill_2 FILLER_6_660 ();
 sg13g2_fill_2 FILLER_6_670 ();
 sg13g2_fill_1 FILLER_6_728 ();
 sg13g2_fill_2 FILLER_6_754 ();
 sg13g2_fill_1 FILLER_6_756 ();
 sg13g2_fill_1 FILLER_6_809 ();
 sg13g2_fill_1 FILLER_6_826 ();
 sg13g2_fill_2 FILLER_6_846 ();
 sg13g2_fill_1 FILLER_6_890 ();
 sg13g2_fill_2 FILLER_6_1006 ();
 sg13g2_fill_2 FILLER_6_1061 ();
 sg13g2_fill_2 FILLER_6_1085 ();
 sg13g2_fill_2 FILLER_6_1147 ();
 sg13g2_fill_2 FILLER_6_1175 ();
 sg13g2_fill_1 FILLER_6_1177 ();
 sg13g2_fill_1 FILLER_6_1205 ();
 sg13g2_fill_1 FILLER_6_1267 ();
 sg13g2_fill_2 FILLER_6_1303 ();
 sg13g2_fill_1 FILLER_6_1305 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_10 ();
 sg13g2_fill_1 FILLER_7_12 ();
 sg13g2_decap_4 FILLER_7_17 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_fill_1 FILLER_7_134 ();
 sg13g2_fill_2 FILLER_7_148 ();
 sg13g2_fill_1 FILLER_7_175 ();
 sg13g2_fill_1 FILLER_7_202 ();
 sg13g2_fill_2 FILLER_7_265 ();
 sg13g2_fill_2 FILLER_7_374 ();
 sg13g2_fill_1 FILLER_7_398 ();
 sg13g2_fill_1 FILLER_7_425 ();
 sg13g2_fill_2 FILLER_7_440 ();
 sg13g2_fill_2 FILLER_7_617 ();
 sg13g2_fill_1 FILLER_7_619 ();
 sg13g2_fill_2 FILLER_7_629 ();
 sg13g2_fill_2 FILLER_7_647 ();
 sg13g2_fill_1 FILLER_7_649 ();
 sg13g2_decap_4 FILLER_7_673 ();
 sg13g2_fill_2 FILLER_7_677 ();
 sg13g2_decap_4 FILLER_7_696 ();
 sg13g2_fill_2 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_746 ();
 sg13g2_decap_8 FILLER_7_753 ();
 sg13g2_fill_2 FILLER_7_760 ();
 sg13g2_decap_4 FILLER_7_775 ();
 sg13g2_fill_1 FILLER_7_779 ();
 sg13g2_fill_1 FILLER_7_785 ();
 sg13g2_decap_4 FILLER_7_790 ();
 sg13g2_decap_4 FILLER_7_809 ();
 sg13g2_fill_2 FILLER_7_813 ();
 sg13g2_fill_2 FILLER_7_820 ();
 sg13g2_decap_8 FILLER_7_831 ();
 sg13g2_fill_2 FILLER_7_838 ();
 sg13g2_fill_1 FILLER_7_840 ();
 sg13g2_decap_4 FILLER_7_854 ();
 sg13g2_fill_2 FILLER_7_865 ();
 sg13g2_fill_1 FILLER_7_1033 ();
 sg13g2_fill_2 FILLER_7_1064 ();
 sg13g2_fill_1 FILLER_7_1066 ();
 sg13g2_fill_1 FILLER_7_1101 ();
 sg13g2_fill_1 FILLER_7_1111 ();
 sg13g2_fill_2 FILLER_7_1121 ();
 sg13g2_fill_1 FILLER_7_1123 ();
 sg13g2_fill_2 FILLER_7_1287 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_85 ();
 sg13g2_fill_2 FILLER_8_95 ();
 sg13g2_fill_2 FILLER_8_106 ();
 sg13g2_decap_4 FILLER_8_148 ();
 sg13g2_fill_1 FILLER_8_152 ();
 sg13g2_fill_2 FILLER_8_159 ();
 sg13g2_fill_1 FILLER_8_196 ();
 sg13g2_fill_1 FILLER_8_253 ();
 sg13g2_fill_2 FILLER_8_294 ();
 sg13g2_fill_2 FILLER_8_335 ();
 sg13g2_fill_1 FILLER_8_354 ();
 sg13g2_fill_2 FILLER_8_412 ();
 sg13g2_fill_1 FILLER_8_440 ();
 sg13g2_fill_1 FILLER_8_477 ();
 sg13g2_fill_1 FILLER_8_500 ();
 sg13g2_fill_2 FILLER_8_520 ();
 sg13g2_fill_2 FILLER_8_558 ();
 sg13g2_fill_2 FILLER_8_565 ();
 sg13g2_fill_1 FILLER_8_567 ();
 sg13g2_fill_2 FILLER_8_580 ();
 sg13g2_fill_1 FILLER_8_582 ();
 sg13g2_fill_1 FILLER_8_592 ();
 sg13g2_fill_2 FILLER_8_611 ();
 sg13g2_fill_1 FILLER_8_647 ();
 sg13g2_fill_2 FILLER_8_678 ();
 sg13g2_fill_1 FILLER_8_680 ();
 sg13g2_fill_2 FILLER_8_698 ();
 sg13g2_fill_2 FILLER_8_704 ();
 sg13g2_fill_1 FILLER_8_711 ();
 sg13g2_fill_1 FILLER_8_722 ();
 sg13g2_decap_8 FILLER_8_727 ();
 sg13g2_decap_8 FILLER_8_734 ();
 sg13g2_decap_8 FILLER_8_741 ();
 sg13g2_decap_4 FILLER_8_748 ();
 sg13g2_fill_1 FILLER_8_752 ();
 sg13g2_fill_2 FILLER_8_761 ();
 sg13g2_fill_2 FILLER_8_805 ();
 sg13g2_fill_1 FILLER_8_807 ();
 sg13g2_fill_2 FILLER_8_831 ();
 sg13g2_fill_1 FILLER_8_876 ();
 sg13g2_fill_2 FILLER_8_1039 ();
 sg13g2_fill_1 FILLER_8_1041 ();
 sg13g2_fill_1 FILLER_8_1156 ();
 sg13g2_fill_2 FILLER_8_1275 ();
 sg13g2_fill_2 FILLER_8_1312 ();
 sg13g2_fill_1 FILLER_8_1314 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_2 ();
 sg13g2_fill_1 FILLER_9_46 ();
 sg13g2_fill_1 FILLER_9_56 ();
 sg13g2_decap_4 FILLER_9_160 ();
 sg13g2_decap_8 FILLER_9_178 ();
 sg13g2_decap_4 FILLER_9_185 ();
 sg13g2_fill_2 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_200 ();
 sg13g2_fill_2 FILLER_9_233 ();
 sg13g2_fill_1 FILLER_9_249 ();
 sg13g2_fill_2 FILLER_9_272 ();
 sg13g2_fill_1 FILLER_9_320 ();
 sg13g2_fill_2 FILLER_9_437 ();
 sg13g2_fill_1 FILLER_9_474 ();
 sg13g2_fill_2 FILLER_9_628 ();
 sg13g2_decap_8 FILLER_9_640 ();
 sg13g2_decap_8 FILLER_9_647 ();
 sg13g2_fill_1 FILLER_9_654 ();
 sg13g2_decap_4 FILLER_9_721 ();
 sg13g2_fill_2 FILLER_9_740 ();
 sg13g2_fill_1 FILLER_9_780 ();
 sg13g2_decap_4 FILLER_9_784 ();
 sg13g2_fill_2 FILLER_9_850 ();
 sg13g2_fill_1 FILLER_9_852 ();
 sg13g2_decap_8 FILLER_9_860 ();
 sg13g2_fill_2 FILLER_9_867 ();
 sg13g2_fill_2 FILLER_9_993 ();
 sg13g2_fill_2 FILLER_9_1008 ();
 sg13g2_fill_1 FILLER_9_1010 ();
 sg13g2_fill_2 FILLER_9_1068 ();
 sg13g2_fill_1 FILLER_9_1070 ();
 sg13g2_fill_2 FILLER_9_1167 ();
 sg13g2_fill_2 FILLER_9_1187 ();
 sg13g2_fill_1 FILLER_9_1189 ();
 sg13g2_fill_2 FILLER_9_1208 ();
 sg13g2_fill_1 FILLER_9_1210 ();
 sg13g2_fill_2 FILLER_9_1286 ();
 sg13g2_fill_1 FILLER_9_1288 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_11 ();
 sg13g2_fill_1 FILLER_10_13 ();
 sg13g2_fill_2 FILLER_10_18 ();
 sg13g2_fill_2 FILLER_10_147 ();
 sg13g2_fill_1 FILLER_10_177 ();
 sg13g2_decap_4 FILLER_10_192 ();
 sg13g2_fill_2 FILLER_10_196 ();
 sg13g2_fill_1 FILLER_10_331 ();
 sg13g2_fill_2 FILLER_10_359 ();
 sg13g2_fill_2 FILLER_10_410 ();
 sg13g2_fill_1 FILLER_10_465 ();
 sg13g2_fill_1 FILLER_10_497 ();
 sg13g2_fill_2 FILLER_10_568 ();
 sg13g2_fill_1 FILLER_10_570 ();
 sg13g2_fill_2 FILLER_10_580 ();
 sg13g2_fill_1 FILLER_10_582 ();
 sg13g2_decap_4 FILLER_10_651 ();
 sg13g2_fill_1 FILLER_10_655 ();
 sg13g2_fill_1 FILLER_10_682 ();
 sg13g2_fill_1 FILLER_10_705 ();
 sg13g2_fill_2 FILLER_10_716 ();
 sg13g2_fill_1 FILLER_10_718 ();
 sg13g2_decap_4 FILLER_10_723 ();
 sg13g2_fill_2 FILLER_10_743 ();
 sg13g2_fill_1 FILLER_10_745 ();
 sg13g2_fill_2 FILLER_10_751 ();
 sg13g2_fill_1 FILLER_10_753 ();
 sg13g2_fill_2 FILLER_10_762 ();
 sg13g2_fill_1 FILLER_10_764 ();
 sg13g2_decap_8 FILLER_10_788 ();
 sg13g2_decap_4 FILLER_10_795 ();
 sg13g2_fill_2 FILLER_10_814 ();
 sg13g2_fill_1 FILLER_10_827 ();
 sg13g2_fill_1 FILLER_10_837 ();
 sg13g2_decap_4 FILLER_10_862 ();
 sg13g2_fill_2 FILLER_10_955 ();
 sg13g2_fill_1 FILLER_10_957 ();
 sg13g2_fill_2 FILLER_10_989 ();
 sg13g2_fill_2 FILLER_10_1130 ();
 sg13g2_fill_1 FILLER_10_1142 ();
 sg13g2_fill_2 FILLER_10_1230 ();
 sg13g2_fill_1 FILLER_10_1314 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_2 ();
 sg13g2_fill_1 FILLER_11_29 ();
 sg13g2_fill_1 FILLER_11_44 ();
 sg13g2_decap_8 FILLER_11_53 ();
 sg13g2_decap_8 FILLER_11_60 ();
 sg13g2_decap_4 FILLER_11_67 ();
 sg13g2_fill_2 FILLER_11_71 ();
 sg13g2_fill_2 FILLER_11_78 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_fill_2 FILLER_11_213 ();
 sg13g2_fill_1 FILLER_11_223 ();
 sg13g2_fill_2 FILLER_11_232 ();
 sg13g2_fill_1 FILLER_11_249 ();
 sg13g2_fill_1 FILLER_11_267 ();
 sg13g2_fill_1 FILLER_11_303 ();
 sg13g2_fill_1 FILLER_11_319 ();
 sg13g2_fill_2 FILLER_11_362 ();
 sg13g2_fill_2 FILLER_11_385 ();
 sg13g2_fill_1 FILLER_11_395 ();
 sg13g2_fill_2 FILLER_11_594 ();
 sg13g2_fill_1 FILLER_11_596 ();
 sg13g2_fill_1 FILLER_11_606 ();
 sg13g2_decap_8 FILLER_11_649 ();
 sg13g2_decap_4 FILLER_11_656 ();
 sg13g2_decap_8 FILLER_11_664 ();
 sg13g2_fill_1 FILLER_11_671 ();
 sg13g2_fill_2 FILLER_11_681 ();
 sg13g2_fill_2 FILLER_11_729 ();
 sg13g2_fill_2 FILLER_11_746 ();
 sg13g2_fill_1 FILLER_11_748 ();
 sg13g2_fill_2 FILLER_11_754 ();
 sg13g2_fill_1 FILLER_11_756 ();
 sg13g2_fill_2 FILLER_11_767 ();
 sg13g2_fill_2 FILLER_11_775 ();
 sg13g2_fill_1 FILLER_11_777 ();
 sg13g2_decap_4 FILLER_11_794 ();
 sg13g2_fill_1 FILLER_11_807 ();
 sg13g2_decap_8 FILLER_11_814 ();
 sg13g2_fill_2 FILLER_11_821 ();
 sg13g2_fill_2 FILLER_11_827 ();
 sg13g2_fill_1 FILLER_11_829 ();
 sg13g2_fill_1 FILLER_11_854 ();
 sg13g2_decap_4 FILLER_11_865 ();
 sg13g2_fill_2 FILLER_11_895 ();
 sg13g2_fill_1 FILLER_11_916 ();
 sg13g2_fill_2 FILLER_11_984 ();
 sg13g2_fill_1 FILLER_11_1012 ();
 sg13g2_fill_1 FILLER_11_1069 ();
 sg13g2_fill_2 FILLER_11_1084 ();
 sg13g2_fill_1 FILLER_11_1178 ();
 sg13g2_fill_2 FILLER_11_1188 ();
 sg13g2_fill_1 FILLER_11_1190 ();
 sg13g2_fill_1 FILLER_11_1204 ();
 sg13g2_fill_1 FILLER_11_1240 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_11 ();
 sg13g2_fill_1 FILLER_12_23 ();
 sg13g2_fill_1 FILLER_12_67 ();
 sg13g2_fill_1 FILLER_12_98 ();
 sg13g2_fill_2 FILLER_12_103 ();
 sg13g2_decap_8 FILLER_12_128 ();
 sg13g2_fill_2 FILLER_12_139 ();
 sg13g2_fill_2 FILLER_12_147 ();
 sg13g2_fill_1 FILLER_12_149 ();
 sg13g2_fill_1 FILLER_12_156 ();
 sg13g2_fill_1 FILLER_12_163 ();
 sg13g2_fill_1 FILLER_12_168 ();
 sg13g2_fill_2 FILLER_12_182 ();
 sg13g2_fill_2 FILLER_12_254 ();
 sg13g2_fill_1 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_262 ();
 sg13g2_decap_4 FILLER_12_269 ();
 sg13g2_fill_2 FILLER_12_276 ();
 sg13g2_fill_1 FILLER_12_278 ();
 sg13g2_decap_8 FILLER_12_283 ();
 sg13g2_fill_2 FILLER_12_290 ();
 sg13g2_fill_2 FILLER_12_317 ();
 sg13g2_fill_1 FILLER_12_417 ();
 sg13g2_fill_1 FILLER_12_431 ();
 sg13g2_fill_2 FILLER_12_504 ();
 sg13g2_fill_2 FILLER_12_562 ();
 sg13g2_fill_1 FILLER_12_564 ();
 sg13g2_fill_2 FILLER_12_701 ();
 sg13g2_fill_1 FILLER_12_726 ();
 sg13g2_fill_2 FILLER_12_749 ();
 sg13g2_fill_2 FILLER_12_762 ();
 sg13g2_fill_1 FILLER_12_764 ();
 sg13g2_fill_1 FILLER_12_824 ();
 sg13g2_fill_2 FILLER_12_830 ();
 sg13g2_decap_4 FILLER_12_845 ();
 sg13g2_fill_2 FILLER_12_849 ();
 sg13g2_fill_1 FILLER_12_877 ();
 sg13g2_fill_2 FILLER_12_888 ();
 sg13g2_fill_2 FILLER_12_895 ();
 sg13g2_fill_2 FILLER_12_932 ();
 sg13g2_fill_1 FILLER_12_957 ();
 sg13g2_fill_1 FILLER_12_1031 ();
 sg13g2_fill_2 FILLER_12_1076 ();
 sg13g2_fill_1 FILLER_12_1122 ();
 sg13g2_fill_2 FILLER_12_1150 ();
 sg13g2_fill_1 FILLER_12_1152 ();
 sg13g2_fill_1 FILLER_12_1266 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_49 ();
 sg13g2_fill_1 FILLER_13_51 ();
 sg13g2_fill_1 FILLER_13_87 ();
 sg13g2_fill_2 FILLER_13_114 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_fill_1 FILLER_13_219 ();
 sg13g2_fill_2 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_248 ();
 sg13g2_fill_2 FILLER_13_314 ();
 sg13g2_fill_1 FILLER_13_320 ();
 sg13g2_fill_1 FILLER_13_330 ();
 sg13g2_fill_1 FILLER_13_529 ();
 sg13g2_fill_1 FILLER_13_681 ();
 sg13g2_fill_2 FILLER_13_773 ();
 sg13g2_fill_1 FILLER_13_775 ();
 sg13g2_fill_1 FILLER_13_780 ();
 sg13g2_decap_8 FILLER_13_790 ();
 sg13g2_fill_2 FILLER_13_797 ();
 sg13g2_decap_8 FILLER_13_817 ();
 sg13g2_decap_8 FILLER_13_824 ();
 sg13g2_fill_2 FILLER_13_831 ();
 sg13g2_fill_2 FILLER_13_842 ();
 sg13g2_fill_1 FILLER_13_848 ();
 sg13g2_fill_2 FILLER_13_869 ();
 sg13g2_fill_2 FILLER_13_906 ();
 sg13g2_fill_2 FILLER_13_956 ();
 sg13g2_fill_1 FILLER_13_967 ();
 sg13g2_fill_1 FILLER_13_1056 ();
 sg13g2_fill_1 FILLER_13_1187 ();
 sg13g2_fill_2 FILLER_13_1205 ();
 sg13g2_fill_1 FILLER_13_1207 ();
 sg13g2_fill_2 FILLER_13_1212 ();
 sg13g2_fill_2 FILLER_13_1223 ();
 sg13g2_fill_2 FILLER_13_1287 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_30 ();
 sg13g2_decap_4 FILLER_14_61 ();
 sg13g2_fill_2 FILLER_14_65 ();
 sg13g2_fill_1 FILLER_14_73 ();
 sg13g2_fill_2 FILLER_14_79 ();
 sg13g2_decap_4 FILLER_14_84 ();
 sg13g2_fill_2 FILLER_14_104 ();
 sg13g2_fill_2 FILLER_14_141 ();
 sg13g2_fill_1 FILLER_14_191 ();
 sg13g2_fill_2 FILLER_14_196 ();
 sg13g2_fill_2 FILLER_14_201 ();
 sg13g2_fill_1 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_fill_1 FILLER_14_227 ();
 sg13g2_fill_2 FILLER_14_242 ();
 sg13g2_fill_1 FILLER_14_304 ();
 sg13g2_fill_1 FILLER_14_350 ();
 sg13g2_fill_1 FILLER_14_416 ();
 sg13g2_fill_1 FILLER_14_452 ();
 sg13g2_fill_1 FILLER_14_467 ();
 sg13g2_fill_1 FILLER_14_620 ();
 sg13g2_fill_2 FILLER_14_626 ();
 sg13g2_fill_1 FILLER_14_628 ();
 sg13g2_fill_2 FILLER_14_648 ();
 sg13g2_fill_2 FILLER_14_694 ();
 sg13g2_fill_1 FILLER_14_696 ();
 sg13g2_fill_1 FILLER_14_703 ();
 sg13g2_decap_8 FILLER_14_708 ();
 sg13g2_decap_4 FILLER_14_715 ();
 sg13g2_fill_1 FILLER_14_719 ();
 sg13g2_fill_2 FILLER_14_729 ();
 sg13g2_fill_2 FILLER_14_762 ();
 sg13g2_fill_1 FILLER_14_764 ();
 sg13g2_fill_1 FILLER_14_777 ();
 sg13g2_fill_1 FILLER_14_783 ();
 sg13g2_fill_1 FILLER_14_815 ();
 sg13g2_fill_1 FILLER_14_845 ();
 sg13g2_fill_1 FILLER_14_851 ();
 sg13g2_fill_2 FILLER_14_857 ();
 sg13g2_fill_1 FILLER_14_867 ();
 sg13g2_decap_8 FILLER_14_873 ();
 sg13g2_fill_2 FILLER_14_880 ();
 sg13g2_decap_8 FILLER_14_886 ();
 sg13g2_fill_2 FILLER_14_934 ();
 sg13g2_fill_1 FILLER_14_948 ();
 sg13g2_fill_2 FILLER_14_1010 ();
 sg13g2_fill_1 FILLER_14_1012 ();
 sg13g2_fill_1 FILLER_14_1071 ();
 sg13g2_fill_2 FILLER_14_1111 ();
 sg13g2_fill_1 FILLER_14_1127 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_17 ();
 sg13g2_fill_2 FILLER_15_24 ();
 sg13g2_fill_1 FILLER_15_61 ();
 sg13g2_fill_2 FILLER_15_88 ();
 sg13g2_decap_4 FILLER_15_116 ();
 sg13g2_decap_4 FILLER_15_123 ();
 sg13g2_decap_4 FILLER_15_161 ();
 sg13g2_fill_1 FILLER_15_165 ();
 sg13g2_decap_4 FILLER_15_207 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_fill_1 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_234 ();
 sg13g2_fill_1 FILLER_15_241 ();
 sg13g2_fill_1 FILLER_15_248 ();
 sg13g2_fill_2 FILLER_15_283 ();
 sg13g2_fill_2 FILLER_15_322 ();
 sg13g2_fill_1 FILLER_15_327 ();
 sg13g2_fill_2 FILLER_15_370 ();
 sg13g2_fill_2 FILLER_15_484 ();
 sg13g2_fill_2 FILLER_15_511 ();
 sg13g2_fill_1 FILLER_15_531 ();
 sg13g2_fill_2 FILLER_15_541 ();
 sg13g2_fill_2 FILLER_15_587 ();
 sg13g2_fill_1 FILLER_15_603 ();
 sg13g2_fill_2 FILLER_15_668 ();
 sg13g2_fill_2 FILLER_15_696 ();
 sg13g2_fill_1 FILLER_15_698 ();
 sg13g2_decap_4 FILLER_15_703 ();
 sg13g2_fill_2 FILLER_15_707 ();
 sg13g2_decap_4 FILLER_15_714 ();
 sg13g2_decap_4 FILLER_15_723 ();
 sg13g2_fill_2 FILLER_15_749 ();
 sg13g2_fill_1 FILLER_15_751 ();
 sg13g2_fill_1 FILLER_15_762 ();
 sg13g2_decap_4 FILLER_15_778 ();
 sg13g2_fill_1 FILLER_15_794 ();
 sg13g2_fill_1 FILLER_15_800 ();
 sg13g2_fill_2 FILLER_15_811 ();
 sg13g2_fill_1 FILLER_15_822 ();
 sg13g2_fill_2 FILLER_15_849 ();
 sg13g2_fill_2 FILLER_15_872 ();
 sg13g2_fill_1 FILLER_15_900 ();
 sg13g2_fill_1 FILLER_15_913 ();
 sg13g2_fill_2 FILLER_15_926 ();
 sg13g2_fill_2 FILLER_15_975 ();
 sg13g2_fill_1 FILLER_15_977 ();
 sg13g2_fill_1 FILLER_15_982 ();
 sg13g2_fill_2 FILLER_15_1035 ();
 sg13g2_fill_1 FILLER_15_1037 ();
 sg13g2_fill_1 FILLER_15_1076 ();
 sg13g2_fill_2 FILLER_15_1177 ();
 sg13g2_fill_2 FILLER_15_1214 ();
 sg13g2_fill_1 FILLER_15_1216 ();
 sg13g2_fill_2 FILLER_15_1235 ();
 sg13g2_fill_1 FILLER_15_1237 ();
 sg13g2_fill_2 FILLER_15_1286 ();
 sg13g2_fill_1 FILLER_15_1288 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_fill_2 FILLER_16_187 ();
 sg13g2_fill_2 FILLER_16_207 ();
 sg13g2_fill_2 FILLER_16_249 ();
 sg13g2_fill_1 FILLER_16_364 ();
 sg13g2_fill_2 FILLER_16_450 ();
 sg13g2_fill_1 FILLER_16_477 ();
 sg13g2_fill_1 FILLER_16_526 ();
 sg13g2_fill_1 FILLER_16_634 ();
 sg13g2_fill_1 FILLER_16_640 ();
 sg13g2_decap_8 FILLER_16_698 ();
 sg13g2_fill_2 FILLER_16_715 ();
 sg13g2_decap_8 FILLER_16_723 ();
 sg13g2_fill_1 FILLER_16_730 ();
 sg13g2_fill_2 FILLER_16_749 ();
 sg13g2_decap_4 FILLER_16_776 ();
 sg13g2_fill_2 FILLER_16_794 ();
 sg13g2_fill_1 FILLER_16_796 ();
 sg13g2_decap_8 FILLER_16_802 ();
 sg13g2_decap_8 FILLER_16_815 ();
 sg13g2_fill_1 FILLER_16_822 ();
 sg13g2_fill_1 FILLER_16_835 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_fill_2 FILLER_16_847 ();
 sg13g2_fill_1 FILLER_16_849 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_4 FILLER_16_871 ();
 sg13g2_fill_1 FILLER_16_884 ();
 sg13g2_fill_2 FILLER_16_889 ();
 sg13g2_fill_1 FILLER_16_891 ();
 sg13g2_fill_2 FILLER_16_989 ();
 sg13g2_fill_1 FILLER_16_991 ();
 sg13g2_fill_1 FILLER_16_1009 ();
 sg13g2_fill_2 FILLER_16_1036 ();
 sg13g2_fill_1 FILLER_16_1038 ();
 sg13g2_fill_2 FILLER_16_1052 ();
 sg13g2_fill_1 FILLER_16_1054 ();
 sg13g2_fill_1 FILLER_16_1102 ();
 sg13g2_fill_1 FILLER_16_1116 ();
 sg13g2_fill_2 FILLER_16_1131 ();
 sg13g2_fill_2 FILLER_16_1198 ();
 sg13g2_fill_1 FILLER_16_1296 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_12 ();
 sg13g2_fill_2 FILLER_17_22 ();
 sg13g2_fill_1 FILLER_17_37 ();
 sg13g2_fill_2 FILLER_17_83 ();
 sg13g2_decap_4 FILLER_17_135 ();
 sg13g2_fill_1 FILLER_17_139 ();
 sg13g2_decap_8 FILLER_17_144 ();
 sg13g2_decap_8 FILLER_17_151 ();
 sg13g2_fill_1 FILLER_17_158 ();
 sg13g2_fill_1 FILLER_17_172 ();
 sg13g2_fill_1 FILLER_17_208 ();
 sg13g2_fill_1 FILLER_17_226 ();
 sg13g2_fill_2 FILLER_17_267 ();
 sg13g2_decap_4 FILLER_17_302 ();
 sg13g2_fill_2 FILLER_17_310 ();
 sg13g2_fill_1 FILLER_17_326 ();
 sg13g2_fill_2 FILLER_17_344 ();
 sg13g2_fill_1 FILLER_17_395 ();
 sg13g2_fill_2 FILLER_17_423 ();
 sg13g2_fill_1 FILLER_17_491 ();
 sg13g2_fill_1 FILLER_17_521 ();
 sg13g2_fill_2 FILLER_17_593 ();
 sg13g2_fill_1 FILLER_17_608 ();
 sg13g2_fill_2 FILLER_17_667 ();
 sg13g2_fill_1 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_691 ();
 sg13g2_decap_4 FILLER_17_698 ();
 sg13g2_fill_1 FILLER_17_702 ();
 sg13g2_fill_2 FILLER_17_708 ();
 sg13g2_decap_8 FILLER_17_719 ();
 sg13g2_fill_1 FILLER_17_739 ();
 sg13g2_fill_2 FILLER_17_748 ();
 sg13g2_fill_1 FILLER_17_750 ();
 sg13g2_fill_1 FILLER_17_770 ();
 sg13g2_fill_2 FILLER_17_795 ();
 sg13g2_fill_1 FILLER_17_797 ();
 sg13g2_fill_2 FILLER_17_856 ();
 sg13g2_fill_2 FILLER_17_882 ();
 sg13g2_decap_8 FILLER_17_889 ();
 sg13g2_decap_8 FILLER_17_896 ();
 sg13g2_fill_1 FILLER_17_903 ();
 sg13g2_decap_4 FILLER_17_909 ();
 sg13g2_fill_1 FILLER_17_917 ();
 sg13g2_fill_1 FILLER_17_948 ();
 sg13g2_fill_2 FILLER_17_1024 ();
 sg13g2_fill_1 FILLER_17_1091 ();
 sg13g2_fill_2 FILLER_17_1105 ();
 sg13g2_fill_1 FILLER_17_1107 ();
 sg13g2_fill_1 FILLER_17_1149 ();
 sg13g2_fill_2 FILLER_17_1251 ();
 sg13g2_fill_1 FILLER_17_1253 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_107 ();
 sg13g2_fill_1 FILLER_18_120 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_fill_2 FILLER_18_160 ();
 sg13g2_fill_1 FILLER_18_162 ();
 sg13g2_fill_1 FILLER_18_173 ();
 sg13g2_fill_2 FILLER_18_202 ();
 sg13g2_fill_1 FILLER_18_204 ();
 sg13g2_fill_2 FILLER_18_293 ();
 sg13g2_fill_1 FILLER_18_316 ();
 sg13g2_fill_2 FILLER_18_357 ();
 sg13g2_fill_2 FILLER_18_416 ();
 sg13g2_fill_2 FILLER_18_567 ();
 sg13g2_fill_1 FILLER_18_578 ();
 sg13g2_fill_2 FILLER_18_610 ();
 sg13g2_fill_1 FILLER_18_612 ();
 sg13g2_fill_2 FILLER_18_641 ();
 sg13g2_fill_2 FILLER_18_674 ();
 sg13g2_fill_2 FILLER_18_739 ();
 sg13g2_decap_4 FILLER_18_756 ();
 sg13g2_fill_1 FILLER_18_760 ();
 sg13g2_decap_8 FILLER_18_773 ();
 sg13g2_fill_2 FILLER_18_780 ();
 sg13g2_fill_1 FILLER_18_782 ();
 sg13g2_decap_8 FILLER_18_804 ();
 sg13g2_fill_2 FILLER_18_811 ();
 sg13g2_fill_1 FILLER_18_824 ();
 sg13g2_fill_2 FILLER_18_830 ();
 sg13g2_fill_2 FILLER_18_843 ();
 sg13g2_fill_1 FILLER_18_845 ();
 sg13g2_decap_8 FILLER_18_870 ();
 sg13g2_fill_2 FILLER_18_877 ();
 sg13g2_decap_8 FILLER_18_905 ();
 sg13g2_fill_2 FILLER_18_922 ();
 sg13g2_fill_2 FILLER_18_937 ();
 sg13g2_fill_1 FILLER_18_973 ();
 sg13g2_fill_1 FILLER_18_997 ();
 sg13g2_fill_1 FILLER_18_1007 ();
 sg13g2_fill_1 FILLER_18_1030 ();
 sg13g2_fill_2 FILLER_18_1049 ();
 sg13g2_fill_1 FILLER_18_1051 ();
 sg13g2_fill_1 FILLER_18_1065 ();
 sg13g2_fill_2 FILLER_18_1127 ();
 sg13g2_fill_1 FILLER_18_1129 ();
 sg13g2_fill_2 FILLER_18_1164 ();
 sg13g2_fill_1 FILLER_18_1197 ();
 sg13g2_fill_2 FILLER_18_1211 ();
 sg13g2_fill_1 FILLER_18_1213 ();
 sg13g2_fill_1 FILLER_18_1275 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_30 ();
 sg13g2_fill_2 FILLER_19_37 ();
 sg13g2_fill_1 FILLER_19_70 ();
 sg13g2_fill_2 FILLER_19_76 ();
 sg13g2_fill_2 FILLER_19_83 ();
 sg13g2_fill_1 FILLER_19_144 ();
 sg13g2_fill_1 FILLER_19_212 ();
 sg13g2_fill_1 FILLER_19_228 ();
 sg13g2_fill_1 FILLER_19_236 ();
 sg13g2_decap_8 FILLER_19_258 ();
 sg13g2_fill_2 FILLER_19_265 ();
 sg13g2_fill_2 FILLER_19_270 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_358 ();
 sg13g2_fill_2 FILLER_19_387 ();
 sg13g2_fill_2 FILLER_19_502 ();
 sg13g2_fill_2 FILLER_19_588 ();
 sg13g2_fill_2 FILLER_19_604 ();
 sg13g2_fill_1 FILLER_19_646 ();
 sg13g2_decap_8 FILLER_19_685 ();
 sg13g2_decap_4 FILLER_19_692 ();
 sg13g2_fill_1 FILLER_19_696 ();
 sg13g2_fill_1 FILLER_19_730 ();
 sg13g2_fill_1 FILLER_19_755 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_fill_2 FILLER_19_792 ();
 sg13g2_fill_1 FILLER_19_814 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_fill_2 FILLER_19_877 ();
 sg13g2_fill_1 FILLER_19_889 ();
 sg13g2_fill_1 FILLER_19_992 ();
 sg13g2_fill_1 FILLER_19_1019 ();
 sg13g2_fill_1 FILLER_19_1050 ();
 sg13g2_fill_2 FILLER_19_1060 ();
 sg13g2_fill_2 FILLER_19_1205 ();
 sg13g2_fill_1 FILLER_19_1225 ();
 sg13g2_fill_2 FILLER_19_1244 ();
 sg13g2_fill_1 FILLER_19_1246 ();
 sg13g2_fill_2 FILLER_19_1286 ();
 sg13g2_fill_1 FILLER_19_1288 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_12 ();
 sg13g2_fill_1 FILLER_20_14 ();
 sg13g2_decap_4 FILLER_20_23 ();
 sg13g2_fill_1 FILLER_20_27 ();
 sg13g2_fill_1 FILLER_20_46 ();
 sg13g2_fill_2 FILLER_20_68 ();
 sg13g2_fill_1 FILLER_20_122 ();
 sg13g2_fill_2 FILLER_20_153 ();
 sg13g2_fill_1 FILLER_20_155 ();
 sg13g2_fill_1 FILLER_20_169 ();
 sg13g2_decap_8 FILLER_20_261 ();
 sg13g2_decap_8 FILLER_20_272 ();
 sg13g2_fill_2 FILLER_20_279 ();
 sg13g2_fill_1 FILLER_20_281 ();
 sg13g2_decap_4 FILLER_20_287 ();
 sg13g2_fill_1 FILLER_20_291 ();
 sg13g2_fill_2 FILLER_20_296 ();
 sg13g2_fill_1 FILLER_20_309 ();
 sg13g2_fill_2 FILLER_20_355 ();
 sg13g2_fill_2 FILLER_20_373 ();
 sg13g2_fill_1 FILLER_20_413 ();
 sg13g2_fill_1 FILLER_20_526 ();
 sg13g2_fill_2 FILLER_20_565 ();
 sg13g2_fill_1 FILLER_20_618 ();
 sg13g2_fill_1 FILLER_20_654 ();
 sg13g2_fill_2 FILLER_20_692 ();
 sg13g2_fill_2 FILLER_20_756 ();
 sg13g2_fill_1 FILLER_20_758 ();
 sg13g2_fill_2 FILLER_20_764 ();
 sg13g2_fill_1 FILLER_20_766 ();
 sg13g2_fill_1 FILLER_20_783 ();
 sg13g2_fill_1 FILLER_20_800 ();
 sg13g2_fill_2 FILLER_20_806 ();
 sg13g2_fill_1 FILLER_20_808 ();
 sg13g2_decap_8 FILLER_20_829 ();
 sg13g2_decap_8 FILLER_20_836 ();
 sg13g2_decap_8 FILLER_20_843 ();
 sg13g2_fill_1 FILLER_20_850 ();
 sg13g2_fill_2 FILLER_20_877 ();
 sg13g2_fill_2 FILLER_20_894 ();
 sg13g2_fill_1 FILLER_20_913 ();
 sg13g2_fill_1 FILLER_20_980 ();
 sg13g2_fill_1 FILLER_20_995 ();
 sg13g2_fill_1 FILLER_20_1013 ();
 sg13g2_fill_1 FILLER_20_1033 ();
 sg13g2_fill_1 FILLER_20_1047 ();
 sg13g2_fill_2 FILLER_20_1087 ();
 sg13g2_fill_1 FILLER_20_1137 ();
 sg13g2_fill_2 FILLER_20_1177 ();
 sg13g2_fill_2 FILLER_20_1265 ();
 sg13g2_fill_1 FILLER_20_1267 ();
 sg13g2_fill_2 FILLER_20_1303 ();
 sg13g2_fill_1 FILLER_20_1305 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_39 ();
 sg13g2_fill_2 FILLER_21_46 ();
 sg13g2_fill_2 FILLER_21_101 ();
 sg13g2_fill_1 FILLER_21_124 ();
 sg13g2_fill_2 FILLER_21_159 ();
 sg13g2_fill_1 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_180 ();
 sg13g2_fill_1 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_219 ();
 sg13g2_fill_2 FILLER_21_226 ();
 sg13g2_decap_4 FILLER_21_233 ();
 sg13g2_fill_1 FILLER_21_237 ();
 sg13g2_decap_8 FILLER_21_242 ();
 sg13g2_fill_2 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_337 ();
 sg13g2_fill_1 FILLER_21_373 ();
 sg13g2_fill_1 FILLER_21_461 ();
 sg13g2_fill_1 FILLER_21_591 ();
 sg13g2_fill_1 FILLER_21_645 ();
 sg13g2_decap_8 FILLER_21_678 ();
 sg13g2_decap_4 FILLER_21_689 ();
 sg13g2_fill_2 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_744 ();
 sg13g2_decap_8 FILLER_21_751 ();
 sg13g2_fill_2 FILLER_21_763 ();
 sg13g2_fill_2 FILLER_21_795 ();
 sg13g2_fill_1 FILLER_21_797 ();
 sg13g2_fill_2 FILLER_21_803 ();
 sg13g2_fill_1 FILLER_21_805 ();
 sg13g2_decap_4 FILLER_21_819 ();
 sg13g2_fill_2 FILLER_21_823 ();
 sg13g2_fill_2 FILLER_21_839 ();
 sg13g2_fill_1 FILLER_21_841 ();
 sg13g2_decap_4 FILLER_21_847 ();
 sg13g2_decap_4 FILLER_21_868 ();
 sg13g2_decap_4 FILLER_21_956 ();
 sg13g2_fill_2 FILLER_21_960 ();
 sg13g2_fill_2 FILLER_21_971 ();
 sg13g2_fill_2 FILLER_21_1031 ();
 sg13g2_fill_1 FILLER_21_1042 ();
 sg13g2_fill_2 FILLER_21_1053 ();
 sg13g2_fill_1 FILLER_21_1055 ();
 sg13g2_fill_1 FILLER_21_1088 ();
 sg13g2_fill_2 FILLER_21_1095 ();
 sg13g2_fill_1 FILLER_21_1097 ();
 sg13g2_fill_1 FILLER_21_1103 ();
 sg13g2_fill_2 FILLER_21_1121 ();
 sg13g2_fill_1 FILLER_21_1123 ();
 sg13g2_fill_2 FILLER_21_1180 ();
 sg13g2_fill_1 FILLER_21_1288 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_4 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_67 ();
 sg13g2_fill_2 FILLER_22_104 ();
 sg13g2_fill_2 FILLER_22_132 ();
 sg13g2_decap_8 FILLER_22_162 ();
 sg13g2_decap_8 FILLER_22_169 ();
 sg13g2_decap_8 FILLER_22_176 ();
 sg13g2_decap_4 FILLER_22_183 ();
 sg13g2_fill_1 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_237 ();
 sg13g2_decap_4 FILLER_22_244 ();
 sg13g2_fill_1 FILLER_22_248 ();
 sg13g2_fill_2 FILLER_22_263 ();
 sg13g2_fill_1 FILLER_22_265 ();
 sg13g2_decap_4 FILLER_22_290 ();
 sg13g2_fill_2 FILLER_22_294 ();
 sg13g2_fill_2 FILLER_22_337 ();
 sg13g2_fill_1 FILLER_22_344 ();
 sg13g2_fill_2 FILLER_22_405 ();
 sg13g2_fill_2 FILLER_22_422 ();
 sg13g2_fill_2 FILLER_22_460 ();
 sg13g2_fill_2 FILLER_22_490 ();
 sg13g2_fill_2 FILLER_22_522 ();
 sg13g2_fill_2 FILLER_22_559 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_fill_1 FILLER_22_705 ();
 sg13g2_decap_8 FILLER_22_745 ();
 sg13g2_fill_1 FILLER_22_752 ();
 sg13g2_decap_4 FILLER_22_757 ();
 sg13g2_fill_1 FILLER_22_761 ();
 sg13g2_fill_1 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_782 ();
 sg13g2_decap_4 FILLER_22_789 ();
 sg13g2_fill_2 FILLER_22_793 ();
 sg13g2_fill_2 FILLER_22_807 ();
 sg13g2_fill_1 FILLER_22_809 ();
 sg13g2_fill_1 FILLER_22_820 ();
 sg13g2_decap_4 FILLER_22_847 ();
 sg13g2_fill_1 FILLER_22_851 ();
 sg13g2_fill_2 FILLER_22_858 ();
 sg13g2_decap_8 FILLER_22_865 ();
 sg13g2_decap_8 FILLER_22_872 ();
 sg13g2_decap_4 FILLER_22_879 ();
 sg13g2_fill_1 FILLER_22_893 ();
 sg13g2_fill_1 FILLER_22_898 ();
 sg13g2_fill_2 FILLER_22_915 ();
 sg13g2_decap_4 FILLER_22_964 ();
 sg13g2_fill_1 FILLER_22_968 ();
 sg13g2_fill_2 FILLER_22_978 ();
 sg13g2_fill_1 FILLER_22_1089 ();
 sg13g2_fill_2 FILLER_22_1104 ();
 sg13g2_fill_1 FILLER_22_1106 ();
 sg13g2_fill_2 FILLER_22_1123 ();
 sg13g2_fill_2 FILLER_22_1135 ();
 sg13g2_fill_1 FILLER_22_1137 ();
 sg13g2_fill_1 FILLER_22_1252 ();
 sg13g2_fill_1 FILLER_22_1314 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_4 ();
 sg13g2_fill_1 FILLER_23_13 ();
 sg13g2_fill_2 FILLER_23_18 ();
 sg13g2_fill_1 FILLER_23_38 ();
 sg13g2_decap_4 FILLER_23_65 ();
 sg13g2_fill_2 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_86 ();
 sg13g2_fill_1 FILLER_23_88 ();
 sg13g2_decap_4 FILLER_23_96 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_221 ();
 sg13g2_fill_2 FILLER_23_228 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_decap_4 FILLER_23_244 ();
 sg13g2_fill_2 FILLER_23_248 ();
 sg13g2_decap_4 FILLER_23_292 ();
 sg13g2_fill_2 FILLER_23_296 ();
 sg13g2_fill_2 FILLER_23_391 ();
 sg13g2_fill_2 FILLER_23_432 ();
 sg13g2_fill_2 FILLER_23_456 ();
 sg13g2_fill_1 FILLER_23_507 ();
 sg13g2_fill_1 FILLER_23_647 ();
 sg13g2_fill_2 FILLER_23_722 ();
 sg13g2_fill_2 FILLER_23_764 ();
 sg13g2_fill_1 FILLER_23_766 ();
 sg13g2_fill_2 FILLER_23_800 ();
 sg13g2_fill_2 FILLER_23_845 ();
 sg13g2_decap_4 FILLER_23_859 ();
 sg13g2_fill_1 FILLER_23_863 ();
 sg13g2_fill_1 FILLER_23_873 ();
 sg13g2_fill_1 FILLER_23_879 ();
 sg13g2_decap_4 FILLER_23_884 ();
 sg13g2_fill_2 FILLER_23_888 ();
 sg13g2_fill_2 FILLER_23_985 ();
 sg13g2_fill_1 FILLER_23_987 ();
 sg13g2_fill_2 FILLER_23_1009 ();
 sg13g2_fill_2 FILLER_23_1015 ();
 sg13g2_fill_1 FILLER_23_1017 ();
 sg13g2_fill_2 FILLER_23_1056 ();
 sg13g2_fill_1 FILLER_23_1058 ();
 sg13g2_fill_2 FILLER_23_1084 ();
 sg13g2_fill_1 FILLER_23_1086 ();
 sg13g2_fill_1 FILLER_23_1093 ();
 sg13g2_fill_2 FILLER_23_1106 ();
 sg13g2_fill_1 FILLER_23_1126 ();
 sg13g2_fill_1 FILLER_23_1145 ();
 sg13g2_fill_2 FILLER_23_1167 ();
 sg13g2_fill_1 FILLER_23_1169 ();
 sg13g2_fill_2 FILLER_23_1264 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_67 ();
 sg13g2_fill_1 FILLER_24_121 ();
 sg13g2_fill_2 FILLER_24_127 ();
 sg13g2_fill_1 FILLER_24_155 ();
 sg13g2_fill_2 FILLER_24_192 ();
 sg13g2_fill_2 FILLER_24_213 ();
 sg13g2_fill_2 FILLER_24_223 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_4 FILLER_24_280 ();
 sg13g2_fill_2 FILLER_24_350 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_fill_1 FILLER_24_466 ();
 sg13g2_fill_1 FILLER_24_499 ();
 sg13g2_fill_2 FILLER_24_531 ();
 sg13g2_fill_1 FILLER_24_614 ();
 sg13g2_fill_2 FILLER_24_669 ();
 sg13g2_fill_1 FILLER_24_671 ();
 sg13g2_fill_1 FILLER_24_681 ();
 sg13g2_fill_1 FILLER_24_716 ();
 sg13g2_fill_2 FILLER_24_731 ();
 sg13g2_fill_1 FILLER_24_733 ();
 sg13g2_fill_2 FILLER_24_782 ();
 sg13g2_fill_1 FILLER_24_811 ();
 sg13g2_fill_1 FILLER_24_820 ();
 sg13g2_fill_1 FILLER_24_914 ();
 sg13g2_fill_1 FILLER_24_921 ();
 sg13g2_decap_8 FILLER_24_993 ();
 sg13g2_fill_2 FILLER_24_1026 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_fill_1 FILLER_24_1033 ();
 sg13g2_fill_2 FILLER_24_1038 ();
 sg13g2_fill_1 FILLER_24_1053 ();
 sg13g2_fill_2 FILLER_24_1058 ();
 sg13g2_fill_2 FILLER_24_1064 ();
 sg13g2_fill_1 FILLER_24_1092 ();
 sg13g2_fill_2 FILLER_24_1136 ();
 sg13g2_fill_1 FILLER_24_1138 ();
 sg13g2_fill_2 FILLER_24_1169 ();
 sg13g2_fill_2 FILLER_24_1223 ();
 sg13g2_fill_2 FILLER_24_1260 ();
 sg13g2_fill_1 FILLER_24_1314 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_94 ();
 sg13g2_decap_4 FILLER_25_101 ();
 sg13g2_fill_1 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_110 ();
 sg13g2_decap_4 FILLER_25_121 ();
 sg13g2_fill_2 FILLER_25_125 ();
 sg13g2_fill_2 FILLER_25_237 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_decap_4 FILLER_25_283 ();
 sg13g2_fill_1 FILLER_25_287 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_fill_1 FILLER_25_474 ();
 sg13g2_fill_2 FILLER_25_510 ();
 sg13g2_fill_1 FILLER_25_521 ();
 sg13g2_fill_1 FILLER_25_576 ();
 sg13g2_fill_2 FILLER_25_590 ();
 sg13g2_fill_1 FILLER_25_605 ();
 sg13g2_fill_1 FILLER_25_637 ();
 sg13g2_fill_1 FILLER_25_666 ();
 sg13g2_fill_2 FILLER_25_745 ();
 sg13g2_fill_1 FILLER_25_747 ();
 sg13g2_fill_2 FILLER_25_788 ();
 sg13g2_fill_1 FILLER_25_814 ();
 sg13g2_decap_8 FILLER_25_837 ();
 sg13g2_fill_2 FILLER_25_844 ();
 sg13g2_decap_4 FILLER_25_851 ();
 sg13g2_decap_8 FILLER_25_864 ();
 sg13g2_decap_4 FILLER_25_871 ();
 sg13g2_fill_1 FILLER_25_875 ();
 sg13g2_fill_2 FILLER_25_1008 ();
 sg13g2_fill_1 FILLER_25_1010 ();
 sg13g2_fill_2 FILLER_25_1020 ();
 sg13g2_fill_1 FILLER_25_1022 ();
 sg13g2_fill_1 FILLER_25_1075 ();
 sg13g2_fill_2 FILLER_25_1106 ();
 sg13g2_fill_1 FILLER_25_1108 ();
 sg13g2_fill_2 FILLER_25_1135 ();
 sg13g2_fill_2 FILLER_25_1241 ();
 sg13g2_fill_2 FILLER_25_1287 ();
 sg13g2_fill_1 FILLER_26_74 ();
 sg13g2_fill_1 FILLER_26_88 ();
 sg13g2_fill_2 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_104 ();
 sg13g2_fill_2 FILLER_26_111 ();
 sg13g2_fill_2 FILLER_26_178 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_fill_2 FILLER_26_253 ();
 sg13g2_fill_1 FILLER_26_255 ();
 sg13g2_fill_2 FILLER_26_265 ();
 sg13g2_fill_1 FILLER_26_267 ();
 sg13g2_decap_8 FILLER_26_285 ();
 sg13g2_fill_2 FILLER_26_318 ();
 sg13g2_fill_1 FILLER_26_364 ();
 sg13g2_fill_2 FILLER_26_374 ();
 sg13g2_fill_2 FILLER_26_416 ();
 sg13g2_fill_2 FILLER_26_474 ();
 sg13g2_fill_1 FILLER_26_554 ();
 sg13g2_fill_2 FILLER_26_585 ();
 sg13g2_decap_8 FILLER_26_669 ();
 sg13g2_fill_1 FILLER_26_676 ();
 sg13g2_fill_2 FILLER_26_686 ();
 sg13g2_fill_1 FILLER_26_688 ();
 sg13g2_fill_2 FILLER_26_693 ();
 sg13g2_fill_2 FILLER_26_717 ();
 sg13g2_fill_2 FILLER_26_728 ();
 sg13g2_fill_1 FILLER_26_829 ();
 sg13g2_decap_4 FILLER_26_846 ();
 sg13g2_fill_2 FILLER_26_857 ();
 sg13g2_fill_1 FILLER_26_902 ();
 sg13g2_fill_1 FILLER_26_1032 ();
 sg13g2_fill_2 FILLER_26_1078 ();
 sg13g2_fill_2 FILLER_26_1084 ();
 sg13g2_fill_1 FILLER_26_1086 ();
 sg13g2_fill_2 FILLER_26_1095 ();
 sg13g2_fill_1 FILLER_26_1097 ();
 sg13g2_fill_2 FILLER_26_1145 ();
 sg13g2_fill_1 FILLER_26_1147 ();
 sg13g2_fill_2 FILLER_26_1152 ();
 sg13g2_fill_1 FILLER_26_1154 ();
 sg13g2_fill_2 FILLER_26_1180 ();
 sg13g2_fill_1 FILLER_26_1182 ();
 sg13g2_fill_1 FILLER_26_1188 ();
 sg13g2_fill_1 FILLER_26_1198 ();
 sg13g2_fill_2 FILLER_26_1303 ();
 sg13g2_fill_1 FILLER_26_1305 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_12 ();
 sg13g2_fill_2 FILLER_27_18 ();
 sg13g2_fill_1 FILLER_27_23 ();
 sg13g2_fill_1 FILLER_27_53 ();
 sg13g2_fill_1 FILLER_27_58 ();
 sg13g2_decap_8 FILLER_27_115 ();
 sg13g2_fill_2 FILLER_27_122 ();
 sg13g2_fill_2 FILLER_27_134 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_fill_2 FILLER_27_156 ();
 sg13g2_fill_2 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_195 ();
 sg13g2_fill_1 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_fill_2 FILLER_27_228 ();
 sg13g2_decap_4 FILLER_27_239 ();
 sg13g2_fill_2 FILLER_27_249 ();
 sg13g2_fill_1 FILLER_27_251 ();
 sg13g2_decap_4 FILLER_27_292 ();
 sg13g2_fill_1 FILLER_27_296 ();
 sg13g2_fill_1 FILLER_27_300 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_fill_2 FILLER_27_326 ();
 sg13g2_fill_2 FILLER_27_343 ();
 sg13g2_fill_2 FILLER_27_384 ();
 sg13g2_fill_1 FILLER_27_391 ();
 sg13g2_fill_2 FILLER_27_451 ();
 sg13g2_fill_2 FILLER_27_482 ();
 sg13g2_fill_2 FILLER_27_545 ();
 sg13g2_fill_1 FILLER_27_565 ();
 sg13g2_fill_1 FILLER_27_596 ();
 sg13g2_fill_2 FILLER_27_601 ();
 sg13g2_fill_1 FILLER_27_603 ();
 sg13g2_decap_8 FILLER_27_648 ();
 sg13g2_decap_8 FILLER_27_655 ();
 sg13g2_fill_1 FILLER_27_662 ();
 sg13g2_fill_2 FILLER_27_689 ();
 sg13g2_fill_2 FILLER_27_696 ();
 sg13g2_fill_1 FILLER_27_698 ();
 sg13g2_fill_2 FILLER_27_803 ();
 sg13g2_fill_2 FILLER_27_848 ();
 sg13g2_fill_2 FILLER_27_865 ();
 sg13g2_fill_1 FILLER_27_867 ();
 sg13g2_fill_1 FILLER_27_892 ();
 sg13g2_fill_2 FILLER_27_945 ();
 sg13g2_fill_1 FILLER_27_947 ();
 sg13g2_fill_2 FILLER_27_981 ();
 sg13g2_fill_1 FILLER_27_983 ();
 sg13g2_fill_2 FILLER_27_1007 ();
 sg13g2_fill_1 FILLER_27_1061 ();
 sg13g2_fill_2 FILLER_27_1067 ();
 sg13g2_fill_1 FILLER_27_1129 ();
 sg13g2_fill_1 FILLER_27_1156 ();
 sg13g2_fill_2 FILLER_28_29 ();
 sg13g2_fill_2 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_96 ();
 sg13g2_fill_1 FILLER_28_113 ();
 sg13g2_fill_2 FILLER_28_136 ();
 sg13g2_fill_1 FILLER_28_138 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_239 ();
 sg13g2_fill_1 FILLER_28_241 ();
 sg13g2_fill_2 FILLER_28_256 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_fill_2 FILLER_28_263 ();
 sg13g2_decap_8 FILLER_28_290 ();
 sg13g2_fill_1 FILLER_28_297 ();
 sg13g2_decap_8 FILLER_28_304 ();
 sg13g2_decap_4 FILLER_28_311 ();
 sg13g2_fill_1 FILLER_28_325 ();
 sg13g2_fill_1 FILLER_28_368 ();
 sg13g2_fill_2 FILLER_28_438 ();
 sg13g2_fill_2 FILLER_28_466 ();
 sg13g2_fill_1 FILLER_28_468 ();
 sg13g2_fill_2 FILLER_28_503 ();
 sg13g2_fill_2 FILLER_28_514 ();
 sg13g2_fill_2 FILLER_28_563 ();
 sg13g2_fill_1 FILLER_28_570 ();
 sg13g2_fill_2 FILLER_28_580 ();
 sg13g2_fill_2 FILLER_28_622 ();
 sg13g2_fill_1 FILLER_28_624 ();
 sg13g2_decap_8 FILLER_28_638 ();
 sg13g2_decap_8 FILLER_28_653 ();
 sg13g2_decap_4 FILLER_28_660 ();
 sg13g2_fill_1 FILLER_28_664 ();
 sg13g2_fill_2 FILLER_28_722 ();
 sg13g2_fill_2 FILLER_28_737 ();
 sg13g2_fill_1 FILLER_28_760 ();
 sg13g2_fill_2 FILLER_28_766 ();
 sg13g2_decap_4 FILLER_28_771 ();
 sg13g2_fill_2 FILLER_28_775 ();
 sg13g2_fill_1 FILLER_28_794 ();
 sg13g2_decap_4 FILLER_28_825 ();
 sg13g2_fill_2 FILLER_28_833 ();
 sg13g2_fill_1 FILLER_28_835 ();
 sg13g2_decap_4 FILLER_28_841 ();
 sg13g2_decap_4 FILLER_28_858 ();
 sg13g2_fill_2 FILLER_28_862 ();
 sg13g2_fill_1 FILLER_28_870 ();
 sg13g2_decap_4 FILLER_28_902 ();
 sg13g2_fill_2 FILLER_28_950 ();
 sg13g2_fill_1 FILLER_28_1013 ();
 sg13g2_decap_8 FILLER_28_1044 ();
 sg13g2_fill_2 FILLER_28_1051 ();
 sg13g2_fill_1 FILLER_28_1053 ();
 sg13g2_fill_2 FILLER_28_1086 ();
 sg13g2_fill_1 FILLER_28_1088 ();
 sg13g2_fill_2 FILLER_28_1117 ();
 sg13g2_fill_1 FILLER_28_1138 ();
 sg13g2_fill_2 FILLER_28_1180 ();
 sg13g2_fill_1 FILLER_28_1182 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_13 ();
 sg13g2_fill_2 FILLER_29_18 ();
 sg13g2_fill_1 FILLER_29_67 ();
 sg13g2_fill_2 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_179 ();
 sg13g2_decap_4 FILLER_29_194 ();
 sg13g2_fill_2 FILLER_29_198 ();
 sg13g2_fill_2 FILLER_29_249 ();
 sg13g2_fill_1 FILLER_29_251 ();
 sg13g2_decap_8 FILLER_29_283 ();
 sg13g2_decap_8 FILLER_29_314 ();
 sg13g2_decap_8 FILLER_29_321 ();
 sg13g2_fill_2 FILLER_29_328 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_fill_2 FILLER_29_375 ();
 sg13g2_fill_1 FILLER_29_381 ();
 sg13g2_fill_1 FILLER_29_445 ();
 sg13g2_fill_1 FILLER_29_464 ();
 sg13g2_fill_1 FILLER_29_489 ();
 sg13g2_fill_1 FILLER_29_515 ();
 sg13g2_fill_1 FILLER_29_523 ();
 sg13g2_fill_2 FILLER_29_531 ();
 sg13g2_fill_2 FILLER_29_612 ();
 sg13g2_fill_1 FILLER_29_640 ();
 sg13g2_decap_4 FILLER_29_661 ();
 sg13g2_fill_2 FILLER_29_686 ();
 sg13g2_fill_1 FILLER_29_693 ();
 sg13g2_fill_2 FILLER_29_703 ();
 sg13g2_fill_1 FILLER_29_751 ();
 sg13g2_fill_1 FILLER_29_756 ();
 sg13g2_decap_8 FILLER_29_792 ();
 sg13g2_fill_2 FILLER_29_799 ();
 sg13g2_fill_1 FILLER_29_862 ();
 sg13g2_decap_4 FILLER_29_868 ();
 sg13g2_fill_1 FILLER_29_892 ();
 sg13g2_fill_2 FILLER_29_919 ();
 sg13g2_fill_2 FILLER_29_995 ();
 sg13g2_fill_2 FILLER_29_1075 ();
 sg13g2_fill_1 FILLER_29_1077 ();
 sg13g2_fill_1 FILLER_29_1288 ();
 sg13g2_fill_2 FILLER_30_34 ();
 sg13g2_fill_2 FILLER_30_55 ();
 sg13g2_fill_1 FILLER_30_73 ();
 sg13g2_fill_2 FILLER_30_93 ();
 sg13g2_fill_1 FILLER_30_125 ();
 sg13g2_fill_2 FILLER_30_134 ();
 sg13g2_fill_1 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_177 ();
 sg13g2_fill_2 FILLER_30_184 ();
 sg13g2_fill_2 FILLER_30_217 ();
 sg13g2_fill_1 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_255 ();
 sg13g2_fill_2 FILLER_30_280 ();
 sg13g2_fill_2 FILLER_30_296 ();
 sg13g2_fill_1 FILLER_30_303 ();
 sg13g2_decap_8 FILLER_30_323 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_decap_4 FILLER_30_393 ();
 sg13g2_fill_2 FILLER_30_481 ();
 sg13g2_fill_1 FILLER_30_483 ();
 sg13g2_fill_2 FILLER_30_495 ();
 sg13g2_fill_2 FILLER_30_505 ();
 sg13g2_fill_1 FILLER_30_518 ();
 sg13g2_fill_1 FILLER_30_527 ();
 sg13g2_fill_1 FILLER_30_533 ();
 sg13g2_fill_2 FILLER_30_562 ();
 sg13g2_fill_2 FILLER_30_577 ();
 sg13g2_fill_2 FILLER_30_611 ();
 sg13g2_fill_2 FILLER_30_631 ();
 sg13g2_fill_1 FILLER_30_633 ();
 sg13g2_fill_2 FILLER_30_642 ();
 sg13g2_fill_2 FILLER_30_650 ();
 sg13g2_fill_1 FILLER_30_657 ();
 sg13g2_fill_1 FILLER_30_684 ();
 sg13g2_fill_1 FILLER_30_711 ();
 sg13g2_fill_1 FILLER_30_718 ();
 sg13g2_fill_2 FILLER_30_730 ();
 sg13g2_fill_1 FILLER_30_741 ();
 sg13g2_fill_1 FILLER_30_768 ();
 sg13g2_fill_1 FILLER_30_800 ();
 sg13g2_decap_8 FILLER_30_832 ();
 sg13g2_fill_2 FILLER_30_839 ();
 sg13g2_fill_1 FILLER_30_841 ();
 sg13g2_fill_1 FILLER_30_857 ();
 sg13g2_fill_1 FILLER_30_875 ();
 sg13g2_fill_2 FILLER_30_913 ();
 sg13g2_fill_1 FILLER_30_915 ();
 sg13g2_fill_2 FILLER_30_931 ();
 sg13g2_fill_2 FILLER_30_946 ();
 sg13g2_fill_1 FILLER_30_948 ();
 sg13g2_fill_1 FILLER_30_969 ();
 sg13g2_fill_2 FILLER_30_992 ();
 sg13g2_fill_2 FILLER_30_1030 ();
 sg13g2_fill_1 FILLER_30_1032 ();
 sg13g2_fill_2 FILLER_30_1042 ();
 sg13g2_fill_1 FILLER_30_1044 ();
 sg13g2_fill_2 FILLER_30_1089 ();
 sg13g2_fill_2 FILLER_30_1128 ();
 sg13g2_fill_2 FILLER_30_1155 ();
 sg13g2_fill_2 FILLER_30_1192 ();
 sg13g2_fill_2 FILLER_30_1217 ();
 sg13g2_fill_1 FILLER_30_1250 ();
 sg13g2_fill_2 FILLER_30_1312 ();
 sg13g2_fill_1 FILLER_30_1314 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_4 ();
 sg13g2_fill_2 FILLER_31_9 ();
 sg13g2_fill_1 FILLER_31_11 ();
 sg13g2_decap_4 FILLER_31_20 ();
 sg13g2_fill_2 FILLER_31_29 ();
 sg13g2_fill_2 FILLER_31_44 ();
 sg13g2_fill_1 FILLER_31_87 ();
 sg13g2_fill_2 FILLER_31_108 ();
 sg13g2_fill_1 FILLER_31_131 ();
 sg13g2_fill_1 FILLER_31_142 ();
 sg13g2_fill_1 FILLER_31_151 ();
 sg13g2_fill_1 FILLER_31_196 ();
 sg13g2_fill_2 FILLER_31_274 ();
 sg13g2_decap_4 FILLER_31_319 ();
 sg13g2_fill_2 FILLER_31_339 ();
 sg13g2_decap_4 FILLER_31_373 ();
 sg13g2_fill_1 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_fill_1 FILLER_31_393 ();
 sg13g2_fill_1 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_432 ();
 sg13g2_fill_2 FILLER_31_444 ();
 sg13g2_fill_1 FILLER_31_446 ();
 sg13g2_fill_1 FILLER_31_469 ();
 sg13g2_fill_2 FILLER_31_523 ();
 sg13g2_fill_1 FILLER_31_531 ();
 sg13g2_fill_2 FILLER_31_561 ();
 sg13g2_decap_8 FILLER_31_594 ();
 sg13g2_fill_1 FILLER_31_601 ();
 sg13g2_decap_8 FILLER_31_606 ();
 sg13g2_fill_1 FILLER_31_613 ();
 sg13g2_fill_2 FILLER_31_620 ();
 sg13g2_fill_1 FILLER_31_622 ();
 sg13g2_fill_2 FILLER_31_649 ();
 sg13g2_fill_2 FILLER_31_686 ();
 sg13g2_fill_1 FILLER_31_688 ();
 sg13g2_fill_1 FILLER_31_705 ();
 sg13g2_fill_1 FILLER_31_760 ();
 sg13g2_decap_8 FILLER_31_767 ();
 sg13g2_fill_1 FILLER_31_779 ();
 sg13g2_fill_1 FILLER_31_789 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_4 FILLER_31_826 ();
 sg13g2_decap_4 FILLER_31_839 ();
 sg13g2_fill_1 FILLER_31_843 ();
 sg13g2_decap_8 FILLER_31_850 ();
 sg13g2_decap_4 FILLER_31_857 ();
 sg13g2_fill_2 FILLER_31_861 ();
 sg13g2_fill_1 FILLER_31_877 ();
 sg13g2_fill_2 FILLER_31_915 ();
 sg13g2_fill_2 FILLER_31_939 ();
 sg13g2_fill_1 FILLER_31_947 ();
 sg13g2_decap_8 FILLER_31_1029 ();
 sg13g2_fill_2 FILLER_31_1036 ();
 sg13g2_fill_2 FILLER_31_1092 ();
 sg13g2_fill_1 FILLER_31_1094 ();
 sg13g2_fill_2 FILLER_31_1114 ();
 sg13g2_fill_2 FILLER_31_1152 ();
 sg13g2_fill_1 FILLER_31_1170 ();
 sg13g2_fill_1 FILLER_31_1197 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_27 ();
 sg13g2_fill_2 FILLER_32_64 ();
 sg13g2_fill_2 FILLER_32_100 ();
 sg13g2_fill_2 FILLER_32_219 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_decap_4 FILLER_32_308 ();
 sg13g2_fill_2 FILLER_32_312 ();
 sg13g2_decap_4 FILLER_32_334 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_350 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_fill_2 FILLER_32_381 ();
 sg13g2_fill_1 FILLER_32_414 ();
 sg13g2_fill_2 FILLER_32_446 ();
 sg13g2_fill_2 FILLER_32_483 ();
 sg13g2_fill_1 FILLER_32_485 ();
 sg13g2_fill_2 FILLER_32_512 ();
 sg13g2_fill_1 FILLER_32_535 ();
 sg13g2_decap_4 FILLER_32_545 ();
 sg13g2_fill_2 FILLER_32_558 ();
 sg13g2_fill_1 FILLER_32_565 ();
 sg13g2_fill_2 FILLER_32_571 ();
 sg13g2_fill_2 FILLER_32_632 ();
 sg13g2_fill_1 FILLER_32_634 ();
 sg13g2_fill_1 FILLER_32_641 ();
 sg13g2_fill_2 FILLER_32_646 ();
 sg13g2_fill_2 FILLER_32_656 ();
 sg13g2_fill_1 FILLER_32_658 ();
 sg13g2_fill_2 FILLER_32_668 ();
 sg13g2_fill_2 FILLER_32_719 ();
 sg13g2_fill_1 FILLER_32_721 ();
 sg13g2_fill_2 FILLER_32_743 ();
 sg13g2_fill_1 FILLER_32_771 ();
 sg13g2_fill_1 FILLER_32_795 ();
 sg13g2_decap_8 FILLER_32_813 ();
 sg13g2_decap_4 FILLER_32_820 ();
 sg13g2_fill_1 FILLER_32_824 ();
 sg13g2_fill_2 FILLER_32_830 ();
 sg13g2_fill_1 FILLER_32_832 ();
 sg13g2_decap_8 FILLER_32_859 ();
 sg13g2_decap_4 FILLER_32_874 ();
 sg13g2_fill_2 FILLER_32_882 ();
 sg13g2_fill_1 FILLER_32_884 ();
 sg13g2_decap_8 FILLER_32_893 ();
 sg13g2_fill_2 FILLER_32_900 ();
 sg13g2_fill_1 FILLER_32_902 ();
 sg13g2_fill_1 FILLER_32_916 ();
 sg13g2_fill_2 FILLER_32_937 ();
 sg13g2_fill_1 FILLER_32_944 ();
 sg13g2_fill_1 FILLER_32_968 ();
 sg13g2_fill_2 FILLER_32_995 ();
 sg13g2_fill_1 FILLER_32_997 ();
 sg13g2_fill_1 FILLER_32_1008 ();
 sg13g2_fill_1 FILLER_32_1114 ();
 sg13g2_fill_1 FILLER_32_1140 ();
 sg13g2_fill_2 FILLER_32_1211 ();
 sg13g2_fill_1 FILLER_32_1213 ();
 sg13g2_fill_1 FILLER_32_1266 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_112 ();
 sg13g2_fill_2 FILLER_33_199 ();
 sg13g2_fill_1 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_233 ();
 sg13g2_fill_1 FILLER_33_244 ();
 sg13g2_decap_8 FILLER_33_289 ();
 sg13g2_fill_2 FILLER_33_296 ();
 sg13g2_fill_1 FILLER_33_298 ();
 sg13g2_decap_4 FILLER_33_312 ();
 sg13g2_fill_2 FILLER_33_316 ();
 sg13g2_decap_4 FILLER_33_323 ();
 sg13g2_fill_2 FILLER_33_363 ();
 sg13g2_fill_1 FILLER_33_377 ();
 sg13g2_fill_1 FILLER_33_425 ();
 sg13g2_decap_4 FILLER_33_435 ();
 sg13g2_fill_2 FILLER_33_439 ();
 sg13g2_fill_1 FILLER_33_471 ();
 sg13g2_fill_1 FILLER_33_481 ();
 sg13g2_fill_2 FILLER_33_492 ();
 sg13g2_fill_1 FILLER_33_499 ();
 sg13g2_decap_4 FILLER_33_508 ();
 sg13g2_fill_2 FILLER_33_527 ();
 sg13g2_fill_2 FILLER_33_560 ();
 sg13g2_decap_8 FILLER_33_602 ();
 sg13g2_decap_8 FILLER_33_609 ();
 sg13g2_fill_1 FILLER_33_616 ();
 sg13g2_fill_2 FILLER_33_632 ();
 sg13g2_fill_2 FILLER_33_640 ();
 sg13g2_fill_1 FILLER_33_652 ();
 sg13g2_decap_4 FILLER_33_664 ();
 sg13g2_fill_2 FILLER_33_676 ();
 sg13g2_decap_8 FILLER_33_695 ();
 sg13g2_decap_8 FILLER_33_702 ();
 sg13g2_fill_2 FILLER_33_709 ();
 sg13g2_fill_2 FILLER_33_716 ();
 sg13g2_fill_1 FILLER_33_718 ();
 sg13g2_fill_1 FILLER_33_745 ();
 sg13g2_fill_1 FILLER_33_773 ();
 sg13g2_fill_1 FILLER_33_786 ();
 sg13g2_fill_2 FILLER_33_799 ();
 sg13g2_decap_4 FILLER_33_825 ();
 sg13g2_fill_2 FILLER_33_850 ();
 sg13g2_fill_1 FILLER_33_852 ();
 sg13g2_fill_1 FILLER_33_879 ();
 sg13g2_fill_2 FILLER_33_949 ();
 sg13g2_fill_1 FILLER_33_986 ();
 sg13g2_decap_8 FILLER_33_1008 ();
 sg13g2_fill_2 FILLER_33_1041 ();
 sg13g2_fill_1 FILLER_33_1043 ();
 sg13g2_fill_2 FILLER_33_1070 ();
 sg13g2_fill_1 FILLER_33_1072 ();
 sg13g2_fill_1 FILLER_33_1079 ();
 sg13g2_fill_1 FILLER_33_1095 ();
 sg13g2_decap_4 FILLER_33_1111 ();
 sg13g2_fill_2 FILLER_33_1155 ();
 sg13g2_fill_1 FILLER_33_1157 ();
 sg13g2_fill_2 FILLER_33_1174 ();
 sg13g2_fill_1 FILLER_33_1176 ();
 sg13g2_fill_2 FILLER_33_1246 ();
 sg13g2_fill_1 FILLER_33_1288 ();
 sg13g2_fill_1 FILLER_34_144 ();
 sg13g2_fill_2 FILLER_34_209 ();
 sg13g2_fill_2 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_247 ();
 sg13g2_fill_1 FILLER_34_274 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_fill_2 FILLER_34_287 ();
 sg13g2_fill_1 FILLER_34_289 ();
 sg13g2_decap_4 FILLER_34_391 ();
 sg13g2_fill_2 FILLER_34_395 ();
 sg13g2_fill_2 FILLER_34_421 ();
 sg13g2_fill_2 FILLER_34_432 ();
 sg13g2_fill_2 FILLER_34_444 ();
 sg13g2_fill_2 FILLER_34_464 ();
 sg13g2_fill_1 FILLER_34_466 ();
 sg13g2_fill_1 FILLER_34_484 ();
 sg13g2_decap_4 FILLER_34_526 ();
 sg13g2_fill_2 FILLER_34_535 ();
 sg13g2_decap_8 FILLER_34_551 ();
 sg13g2_fill_1 FILLER_34_558 ();
 sg13g2_fill_1 FILLER_34_582 ();
 sg13g2_fill_2 FILLER_34_623 ();
 sg13g2_fill_1 FILLER_34_625 ();
 sg13g2_fill_2 FILLER_34_701 ();
 sg13g2_fill_1 FILLER_34_703 ();
 sg13g2_decap_4 FILLER_34_709 ();
 sg13g2_fill_1 FILLER_34_713 ();
 sg13g2_decap_8 FILLER_34_776 ();
 sg13g2_fill_1 FILLER_34_783 ();
 sg13g2_decap_4 FILLER_34_790 ();
 sg13g2_fill_1 FILLER_34_794 ();
 sg13g2_fill_2 FILLER_34_805 ();
 sg13g2_fill_1 FILLER_34_807 ();
 sg13g2_fill_1 FILLER_34_824 ();
 sg13g2_fill_2 FILLER_34_838 ();
 sg13g2_decap_8 FILLER_34_854 ();
 sg13g2_decap_8 FILLER_34_874 ();
 sg13g2_decap_4 FILLER_34_881 ();
 sg13g2_decap_8 FILLER_34_889 ();
 sg13g2_decap_4 FILLER_34_896 ();
 sg13g2_fill_2 FILLER_34_900 ();
 sg13g2_fill_1 FILLER_34_940 ();
 sg13g2_fill_1 FILLER_34_970 ();
 sg13g2_decap_4 FILLER_34_984 ();
 sg13g2_fill_1 FILLER_34_988 ();
 sg13g2_fill_1 FILLER_34_999 ();
 sg13g2_decap_8 FILLER_34_1026 ();
 sg13g2_decap_4 FILLER_34_1033 ();
 sg13g2_fill_1 FILLER_34_1037 ();
 sg13g2_decap_4 FILLER_34_1072 ();
 sg13g2_fill_2 FILLER_34_1112 ();
 sg13g2_decap_8 FILLER_34_1119 ();
 sg13g2_fill_1 FILLER_34_1126 ();
 sg13g2_fill_2 FILLER_34_1132 ();
 sg13g2_fill_2 FILLER_34_1145 ();
 sg13g2_fill_1 FILLER_34_1153 ();
 sg13g2_fill_2 FILLER_34_1168 ();
 sg13g2_fill_1 FILLER_34_1262 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_22 ();
 sg13g2_fill_1 FILLER_35_70 ();
 sg13g2_fill_1 FILLER_35_79 ();
 sg13g2_fill_2 FILLER_35_270 ();
 sg13g2_fill_2 FILLER_35_298 ();
 sg13g2_fill_1 FILLER_35_300 ();
 sg13g2_fill_2 FILLER_35_337 ();
 sg13g2_fill_1 FILLER_35_370 ();
 sg13g2_fill_2 FILLER_35_380 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_409 ();
 sg13g2_decap_4 FILLER_35_416 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_fill_2 FILLER_35_443 ();
 sg13g2_fill_1 FILLER_35_485 ();
 sg13g2_decap_8 FILLER_35_500 ();
 sg13g2_decap_8 FILLER_35_507 ();
 sg13g2_decap_4 FILLER_35_514 ();
 sg13g2_fill_1 FILLER_35_518 ();
 sg13g2_fill_2 FILLER_35_524 ();
 sg13g2_fill_1 FILLER_35_536 ();
 sg13g2_fill_1 FILLER_35_558 ();
 sg13g2_fill_2 FILLER_35_582 ();
 sg13g2_decap_8 FILLER_35_599 ();
 sg13g2_fill_2 FILLER_35_606 ();
 sg13g2_decap_8 FILLER_35_612 ();
 sg13g2_fill_2 FILLER_35_619 ();
 sg13g2_fill_2 FILLER_35_631 ();
 sg13g2_decap_4 FILLER_35_704 ();
 sg13g2_fill_1 FILLER_35_732 ();
 sg13g2_decap_8 FILLER_35_750 ();
 sg13g2_fill_1 FILLER_35_775 ();
 sg13g2_decap_8 FILLER_35_780 ();
 sg13g2_decap_8 FILLER_35_787 ();
 sg13g2_decap_4 FILLER_35_794 ();
 sg13g2_fill_1 FILLER_35_798 ();
 sg13g2_fill_2 FILLER_35_803 ();
 sg13g2_decap_8 FILLER_35_856 ();
 sg13g2_decap_4 FILLER_35_872 ();
 sg13g2_fill_2 FILLER_35_876 ();
 sg13g2_decap_8 FILLER_35_883 ();
 sg13g2_decap_8 FILLER_35_890 ();
 sg13g2_fill_1 FILLER_35_897 ();
 sg13g2_fill_2 FILLER_35_907 ();
 sg13g2_fill_1 FILLER_35_909 ();
 sg13g2_fill_2 FILLER_35_987 ();
 sg13g2_fill_2 FILLER_35_996 ();
 sg13g2_fill_1 FILLER_35_998 ();
 sg13g2_fill_2 FILLER_35_1008 ();
 sg13g2_fill_1 FILLER_35_1010 ();
 sg13g2_fill_2 FILLER_35_1015 ();
 sg13g2_fill_2 FILLER_35_1030 ();
 sg13g2_fill_1 FILLER_35_1041 ();
 sg13g2_fill_1 FILLER_35_1051 ();
 sg13g2_decap_4 FILLER_35_1078 ();
 sg13g2_fill_1 FILLER_35_1082 ();
 sg13g2_fill_2 FILLER_35_1095 ();
 sg13g2_decap_8 FILLER_35_1116 ();
 sg13g2_fill_1 FILLER_35_1123 ();
 sg13g2_fill_2 FILLER_35_1134 ();
 sg13g2_fill_1 FILLER_35_1136 ();
 sg13g2_fill_2 FILLER_35_1147 ();
 sg13g2_fill_1 FILLER_35_1149 ();
 sg13g2_fill_2 FILLER_35_1175 ();
 sg13g2_fill_1 FILLER_35_1177 ();
 sg13g2_fill_2 FILLER_35_1194 ();
 sg13g2_fill_2 FILLER_35_1226 ();
 sg13g2_fill_1 FILLER_35_1228 ();
 sg13g2_fill_2 FILLER_35_1259 ();
 sg13g2_fill_2 FILLER_35_1287 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_39 ();
 sg13g2_fill_2 FILLER_36_73 ();
 sg13g2_fill_1 FILLER_36_106 ();
 sg13g2_fill_1 FILLER_36_120 ();
 sg13g2_fill_2 FILLER_36_144 ();
 sg13g2_fill_2 FILLER_36_259 ();
 sg13g2_fill_2 FILLER_36_287 ();
 sg13g2_fill_2 FILLER_36_302 ();
 sg13g2_fill_1 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_325 ();
 sg13g2_fill_1 FILLER_36_364 ();
 sg13g2_fill_1 FILLER_36_384 ();
 sg13g2_fill_1 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_437 ();
 sg13g2_fill_1 FILLER_36_439 ();
 sg13g2_fill_2 FILLER_36_469 ();
 sg13g2_fill_2 FILLER_36_489 ();
 sg13g2_fill_1 FILLER_36_496 ();
 sg13g2_decap_4 FILLER_36_507 ();
 sg13g2_decap_8 FILLER_36_516 ();
 sg13g2_fill_2 FILLER_36_531 ();
 sg13g2_fill_1 FILLER_36_533 ();
 sg13g2_decap_4 FILLER_36_590 ();
 sg13g2_fill_2 FILLER_36_631 ();
 sg13g2_fill_1 FILLER_36_667 ();
 sg13g2_fill_1 FILLER_36_676 ();
 sg13g2_fill_2 FILLER_36_685 ();
 sg13g2_decap_8 FILLER_36_744 ();
 sg13g2_decap_8 FILLER_36_751 ();
 sg13g2_decap_4 FILLER_36_758 ();
 sg13g2_fill_1 FILLER_36_762 ();
 sg13g2_decap_8 FILLER_36_786 ();
 sg13g2_decap_4 FILLER_36_793 ();
 sg13g2_fill_1 FILLER_36_797 ();
 sg13g2_decap_4 FILLER_36_803 ();
 sg13g2_fill_2 FILLER_36_807 ();
 sg13g2_fill_2 FILLER_36_825 ();
 sg13g2_fill_2 FILLER_36_878 ();
 sg13g2_fill_1 FILLER_36_880 ();
 sg13g2_fill_1 FILLER_36_926 ();
 sg13g2_decap_4 FILLER_36_947 ();
 sg13g2_fill_2 FILLER_36_955 ();
 sg13g2_fill_1 FILLER_36_973 ();
 sg13g2_fill_2 FILLER_36_983 ();
 sg13g2_fill_1 FILLER_36_991 ();
 sg13g2_fill_1 FILLER_36_1004 ();
 sg13g2_fill_2 FILLER_36_1031 ();
 sg13g2_fill_2 FILLER_36_1044 ();
 sg13g2_fill_1 FILLER_36_1046 ();
 sg13g2_fill_2 FILLER_36_1056 ();
 sg13g2_fill_2 FILLER_36_1071 ();
 sg13g2_fill_1 FILLER_36_1073 ();
 sg13g2_decap_8 FILLER_36_1085 ();
 sg13g2_decap_4 FILLER_36_1092 ();
 sg13g2_fill_2 FILLER_36_1096 ();
 sg13g2_decap_8 FILLER_36_1145 ();
 sg13g2_decap_4 FILLER_36_1152 ();
 sg13g2_fill_1 FILLER_36_1206 ();
 sg13g2_fill_2 FILLER_36_1211 ();
 sg13g2_fill_2 FILLER_36_1243 ();
 sg13g2_fill_2 FILLER_36_1280 ();
 sg13g2_fill_2 FILLER_36_1312 ();
 sg13g2_fill_1 FILLER_36_1314 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_16 ();
 sg13g2_decap_8 FILLER_37_26 ();
 sg13g2_decap_4 FILLER_37_33 ();
 sg13g2_decap_4 FILLER_37_40 ();
 sg13g2_fill_2 FILLER_37_44 ();
 sg13g2_decap_4 FILLER_37_55 ();
 sg13g2_decap_4 FILLER_37_72 ();
 sg13g2_fill_2 FILLER_37_84 ();
 sg13g2_fill_2 FILLER_37_138 ();
 sg13g2_fill_1 FILLER_37_171 ();
 sg13g2_fill_2 FILLER_37_234 ();
 sg13g2_fill_1 FILLER_37_326 ();
 sg13g2_fill_1 FILLER_37_351 ();
 sg13g2_fill_2 FILLER_37_357 ();
 sg13g2_fill_1 FILLER_37_395 ();
 sg13g2_fill_1 FILLER_37_427 ();
 sg13g2_fill_1 FILLER_37_442 ();
 sg13g2_decap_4 FILLER_37_493 ();
 sg13g2_fill_2 FILLER_37_501 ();
 sg13g2_fill_1 FILLER_37_503 ();
 sg13g2_fill_1 FILLER_37_537 ();
 sg13g2_fill_2 FILLER_37_585 ();
 sg13g2_decap_4 FILLER_37_612 ();
 sg13g2_fill_1 FILLER_37_616 ();
 sg13g2_decap_8 FILLER_37_622 ();
 sg13g2_fill_1 FILLER_37_629 ();
 sg13g2_decap_8 FILLER_37_693 ();
 sg13g2_fill_2 FILLER_37_700 ();
 sg13g2_fill_1 FILLER_37_702 ();
 sg13g2_decap_4 FILLER_37_707 ();
 sg13g2_fill_1 FILLER_37_730 ();
 sg13g2_decap_8 FILLER_37_739 ();
 sg13g2_fill_1 FILLER_37_746 ();
 sg13g2_fill_2 FILLER_37_773 ();
 sg13g2_fill_1 FILLER_37_780 ();
 sg13g2_decap_4 FILLER_37_813 ();
 sg13g2_fill_1 FILLER_37_817 ();
 sg13g2_fill_2 FILLER_37_837 ();
 sg13g2_fill_1 FILLER_37_839 ();
 sg13g2_fill_2 FILLER_37_930 ();
 sg13g2_fill_1 FILLER_37_932 ();
 sg13g2_decap_4 FILLER_37_943 ();
 sg13g2_fill_1 FILLER_37_966 ();
 sg13g2_decap_8 FILLER_37_990 ();
 sg13g2_decap_4 FILLER_37_997 ();
 sg13g2_decap_8 FILLER_37_1008 ();
 sg13g2_fill_1 FILLER_37_1028 ();
 sg13g2_fill_2 FILLER_37_1047 ();
 sg13g2_decap_8 FILLER_37_1057 ();
 sg13g2_fill_1 FILLER_37_1078 ();
 sg13g2_fill_1 FILLER_37_1124 ();
 sg13g2_fill_1 FILLER_37_1135 ();
 sg13g2_fill_1 FILLER_37_1151 ();
 sg13g2_decap_4 FILLER_37_1157 ();
 sg13g2_fill_1 FILLER_37_1173 ();
 sg13g2_fill_2 FILLER_37_1184 ();
 sg13g2_fill_1 FILLER_37_1186 ();
 sg13g2_fill_2 FILLER_37_1195 ();
 sg13g2_fill_2 FILLER_37_1215 ();
 sg13g2_fill_1 FILLER_37_1217 ();
 sg13g2_fill_2 FILLER_37_1231 ();
 sg13g2_fill_1 FILLER_37_1233 ();
 sg13g2_fill_1 FILLER_37_1265 ();
 sg13g2_fill_1 FILLER_37_1284 ();
 sg13g2_fill_2 FILLER_37_1294 ();
 sg13g2_fill_1 FILLER_37_1296 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_1 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_45 ();
 sg13g2_fill_2 FILLER_38_53 ();
 sg13g2_decap_4 FILLER_38_64 ();
 sg13g2_fill_1 FILLER_38_68 ();
 sg13g2_fill_2 FILLER_38_78 ();
 sg13g2_fill_1 FILLER_38_80 ();
 sg13g2_fill_2 FILLER_38_122 ();
 sg13g2_fill_2 FILLER_38_172 ();
 sg13g2_fill_1 FILLER_38_181 ();
 sg13g2_fill_2 FILLER_38_204 ();
 sg13g2_fill_1 FILLER_38_220 ();
 sg13g2_fill_1 FILLER_38_229 ();
 sg13g2_fill_2 FILLER_38_235 ();
 sg13g2_fill_1 FILLER_38_237 ();
 sg13g2_fill_2 FILLER_38_245 ();
 sg13g2_fill_1 FILLER_38_251 ();
 sg13g2_fill_1 FILLER_38_265 ();
 sg13g2_fill_1 FILLER_38_288 ();
 sg13g2_fill_1 FILLER_38_322 ();
 sg13g2_fill_1 FILLER_38_338 ();
 sg13g2_fill_1 FILLER_38_352 ();
 sg13g2_fill_1 FILLER_38_440 ();
 sg13g2_fill_2 FILLER_38_474 ();
 sg13g2_fill_2 FILLER_38_575 ();
 sg13g2_decap_4 FILLER_38_605 ();
 sg13g2_fill_2 FILLER_38_609 ();
 sg13g2_decap_8 FILLER_38_615 ();
 sg13g2_decap_8 FILLER_38_622 ();
 sg13g2_decap_8 FILLER_38_629 ();
 sg13g2_decap_8 FILLER_38_636 ();
 sg13g2_fill_1 FILLER_38_643 ();
 sg13g2_fill_2 FILLER_38_648 ();
 sg13g2_fill_1 FILLER_38_653 ();
 sg13g2_fill_1 FILLER_38_680 ();
 sg13g2_fill_2 FILLER_38_704 ();
 sg13g2_fill_1 FILLER_38_726 ();
 sg13g2_fill_2 FILLER_38_756 ();
 sg13g2_decap_8 FILLER_38_762 ();
 sg13g2_fill_1 FILLER_38_769 ();
 sg13g2_decap_8 FILLER_38_788 ();
 sg13g2_fill_2 FILLER_38_795 ();
 sg13g2_fill_1 FILLER_38_797 ();
 sg13g2_fill_1 FILLER_38_802 ();
 sg13g2_fill_1 FILLER_38_808 ();
 sg13g2_fill_2 FILLER_38_841 ();
 sg13g2_fill_1 FILLER_38_843 ();
 sg13g2_fill_2 FILLER_38_854 ();
 sg13g2_fill_1 FILLER_38_856 ();
 sg13g2_decap_8 FILLER_38_861 ();
 sg13g2_fill_2 FILLER_38_868 ();
 sg13g2_decap_4 FILLER_38_892 ();
 sg13g2_fill_1 FILLER_38_904 ();
 sg13g2_fill_1 FILLER_38_914 ();
 sg13g2_decap_8 FILLER_38_939 ();
 sg13g2_fill_2 FILLER_38_946 ();
 sg13g2_fill_2 FILLER_38_958 ();
 sg13g2_fill_2 FILLER_38_967 ();
 sg13g2_fill_1 FILLER_38_969 ();
 sg13g2_fill_1 FILLER_38_1006 ();
 sg13g2_fill_1 FILLER_38_1029 ();
 sg13g2_decap_4 FILLER_38_1036 ();
 sg13g2_fill_2 FILLER_38_1040 ();
 sg13g2_decap_8 FILLER_38_1068 ();
 sg13g2_decap_8 FILLER_38_1075 ();
 sg13g2_fill_1 FILLER_38_1082 ();
 sg13g2_fill_1 FILLER_38_1092 ();
 sg13g2_fill_1 FILLER_38_1121 ();
 sg13g2_fill_2 FILLER_38_1131 ();
 sg13g2_fill_1 FILLER_38_1133 ();
 sg13g2_fill_1 FILLER_38_1139 ();
 sg13g2_fill_2 FILLER_38_1156 ();
 sg13g2_fill_1 FILLER_38_1158 ();
 sg13g2_decap_8 FILLER_38_1175 ();
 sg13g2_decap_4 FILLER_38_1182 ();
 sg13g2_fill_2 FILLER_38_1273 ();
 sg13g2_fill_1 FILLER_38_1275 ();
 sg13g2_fill_2 FILLER_39_13 ();
 sg13g2_fill_1 FILLER_39_15 ();
 sg13g2_fill_2 FILLER_39_77 ();
 sg13g2_fill_1 FILLER_39_118 ();
 sg13g2_fill_2 FILLER_39_133 ();
 sg13g2_fill_2 FILLER_39_139 ();
 sg13g2_fill_2 FILLER_39_269 ();
 sg13g2_fill_1 FILLER_39_271 ();
 sg13g2_decap_8 FILLER_39_321 ();
 sg13g2_decap_4 FILLER_39_328 ();
 sg13g2_fill_2 FILLER_39_332 ();
 sg13g2_decap_4 FILLER_39_344 ();
 sg13g2_fill_1 FILLER_39_348 ();
 sg13g2_fill_1 FILLER_39_375 ();
 sg13g2_fill_1 FILLER_39_443 ();
 sg13g2_fill_1 FILLER_39_466 ();
 sg13g2_fill_2 FILLER_39_506 ();
 sg13g2_fill_2 FILLER_39_543 ();
 sg13g2_fill_2 FILLER_39_571 ();
 sg13g2_fill_1 FILLER_39_573 ();
 sg13g2_fill_1 FILLER_39_626 ();
 sg13g2_decap_4 FILLER_39_672 ();
 sg13g2_fill_2 FILLER_39_710 ();
 sg13g2_decap_4 FILLER_39_720 ();
 sg13g2_fill_2 FILLER_39_724 ();
 sg13g2_decap_8 FILLER_39_747 ();
 sg13g2_decap_8 FILLER_39_768 ();
 sg13g2_fill_2 FILLER_39_775 ();
 sg13g2_fill_1 FILLER_39_777 ();
 sg13g2_decap_8 FILLER_39_783 ();
 sg13g2_decap_8 FILLER_39_790 ();
 sg13g2_fill_1 FILLER_39_797 ();
 sg13g2_decap_8 FILLER_39_807 ();
 sg13g2_fill_2 FILLER_39_814 ();
 sg13g2_fill_1 FILLER_39_816 ();
 sg13g2_decap_4 FILLER_39_825 ();
 sg13g2_decap_4 FILLER_39_836 ();
 sg13g2_decap_4 FILLER_39_844 ();
 sg13g2_fill_2 FILLER_39_851 ();
 sg13g2_decap_4 FILLER_39_880 ();
 sg13g2_fill_2 FILLER_39_945 ();
 sg13g2_fill_1 FILLER_39_947 ();
 sg13g2_fill_1 FILLER_39_956 ();
 sg13g2_decap_4 FILLER_39_962 ();
 sg13g2_fill_2 FILLER_39_989 ();
 sg13g2_decap_8 FILLER_39_1037 ();
 sg13g2_decap_8 FILLER_39_1044 ();
 sg13g2_fill_2 FILLER_39_1051 ();
 sg13g2_decap_8 FILLER_39_1057 ();
 sg13g2_decap_8 FILLER_39_1064 ();
 sg13g2_decap_8 FILLER_39_1071 ();
 sg13g2_decap_8 FILLER_39_1078 ();
 sg13g2_fill_1 FILLER_39_1085 ();
 sg13g2_fill_2 FILLER_39_1129 ();
 sg13g2_fill_1 FILLER_39_1131 ();
 sg13g2_fill_1 FILLER_39_1165 ();
 sg13g2_fill_2 FILLER_39_1202 ();
 sg13g2_fill_1 FILLER_39_1256 ();
 sg13g2_fill_2 FILLER_39_1313 ();
 sg13g2_decap_4 FILLER_40_92 ();
 sg13g2_fill_2 FILLER_40_96 ();
 sg13g2_fill_2 FILLER_40_138 ();
 sg13g2_fill_1 FILLER_40_207 ();
 sg13g2_fill_2 FILLER_40_216 ();
 sg13g2_fill_2 FILLER_40_223 ();
 sg13g2_fill_2 FILLER_40_248 ();
 sg13g2_fill_1 FILLER_40_250 ();
 sg13g2_fill_2 FILLER_40_273 ();
 sg13g2_fill_1 FILLER_40_275 ();
 sg13g2_decap_4 FILLER_40_332 ();
 sg13g2_fill_2 FILLER_40_346 ();
 sg13g2_decap_8 FILLER_40_365 ();
 sg13g2_fill_2 FILLER_40_372 ();
 sg13g2_fill_1 FILLER_40_459 ();
 sg13g2_fill_1 FILLER_40_475 ();
 sg13g2_fill_2 FILLER_40_494 ();
 sg13g2_fill_2 FILLER_40_509 ();
 sg13g2_decap_4 FILLER_40_568 ();
 sg13g2_fill_1 FILLER_40_572 ();
 sg13g2_decap_4 FILLER_40_599 ();
 sg13g2_fill_1 FILLER_40_603 ();
 sg13g2_fill_2 FILLER_40_641 ();
 sg13g2_fill_2 FILLER_40_647 ();
 sg13g2_decap_4 FILLER_40_653 ();
 sg13g2_fill_1 FILLER_40_657 ();
 sg13g2_fill_2 FILLER_40_687 ();
 sg13g2_decap_4 FILLER_40_708 ();
 sg13g2_fill_1 FILLER_40_712 ();
 sg13g2_decap_8 FILLER_40_721 ();
 sg13g2_fill_2 FILLER_40_728 ();
 sg13g2_fill_1 FILLER_40_730 ();
 sg13g2_fill_2 FILLER_40_744 ();
 sg13g2_decap_4 FILLER_40_776 ();
 sg13g2_fill_2 FILLER_40_819 ();
 sg13g2_decap_8 FILLER_40_842 ();
 sg13g2_decap_8 FILLER_40_849 ();
 sg13g2_decap_4 FILLER_40_856 ();
 sg13g2_fill_1 FILLER_40_860 ();
 sg13g2_fill_1 FILLER_40_871 ();
 sg13g2_fill_2 FILLER_40_876 ();
 sg13g2_fill_1 FILLER_40_878 ();
 sg13g2_fill_2 FILLER_40_895 ();
 sg13g2_fill_1 FILLER_40_897 ();
 sg13g2_fill_1 FILLER_40_926 ();
 sg13g2_fill_1 FILLER_40_963 ();
 sg13g2_fill_1 FILLER_40_984 ();
 sg13g2_fill_2 FILLER_40_994 ();
 sg13g2_decap_4 FILLER_40_1026 ();
 sg13g2_fill_2 FILLER_40_1030 ();
 sg13g2_decap_8 FILLER_40_1054 ();
 sg13g2_decap_4 FILLER_40_1061 ();
 sg13g2_decap_8 FILLER_40_1083 ();
 sg13g2_fill_1 FILLER_40_1090 ();
 sg13g2_fill_2 FILLER_40_1127 ();
 sg13g2_fill_2 FILLER_40_1155 ();
 sg13g2_fill_1 FILLER_40_1157 ();
 sg13g2_decap_8 FILLER_40_1173 ();
 sg13g2_decap_8 FILLER_40_1180 ();
 sg13g2_fill_1 FILLER_40_1191 ();
 sg13g2_fill_2 FILLER_40_1249 ();
 sg13g2_fill_1 FILLER_40_1251 ();
 sg13g2_fill_2 FILLER_40_1265 ();
 sg13g2_fill_1 FILLER_40_1267 ();
 sg13g2_fill_2 FILLER_40_1312 ();
 sg13g2_fill_1 FILLER_40_1314 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_25 ();
 sg13g2_fill_2 FILLER_41_75 ();
 sg13g2_fill_1 FILLER_41_77 ();
 sg13g2_fill_2 FILLER_41_88 ();
 sg13g2_decap_4 FILLER_41_101 ();
 sg13g2_fill_1 FILLER_41_105 ();
 sg13g2_fill_1 FILLER_41_162 ();
 sg13g2_fill_2 FILLER_41_172 ();
 sg13g2_fill_2 FILLER_41_199 ();
 sg13g2_fill_1 FILLER_41_211 ();
 sg13g2_decap_4 FILLER_41_218 ();
 sg13g2_fill_1 FILLER_41_222 ();
 sg13g2_decap_8 FILLER_41_227 ();
 sg13g2_fill_1 FILLER_41_234 ();
 sg13g2_fill_1 FILLER_41_261 ();
 sg13g2_fill_2 FILLER_41_277 ();
 sg13g2_fill_1 FILLER_41_279 ();
 sg13g2_fill_2 FILLER_41_288 ();
 sg13g2_fill_1 FILLER_41_290 ();
 sg13g2_fill_2 FILLER_41_300 ();
 sg13g2_fill_1 FILLER_41_316 ();
 sg13g2_fill_1 FILLER_41_350 ();
 sg13g2_fill_2 FILLER_41_369 ();
 sg13g2_fill_1 FILLER_41_371 ();
 sg13g2_fill_1 FILLER_41_376 ();
 sg13g2_fill_1 FILLER_41_387 ();
 sg13g2_fill_2 FILLER_41_398 ();
 sg13g2_fill_1 FILLER_41_417 ();
 sg13g2_fill_2 FILLER_41_451 ();
 sg13g2_fill_2 FILLER_41_476 ();
 sg13g2_decap_8 FILLER_41_535 ();
 sg13g2_decap_8 FILLER_41_542 ();
 sg13g2_fill_1 FILLER_41_678 ();
 sg13g2_decap_8 FILLER_41_713 ();
 sg13g2_fill_2 FILLER_41_720 ();
 sg13g2_decap_8 FILLER_41_732 ();
 sg13g2_decap_4 FILLER_41_739 ();
 sg13g2_decap_8 FILLER_41_751 ();
 sg13g2_decap_8 FILLER_41_758 ();
 sg13g2_fill_1 FILLER_41_781 ();
 sg13g2_fill_2 FILLER_41_787 ();
 sg13g2_fill_1 FILLER_41_789 ();
 sg13g2_decap_8 FILLER_41_809 ();
 sg13g2_fill_1 FILLER_41_816 ();
 sg13g2_decap_4 FILLER_41_823 ();
 sg13g2_fill_2 FILLER_41_827 ();
 sg13g2_fill_2 FILLER_41_838 ();
 sg13g2_fill_2 FILLER_41_844 ();
 sg13g2_fill_1 FILLER_41_846 ();
 sg13g2_decap_8 FILLER_41_877 ();
 sg13g2_fill_2 FILLER_41_884 ();
 sg13g2_fill_1 FILLER_41_886 ();
 sg13g2_fill_2 FILLER_41_948 ();
 sg13g2_fill_1 FILLER_41_950 ();
 sg13g2_decap_8 FILLER_41_976 ();
 sg13g2_fill_2 FILLER_41_983 ();
 sg13g2_fill_1 FILLER_41_995 ();
 sg13g2_fill_2 FILLER_41_1010 ();
 sg13g2_fill_2 FILLER_41_1087 ();
 sg13g2_fill_2 FILLER_41_1097 ();
 sg13g2_fill_1 FILLER_41_1103 ();
 sg13g2_decap_8 FILLER_41_1114 ();
 sg13g2_decap_4 FILLER_41_1121 ();
 sg13g2_decap_8 FILLER_41_1154 ();
 sg13g2_fill_1 FILLER_41_1161 ();
 sg13g2_fill_2 FILLER_41_1166 ();
 sg13g2_fill_1 FILLER_41_1168 ();
 sg13g2_fill_1 FILLER_41_1221 ();
 sg13g2_fill_2 FILLER_41_1287 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_30 ();
 sg13g2_fill_1 FILLER_42_34 ();
 sg13g2_fill_1 FILLER_42_44 ();
 sg13g2_fill_2 FILLER_42_71 ();
 sg13g2_fill_2 FILLER_42_196 ();
 sg13g2_fill_1 FILLER_42_198 ();
 sg13g2_fill_2 FILLER_42_250 ();
 sg13g2_fill_1 FILLER_42_272 ();
 sg13g2_fill_2 FILLER_42_289 ();
 sg13g2_fill_1 FILLER_42_291 ();
 sg13g2_fill_2 FILLER_42_296 ();
 sg13g2_fill_2 FILLER_42_307 ();
 sg13g2_fill_1 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_354 ();
 sg13g2_fill_1 FILLER_42_361 ();
 sg13g2_fill_2 FILLER_42_450 ();
 sg13g2_fill_1 FILLER_42_471 ();
 sg13g2_fill_2 FILLER_42_476 ();
 sg13g2_fill_1 FILLER_42_511 ();
 sg13g2_fill_2 FILLER_42_554 ();
 sg13g2_fill_1 FILLER_42_556 ();
 sg13g2_decap_8 FILLER_42_570 ();
 sg13g2_fill_2 FILLER_42_577 ();
 sg13g2_fill_2 FILLER_42_583 ();
 sg13g2_fill_1 FILLER_42_585 ();
 sg13g2_decap_4 FILLER_42_590 ();
 sg13g2_fill_1 FILLER_42_610 ();
 sg13g2_fill_2 FILLER_42_620 ();
 sg13g2_fill_1 FILLER_42_639 ();
 sg13g2_fill_2 FILLER_42_659 ();
 sg13g2_fill_1 FILLER_42_661 ();
 sg13g2_fill_2 FILLER_42_670 ();
 sg13g2_decap_8 FILLER_42_725 ();
 sg13g2_decap_4 FILLER_42_732 ();
 sg13g2_fill_2 FILLER_42_781 ();
 sg13g2_fill_2 FILLER_42_800 ();
 sg13g2_fill_1 FILLER_42_802 ();
 sg13g2_decap_8 FILLER_42_868 ();
 sg13g2_decap_8 FILLER_42_875 ();
 sg13g2_fill_1 FILLER_42_901 ();
 sg13g2_fill_2 FILLER_42_965 ();
 sg13g2_fill_2 FILLER_42_1016 ();
 sg13g2_fill_1 FILLER_42_1018 ();
 sg13g2_decap_4 FILLER_42_1027 ();
 sg13g2_fill_1 FILLER_42_1031 ();
 sg13g2_fill_1 FILLER_42_1055 ();
 sg13g2_decap_4 FILLER_42_1082 ();
 sg13g2_fill_1 FILLER_42_1150 ();
 sg13g2_fill_1 FILLER_42_1190 ();
 sg13g2_fill_1 FILLER_42_1226 ();
 sg13g2_fill_2 FILLER_42_1257 ();
 sg13g2_fill_1 FILLER_42_1259 ();
 sg13g2_fill_2 FILLER_42_1286 ();
 sg13g2_fill_1 FILLER_42_1288 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_21 ();
 sg13g2_fill_2 FILLER_43_31 ();
 sg13g2_fill_2 FILLER_43_76 ();
 sg13g2_fill_1 FILLER_43_78 ();
 sg13g2_fill_2 FILLER_43_132 ();
 sg13g2_fill_2 FILLER_43_150 ();
 sg13g2_fill_2 FILLER_43_174 ();
 sg13g2_fill_2 FILLER_43_270 ();
 sg13g2_decap_8 FILLER_43_317 ();
 sg13g2_decap_4 FILLER_43_324 ();
 sg13g2_decap_8 FILLER_43_349 ();
 sg13g2_fill_2 FILLER_43_356 ();
 sg13g2_decap_8 FILLER_43_362 ();
 sg13g2_decap_8 FILLER_43_369 ();
 sg13g2_decap_8 FILLER_43_376 ();
 sg13g2_fill_2 FILLER_43_383 ();
 sg13g2_fill_2 FILLER_43_416 ();
 sg13g2_fill_1 FILLER_43_418 ();
 sg13g2_fill_1 FILLER_43_479 ();
 sg13g2_decap_8 FILLER_43_492 ();
 sg13g2_decap_8 FILLER_43_499 ();
 sg13g2_decap_8 FILLER_43_512 ();
 sg13g2_fill_2 FILLER_43_519 ();
 sg13g2_decap_8 FILLER_43_536 ();
 sg13g2_fill_2 FILLER_43_543 ();
 sg13g2_decap_8 FILLER_43_549 ();
 sg13g2_fill_2 FILLER_43_556 ();
 sg13g2_decap_4 FILLER_43_570 ();
 sg13g2_fill_2 FILLER_43_587 ();
 sg13g2_fill_1 FILLER_43_614 ();
 sg13g2_decap_4 FILLER_43_651 ();
 sg13g2_fill_1 FILLER_43_655 ();
 sg13g2_fill_1 FILLER_43_685 ();
 sg13g2_fill_2 FILLER_43_691 ();
 sg13g2_fill_1 FILLER_43_735 ();
 sg13g2_decap_4 FILLER_43_759 ();
 sg13g2_fill_2 FILLER_43_763 ();
 sg13g2_fill_1 FILLER_43_769 ();
 sg13g2_fill_1 FILLER_43_778 ();
 sg13g2_fill_2 FILLER_43_789 ();
 sg13g2_fill_2 FILLER_43_797 ();
 sg13g2_fill_1 FILLER_43_819 ();
 sg13g2_fill_2 FILLER_43_823 ();
 sg13g2_fill_1 FILLER_43_825 ();
 sg13g2_fill_2 FILLER_43_835 ();
 sg13g2_fill_1 FILLER_43_926 ();
 sg13g2_decap_8 FILLER_43_961 ();
 sg13g2_fill_2 FILLER_43_968 ();
 sg13g2_fill_1 FILLER_43_970 ();
 sg13g2_fill_1 FILLER_43_984 ();
 sg13g2_fill_2 FILLER_43_994 ();
 sg13g2_fill_1 FILLER_43_1001 ();
 sg13g2_decap_4 FILLER_43_1025 ();
 sg13g2_fill_2 FILLER_43_1042 ();
 sg13g2_fill_1 FILLER_43_1044 ();
 sg13g2_decap_4 FILLER_43_1062 ();
 sg13g2_decap_8 FILLER_43_1070 ();
 sg13g2_fill_2 FILLER_43_1077 ();
 sg13g2_fill_2 FILLER_43_1120 ();
 sg13g2_fill_1 FILLER_43_1130 ();
 sg13g2_fill_2 FILLER_43_1168 ();
 sg13g2_fill_1 FILLER_43_1170 ();
 sg13g2_fill_1 FILLER_43_1175 ();
 sg13g2_fill_2 FILLER_43_1242 ();
 sg13g2_fill_1 FILLER_43_1244 ();
 sg13g2_fill_1 FILLER_43_1280 ();
 sg13g2_fill_2 FILLER_43_1312 ();
 sg13g2_fill_1 FILLER_43_1314 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_30 ();
 sg13g2_fill_2 FILLER_44_252 ();
 sg13g2_fill_2 FILLER_44_274 ();
 sg13g2_fill_1 FILLER_44_291 ();
 sg13g2_fill_2 FILLER_44_360 ();
 sg13g2_fill_1 FILLER_44_366 ();
 sg13g2_decap_8 FILLER_44_383 ();
 sg13g2_fill_2 FILLER_44_390 ();
 sg13g2_fill_1 FILLER_44_392 ();
 sg13g2_fill_2 FILLER_44_405 ();
 sg13g2_fill_1 FILLER_44_407 ();
 sg13g2_fill_1 FILLER_44_412 ();
 sg13g2_fill_2 FILLER_44_453 ();
 sg13g2_fill_2 FILLER_44_495 ();
 sg13g2_fill_1 FILLER_44_569 ();
 sg13g2_fill_1 FILLER_44_605 ();
 sg13g2_fill_2 FILLER_44_620 ();
 sg13g2_fill_2 FILLER_44_630 ();
 sg13g2_fill_1 FILLER_44_632 ();
 sg13g2_fill_1 FILLER_44_708 ();
 sg13g2_fill_2 FILLER_44_717 ();
 sg13g2_decap_8 FILLER_44_745 ();
 sg13g2_fill_1 FILLER_44_752 ();
 sg13g2_decap_4 FILLER_44_808 ();
 sg13g2_fill_1 FILLER_44_812 ();
 sg13g2_fill_1 FILLER_44_823 ();
 sg13g2_fill_2 FILLER_44_844 ();
 sg13g2_fill_2 FILLER_44_875 ();
 sg13g2_fill_2 FILLER_44_900 ();
 sg13g2_decap_8 FILLER_44_969 ();
 sg13g2_decap_8 FILLER_44_976 ();
 sg13g2_fill_1 FILLER_44_983 ();
 sg13g2_fill_1 FILLER_44_996 ();
 sg13g2_decap_8 FILLER_44_1005 ();
 sg13g2_fill_1 FILLER_44_1012 ();
 sg13g2_fill_2 FILLER_44_1017 ();
 sg13g2_fill_1 FILLER_44_1019 ();
 sg13g2_decap_8 FILLER_44_1025 ();
 sg13g2_decap_4 FILLER_44_1032 ();
 sg13g2_fill_1 FILLER_44_1036 ();
 sg13g2_fill_2 FILLER_44_1102 ();
 sg13g2_fill_1 FILLER_44_1132 ();
 sg13g2_fill_1 FILLER_44_1195 ();
 sg13g2_fill_2 FILLER_44_1200 ();
 sg13g2_fill_1 FILLER_44_1202 ();
 sg13g2_fill_2 FILLER_44_1229 ();
 sg13g2_fill_1 FILLER_44_1288 ();
 sg13g2_fill_2 FILLER_45_33 ();
 sg13g2_fill_2 FILLER_45_49 ();
 sg13g2_fill_1 FILLER_45_149 ();
 sg13g2_fill_1 FILLER_45_177 ();
 sg13g2_fill_2 FILLER_45_202 ();
 sg13g2_fill_1 FILLER_45_235 ();
 sg13g2_fill_1 FILLER_45_365 ();
 sg13g2_fill_2 FILLER_45_389 ();
 sg13g2_fill_1 FILLER_45_402 ();
 sg13g2_fill_1 FILLER_45_413 ();
 sg13g2_fill_1 FILLER_45_436 ();
 sg13g2_fill_2 FILLER_45_463 ();
 sg13g2_fill_2 FILLER_45_474 ();
 sg13g2_fill_1 FILLER_45_476 ();
 sg13g2_fill_2 FILLER_45_519 ();
 sg13g2_fill_1 FILLER_45_537 ();
 sg13g2_decap_4 FILLER_45_548 ();
 sg13g2_fill_1 FILLER_45_576 ();
 sg13g2_fill_1 FILLER_45_596 ();
 sg13g2_fill_1 FILLER_45_616 ();
 sg13g2_decap_8 FILLER_45_657 ();
 sg13g2_decap_8 FILLER_45_705 ();
 sg13g2_decap_4 FILLER_45_712 ();
 sg13g2_fill_2 FILLER_45_716 ();
 sg13g2_fill_1 FILLER_45_779 ();
 sg13g2_fill_1 FILLER_45_799 ();
 sg13g2_fill_1 FILLER_45_812 ();
 sg13g2_fill_1 FILLER_45_820 ();
 sg13g2_fill_2 FILLER_45_833 ();
 sg13g2_fill_1 FILLER_45_849 ();
 sg13g2_fill_1 FILLER_45_855 ();
 sg13g2_fill_2 FILLER_45_865 ();
 sg13g2_fill_1 FILLER_45_867 ();
 sg13g2_fill_1 FILLER_45_876 ();
 sg13g2_fill_1 FILLER_45_884 ();
 sg13g2_fill_2 FILLER_45_951 ();
 sg13g2_fill_1 FILLER_45_953 ();
 sg13g2_decap_8 FILLER_45_963 ();
 sg13g2_decap_4 FILLER_45_970 ();
 sg13g2_fill_2 FILLER_45_974 ();
 sg13g2_fill_2 FILLER_45_986 ();
 sg13g2_fill_1 FILLER_45_1014 ();
 sg13g2_fill_2 FILLER_45_1020 ();
 sg13g2_fill_2 FILLER_45_1042 ();
 sg13g2_fill_1 FILLER_45_1044 ();
 sg13g2_fill_2 FILLER_45_1095 ();
 sg13g2_fill_2 FILLER_45_1137 ();
 sg13g2_fill_2 FILLER_45_1257 ();
 sg13g2_fill_1 FILLER_45_1259 ();
 sg13g2_fill_2 FILLER_45_1312 ();
 sg13g2_fill_1 FILLER_45_1314 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_9 ();
 sg13g2_fill_2 FILLER_46_65 ();
 sg13g2_fill_1 FILLER_46_76 ();
 sg13g2_fill_2 FILLER_46_85 ();
 sg13g2_fill_1 FILLER_46_100 ();
 sg13g2_fill_2 FILLER_46_117 ();
 sg13g2_fill_1 FILLER_46_119 ();
 sg13g2_fill_2 FILLER_46_127 ();
 sg13g2_decap_8 FILLER_46_155 ();
 sg13g2_fill_1 FILLER_46_162 ();
 sg13g2_fill_2 FILLER_46_189 ();
 sg13g2_fill_1 FILLER_46_191 ();
 sg13g2_fill_1 FILLER_46_253 ();
 sg13g2_fill_2 FILLER_46_259 ();
 sg13g2_fill_1 FILLER_46_309 ();
 sg13g2_decap_8 FILLER_46_314 ();
 sg13g2_decap_8 FILLER_46_321 ();
 sg13g2_fill_2 FILLER_46_328 ();
 sg13g2_fill_1 FILLER_46_330 ();
 sg13g2_fill_2 FILLER_46_335 ();
 sg13g2_fill_1 FILLER_46_359 ();
 sg13g2_fill_2 FILLER_46_373 ();
 sg13g2_decap_8 FILLER_46_384 ();
 sg13g2_decap_4 FILLER_46_391 ();
 sg13g2_fill_1 FILLER_46_395 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_fill_2 FILLER_46_417 ();
 sg13g2_fill_1 FILLER_46_419 ();
 sg13g2_fill_1 FILLER_46_446 ();
 sg13g2_fill_2 FILLER_46_454 ();
 sg13g2_fill_1 FILLER_46_456 ();
 sg13g2_fill_2 FILLER_46_501 ();
 sg13g2_fill_2 FILLER_46_529 ();
 sg13g2_decap_8 FILLER_46_554 ();
 sg13g2_decap_8 FILLER_46_561 ();
 sg13g2_fill_2 FILLER_46_573 ();
 sg13g2_fill_1 FILLER_46_601 ();
 sg13g2_fill_1 FILLER_46_640 ();
 sg13g2_decap_8 FILLER_46_689 ();
 sg13g2_decap_4 FILLER_46_696 ();
 sg13g2_fill_2 FILLER_46_700 ();
 sg13g2_fill_1 FILLER_46_706 ();
 sg13g2_decap_4 FILLER_46_733 ();
 sg13g2_fill_2 FILLER_46_737 ();
 sg13g2_decap_8 FILLER_46_743 ();
 sg13g2_decap_4 FILLER_46_750 ();
 sg13g2_fill_2 FILLER_46_754 ();
 sg13g2_fill_2 FILLER_46_774 ();
 sg13g2_fill_1 FILLER_46_806 ();
 sg13g2_decap_8 FILLER_46_821 ();
 sg13g2_fill_1 FILLER_46_828 ();
 sg13g2_decap_8 FILLER_46_833 ();
 sg13g2_fill_1 FILLER_46_854 ();
 sg13g2_fill_1 FILLER_46_881 ();
 sg13g2_decap_8 FILLER_46_886 ();
 sg13g2_fill_1 FILLER_46_893 ();
 sg13g2_fill_2 FILLER_46_898 ();
 sg13g2_fill_1 FILLER_46_900 ();
 sg13g2_fill_1 FILLER_46_905 ();
 sg13g2_fill_2 FILLER_46_931 ();
 sg13g2_fill_1 FILLER_46_933 ();
 sg13g2_fill_1 FILLER_46_957 ();
 sg13g2_fill_2 FILLER_46_963 ();
 sg13g2_fill_1 FILLER_46_965 ();
 sg13g2_decap_8 FILLER_46_1015 ();
 sg13g2_fill_1 FILLER_46_1022 ();
 sg13g2_fill_2 FILLER_46_1027 ();
 sg13g2_fill_1 FILLER_46_1029 ();
 sg13g2_fill_1 FILLER_46_1045 ();
 sg13g2_fill_2 FILLER_46_1076 ();
 sg13g2_fill_2 FILLER_46_1134 ();
 sg13g2_decap_8 FILLER_46_1151 ();
 sg13g2_fill_2 FILLER_46_1158 ();
 sg13g2_decap_4 FILLER_46_1164 ();
 sg13g2_fill_1 FILLER_46_1216 ();
 sg13g2_fill_1 FILLER_46_1226 ();
 sg13g2_fill_2 FILLER_46_1240 ();
 sg13g2_fill_1 FILLER_46_1242 ();
 sg13g2_fill_2 FILLER_46_1278 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_2 ();
 sg13g2_fill_1 FILLER_47_29 ();
 sg13g2_decap_8 FILLER_47_34 ();
 sg13g2_fill_1 FILLER_47_41 ();
 sg13g2_fill_2 FILLER_47_68 ();
 sg13g2_decap_4 FILLER_47_96 ();
 sg13g2_fill_2 FILLER_47_126 ();
 sg13g2_decap_4 FILLER_47_166 ();
 sg13g2_fill_2 FILLER_47_194 ();
 sg13g2_fill_1 FILLER_47_250 ();
 sg13g2_fill_2 FILLER_47_274 ();
 sg13g2_fill_1 FILLER_47_375 ();
 sg13g2_fill_2 FILLER_47_388 ();
 sg13g2_fill_2 FILLER_47_401 ();
 sg13g2_fill_1 FILLER_47_403 ();
 sg13g2_fill_1 FILLER_47_440 ();
 sg13g2_decap_4 FILLER_47_450 ();
 sg13g2_fill_1 FILLER_47_454 ();
 sg13g2_fill_1 FILLER_47_465 ();
 sg13g2_fill_1 FILLER_47_510 ();
 sg13g2_fill_1 FILLER_47_515 ();
 sg13g2_fill_2 FILLER_47_531 ();
 sg13g2_fill_1 FILLER_47_533 ();
 sg13g2_decap_4 FILLER_47_545 ();
 sg13g2_fill_2 FILLER_47_560 ();
 sg13g2_decap_8 FILLER_47_617 ();
 sg13g2_fill_1 FILLER_47_624 ();
 sg13g2_decap_8 FILLER_47_631 ();
 sg13g2_fill_2 FILLER_47_638 ();
 sg13g2_decap_8 FILLER_47_663 ();
 sg13g2_decap_4 FILLER_47_670 ();
 sg13g2_fill_1 FILLER_47_674 ();
 sg13g2_fill_2 FILLER_47_701 ();
 sg13g2_decap_8 FILLER_47_721 ();
 sg13g2_fill_1 FILLER_47_728 ();
 sg13g2_decap_4 FILLER_47_760 ();
 sg13g2_fill_1 FILLER_47_764 ();
 sg13g2_fill_1 FILLER_47_783 ();
 sg13g2_fill_2 FILLER_47_818 ();
 sg13g2_fill_1 FILLER_47_820 ();
 sg13g2_decap_4 FILLER_47_860 ();
 sg13g2_fill_2 FILLER_47_864 ();
 sg13g2_fill_1 FILLER_47_874 ();
 sg13g2_decap_4 FILLER_47_879 ();
 sg13g2_decap_4 FILLER_47_909 ();
 sg13g2_fill_2 FILLER_47_921 ();
 sg13g2_fill_1 FILLER_47_923 ();
 sg13g2_decap_4 FILLER_47_953 ();
 sg13g2_decap_4 FILLER_47_968 ();
 sg13g2_fill_1 FILLER_47_984 ();
 sg13g2_fill_2 FILLER_47_1001 ();
 sg13g2_fill_1 FILLER_47_1028 ();
 sg13g2_decap_8 FILLER_47_1049 ();
 sg13g2_fill_2 FILLER_47_1056 ();
 sg13g2_fill_1 FILLER_47_1058 ();
 sg13g2_decap_4 FILLER_47_1067 ();
 sg13g2_fill_2 FILLER_47_1071 ();
 sg13g2_decap_4 FILLER_47_1081 ();
 sg13g2_fill_2 FILLER_47_1085 ();
 sg13g2_fill_2 FILLER_47_1139 ();
 sg13g2_fill_1 FILLER_47_1141 ();
 sg13g2_fill_2 FILLER_47_1199 ();
 sg13g2_fill_1 FILLER_47_1314 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_29 ();
 sg13g2_fill_1 FILLER_48_31 ();
 sg13g2_fill_2 FILLER_48_41 ();
 sg13g2_fill_2 FILLER_48_69 ();
 sg13g2_fill_2 FILLER_48_97 ();
 sg13g2_fill_2 FILLER_48_172 ();
 sg13g2_fill_1 FILLER_48_267 ();
 sg13g2_fill_1 FILLER_48_273 ();
 sg13g2_fill_1 FILLER_48_298 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_333 ();
 sg13g2_decap_4 FILLER_48_340 ();
 sg13g2_fill_1 FILLER_48_344 ();
 sg13g2_fill_2 FILLER_48_358 ();
 sg13g2_fill_1 FILLER_48_360 ();
 sg13g2_decap_8 FILLER_48_366 ();
 sg13g2_decap_4 FILLER_48_373 ();
 sg13g2_fill_2 FILLER_48_377 ();
 sg13g2_decap_4 FILLER_48_385 ();
 sg13g2_fill_2 FILLER_48_400 ();
 sg13g2_fill_1 FILLER_48_402 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_fill_2 FILLER_48_428 ();
 sg13g2_fill_1 FILLER_48_430 ();
 sg13g2_fill_1 FILLER_48_524 ();
 sg13g2_fill_2 FILLER_48_532 ();
 sg13g2_fill_2 FILLER_48_545 ();
 sg13g2_fill_1 FILLER_48_547 ();
 sg13g2_decap_8 FILLER_48_566 ();
 sg13g2_fill_1 FILLER_48_579 ();
 sg13g2_fill_2 FILLER_48_602 ();
 sg13g2_fill_2 FILLER_48_609 ();
 sg13g2_fill_1 FILLER_48_611 ();
 sg13g2_fill_1 FILLER_48_616 ();
 sg13g2_decap_4 FILLER_48_680 ();
 sg13g2_fill_2 FILLER_48_684 ();
 sg13g2_decap_4 FILLER_48_690 ();
 sg13g2_fill_2 FILLER_48_694 ();
 sg13g2_fill_2 FILLER_48_723 ();
 sg13g2_fill_1 FILLER_48_730 ();
 sg13g2_fill_1 FILLER_48_773 ();
 sg13g2_fill_2 FILLER_48_816 ();
 sg13g2_fill_1 FILLER_48_818 ();
 sg13g2_fill_2 FILLER_48_827 ();
 sg13g2_fill_1 FILLER_48_829 ();
 sg13g2_decap_4 FILLER_48_853 ();
 sg13g2_fill_2 FILLER_48_857 ();
 sg13g2_fill_1 FILLER_48_885 ();
 sg13g2_fill_2 FILLER_48_903 ();
 sg13g2_fill_2 FILLER_48_954 ();
 sg13g2_fill_2 FILLER_48_974 ();
 sg13g2_fill_1 FILLER_48_976 ();
 sg13g2_fill_1 FILLER_48_986 ();
 sg13g2_fill_2 FILLER_48_991 ();
 sg13g2_fill_1 FILLER_48_993 ();
 sg13g2_decap_8 FILLER_48_999 ();
 sg13g2_decap_8 FILLER_48_1006 ();
 sg13g2_fill_1 FILLER_48_1029 ();
 sg13g2_fill_2 FILLER_48_1040 ();
 sg13g2_fill_2 FILLER_48_1046 ();
 sg13g2_fill_2 FILLER_48_1053 ();
 sg13g2_fill_1 FILLER_48_1055 ();
 sg13g2_fill_1 FILLER_48_1061 ();
 sg13g2_fill_1 FILLER_48_1075 ();
 sg13g2_fill_1 FILLER_48_1084 ();
 sg13g2_fill_2 FILLER_48_1090 ();
 sg13g2_fill_2 FILLER_48_1108 ();
 sg13g2_fill_2 FILLER_48_1136 ();
 sg13g2_fill_1 FILLER_48_1138 ();
 sg13g2_decap_8 FILLER_48_1144 ();
 sg13g2_fill_2 FILLER_48_1185 ();
 sg13g2_fill_1 FILLER_48_1187 ();
 sg13g2_fill_1 FILLER_48_1250 ();
 sg13g2_fill_2 FILLER_48_1286 ();
 sg13g2_fill_1 FILLER_48_1288 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_16 ();
 sg13g2_fill_1 FILLER_49_18 ();
 sg13g2_fill_1 FILLER_49_111 ();
 sg13g2_decap_4 FILLER_49_156 ();
 sg13g2_fill_1 FILLER_49_160 ();
 sg13g2_fill_1 FILLER_49_210 ();
 sg13g2_fill_2 FILLER_49_220 ();
 sg13g2_fill_1 FILLER_49_227 ();
 sg13g2_fill_1 FILLER_49_386 ();
 sg13g2_fill_2 FILLER_49_401 ();
 sg13g2_fill_1 FILLER_49_403 ();
 sg13g2_fill_1 FILLER_49_413 ();
 sg13g2_fill_2 FILLER_49_434 ();
 sg13g2_fill_1 FILLER_49_450 ();
 sg13g2_fill_2 FILLER_49_460 ();
 sg13g2_fill_1 FILLER_49_472 ();
 sg13g2_fill_2 FILLER_49_478 ();
 sg13g2_fill_2 FILLER_49_506 ();
 sg13g2_fill_2 FILLER_49_541 ();
 sg13g2_fill_1 FILLER_49_561 ();
 sg13g2_fill_1 FILLER_49_578 ();
 sg13g2_fill_1 FILLER_49_592 ();
 sg13g2_decap_4 FILLER_49_597 ();
 sg13g2_fill_1 FILLER_49_633 ();
 sg13g2_fill_2 FILLER_49_658 ();
 sg13g2_fill_2 FILLER_49_686 ();
 sg13g2_fill_1 FILLER_49_688 ();
 sg13g2_fill_2 FILLER_49_749 ();
 sg13g2_decap_8 FILLER_49_761 ();
 sg13g2_decap_4 FILLER_49_768 ();
 sg13g2_decap_4 FILLER_49_777 ();
 sg13g2_fill_1 FILLER_49_831 ();
 sg13g2_fill_2 FILLER_49_875 ();
 sg13g2_decap_8 FILLER_49_922 ();
 sg13g2_fill_1 FILLER_49_938 ();
 sg13g2_fill_2 FILLER_49_949 ();
 sg13g2_fill_1 FILLER_49_974 ();
 sg13g2_fill_1 FILLER_49_989 ();
 sg13g2_fill_2 FILLER_49_1021 ();
 sg13g2_fill_1 FILLER_49_1023 ();
 sg13g2_fill_2 FILLER_49_1033 ();
 sg13g2_fill_2 FILLER_49_1068 ();
 sg13g2_fill_1 FILLER_49_1083 ();
 sg13g2_decap_4 FILLER_49_1096 ();
 sg13g2_decap_4 FILLER_49_1116 ();
 sg13g2_fill_1 FILLER_49_1124 ();
 sg13g2_fill_2 FILLER_49_1208 ();
 sg13g2_fill_1 FILLER_49_1210 ();
 sg13g2_fill_1 FILLER_49_1267 ();
 sg13g2_decap_4 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_4 ();
 sg13g2_fill_2 FILLER_50_70 ();
 sg13g2_fill_2 FILLER_50_77 ();
 sg13g2_fill_1 FILLER_50_79 ();
 sg13g2_fill_1 FILLER_50_97 ();
 sg13g2_fill_1 FILLER_50_157 ();
 sg13g2_decap_8 FILLER_50_163 ();
 sg13g2_decap_4 FILLER_50_170 ();
 sg13g2_fill_2 FILLER_50_231 ();
 sg13g2_fill_1 FILLER_50_272 ();
 sg13g2_decap_4 FILLER_50_304 ();
 sg13g2_fill_1 FILLER_50_318 ();
 sg13g2_fill_2 FILLER_50_336 ();
 sg13g2_fill_2 FILLER_50_359 ();
 sg13g2_decap_4 FILLER_50_364 ();
 sg13g2_fill_1 FILLER_50_368 ();
 sg13g2_fill_1 FILLER_50_382 ();
 sg13g2_fill_2 FILLER_50_392 ();
 sg13g2_fill_2 FILLER_50_419 ();
 sg13g2_fill_1 FILLER_50_421 ();
 sg13g2_fill_2 FILLER_50_464 ();
 sg13g2_fill_1 FILLER_50_496 ();
 sg13g2_fill_2 FILLER_50_509 ();
 sg13g2_fill_1 FILLER_50_522 ();
 sg13g2_decap_4 FILLER_50_544 ();
 sg13g2_fill_2 FILLER_50_548 ();
 sg13g2_fill_1 FILLER_50_574 ();
 sg13g2_fill_2 FILLER_50_580 ();
 sg13g2_decap_8 FILLER_50_617 ();
 sg13g2_fill_1 FILLER_50_624 ();
 sg13g2_decap_8 FILLER_50_631 ();
 sg13g2_fill_1 FILLER_50_643 ();
 sg13g2_fill_2 FILLER_50_649 ();
 sg13g2_decap_4 FILLER_50_668 ();
 sg13g2_fill_2 FILLER_50_685 ();
 sg13g2_fill_1 FILLER_50_687 ();
 sg13g2_fill_2 FILLER_50_692 ();
 sg13g2_fill_1 FILLER_50_694 ();
 sg13g2_decap_4 FILLER_50_733 ();
 sg13g2_decap_4 FILLER_50_766 ();
 sg13g2_fill_2 FILLER_50_770 ();
 sg13g2_fill_2 FILLER_50_799 ();
 sg13g2_fill_1 FILLER_50_801 ();
 sg13g2_fill_1 FILLER_50_819 ();
 sg13g2_fill_1 FILLER_50_825 ();
 sg13g2_decap_4 FILLER_50_839 ();
 sg13g2_fill_1 FILLER_50_843 ();
 sg13g2_fill_1 FILLER_50_852 ();
 sg13g2_fill_2 FILLER_50_909 ();
 sg13g2_fill_1 FILLER_50_916 ();
 sg13g2_decap_8 FILLER_50_930 ();
 sg13g2_fill_2 FILLER_50_937 ();
 sg13g2_fill_1 FILLER_50_939 ();
 sg13g2_decap_4 FILLER_50_992 ();
 sg13g2_fill_2 FILLER_50_996 ();
 sg13g2_decap_4 FILLER_50_1011 ();
 sg13g2_fill_1 FILLER_50_1015 ();
 sg13g2_fill_2 FILLER_50_1031 ();
 sg13g2_fill_2 FILLER_50_1056 ();
 sg13g2_fill_1 FILLER_50_1058 ();
 sg13g2_fill_2 FILLER_50_1064 ();
 sg13g2_decap_4 FILLER_50_1101 ();
 sg13g2_decap_8 FILLER_50_1123 ();
 sg13g2_decap_4 FILLER_50_1130 ();
 sg13g2_fill_2 FILLER_50_1134 ();
 sg13g2_fill_1 FILLER_50_1159 ();
 sg13g2_fill_2 FILLER_50_1164 ();
 sg13g2_fill_2 FILLER_50_1244 ();
 sg13g2_fill_1 FILLER_50_1246 ();
 sg13g2_fill_2 FILLER_50_1287 ();
 sg13g2_fill_1 FILLER_51_21 ();
 sg13g2_fill_2 FILLER_51_40 ();
 sg13g2_fill_2 FILLER_51_60 ();
 sg13g2_fill_2 FILLER_51_114 ();
 sg13g2_fill_1 FILLER_51_116 ();
 sg13g2_fill_1 FILLER_51_210 ();
 sg13g2_fill_2 FILLER_51_216 ();
 sg13g2_fill_2 FILLER_51_223 ();
 sg13g2_fill_1 FILLER_51_265 ();
 sg13g2_fill_2 FILLER_51_280 ();
 sg13g2_fill_2 FILLER_51_287 ();
 sg13g2_decap_4 FILLER_51_297 ();
 sg13g2_fill_1 FILLER_51_301 ();
 sg13g2_fill_2 FILLER_51_340 ();
 sg13g2_fill_2 FILLER_51_378 ();
 sg13g2_fill_1 FILLER_51_386 ();
 sg13g2_fill_2 FILLER_51_412 ();
 sg13g2_fill_1 FILLER_51_419 ();
 sg13g2_fill_1 FILLER_51_434 ();
 sg13g2_fill_2 FILLER_51_492 ();
 sg13g2_fill_1 FILLER_51_494 ();
 sg13g2_decap_8 FILLER_51_507 ();
 sg13g2_fill_2 FILLER_51_545 ();
 sg13g2_fill_2 FILLER_51_569 ();
 sg13g2_decap_4 FILLER_51_608 ();
 sg13g2_fill_2 FILLER_51_708 ();
 sg13g2_fill_2 FILLER_51_717 ();
 sg13g2_fill_1 FILLER_51_736 ();
 sg13g2_decap_4 FILLER_51_763 ();
 sg13g2_decap_8 FILLER_51_772 ();
 sg13g2_decap_8 FILLER_51_779 ();
 sg13g2_decap_8 FILLER_51_791 ();
 sg13g2_fill_2 FILLER_51_798 ();
 sg13g2_fill_2 FILLER_51_813 ();
 sg13g2_fill_1 FILLER_51_815 ();
 sg13g2_decap_8 FILLER_51_824 ();
 sg13g2_fill_2 FILLER_51_844 ();
 sg13g2_fill_2 FILLER_51_911 ();
 sg13g2_decap_8 FILLER_51_930 ();
 sg13g2_fill_2 FILLER_51_937 ();
 sg13g2_decap_4 FILLER_51_947 ();
 sg13g2_fill_1 FILLER_51_951 ();
 sg13g2_fill_2 FILLER_51_974 ();
 sg13g2_decap_4 FILLER_51_1024 ();
 sg13g2_fill_2 FILLER_51_1028 ();
 sg13g2_fill_2 FILLER_51_1112 ();
 sg13g2_decap_8 FILLER_51_1135 ();
 sg13g2_fill_2 FILLER_51_1142 ();
 sg13g2_fill_1 FILLER_51_1148 ();
 sg13g2_fill_1 FILLER_51_1206 ();
 sg13g2_fill_1 FILLER_51_1268 ();
 sg13g2_fill_2 FILLER_51_1313 ();
 sg13g2_fill_1 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_39 ();
 sg13g2_fill_2 FILLER_52_71 ();
 sg13g2_decap_4 FILLER_52_77 ();
 sg13g2_fill_1 FILLER_52_81 ();
 sg13g2_decap_4 FILLER_52_113 ();
 sg13g2_fill_2 FILLER_52_117 ();
 sg13g2_fill_1 FILLER_52_132 ();
 sg13g2_decap_8 FILLER_52_149 ();
 sg13g2_decap_8 FILLER_52_156 ();
 sg13g2_decap_8 FILLER_52_163 ();
 sg13g2_fill_2 FILLER_52_174 ();
 sg13g2_fill_1 FILLER_52_218 ();
 sg13g2_fill_1 FILLER_52_228 ();
 sg13g2_decap_4 FILLER_52_287 ();
 sg13g2_fill_1 FILLER_52_291 ();
 sg13g2_decap_8 FILLER_52_297 ();
 sg13g2_decap_8 FILLER_52_304 ();
 sg13g2_decap_8 FILLER_52_311 ();
 sg13g2_decap_8 FILLER_52_318 ();
 sg13g2_decap_4 FILLER_52_325 ();
 sg13g2_fill_1 FILLER_52_329 ();
 sg13g2_fill_1 FILLER_52_349 ();
 sg13g2_fill_2 FILLER_52_394 ();
 sg13g2_fill_2 FILLER_52_414 ();
 sg13g2_fill_1 FILLER_52_416 ();
 sg13g2_fill_1 FILLER_52_442 ();
 sg13g2_fill_2 FILLER_52_468 ();
 sg13g2_fill_1 FILLER_52_470 ();
 sg13g2_fill_2 FILLER_52_508 ();
 sg13g2_decap_4 FILLER_52_529 ();
 sg13g2_fill_2 FILLER_52_533 ();
 sg13g2_decap_4 FILLER_52_575 ();
 sg13g2_fill_2 FILLER_52_579 ();
 sg13g2_fill_1 FILLER_52_585 ();
 sg13g2_decap_4 FILLER_52_607 ();
 sg13g2_fill_2 FILLER_52_621 ();
 sg13g2_fill_1 FILLER_52_623 ();
 sg13g2_decap_4 FILLER_52_628 ();
 sg13g2_fill_1 FILLER_52_640 ();
 sg13g2_fill_2 FILLER_52_645 ();
 sg13g2_fill_1 FILLER_52_690 ();
 sg13g2_fill_2 FILLER_52_751 ();
 sg13g2_fill_1 FILLER_52_753 ();
 sg13g2_decap_4 FILLER_52_759 ();
 sg13g2_fill_1 FILLER_52_763 ();
 sg13g2_fill_2 FILLER_52_781 ();
 sg13g2_fill_1 FILLER_52_783 ();
 sg13g2_fill_1 FILLER_52_804 ();
 sg13g2_fill_2 FILLER_52_838 ();
 sg13g2_fill_1 FILLER_52_840 ();
 sg13g2_decap_4 FILLER_52_844 ();
 sg13g2_fill_2 FILLER_52_848 ();
 sg13g2_fill_2 FILLER_52_867 ();
 sg13g2_fill_1 FILLER_52_914 ();
 sg13g2_decap_8 FILLER_52_927 ();
 sg13g2_decap_4 FILLER_52_1047 ();
 sg13g2_fill_2 FILLER_52_1051 ();
 sg13g2_fill_2 FILLER_52_1072 ();
 sg13g2_decap_4 FILLER_52_1100 ();
 sg13g2_fill_2 FILLER_52_1130 ();
 sg13g2_fill_1 FILLER_52_1132 ();
 sg13g2_decap_4 FILLER_52_1159 ();
 sg13g2_fill_2 FILLER_52_1184 ();
 sg13g2_fill_1 FILLER_52_1248 ();
 sg13g2_fill_1 FILLER_52_1288 ();
 sg13g2_decap_4 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_17 ();
 sg13g2_fill_2 FILLER_53_25 ();
 sg13g2_fill_2 FILLER_53_68 ();
 sg13g2_decap_4 FILLER_53_151 ();
 sg13g2_fill_1 FILLER_53_193 ();
 sg13g2_fill_1 FILLER_53_255 ();
 sg13g2_fill_1 FILLER_53_265 ();
 sg13g2_fill_1 FILLER_53_306 ();
 sg13g2_fill_2 FILLER_53_311 ();
 sg13g2_fill_1 FILLER_53_313 ();
 sg13g2_fill_1 FILLER_53_356 ();
 sg13g2_decap_8 FILLER_53_386 ();
 sg13g2_fill_2 FILLER_53_393 ();
 sg13g2_fill_2 FILLER_53_431 ();
 sg13g2_fill_1 FILLER_53_433 ();
 sg13g2_fill_1 FILLER_53_460 ();
 sg13g2_decap_4 FILLER_53_495 ();
 sg13g2_decap_4 FILLER_53_505 ();
 sg13g2_fill_1 FILLER_53_509 ();
 sg13g2_decap_8 FILLER_53_515 ();
 sg13g2_decap_8 FILLER_53_522 ();
 sg13g2_fill_2 FILLER_53_529 ();
 sg13g2_fill_2 FILLER_53_594 ();
 sg13g2_fill_1 FILLER_53_596 ();
 sg13g2_fill_1 FILLER_53_617 ();
 sg13g2_fill_2 FILLER_53_628 ();
 sg13g2_fill_1 FILLER_53_630 ();
 sg13g2_decap_4 FILLER_53_651 ();
 sg13g2_fill_2 FILLER_53_721 ();
 sg13g2_fill_1 FILLER_53_723 ();
 sg13g2_fill_2 FILLER_53_746 ();
 sg13g2_fill_1 FILLER_53_752 ();
 sg13g2_fill_2 FILLER_53_805 ();
 sg13g2_fill_1 FILLER_53_807 ();
 sg13g2_fill_1 FILLER_53_813 ();
 sg13g2_fill_1 FILLER_53_836 ();
 sg13g2_fill_2 FILLER_53_850 ();
 sg13g2_fill_1 FILLER_53_852 ();
 sg13g2_fill_1 FILLER_53_871 ();
 sg13g2_decap_8 FILLER_53_907 ();
 sg13g2_decap_4 FILLER_53_940 ();
 sg13g2_fill_1 FILLER_53_944 ();
 sg13g2_decap_8 FILLER_53_953 ();
 sg13g2_fill_2 FILLER_53_960 ();
 sg13g2_fill_1 FILLER_53_962 ();
 sg13g2_fill_2 FILLER_53_1063 ();
 sg13g2_fill_1 FILLER_53_1065 ();
 sg13g2_fill_1 FILLER_53_1096 ();
 sg13g2_fill_1 FILLER_53_1119 ();
 sg13g2_fill_2 FILLER_53_1134 ();
 sg13g2_fill_1 FILLER_53_1136 ();
 sg13g2_fill_2 FILLER_53_1268 ();
 sg13g2_fill_1 FILLER_53_1314 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_2 ();
 sg13g2_fill_1 FILLER_54_39 ();
 sg13g2_fill_2 FILLER_54_45 ();
 sg13g2_fill_1 FILLER_54_77 ();
 sg13g2_fill_2 FILLER_54_94 ();
 sg13g2_fill_1 FILLER_54_113 ();
 sg13g2_fill_1 FILLER_54_123 ();
 sg13g2_fill_2 FILLER_54_161 ();
 sg13g2_fill_1 FILLER_54_238 ();
 sg13g2_fill_1 FILLER_54_349 ();
 sg13g2_fill_1 FILLER_54_355 ();
 sg13g2_fill_1 FILLER_54_361 ();
 sg13g2_fill_2 FILLER_54_371 ();
 sg13g2_decap_8 FILLER_54_382 ();
 sg13g2_decap_8 FILLER_54_389 ();
 sg13g2_decap_4 FILLER_54_426 ();
 sg13g2_fill_1 FILLER_54_458 ();
 sg13g2_fill_2 FILLER_54_474 ();
 sg13g2_decap_8 FILLER_54_480 ();
 sg13g2_decap_8 FILLER_54_487 ();
 sg13g2_fill_1 FILLER_54_500 ();
 sg13g2_decap_4 FILLER_54_513 ();
 sg13g2_fill_1 FILLER_54_517 ();
 sg13g2_fill_1 FILLER_54_560 ();
 sg13g2_fill_1 FILLER_54_586 ();
 sg13g2_fill_2 FILLER_54_600 ();
 sg13g2_fill_1 FILLER_54_610 ();
 sg13g2_decap_8 FILLER_54_624 ();
 sg13g2_decap_4 FILLER_54_631 ();
 sg13g2_fill_1 FILLER_54_657 ();
 sg13g2_decap_8 FILLER_54_662 ();
 sg13g2_decap_8 FILLER_54_669 ();
 sg13g2_fill_2 FILLER_54_676 ();
 sg13g2_fill_1 FILLER_54_701 ();
 sg13g2_fill_1 FILLER_54_715 ();
 sg13g2_decap_8 FILLER_54_750 ();
 sg13g2_decap_4 FILLER_54_757 ();
 sg13g2_decap_8 FILLER_54_766 ();
 sg13g2_fill_2 FILLER_54_773 ();
 sg13g2_fill_1 FILLER_54_775 ();
 sg13g2_decap_4 FILLER_54_780 ();
 sg13g2_fill_1 FILLER_54_789 ();
 sg13g2_fill_1 FILLER_54_795 ();
 sg13g2_fill_2 FILLER_54_800 ();
 sg13g2_fill_1 FILLER_54_802 ();
 sg13g2_fill_1 FILLER_54_841 ();
 sg13g2_fill_1 FILLER_54_847 ();
 sg13g2_fill_1 FILLER_54_852 ();
 sg13g2_decap_4 FILLER_54_891 ();
 sg13g2_fill_1 FILLER_54_895 ();
 sg13g2_fill_1 FILLER_54_909 ();
 sg13g2_decap_4 FILLER_54_930 ();
 sg13g2_fill_1 FILLER_54_964 ();
 sg13g2_fill_2 FILLER_54_1008 ();
 sg13g2_fill_1 FILLER_54_1010 ();
 sg13g2_fill_1 FILLER_54_1034 ();
 sg13g2_decap_4 FILLER_54_1114 ();
 sg13g2_fill_1 FILLER_54_1118 ();
 sg13g2_fill_2 FILLER_54_1123 ();
 sg13g2_decap_4 FILLER_54_1151 ();
 sg13g2_fill_1 FILLER_54_1155 ();
 sg13g2_fill_2 FILLER_54_1186 ();
 sg13g2_fill_1 FILLER_54_1188 ();
 sg13g2_fill_1 FILLER_54_1219 ();
 sg13g2_fill_2 FILLER_54_1251 ();
 sg13g2_fill_1 FILLER_54_1253 ();
 sg13g2_decap_4 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_4 ();
 sg13g2_fill_2 FILLER_55_18 ();
 sg13g2_fill_1 FILLER_55_84 ();
 sg13g2_fill_2 FILLER_55_120 ();
 sg13g2_decap_4 FILLER_55_176 ();
 sg13g2_fill_2 FILLER_55_180 ();
 sg13g2_fill_1 FILLER_55_194 ();
 sg13g2_fill_1 FILLER_55_223 ();
 sg13g2_fill_2 FILLER_55_255 ();
 sg13g2_fill_1 FILLER_55_262 ();
 sg13g2_fill_2 FILLER_55_296 ();
 sg13g2_fill_2 FILLER_55_396 ();
 sg13g2_fill_1 FILLER_55_473 ();
 sg13g2_fill_2 FILLER_55_500 ();
 sg13g2_decap_8 FILLER_55_528 ();
 sg13g2_decap_8 FILLER_55_535 ();
 sg13g2_decap_8 FILLER_55_542 ();
 sg13g2_decap_8 FILLER_55_549 ();
 sg13g2_decap_8 FILLER_55_556 ();
 sg13g2_decap_8 FILLER_55_563 ();
 sg13g2_fill_2 FILLER_55_570 ();
 sg13g2_fill_1 FILLER_55_572 ();
 sg13g2_fill_2 FILLER_55_581 ();
 sg13g2_fill_1 FILLER_55_596 ();
 sg13g2_decap_4 FILLER_55_604 ();
 sg13g2_fill_1 FILLER_55_608 ();
 sg13g2_fill_1 FILLER_55_635 ();
 sg13g2_fill_2 FILLER_55_729 ();
 sg13g2_fill_1 FILLER_55_731 ();
 sg13g2_fill_1 FILLER_55_773 ();
 sg13g2_decap_4 FILLER_55_809 ();
 sg13g2_fill_1 FILLER_55_813 ();
 sg13g2_fill_1 FILLER_55_904 ();
 sg13g2_fill_2 FILLER_55_915 ();
 sg13g2_fill_1 FILLER_55_917 ();
 sg13g2_decap_8 FILLER_55_937 ();
 sg13g2_fill_2 FILLER_55_964 ();
 sg13g2_fill_1 FILLER_55_983 ();
 sg13g2_decap_4 FILLER_55_989 ();
 sg13g2_fill_2 FILLER_55_993 ();
 sg13g2_fill_2 FILLER_55_998 ();
 sg13g2_fill_1 FILLER_55_1000 ();
 sg13g2_fill_2 FILLER_55_1037 ();
 sg13g2_fill_1 FILLER_55_1039 ();
 sg13g2_fill_2 FILLER_55_1050 ();
 sg13g2_fill_1 FILLER_55_1072 ();
 sg13g2_fill_2 FILLER_55_1081 ();
 sg13g2_fill_1 FILLER_55_1083 ();
 sg13g2_fill_2 FILLER_55_1109 ();
 sg13g2_fill_1 FILLER_55_1127 ();
 sg13g2_decap_4 FILLER_55_1142 ();
 sg13g2_fill_2 FILLER_55_1156 ();
 sg13g2_fill_2 FILLER_55_1236 ();
 sg13g2_fill_1 FILLER_55_1273 ();
 sg13g2_fill_2 FILLER_55_1313 ();
 sg13g2_fill_1 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_58 ();
 sg13g2_fill_1 FILLER_56_95 ();
 sg13g2_fill_1 FILLER_56_136 ();
 sg13g2_fill_2 FILLER_56_207 ();
 sg13g2_fill_1 FILLER_56_209 ();
 sg13g2_fill_1 FILLER_56_224 ();
 sg13g2_fill_2 FILLER_56_304 ();
 sg13g2_fill_1 FILLER_56_366 ();
 sg13g2_fill_2 FILLER_56_372 ();
 sg13g2_fill_2 FILLER_56_387 ();
 sg13g2_fill_1 FILLER_56_389 ();
 sg13g2_decap_8 FILLER_56_399 ();
 sg13g2_decap_8 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_413 ();
 sg13g2_fill_2 FILLER_56_429 ();
 sg13g2_fill_1 FILLER_56_436 ();
 sg13g2_decap_4 FILLER_56_444 ();
 sg13g2_fill_1 FILLER_56_461 ();
 sg13g2_fill_1 FILLER_56_468 ();
 sg13g2_fill_2 FILLER_56_483 ();
 sg13g2_fill_1 FILLER_56_485 ();
 sg13g2_decap_8 FILLER_56_524 ();
 sg13g2_fill_1 FILLER_56_531 ();
 sg13g2_decap_8 FILLER_56_563 ();
 sg13g2_decap_8 FILLER_56_570 ();
 sg13g2_fill_2 FILLER_56_577 ();
 sg13g2_fill_1 FILLER_56_612 ();
 sg13g2_fill_2 FILLER_56_617 ();
 sg13g2_fill_1 FILLER_56_619 ();
 sg13g2_fill_2 FILLER_56_624 ();
 sg13g2_fill_1 FILLER_56_626 ();
 sg13g2_fill_1 FILLER_56_668 ();
 sg13g2_fill_2 FILLER_56_696 ();
 sg13g2_fill_1 FILLER_56_703 ();
 sg13g2_fill_2 FILLER_56_721 ();
 sg13g2_fill_1 FILLER_56_723 ();
 sg13g2_fill_1 FILLER_56_754 ();
 sg13g2_decap_4 FILLER_56_781 ();
 sg13g2_fill_2 FILLER_56_785 ();
 sg13g2_fill_1 FILLER_56_805 ();
 sg13g2_fill_2 FILLER_56_818 ();
 sg13g2_fill_2 FILLER_56_832 ();
 sg13g2_decap_8 FILLER_56_842 ();
 sg13g2_decap_4 FILLER_56_849 ();
 sg13g2_fill_2 FILLER_56_853 ();
 sg13g2_fill_2 FILLER_56_876 ();
 sg13g2_fill_1 FILLER_56_913 ();
 sg13g2_fill_2 FILLER_56_943 ();
 sg13g2_decap_4 FILLER_56_986 ();
 sg13g2_fill_2 FILLER_56_990 ();
 sg13g2_decap_8 FILLER_56_997 ();
 sg13g2_fill_1 FILLER_56_1004 ();
 sg13g2_fill_2 FILLER_56_1015 ();
 sg13g2_decap_4 FILLER_56_1021 ();
 sg13g2_fill_1 FILLER_56_1025 ();
 sg13g2_fill_2 FILLER_56_1078 ();
 sg13g2_fill_1 FILLER_56_1080 ();
 sg13g2_fill_2 FILLER_56_1094 ();
 sg13g2_fill_1 FILLER_56_1096 ();
 sg13g2_fill_2 FILLER_56_1118 ();
 sg13g2_fill_2 FILLER_56_1151 ();
 sg13g2_fill_1 FILLER_56_1165 ();
 sg13g2_fill_2 FILLER_56_1223 ();
 sg13g2_fill_2 FILLER_56_1287 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_65 ();
 sg13g2_fill_1 FILLER_57_72 ();
 sg13g2_fill_2 FILLER_57_121 ();
 sg13g2_fill_1 FILLER_57_149 ();
 sg13g2_fill_2 FILLER_57_159 ();
 sg13g2_fill_1 FILLER_57_201 ();
 sg13g2_fill_1 FILLER_57_240 ();
 sg13g2_fill_2 FILLER_57_257 ();
 sg13g2_fill_2 FILLER_57_264 ();
 sg13g2_decap_4 FILLER_57_327 ();
 sg13g2_fill_1 FILLER_57_331 ();
 sg13g2_fill_1 FILLER_57_341 ();
 sg13g2_decap_4 FILLER_57_416 ();
 sg13g2_decap_8 FILLER_57_424 ();
 sg13g2_fill_1 FILLER_57_431 ();
 sg13g2_fill_1 FILLER_57_467 ();
 sg13g2_decap_4 FILLER_57_476 ();
 sg13g2_fill_2 FILLER_57_494 ();
 sg13g2_fill_2 FILLER_57_515 ();
 sg13g2_decap_4 FILLER_57_585 ();
 sg13g2_fill_2 FILLER_57_589 ();
 sg13g2_decap_8 FILLER_57_598 ();
 sg13g2_decap_8 FILLER_57_605 ();
 sg13g2_decap_8 FILLER_57_612 ();
 sg13g2_fill_2 FILLER_57_619 ();
 sg13g2_fill_2 FILLER_57_666 ();
 sg13g2_fill_1 FILLER_57_668 ();
 sg13g2_fill_2 FILLER_57_723 ();
 sg13g2_decap_8 FILLER_57_740 ();
 sg13g2_decap_8 FILLER_57_747 ();
 sg13g2_fill_2 FILLER_57_754 ();
 sg13g2_fill_1 FILLER_57_756 ();
 sg13g2_decap_4 FILLER_57_774 ();
 sg13g2_fill_1 FILLER_57_855 ();
 sg13g2_fill_1 FILLER_57_865 ();
 sg13g2_fill_1 FILLER_57_881 ();
 sg13g2_fill_1 FILLER_57_910 ();
 sg13g2_fill_1 FILLER_57_916 ();
 sg13g2_decap_4 FILLER_57_927 ();
 sg13g2_decap_4 FILLER_57_948 ();
 sg13g2_fill_1 FILLER_57_952 ();
 sg13g2_decap_4 FILLER_57_970 ();
 sg13g2_fill_1 FILLER_57_1005 ();
 sg13g2_decap_8 FILLER_57_1030 ();
 sg13g2_decap_8 FILLER_57_1041 ();
 sg13g2_fill_1 FILLER_57_1048 ();
 sg13g2_decap_4 FILLER_57_1067 ();
 sg13g2_fill_1 FILLER_57_1071 ();
 sg13g2_fill_2 FILLER_57_1101 ();
 sg13g2_fill_1 FILLER_57_1103 ();
 sg13g2_fill_2 FILLER_57_1117 ();
 sg13g2_fill_1 FILLER_57_1119 ();
 sg13g2_decap_4 FILLER_57_1129 ();
 sg13g2_fill_2 FILLER_57_1242 ();
 sg13g2_fill_1 FILLER_57_1249 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_28 ();
 sg13g2_fill_1 FILLER_58_131 ();
 sg13g2_fill_1 FILLER_58_181 ();
 sg13g2_fill_2 FILLER_58_191 ();
 sg13g2_fill_2 FILLER_58_216 ();
 sg13g2_fill_1 FILLER_58_304 ();
 sg13g2_fill_1 FILLER_58_335 ();
 sg13g2_fill_2 FILLER_58_375 ();
 sg13g2_fill_1 FILLER_58_377 ();
 sg13g2_decap_4 FILLER_58_382 ();
 sg13g2_fill_1 FILLER_58_386 ();
 sg13g2_decap_4 FILLER_58_392 ();
 sg13g2_fill_1 FILLER_58_396 ();
 sg13g2_fill_1 FILLER_58_414 ();
 sg13g2_fill_2 FILLER_58_439 ();
 sg13g2_fill_1 FILLER_58_475 ();
 sg13g2_fill_2 FILLER_58_507 ();
 sg13g2_fill_1 FILLER_58_514 ();
 sg13g2_decap_4 FILLER_58_539 ();
 sg13g2_fill_1 FILLER_58_543 ();
 sg13g2_fill_1 FILLER_58_565 ();
 sg13g2_fill_1 FILLER_58_655 ();
 sg13g2_fill_1 FILLER_58_665 ();
 sg13g2_fill_1 FILLER_58_699 ();
 sg13g2_decap_4 FILLER_58_708 ();
 sg13g2_fill_2 FILLER_58_712 ();
 sg13g2_decap_8 FILLER_58_734 ();
 sg13g2_decap_4 FILLER_58_750 ();
 sg13g2_fill_2 FILLER_58_754 ();
 sg13g2_fill_2 FILLER_58_761 ();
 sg13g2_fill_2 FILLER_58_771 ();
 sg13g2_fill_1 FILLER_58_773 ();
 sg13g2_decap_4 FILLER_58_779 ();
 sg13g2_fill_2 FILLER_58_783 ();
 sg13g2_fill_2 FILLER_58_950 ();
 sg13g2_fill_1 FILLER_58_952 ();
 sg13g2_fill_1 FILLER_58_968 ();
 sg13g2_fill_1 FILLER_58_975 ();
 sg13g2_fill_2 FILLER_58_989 ();
 sg13g2_fill_1 FILLER_58_991 ();
 sg13g2_decap_8 FILLER_58_1010 ();
 sg13g2_decap_8 FILLER_58_1041 ();
 sg13g2_decap_8 FILLER_58_1048 ();
 sg13g2_decap_8 FILLER_58_1055 ();
 sg13g2_fill_2 FILLER_58_1062 ();
 sg13g2_decap_8 FILLER_58_1068 ();
 sg13g2_fill_2 FILLER_58_1075 ();
 sg13g2_fill_2 FILLER_58_1081 ();
 sg13g2_fill_1 FILLER_58_1083 ();
 sg13g2_decap_4 FILLER_58_1093 ();
 sg13g2_decap_8 FILLER_58_1137 ();
 sg13g2_decap_8 FILLER_58_1148 ();
 sg13g2_fill_2 FILLER_58_1155 ();
 sg13g2_fill_1 FILLER_58_1157 ();
 sg13g2_fill_2 FILLER_58_1166 ();
 sg13g2_fill_1 FILLER_58_1177 ();
 sg13g2_fill_1 FILLER_58_1191 ();
 sg13g2_fill_2 FILLER_58_1218 ();
 sg13g2_fill_2 FILLER_58_1278 ();
 sg13g2_fill_1 FILLER_58_1280 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_20 ();
 sg13g2_fill_2 FILLER_59_42 ();
 sg13g2_fill_1 FILLER_59_44 ();
 sg13g2_fill_2 FILLER_59_49 ();
 sg13g2_fill_1 FILLER_59_164 ();
 sg13g2_fill_2 FILLER_59_182 ();
 sg13g2_fill_1 FILLER_59_212 ();
 sg13g2_fill_1 FILLER_59_232 ();
 sg13g2_fill_2 FILLER_59_246 ();
 sg13g2_fill_1 FILLER_59_312 ();
 sg13g2_fill_2 FILLER_59_323 ();
 sg13g2_fill_1 FILLER_59_325 ();
 sg13g2_fill_2 FILLER_59_341 ();
 sg13g2_fill_2 FILLER_59_353 ();
 sg13g2_fill_1 FILLER_59_355 ();
 sg13g2_fill_1 FILLER_59_488 ();
 sg13g2_fill_1 FILLER_59_503 ();
 sg13g2_fill_2 FILLER_59_533 ();
 sg13g2_fill_1 FILLER_59_535 ();
 sg13g2_fill_2 FILLER_59_588 ();
 sg13g2_fill_1 FILLER_59_590 ();
 sg13g2_fill_1 FILLER_59_615 ();
 sg13g2_decap_4 FILLER_59_712 ();
 sg13g2_fill_2 FILLER_59_716 ();
 sg13g2_fill_2 FILLER_59_723 ();
 sg13g2_fill_1 FILLER_59_755 ();
 sg13g2_decap_4 FILLER_59_764 ();
 sg13g2_decap_8 FILLER_59_786 ();
 sg13g2_fill_1 FILLER_59_793 ();
 sg13g2_fill_1 FILLER_59_799 ();
 sg13g2_fill_2 FILLER_59_839 ();
 sg13g2_fill_1 FILLER_59_841 ();
 sg13g2_decap_8 FILLER_59_865 ();
 sg13g2_decap_8 FILLER_59_872 ();
 sg13g2_decap_8 FILLER_59_879 ();
 sg13g2_decap_8 FILLER_59_886 ();
 sg13g2_decap_4 FILLER_59_893 ();
 sg13g2_fill_2 FILLER_59_897 ();
 sg13g2_fill_2 FILLER_59_908 ();
 sg13g2_decap_4 FILLER_59_925 ();
 sg13g2_fill_2 FILLER_59_929 ();
 sg13g2_decap_4 FILLER_59_935 ();
 sg13g2_fill_1 FILLER_59_939 ();
 sg13g2_fill_2 FILLER_59_964 ();
 sg13g2_decap_8 FILLER_59_1014 ();
 sg13g2_fill_1 FILLER_59_1021 ();
 sg13g2_decap_8 FILLER_59_1039 ();
 sg13g2_decap_8 FILLER_59_1046 ();
 sg13g2_decap_8 FILLER_59_1053 ();
 sg13g2_decap_8 FILLER_59_1060 ();
 sg13g2_fill_1 FILLER_59_1067 ();
 sg13g2_decap_4 FILLER_59_1097 ();
 sg13g2_fill_1 FILLER_59_1101 ();
 sg13g2_decap_8 FILLER_59_1111 ();
 sg13g2_fill_2 FILLER_59_1136 ();
 sg13g2_fill_1 FILLER_59_1212 ();
 sg13g2_fill_2 FILLER_59_1304 ();
 sg13g2_fill_1 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_64 ();
 sg13g2_fill_1 FILLER_60_66 ();
 sg13g2_fill_2 FILLER_60_102 ();
 sg13g2_fill_1 FILLER_60_121 ();
 sg13g2_fill_2 FILLER_60_146 ();
 sg13g2_fill_1 FILLER_60_148 ();
 sg13g2_decap_4 FILLER_60_157 ();
 sg13g2_fill_1 FILLER_60_253 ();
 sg13g2_fill_2 FILLER_60_264 ();
 sg13g2_fill_2 FILLER_60_290 ();
 sg13g2_fill_2 FILLER_60_314 ();
 sg13g2_fill_2 FILLER_60_326 ();
 sg13g2_fill_1 FILLER_60_333 ();
 sg13g2_fill_1 FILLER_60_350 ();
 sg13g2_fill_1 FILLER_60_382 ();
 sg13g2_decap_8 FILLER_60_401 ();
 sg13g2_decap_8 FILLER_60_412 ();
 sg13g2_fill_2 FILLER_60_419 ();
 sg13g2_decap_8 FILLER_60_425 ();
 sg13g2_fill_2 FILLER_60_463 ();
 sg13g2_fill_1 FILLER_60_465 ();
 sg13g2_fill_2 FILLER_60_475 ();
 sg13g2_fill_1 FILLER_60_477 ();
 sg13g2_fill_2 FILLER_60_514 ();
 sg13g2_fill_2 FILLER_60_636 ();
 sg13g2_fill_1 FILLER_60_638 ();
 sg13g2_fill_2 FILLER_60_654 ();
 sg13g2_fill_1 FILLER_60_656 ();
 sg13g2_fill_1 FILLER_60_680 ();
 sg13g2_fill_1 FILLER_60_704 ();
 sg13g2_fill_2 FILLER_60_728 ();
 sg13g2_fill_1 FILLER_60_730 ();
 sg13g2_decap_8 FILLER_60_750 ();
 sg13g2_fill_1 FILLER_60_818 ();
 sg13g2_decap_4 FILLER_60_837 ();
 sg13g2_decap_4 FILLER_60_880 ();
 sg13g2_fill_1 FILLER_60_947 ();
 sg13g2_fill_1 FILLER_60_977 ();
 sg13g2_fill_2 FILLER_60_988 ();
 sg13g2_fill_2 FILLER_60_994 ();
 sg13g2_fill_2 FILLER_60_1028 ();
 sg13g2_decap_8 FILLER_60_1051 ();
 sg13g2_fill_2 FILLER_60_1058 ();
 sg13g2_fill_1 FILLER_60_1060 ();
 sg13g2_fill_1 FILLER_60_1081 ();
 sg13g2_decap_8 FILLER_60_1091 ();
 sg13g2_decap_4 FILLER_60_1098 ();
 sg13g2_fill_1 FILLER_60_1102 ();
 sg13g2_fill_2 FILLER_60_1131 ();
 sg13g2_fill_1 FILLER_60_1133 ();
 sg13g2_fill_2 FILLER_60_1144 ();
 sg13g2_fill_2 FILLER_60_1254 ();
 sg13g2_fill_1 FILLER_60_1256 ();
 sg13g2_fill_1 FILLER_60_1314 ();
 sg13g2_fill_2 FILLER_61_40 ();
 sg13g2_fill_1 FILLER_61_42 ();
 sg13g2_decap_4 FILLER_61_73 ();
 sg13g2_fill_2 FILLER_61_77 ();
 sg13g2_fill_2 FILLER_61_214 ();
 sg13g2_fill_2 FILLER_61_220 ();
 sg13g2_fill_1 FILLER_61_222 ();
 sg13g2_fill_2 FILLER_61_325 ();
 sg13g2_fill_1 FILLER_61_357 ();
 sg13g2_decap_8 FILLER_61_389 ();
 sg13g2_decap_4 FILLER_61_396 ();
 sg13g2_fill_1 FILLER_61_400 ();
 sg13g2_decap_8 FILLER_61_405 ();
 sg13g2_fill_2 FILLER_61_412 ();
 sg13g2_decap_4 FILLER_61_419 ();
 sg13g2_fill_1 FILLER_61_423 ();
 sg13g2_fill_1 FILLER_61_449 ();
 sg13g2_fill_1 FILLER_61_480 ();
 sg13g2_fill_1 FILLER_61_490 ();
 sg13g2_fill_2 FILLER_61_519 ();
 sg13g2_fill_2 FILLER_61_535 ();
 sg13g2_decap_4 FILLER_61_541 ();
 sg13g2_decap_8 FILLER_61_575 ();
 sg13g2_decap_4 FILLER_61_582 ();
 sg13g2_fill_2 FILLER_61_594 ();
 sg13g2_fill_2 FILLER_61_695 ();
 sg13g2_fill_1 FILLER_61_697 ();
 sg13g2_decap_4 FILLER_61_702 ();
 sg13g2_fill_1 FILLER_61_706 ();
 sg13g2_decap_8 FILLER_61_711 ();
 sg13g2_fill_1 FILLER_61_718 ();
 sg13g2_fill_1 FILLER_61_727 ();
 sg13g2_fill_2 FILLER_61_733 ();
 sg13g2_decap_4 FILLER_61_752 ();
 sg13g2_decap_8 FILLER_61_764 ();
 sg13g2_fill_1 FILLER_61_771 ();
 sg13g2_fill_2 FILLER_61_781 ();
 sg13g2_fill_1 FILLER_61_783 ();
 sg13g2_fill_2 FILLER_61_789 ();
 sg13g2_decap_8 FILLER_61_796 ();
 sg13g2_fill_1 FILLER_61_803 ();
 sg13g2_decap_8 FILLER_61_809 ();
 sg13g2_fill_2 FILLER_61_816 ();
 sg13g2_fill_1 FILLER_61_834 ();
 sg13g2_decap_4 FILLER_61_861 ();
 sg13g2_fill_2 FILLER_61_869 ();
 sg13g2_fill_1 FILLER_61_871 ();
 sg13g2_fill_1 FILLER_61_908 ();
 sg13g2_decap_4 FILLER_61_957 ();
 sg13g2_fill_1 FILLER_61_961 ();
 sg13g2_decap_8 FILLER_61_983 ();
 sg13g2_decap_4 FILLER_61_990 ();
 sg13g2_fill_1 FILLER_61_994 ();
 sg13g2_fill_2 FILLER_61_1022 ();
 sg13g2_fill_1 FILLER_61_1032 ();
 sg13g2_decap_8 FILLER_61_1042 ();
 sg13g2_decap_8 FILLER_61_1049 ();
 sg13g2_fill_2 FILLER_61_1056 ();
 sg13g2_fill_1 FILLER_61_1067 ();
 sg13g2_decap_4 FILLER_61_1073 ();
 sg13g2_decap_8 FILLER_61_1101 ();
 sg13g2_fill_2 FILLER_61_1108 ();
 sg13g2_decap_8 FILLER_61_1132 ();
 sg13g2_fill_1 FILLER_61_1139 ();
 sg13g2_fill_2 FILLER_61_1287 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_56 ();
 sg13g2_decap_4 FILLER_62_74 ();
 sg13g2_fill_2 FILLER_62_139 ();
 sg13g2_fill_2 FILLER_62_146 ();
 sg13g2_fill_2 FILLER_62_165 ();
 sg13g2_fill_2 FILLER_62_233 ();
 sg13g2_fill_1 FILLER_62_270 ();
 sg13g2_fill_1 FILLER_62_279 ();
 sg13g2_decap_4 FILLER_62_296 ();
 sg13g2_fill_1 FILLER_62_300 ();
 sg13g2_fill_2 FILLER_62_304 ();
 sg13g2_fill_1 FILLER_62_306 ();
 sg13g2_fill_2 FILLER_62_312 ();
 sg13g2_fill_1 FILLER_62_314 ();
 sg13g2_fill_1 FILLER_62_326 ();
 sg13g2_fill_2 FILLER_62_332 ();
 sg13g2_fill_1 FILLER_62_340 ();
 sg13g2_fill_2 FILLER_62_345 ();
 sg13g2_decap_8 FILLER_62_357 ();
 sg13g2_decap_4 FILLER_62_364 ();
 sg13g2_fill_2 FILLER_62_368 ();
 sg13g2_fill_1 FILLER_62_378 ();
 sg13g2_fill_2 FILLER_62_383 ();
 sg13g2_fill_1 FILLER_62_520 ();
 sg13g2_fill_2 FILLER_62_530 ();
 sg13g2_fill_1 FILLER_62_532 ();
 sg13g2_decap_8 FILLER_62_537 ();
 sg13g2_decap_4 FILLER_62_544 ();
 sg13g2_fill_2 FILLER_62_560 ();
 sg13g2_fill_1 FILLER_62_562 ();
 sg13g2_decap_8 FILLER_62_593 ();
 sg13g2_fill_2 FILLER_62_600 ();
 sg13g2_fill_1 FILLER_62_602 ();
 sg13g2_fill_2 FILLER_62_631 ();
 sg13g2_fill_1 FILLER_62_637 ();
 sg13g2_fill_1 FILLER_62_664 ();
 sg13g2_fill_1 FILLER_62_704 ();
 sg13g2_decap_4 FILLER_62_715 ();
 sg13g2_fill_2 FILLER_62_719 ();
 sg13g2_fill_1 FILLER_62_726 ();
 sg13g2_decap_4 FILLER_62_735 ();
 sg13g2_fill_1 FILLER_62_739 ();
 sg13g2_fill_2 FILLER_62_752 ();
 sg13g2_fill_1 FILLER_62_754 ();
 sg13g2_decap_4 FILLER_62_833 ();
 sg13g2_fill_2 FILLER_62_871 ();
 sg13g2_fill_1 FILLER_62_882 ();
 sg13g2_decap_8 FILLER_62_978 ();
 sg13g2_decap_8 FILLER_62_985 ();
 sg13g2_fill_1 FILLER_62_992 ();
 sg13g2_decap_8 FILLER_62_998 ();
 sg13g2_fill_1 FILLER_62_1005 ();
 sg13g2_decap_8 FILLER_62_1011 ();
 sg13g2_decap_8 FILLER_62_1018 ();
 sg13g2_fill_2 FILLER_62_1025 ();
 sg13g2_fill_1 FILLER_62_1052 ();
 sg13g2_fill_1 FILLER_62_1073 ();
 sg13g2_decap_4 FILLER_62_1086 ();
 sg13g2_decap_4 FILLER_62_1099 ();
 sg13g2_fill_1 FILLER_62_1103 ();
 sg13g2_fill_1 FILLER_62_1112 ();
 sg13g2_fill_1 FILLER_62_1116 ();
 sg13g2_fill_2 FILLER_62_1121 ();
 sg13g2_fill_1 FILLER_62_1149 ();
 sg13g2_fill_2 FILLER_62_1175 ();
 sg13g2_fill_2 FILLER_62_1247 ();
 sg13g2_fill_1 FILLER_62_1288 ();
 sg13g2_fill_2 FILLER_63_93 ();
 sg13g2_fill_2 FILLER_63_130 ();
 sg13g2_fill_1 FILLER_63_145 ();
 sg13g2_fill_1 FILLER_63_205 ();
 sg13g2_fill_1 FILLER_63_215 ();
 sg13g2_fill_2 FILLER_63_230 ();
 sg13g2_fill_1 FILLER_63_232 ();
 sg13g2_fill_1 FILLER_63_252 ();
 sg13g2_fill_2 FILLER_63_272 ();
 sg13g2_fill_1 FILLER_63_320 ();
 sg13g2_fill_1 FILLER_63_350 ();
 sg13g2_decap_4 FILLER_63_360 ();
 sg13g2_fill_1 FILLER_63_390 ();
 sg13g2_fill_2 FILLER_63_417 ();
 sg13g2_decap_4 FILLER_63_423 ();
 sg13g2_decap_8 FILLER_63_431 ();
 sg13g2_decap_4 FILLER_63_465 ();
 sg13g2_fill_2 FILLER_63_505 ();
 sg13g2_fill_1 FILLER_63_507 ();
 sg13g2_fill_2 FILLER_63_514 ();
 sg13g2_fill_1 FILLER_63_526 ();
 sg13g2_fill_2 FILLER_63_538 ();
 sg13g2_fill_1 FILLER_63_545 ();
 sg13g2_fill_1 FILLER_63_564 ();
 sg13g2_fill_1 FILLER_63_709 ();
 sg13g2_fill_1 FILLER_63_719 ();
 sg13g2_decap_8 FILLER_63_728 ();
 sg13g2_decap_4 FILLER_63_735 ();
 sg13g2_fill_1 FILLER_63_739 ();
 sg13g2_decap_4 FILLER_63_750 ();
 sg13g2_fill_1 FILLER_63_754 ();
 sg13g2_fill_2 FILLER_63_770 ();
 sg13g2_fill_2 FILLER_63_776 ();
 sg13g2_fill_1 FILLER_63_778 ();
 sg13g2_fill_2 FILLER_63_833 ();
 sg13g2_decap_8 FILLER_63_849 ();
 sg13g2_decap_4 FILLER_63_860 ();
 sg13g2_fill_1 FILLER_63_899 ();
 sg13g2_fill_1 FILLER_63_955 ();
 sg13g2_fill_1 FILLER_63_985 ();
 sg13g2_decap_4 FILLER_63_999 ();
 sg13g2_fill_2 FILLER_63_1028 ();
 sg13g2_decap_8 FILLER_63_1047 ();
 sg13g2_decap_4 FILLER_63_1054 ();
 sg13g2_decap_4 FILLER_63_1067 ();
 sg13g2_fill_1 FILLER_63_1071 ();
 sg13g2_fill_2 FILLER_63_1089 ();
 sg13g2_fill_1 FILLER_63_1091 ();
 sg13g2_fill_1 FILLER_63_1115 ();
 sg13g2_decap_4 FILLER_63_1129 ();
 sg13g2_fill_1 FILLER_63_1133 ();
 sg13g2_decap_4 FILLER_63_1138 ();
 sg13g2_fill_1 FILLER_63_1204 ();
 sg13g2_fill_2 FILLER_63_1266 ();
 sg13g2_fill_1 FILLER_63_1268 ();
 sg13g2_fill_2 FILLER_63_1295 ();
 sg13g2_fill_1 FILLER_64_33 ();
 sg13g2_fill_2 FILLER_64_60 ();
 sg13g2_fill_2 FILLER_64_76 ();
 sg13g2_decap_4 FILLER_64_89 ();
 sg13g2_fill_2 FILLER_64_93 ();
 sg13g2_fill_2 FILLER_64_116 ();
 sg13g2_fill_1 FILLER_64_156 ();
 sg13g2_decap_4 FILLER_64_164 ();
 sg13g2_fill_2 FILLER_64_194 ();
 sg13g2_fill_2 FILLER_64_249 ();
 sg13g2_fill_1 FILLER_64_251 ();
 sg13g2_fill_1 FILLER_64_278 ();
 sg13g2_fill_1 FILLER_64_298 ();
 sg13g2_fill_1 FILLER_64_315 ();
 sg13g2_fill_2 FILLER_64_324 ();
 sg13g2_decap_8 FILLER_64_399 ();
 sg13g2_fill_2 FILLER_64_406 ();
 sg13g2_decap_8 FILLER_64_434 ();
 sg13g2_fill_2 FILLER_64_441 ();
 sg13g2_fill_2 FILLER_64_469 ();
 sg13g2_fill_2 FILLER_64_514 ();
 sg13g2_fill_2 FILLER_64_522 ();
 sg13g2_fill_1 FILLER_64_524 ();
 sg13g2_fill_2 FILLER_64_539 ();
 sg13g2_fill_1 FILLER_64_541 ();
 sg13g2_decap_8 FILLER_64_567 ();
 sg13g2_fill_1 FILLER_64_574 ();
 sg13g2_decap_4 FILLER_64_600 ();
 sg13g2_fill_2 FILLER_64_618 ();
 sg13g2_fill_1 FILLER_64_620 ();
 sg13g2_fill_2 FILLER_64_660 ();
 sg13g2_fill_1 FILLER_64_662 ();
 sg13g2_fill_1 FILLER_64_702 ();
 sg13g2_fill_2 FILLER_64_716 ();
 sg13g2_fill_1 FILLER_64_718 ();
 sg13g2_decap_8 FILLER_64_745 ();
 sg13g2_fill_2 FILLER_64_752 ();
 sg13g2_decap_8 FILLER_64_758 ();
 sg13g2_fill_2 FILLER_64_765 ();
 sg13g2_fill_1 FILLER_64_778 ();
 sg13g2_fill_2 FILLER_64_783 ();
 sg13g2_fill_1 FILLER_64_793 ();
 sg13g2_decap_8 FILLER_64_803 ();
 sg13g2_fill_2 FILLER_64_810 ();
 sg13g2_fill_1 FILLER_64_812 ();
 sg13g2_fill_2 FILLER_64_817 ();
 sg13g2_fill_2 FILLER_64_848 ();
 sg13g2_fill_1 FILLER_64_850 ();
 sg13g2_fill_2 FILLER_64_871 ();
 sg13g2_fill_2 FILLER_64_913 ();
 sg13g2_fill_2 FILLER_64_951 ();
 sg13g2_fill_1 FILLER_64_953 ();
 sg13g2_fill_1 FILLER_64_979 ();
 sg13g2_fill_2 FILLER_64_1017 ();
 sg13g2_fill_1 FILLER_64_1019 ();
 sg13g2_fill_1 FILLER_64_1030 ();
 sg13g2_decap_8 FILLER_64_1039 ();
 sg13g2_decap_8 FILLER_64_1046 ();
 sg13g2_fill_2 FILLER_64_1053 ();
 sg13g2_fill_1 FILLER_64_1055 ();
 sg13g2_fill_2 FILLER_64_1069 ();
 sg13g2_fill_1 FILLER_64_1071 ();
 sg13g2_fill_2 FILLER_64_1077 ();
 sg13g2_fill_1 FILLER_64_1079 ();
 sg13g2_decap_8 FILLER_64_1085 ();
 sg13g2_fill_2 FILLER_64_1096 ();
 sg13g2_fill_1 FILLER_64_1098 ();
 sg13g2_fill_1 FILLER_64_1104 ();
 sg13g2_fill_2 FILLER_64_1148 ();
 sg13g2_fill_2 FILLER_64_1187 ();
 sg13g2_fill_2 FILLER_64_1233 ();
 sg13g2_fill_1 FILLER_64_1235 ();
 sg13g2_fill_2 FILLER_64_1245 ();
 sg13g2_fill_1 FILLER_64_1247 ();
 sg13g2_fill_2 FILLER_64_1304 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_8 ();
 sg13g2_fill_1 FILLER_65_27 ();
 sg13g2_fill_1 FILLER_65_45 ();
 sg13g2_fill_1 FILLER_65_82 ();
 sg13g2_fill_2 FILLER_65_92 ();
 sg13g2_decap_8 FILLER_65_97 ();
 sg13g2_decap_8 FILLER_65_104 ();
 sg13g2_decap_4 FILLER_65_173 ();
 sg13g2_fill_2 FILLER_65_177 ();
 sg13g2_decap_4 FILLER_65_183 ();
 sg13g2_fill_1 FILLER_65_187 ();
 sg13g2_fill_2 FILLER_65_217 ();
 sg13g2_fill_2 FILLER_65_306 ();
 sg13g2_fill_1 FILLER_65_313 ();
 sg13g2_decap_4 FILLER_65_360 ();
 sg13g2_fill_2 FILLER_65_364 ();
 sg13g2_fill_1 FILLER_65_376 ();
 sg13g2_decap_8 FILLER_65_417 ();
 sg13g2_decap_4 FILLER_65_424 ();
 sg13g2_fill_1 FILLER_65_428 ();
 sg13g2_fill_1 FILLER_65_460 ();
 sg13g2_fill_2 FILLER_65_523 ();
 sg13g2_fill_1 FILLER_65_549 ();
 sg13g2_fill_1 FILLER_65_559 ();
 sg13g2_fill_1 FILLER_65_565 ();
 sg13g2_fill_1 FILLER_65_574 ();
 sg13g2_fill_2 FILLER_65_586 ();
 sg13g2_fill_1 FILLER_65_588 ();
 sg13g2_fill_1 FILLER_65_667 ();
 sg13g2_fill_2 FILLER_65_689 ();
 sg13g2_fill_2 FILLER_65_717 ();
 sg13g2_decap_8 FILLER_65_723 ();
 sg13g2_decap_4 FILLER_65_734 ();
 sg13g2_decap_4 FILLER_65_798 ();
 sg13g2_fill_1 FILLER_65_837 ();
 sg13g2_fill_2 FILLER_65_847 ();
 sg13g2_fill_2 FILLER_65_914 ();
 sg13g2_fill_1 FILLER_65_916 ();
 sg13g2_fill_2 FILLER_65_935 ();
 sg13g2_fill_1 FILLER_65_937 ();
 sg13g2_fill_2 FILLER_65_953 ();
 sg13g2_decap_4 FILLER_65_985 ();
 sg13g2_decap_8 FILLER_65_999 ();
 sg13g2_fill_1 FILLER_65_1020 ();
 sg13g2_fill_2 FILLER_65_1026 ();
 sg13g2_fill_2 FILLER_65_1071 ();
 sg13g2_fill_1 FILLER_65_1073 ();
 sg13g2_fill_2 FILLER_65_1269 ();
 sg13g2_fill_1 FILLER_65_1271 ();
 sg13g2_fill_2 FILLER_65_1286 ();
 sg13g2_fill_1 FILLER_65_1288 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_47 ();
 sg13g2_fill_1 FILLER_66_244 ();
 sg13g2_fill_2 FILLER_66_253 ();
 sg13g2_fill_1 FILLER_66_315 ();
 sg13g2_fill_1 FILLER_66_411 ();
 sg13g2_decap_8 FILLER_66_438 ();
 sg13g2_fill_2 FILLER_66_449 ();
 sg13g2_fill_1 FILLER_66_451 ();
 sg13g2_fill_2 FILLER_66_470 ();
 sg13g2_fill_2 FILLER_66_503 ();
 sg13g2_fill_2 FILLER_66_510 ();
 sg13g2_fill_1 FILLER_66_512 ();
 sg13g2_fill_1 FILLER_66_526 ();
 sg13g2_fill_2 FILLER_66_541 ();
 sg13g2_fill_2 FILLER_66_549 ();
 sg13g2_fill_1 FILLER_66_551 ();
 sg13g2_decap_4 FILLER_66_574 ();
 sg13g2_fill_1 FILLER_66_578 ();
 sg13g2_decap_8 FILLER_66_612 ();
 sg13g2_decap_8 FILLER_66_619 ();
 sg13g2_fill_2 FILLER_66_626 ();
 sg13g2_decap_4 FILLER_66_632 ();
 sg13g2_fill_1 FILLER_66_636 ();
 sg13g2_fill_2 FILLER_66_680 ();
 sg13g2_fill_1 FILLER_66_682 ();
 sg13g2_fill_1 FILLER_66_706 ();
 sg13g2_fill_1 FILLER_66_728 ();
 sg13g2_fill_1 FILLER_66_745 ();
 sg13g2_fill_2 FILLER_66_772 ();
 sg13g2_fill_1 FILLER_66_788 ();
 sg13g2_fill_1 FILLER_66_793 ();
 sg13g2_fill_2 FILLER_66_854 ();
 sg13g2_fill_1 FILLER_66_884 ();
 sg13g2_fill_1 FILLER_66_921 ();
 sg13g2_fill_1 FILLER_66_952 ();
 sg13g2_decap_8 FILLER_66_974 ();
 sg13g2_fill_1 FILLER_66_981 ();
 sg13g2_decap_4 FILLER_66_1004 ();
 sg13g2_fill_1 FILLER_66_1025 ();
 sg13g2_fill_2 FILLER_66_1045 ();
 sg13g2_fill_1 FILLER_66_1047 ();
 sg13g2_fill_2 FILLER_66_1057 ();
 sg13g2_fill_1 FILLER_66_1081 ();
 sg13g2_decap_8 FILLER_66_1087 ();
 sg13g2_decap_4 FILLER_66_1094 ();
 sg13g2_fill_1 FILLER_66_1098 ();
 sg13g2_fill_1 FILLER_66_1103 ();
 sg13g2_fill_2 FILLER_66_1107 ();
 sg13g2_fill_1 FILLER_66_1109 ();
 sg13g2_decap_8 FILLER_66_1119 ();
 sg13g2_decap_8 FILLER_66_1126 ();
 sg13g2_decap_4 FILLER_66_1133 ();
 sg13g2_fill_1 FILLER_66_1137 ();
 sg13g2_fill_2 FILLER_66_1210 ();
 sg13g2_fill_1 FILLER_66_1234 ();
 sg13g2_fill_2 FILLER_66_1287 ();
 sg13g2_decap_4 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_4 ();
 sg13g2_fill_1 FILLER_67_21 ();
 sg13g2_fill_1 FILLER_67_79 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_fill_2 FILLER_67_91 ();
 sg13g2_fill_2 FILLER_67_96 ();
 sg13g2_fill_1 FILLER_67_98 ();
 sg13g2_fill_2 FILLER_67_155 ();
 sg13g2_fill_1 FILLER_67_157 ();
 sg13g2_fill_1 FILLER_67_162 ();
 sg13g2_fill_1 FILLER_67_211 ();
 sg13g2_fill_2 FILLER_67_217 ();
 sg13g2_fill_2 FILLER_67_254 ();
 sg13g2_fill_1 FILLER_67_256 ();
 sg13g2_decap_8 FILLER_67_298 ();
 sg13g2_decap_4 FILLER_67_305 ();
 sg13g2_fill_1 FILLER_67_309 ();
 sg13g2_decap_8 FILLER_67_313 ();
 sg13g2_fill_2 FILLER_67_320 ();
 sg13g2_fill_1 FILLER_67_322 ();
 sg13g2_fill_1 FILLER_67_338 ();
 sg13g2_fill_2 FILLER_67_351 ();
 sg13g2_fill_1 FILLER_67_367 ();
 sg13g2_fill_2 FILLER_67_398 ();
 sg13g2_fill_1 FILLER_67_427 ();
 sg13g2_decap_8 FILLER_67_454 ();
 sg13g2_decap_4 FILLER_67_461 ();
 sg13g2_fill_1 FILLER_67_491 ();
 sg13g2_fill_1 FILLER_67_501 ();
 sg13g2_fill_2 FILLER_67_536 ();
 sg13g2_fill_1 FILLER_67_550 ();
 sg13g2_fill_1 FILLER_67_577 ();
 sg13g2_decap_4 FILLER_67_622 ();
 sg13g2_fill_1 FILLER_67_626 ();
 sg13g2_decap_8 FILLER_67_631 ();
 sg13g2_fill_1 FILLER_67_638 ();
 sg13g2_fill_1 FILLER_67_683 ();
 sg13g2_fill_2 FILLER_67_754 ();
 sg13g2_fill_1 FILLER_67_830 ();
 sg13g2_fill_1 FILLER_67_876 ();
 sg13g2_fill_2 FILLER_67_893 ();
 sg13g2_fill_2 FILLER_67_936 ();
 sg13g2_decap_8 FILLER_67_981 ();
 sg13g2_fill_2 FILLER_67_988 ();
 sg13g2_decap_4 FILLER_67_1000 ();
 sg13g2_fill_2 FILLER_67_1004 ();
 sg13g2_fill_2 FILLER_67_1028 ();
 sg13g2_fill_1 FILLER_67_1030 ();
 sg13g2_decap_8 FILLER_67_1045 ();
 sg13g2_fill_1 FILLER_67_1052 ();
 sg13g2_fill_2 FILLER_67_1073 ();
 sg13g2_fill_2 FILLER_67_1099 ();
 sg13g2_decap_8 FILLER_67_1147 ();
 sg13g2_fill_2 FILLER_67_1162 ();
 sg13g2_fill_1 FILLER_67_1164 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_fill_2 FILLER_68_29 ();
 sg13g2_fill_1 FILLER_68_31 ();
 sg13g2_fill_2 FILLER_68_137 ();
 sg13g2_fill_2 FILLER_68_171 ();
 sg13g2_fill_1 FILLER_68_244 ();
 sg13g2_fill_2 FILLER_68_269 ();
 sg13g2_fill_1 FILLER_68_271 ();
 sg13g2_fill_2 FILLER_68_290 ();
 sg13g2_decap_8 FILLER_68_298 ();
 sg13g2_fill_1 FILLER_68_368 ();
 sg13g2_fill_2 FILLER_68_429 ();
 sg13g2_decap_4 FILLER_68_465 ();
 sg13g2_fill_2 FILLER_68_469 ();
 sg13g2_fill_2 FILLER_68_540 ();
 sg13g2_fill_1 FILLER_68_568 ();
 sg13g2_fill_2 FILLER_68_593 ();
 sg13g2_fill_2 FILLER_68_686 ();
 sg13g2_fill_1 FILLER_68_688 ();
 sg13g2_fill_1 FILLER_68_730 ();
 sg13g2_fill_2 FILLER_68_762 ();
 sg13g2_fill_1 FILLER_68_769 ();
 sg13g2_fill_1 FILLER_68_789 ();
 sg13g2_fill_1 FILLER_68_818 ();
 sg13g2_fill_2 FILLER_68_925 ();
 sg13g2_fill_1 FILLER_68_927 ();
 sg13g2_decap_4 FILLER_68_979 ();
 sg13g2_fill_2 FILLER_68_983 ();
 sg13g2_fill_2 FILLER_68_1011 ();
 sg13g2_fill_1 FILLER_68_1018 ();
 sg13g2_decap_8 FILLER_68_1028 ();
 sg13g2_decap_8 FILLER_68_1035 ();
 sg13g2_decap_4 FILLER_68_1042 ();
 sg13g2_fill_2 FILLER_68_1046 ();
 sg13g2_fill_2 FILLER_68_1052 ();
 sg13g2_fill_2 FILLER_68_1059 ();
 sg13g2_fill_1 FILLER_68_1061 ();
 sg13g2_fill_2 FILLER_68_1067 ();
 sg13g2_fill_1 FILLER_68_1069 ();
 sg13g2_fill_2 FILLER_68_1074 ();
 sg13g2_fill_1 FILLER_68_1076 ();
 sg13g2_decap_4 FILLER_68_1086 ();
 sg13g2_decap_4 FILLER_68_1094 ();
 sg13g2_fill_1 FILLER_68_1098 ();
 sg13g2_fill_1 FILLER_68_1134 ();
 sg13g2_fill_1 FILLER_68_1171 ();
 sg13g2_fill_2 FILLER_68_1185 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_187 ();
 sg13g2_fill_1 FILLER_69_198 ();
 sg13g2_fill_2 FILLER_69_203 ();
 sg13g2_fill_2 FILLER_69_210 ();
 sg13g2_fill_1 FILLER_69_252 ();
 sg13g2_fill_1 FILLER_69_284 ();
 sg13g2_fill_2 FILLER_69_381 ();
 sg13g2_fill_1 FILLER_69_404 ();
 sg13g2_fill_2 FILLER_69_446 ();
 sg13g2_fill_1 FILLER_69_448 ();
 sg13g2_fill_2 FILLER_69_458 ();
 sg13g2_decap_4 FILLER_69_464 ();
 sg13g2_fill_1 FILLER_69_468 ();
 sg13g2_decap_4 FILLER_69_476 ();
 sg13g2_fill_2 FILLER_69_506 ();
 sg13g2_fill_1 FILLER_69_508 ();
 sg13g2_fill_1 FILLER_69_525 ();
 sg13g2_fill_1 FILLER_69_531 ();
 sg13g2_fill_1 FILLER_69_549 ();
 sg13g2_decap_4 FILLER_69_556 ();
 sg13g2_decap_8 FILLER_69_576 ();
 sg13g2_decap_4 FILLER_69_588 ();
 sg13g2_fill_1 FILLER_69_592 ();
 sg13g2_fill_2 FILLER_69_605 ();
 sg13g2_fill_2 FILLER_69_611 ();
 sg13g2_fill_2 FILLER_69_617 ();
 sg13g2_fill_1 FILLER_69_652 ();
 sg13g2_fill_2 FILLER_69_663 ();
 sg13g2_fill_1 FILLER_69_743 ();
 sg13g2_fill_2 FILLER_69_791 ();
 sg13g2_fill_2 FILLER_69_916 ();
 sg13g2_fill_1 FILLER_69_918 ();
 sg13g2_fill_2 FILLER_69_964 ();
 sg13g2_decap_4 FILLER_69_987 ();
 sg13g2_fill_1 FILLER_69_991 ();
 sg13g2_fill_2 FILLER_69_997 ();
 sg13g2_fill_1 FILLER_69_999 ();
 sg13g2_fill_2 FILLER_69_1043 ();
 sg13g2_fill_1 FILLER_69_1045 ();
 sg13g2_fill_2 FILLER_69_1066 ();
 sg13g2_fill_1 FILLER_69_1068 ();
 sg13g2_fill_1 FILLER_69_1077 ();
 sg13g2_fill_2 FILLER_69_1086 ();
 sg13g2_fill_1 FILLER_69_1096 ();
 sg13g2_fill_2 FILLER_69_1105 ();
 sg13g2_decap_8 FILLER_69_1120 ();
 sg13g2_fill_2 FILLER_69_1127 ();
 sg13g2_decap_4 FILLER_69_1133 ();
 sg13g2_fill_2 FILLER_69_1137 ();
 sg13g2_fill_1 FILLER_69_1166 ();
 sg13g2_fill_2 FILLER_69_1228 ();
 sg13g2_fill_2 FILLER_69_1287 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_40 ();
 sg13g2_fill_2 FILLER_70_125 ();
 sg13g2_fill_2 FILLER_70_153 ();
 sg13g2_fill_2 FILLER_70_181 ();
 sg13g2_fill_2 FILLER_70_201 ();
 sg13g2_fill_2 FILLER_70_207 ();
 sg13g2_fill_1 FILLER_70_231 ();
 sg13g2_fill_2 FILLER_70_245 ();
 sg13g2_fill_2 FILLER_70_252 ();
 sg13g2_fill_1 FILLER_70_267 ();
 sg13g2_fill_2 FILLER_70_323 ();
 sg13g2_fill_1 FILLER_70_357 ();
 sg13g2_fill_1 FILLER_70_362 ();
 sg13g2_fill_2 FILLER_70_394 ();
 sg13g2_fill_2 FILLER_70_526 ();
 sg13g2_fill_2 FILLER_70_534 ();
 sg13g2_decap_4 FILLER_70_553 ();
 sg13g2_fill_2 FILLER_70_557 ();
 sg13g2_fill_2 FILLER_70_573 ();
 sg13g2_fill_1 FILLER_70_584 ();
 sg13g2_decap_4 FILLER_70_611 ();
 sg13g2_fill_1 FILLER_70_615 ();
 sg13g2_fill_1 FILLER_70_624 ();
 sg13g2_fill_1 FILLER_70_634 ();
 sg13g2_fill_1 FILLER_70_644 ();
 sg13g2_fill_2 FILLER_70_658 ();
 sg13g2_fill_2 FILLER_70_694 ();
 sg13g2_fill_1 FILLER_70_809 ();
 sg13g2_fill_2 FILLER_70_844 ();
 sg13g2_fill_1 FILLER_70_846 ();
 sg13g2_fill_1 FILLER_70_874 ();
 sg13g2_fill_1 FILLER_70_931 ();
 sg13g2_fill_2 FILLER_70_966 ();
 sg13g2_decap_8 FILLER_70_994 ();
 sg13g2_fill_1 FILLER_70_1001 ();
 sg13g2_decap_8 FILLER_70_1029 ();
 sg13g2_decap_4 FILLER_70_1036 ();
 sg13g2_fill_2 FILLER_70_1040 ();
 sg13g2_decap_4 FILLER_70_1051 ();
 sg13g2_fill_1 FILLER_70_1068 ();
 sg13g2_decap_8 FILLER_70_1082 ();
 sg13g2_decap_8 FILLER_70_1089 ();
 sg13g2_fill_2 FILLER_70_1096 ();
 sg13g2_fill_1 FILLER_70_1098 ();
 sg13g2_fill_2 FILLER_70_1104 ();
 sg13g2_decap_4 FILLER_70_1114 ();
 sg13g2_fill_1 FILLER_70_1118 ();
 sg13g2_fill_2 FILLER_70_1145 ();
 sg13g2_fill_1 FILLER_70_1147 ();
 sg13g2_fill_2 FILLER_70_1191 ();
 sg13g2_fill_1 FILLER_70_1206 ();
 sg13g2_fill_2 FILLER_70_1269 ();
 sg13g2_fill_2 FILLER_70_1297 ();
 sg13g2_fill_1 FILLER_70_1299 ();
 sg13g2_fill_2 FILLER_70_1313 ();
 sg13g2_fill_1 FILLER_71_90 ();
 sg13g2_fill_1 FILLER_71_121 ();
 sg13g2_fill_2 FILLER_71_127 ();
 sg13g2_fill_1 FILLER_71_135 ();
 sg13g2_fill_1 FILLER_71_140 ();
 sg13g2_fill_1 FILLER_71_149 ();
 sg13g2_fill_2 FILLER_71_176 ();
 sg13g2_fill_2 FILLER_71_247 ();
 sg13g2_fill_1 FILLER_71_249 ();
 sg13g2_fill_2 FILLER_71_255 ();
 sg13g2_fill_1 FILLER_71_266 ();
 sg13g2_fill_1 FILLER_71_363 ();
 sg13g2_fill_2 FILLER_71_378 ();
 sg13g2_fill_2 FILLER_71_389 ();
 sg13g2_fill_1 FILLER_71_432 ();
 sg13g2_fill_1 FILLER_71_459 ();
 sg13g2_fill_2 FILLER_71_469 ();
 sg13g2_fill_2 FILLER_71_476 ();
 sg13g2_fill_2 FILLER_71_492 ();
 sg13g2_fill_1 FILLER_71_528 ();
 sg13g2_fill_1 FILLER_71_544 ();
 sg13g2_fill_1 FILLER_71_588 ();
 sg13g2_fill_1 FILLER_71_597 ();
 sg13g2_fill_1 FILLER_71_608 ();
 sg13g2_decap_4 FILLER_71_614 ();
 sg13g2_decap_8 FILLER_71_632 ();
 sg13g2_fill_1 FILLER_71_643 ();
 sg13g2_fill_1 FILLER_71_712 ();
 sg13g2_fill_1 FILLER_71_744 ();
 sg13g2_fill_2 FILLER_71_771 ();
 sg13g2_fill_2 FILLER_71_791 ();
 sg13g2_fill_2 FILLER_71_830 ();
 sg13g2_fill_2 FILLER_71_862 ();
 sg13g2_fill_2 FILLER_71_875 ();
 sg13g2_fill_1 FILLER_71_877 ();
 sg13g2_fill_1 FILLER_71_921 ();
 sg13g2_fill_2 FILLER_71_959 ();
 sg13g2_fill_1 FILLER_71_961 ();
 sg13g2_fill_1 FILLER_71_987 ();
 sg13g2_decap_4 FILLER_71_997 ();
 sg13g2_fill_2 FILLER_71_1001 ();
 sg13g2_fill_2 FILLER_71_1007 ();
 sg13g2_decap_8 FILLER_71_1027 ();
 sg13g2_fill_2 FILLER_71_1054 ();
 sg13g2_fill_1 FILLER_71_1056 ();
 sg13g2_fill_2 FILLER_71_1069 ();
 sg13g2_fill_1 FILLER_71_1088 ();
 sg13g2_fill_1 FILLER_71_1101 ();
 sg13g2_decap_8 FILLER_71_1123 ();
 sg13g2_decap_4 FILLER_71_1130 ();
 sg13g2_fill_1 FILLER_71_1134 ();
 sg13g2_fill_2 FILLER_71_1138 ();
 sg13g2_fill_1 FILLER_71_1140 ();
 sg13g2_fill_1 FILLER_71_1154 ();
 sg13g2_fill_2 FILLER_71_1224 ();
 sg13g2_fill_2 FILLER_71_1304 ();
 sg13g2_fill_2 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_93 ();
 sg13g2_fill_2 FILLER_72_114 ();
 sg13g2_fill_1 FILLER_72_161 ();
 sg13g2_fill_2 FILLER_72_181 ();
 sg13g2_fill_1 FILLER_72_194 ();
 sg13g2_fill_2 FILLER_72_201 ();
 sg13g2_fill_1 FILLER_72_216 ();
 sg13g2_fill_2 FILLER_72_227 ();
 sg13g2_fill_1 FILLER_72_242 ();
 sg13g2_fill_1 FILLER_72_302 ();
 sg13g2_fill_2 FILLER_72_311 ();
 sg13g2_fill_1 FILLER_72_437 ();
 sg13g2_fill_1 FILLER_72_448 ();
 sg13g2_decap_4 FILLER_72_475 ();
 sg13g2_fill_2 FILLER_72_531 ();
 sg13g2_fill_2 FILLER_72_557 ();
 sg13g2_fill_2 FILLER_72_564 ();
 sg13g2_fill_1 FILLER_72_570 ();
 sg13g2_decap_4 FILLER_72_586 ();
 sg13g2_fill_2 FILLER_72_594 ();
 sg13g2_fill_2 FILLER_72_609 ();
 sg13g2_fill_1 FILLER_72_611 ();
 sg13g2_fill_1 FILLER_72_621 ();
 sg13g2_fill_1 FILLER_72_687 ();
 sg13g2_fill_1 FILLER_72_778 ();
 sg13g2_fill_1 FILLER_72_810 ();
 sg13g2_fill_1 FILLER_72_853 ();
 sg13g2_fill_1 FILLER_72_865 ();
 sg13g2_fill_2 FILLER_72_928 ();
 sg13g2_fill_1 FILLER_72_930 ();
 sg13g2_fill_2 FILLER_72_966 ();
 sg13g2_fill_1 FILLER_72_968 ();
 sg13g2_decap_4 FILLER_72_1032 ();
 sg13g2_fill_1 FILLER_72_1036 ();
 sg13g2_decap_4 FILLER_72_1048 ();
 sg13g2_fill_1 FILLER_72_1081 ();
 sg13g2_decap_4 FILLER_72_1094 ();
 sg13g2_fill_1 FILLER_72_1102 ();
 sg13g2_decap_4 FILLER_72_1108 ();
 sg13g2_fill_1 FILLER_72_1112 ();
 sg13g2_fill_2 FILLER_72_1126 ();
 sg13g2_fill_1 FILLER_72_1128 ();
 sg13g2_fill_2 FILLER_72_1156 ();
 sg13g2_fill_1 FILLER_72_1158 ();
 sg13g2_fill_2 FILLER_72_1168 ();
 sg13g2_fill_1 FILLER_72_1170 ();
 sg13g2_fill_2 FILLER_72_1245 ();
 sg13g2_fill_2 FILLER_72_1286 ();
 sg13g2_fill_1 FILLER_72_1288 ();
 sg13g2_fill_1 FILLER_73_117 ();
 sg13g2_fill_2 FILLER_73_199 ();
 sg13g2_fill_1 FILLER_73_214 ();
 sg13g2_fill_2 FILLER_73_298 ();
 sg13g2_fill_2 FILLER_73_319 ();
 sg13g2_fill_2 FILLER_73_392 ();
 sg13g2_fill_1 FILLER_73_410 ();
 sg13g2_fill_2 FILLER_73_442 ();
 sg13g2_fill_1 FILLER_73_478 ();
 sg13g2_decap_8 FILLER_73_484 ();
 sg13g2_fill_2 FILLER_73_491 ();
 sg13g2_decap_8 FILLER_73_506 ();
 sg13g2_fill_1 FILLER_73_530 ();
 sg13g2_fill_1 FILLER_73_553 ();
 sg13g2_fill_1 FILLER_73_624 ();
 sg13g2_fill_2 FILLER_73_656 ();
 sg13g2_fill_1 FILLER_73_733 ();
 sg13g2_fill_1 FILLER_73_782 ();
 sg13g2_fill_2 FILLER_73_816 ();
 sg13g2_fill_1 FILLER_73_837 ();
 sg13g2_fill_1 FILLER_73_920 ();
 sg13g2_fill_1 FILLER_73_941 ();
 sg13g2_fill_1 FILLER_73_968 ();
 sg13g2_fill_2 FILLER_73_974 ();
 sg13g2_fill_1 FILLER_73_976 ();
 sg13g2_decap_4 FILLER_73_1027 ();
 sg13g2_fill_1 FILLER_73_1031 ();
 sg13g2_fill_1 FILLER_73_1046 ();
 sg13g2_decap_4 FILLER_73_1064 ();
 sg13g2_decap_4 FILLER_73_1077 ();
 sg13g2_fill_1 FILLER_73_1081 ();
 sg13g2_fill_1 FILLER_73_1103 ();
 sg13g2_fill_1 FILLER_73_1117 ();
 sg13g2_fill_2 FILLER_73_1144 ();
 sg13g2_fill_1 FILLER_73_1206 ();
 sg13g2_fill_2 FILLER_73_1312 ();
 sg13g2_fill_1 FILLER_73_1314 ();
 sg13g2_fill_1 FILLER_74_82 ();
 sg13g2_fill_1 FILLER_74_113 ();
 sg13g2_fill_1 FILLER_74_153 ();
 sg13g2_fill_1 FILLER_74_167 ();
 sg13g2_fill_2 FILLER_74_194 ();
 sg13g2_fill_2 FILLER_74_322 ();
 sg13g2_fill_1 FILLER_74_334 ();
 sg13g2_fill_1 FILLER_74_394 ();
 sg13g2_fill_2 FILLER_74_435 ();
 sg13g2_fill_1 FILLER_74_437 ();
 sg13g2_fill_1 FILLER_74_447 ();
 sg13g2_fill_2 FILLER_74_475 ();
 sg13g2_fill_1 FILLER_74_477 ();
 sg13g2_decap_4 FILLER_74_482 ();
 sg13g2_fill_2 FILLER_74_486 ();
 sg13g2_decap_8 FILLER_74_494 ();
 sg13g2_fill_2 FILLER_74_524 ();
 sg13g2_fill_1 FILLER_74_584 ();
 sg13g2_fill_1 FILLER_74_602 ();
 sg13g2_decap_4 FILLER_74_613 ();
 sg13g2_fill_1 FILLER_74_617 ();
 sg13g2_fill_2 FILLER_74_629 ();
 sg13g2_decap_4 FILLER_74_654 ();
 sg13g2_fill_2 FILLER_74_717 ();
 sg13g2_fill_1 FILLER_74_848 ();
 sg13g2_fill_1 FILLER_74_900 ();
 sg13g2_fill_1 FILLER_74_973 ();
 sg13g2_fill_1 FILLER_74_988 ();
 sg13g2_fill_2 FILLER_74_1028 ();
 sg13g2_fill_1 FILLER_74_1030 ();
 sg13g2_fill_1 FILLER_74_1069 ();
 sg13g2_decap_8 FILLER_74_1082 ();
 sg13g2_decap_8 FILLER_74_1089 ();
 sg13g2_fill_2 FILLER_74_1096 ();
 sg13g2_fill_1 FILLER_74_1098 ();
 sg13g2_fill_2 FILLER_74_1112 ();
 sg13g2_decap_4 FILLER_74_1122 ();
 sg13g2_fill_2 FILLER_74_1126 ();
 sg13g2_fill_1 FILLER_74_1202 ();
 sg13g2_fill_2 FILLER_74_1207 ();
 sg13g2_fill_1 FILLER_74_1209 ();
 sg13g2_fill_2 FILLER_75_30 ();
 sg13g2_fill_1 FILLER_75_62 ();
 sg13g2_fill_2 FILLER_75_102 ();
 sg13g2_fill_1 FILLER_75_113 ();
 sg13g2_fill_1 FILLER_75_188 ();
 sg13g2_fill_1 FILLER_75_260 ();
 sg13g2_fill_2 FILLER_75_282 ();
 sg13g2_fill_1 FILLER_75_323 ();
 sg13g2_fill_2 FILLER_75_338 ();
 sg13g2_fill_2 FILLER_75_383 ();
 sg13g2_fill_2 FILLER_75_439 ();
 sg13g2_fill_1 FILLER_75_441 ();
 sg13g2_fill_1 FILLER_75_492 ();
 sg13g2_fill_1 FILLER_75_541 ();
 sg13g2_decap_8 FILLER_75_648 ();
 sg13g2_decap_4 FILLER_75_655 ();
 sg13g2_fill_1 FILLER_75_667 ();
 sg13g2_fill_2 FILLER_75_681 ();
 sg13g2_fill_1 FILLER_75_714 ();
 sg13g2_fill_2 FILLER_75_733 ();
 sg13g2_fill_2 FILLER_75_752 ();
 sg13g2_fill_2 FILLER_75_797 ();
 sg13g2_fill_2 FILLER_75_865 ();
 sg13g2_fill_2 FILLER_75_878 ();
 sg13g2_fill_2 FILLER_75_919 ();
 sg13g2_fill_1 FILLER_75_926 ();
 sg13g2_fill_1 FILLER_75_946 ();
 sg13g2_fill_2 FILLER_75_987 ();
 sg13g2_fill_1 FILLER_75_1009 ();
 sg13g2_fill_2 FILLER_75_1027 ();
 sg13g2_fill_2 FILLER_75_1053 ();
 sg13g2_fill_1 FILLER_75_1055 ();
 sg13g2_fill_2 FILLER_75_1069 ();
 sg13g2_decap_4 FILLER_75_1084 ();
 sg13g2_decap_8 FILLER_75_1100 ();
 sg13g2_fill_1 FILLER_75_1107 ();
 sg13g2_fill_2 FILLER_75_1157 ();
 sg13g2_fill_2 FILLER_75_1229 ();
 sg13g2_fill_2 FILLER_75_1266 ();
 sg13g2_fill_1 FILLER_75_1273 ();
 sg13g2_fill_2 FILLER_75_1304 ();
 sg13g2_fill_1 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_22 ();
 sg13g2_fill_2 FILLER_76_68 ();
 sg13g2_fill_1 FILLER_76_70 ();
 sg13g2_fill_1 FILLER_76_98 ();
 sg13g2_fill_1 FILLER_76_137 ();
 sg13g2_fill_1 FILLER_76_196 ();
 sg13g2_fill_2 FILLER_76_328 ();
 sg13g2_fill_2 FILLER_76_356 ();
 sg13g2_fill_1 FILLER_76_403 ();
 sg13g2_fill_1 FILLER_76_435 ();
 sg13g2_fill_2 FILLER_76_462 ();
 sg13g2_fill_1 FILLER_76_481 ();
 sg13g2_fill_2 FILLER_76_487 ();
 sg13g2_fill_2 FILLER_76_506 ();
 sg13g2_fill_2 FILLER_76_538 ();
 sg13g2_fill_1 FILLER_76_540 ();
 sg13g2_fill_1 FILLER_76_576 ();
 sg13g2_fill_2 FILLER_76_597 ();
 sg13g2_fill_1 FILLER_76_618 ();
 sg13g2_fill_1 FILLER_76_623 ();
 sg13g2_fill_2 FILLER_76_629 ();
 sg13g2_fill_1 FILLER_76_647 ();
 sg13g2_fill_1 FILLER_76_674 ();
 sg13g2_fill_2 FILLER_76_684 ();
 sg13g2_fill_1 FILLER_76_783 ();
 sg13g2_fill_2 FILLER_76_803 ();
 sg13g2_fill_1 FILLER_76_837 ();
 sg13g2_fill_2 FILLER_76_847 ();
 sg13g2_fill_1 FILLER_76_933 ();
 sg13g2_fill_1 FILLER_76_1001 ();
 sg13g2_fill_1 FILLER_76_1047 ();
 sg13g2_decap_8 FILLER_76_1084 ();
 sg13g2_fill_2 FILLER_76_1091 ();
 sg13g2_fill_1 FILLER_76_1093 ();
 sg13g2_fill_2 FILLER_76_1107 ();
 sg13g2_fill_1 FILLER_76_1109 ();
 sg13g2_decap_8 FILLER_76_1120 ();
 sg13g2_fill_1 FILLER_76_1127 ();
 sg13g2_fill_1 FILLER_76_1136 ();
 sg13g2_fill_1 FILLER_76_1154 ();
 sg13g2_fill_1 FILLER_76_1194 ();
 sg13g2_fill_2 FILLER_76_1213 ();
 sg13g2_fill_1 FILLER_76_1215 ();
 sg13g2_fill_2 FILLER_76_1247 ();
 sg13g2_fill_1 FILLER_76_1249 ();
 sg13g2_fill_1 FILLER_77_26 ();
 sg13g2_fill_2 FILLER_77_178 ();
 sg13g2_fill_2 FILLER_77_204 ();
 sg13g2_fill_1 FILLER_77_216 ();
 sg13g2_fill_1 FILLER_77_235 ();
 sg13g2_fill_1 FILLER_77_428 ();
 sg13g2_fill_1 FILLER_77_448 ();
 sg13g2_fill_2 FILLER_77_473 ();
 sg13g2_fill_2 FILLER_77_512 ();
 sg13g2_fill_1 FILLER_77_551 ();
 sg13g2_fill_1 FILLER_77_556 ();
 sg13g2_fill_2 FILLER_77_585 ();
 sg13g2_fill_1 FILLER_77_668 ();
 sg13g2_fill_2 FILLER_77_706 ();
 sg13g2_fill_1 FILLER_77_708 ();
 sg13g2_fill_1 FILLER_77_783 ();
 sg13g2_fill_1 FILLER_77_866 ();
 sg13g2_fill_2 FILLER_77_903 ();
 sg13g2_fill_1 FILLER_77_905 ();
 sg13g2_fill_1 FILLER_77_916 ();
 sg13g2_fill_2 FILLER_77_935 ();
 sg13g2_fill_1 FILLER_77_937 ();
 sg13g2_fill_1 FILLER_77_952 ();
 sg13g2_fill_1 FILLER_77_1068 ();
 sg13g2_fill_1 FILLER_77_1079 ();
 sg13g2_fill_2 FILLER_77_1105 ();
 sg13g2_fill_1 FILLER_77_1107 ();
 sg13g2_fill_1 FILLER_77_1116 ();
 sg13g2_fill_1 FILLER_77_1143 ();
 sg13g2_fill_1 FILLER_77_1179 ();
 sg13g2_fill_2 FILLER_77_1276 ();
 sg13g2_fill_2 FILLER_77_1313 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_2 ();
 sg13g2_fill_2 FILLER_78_22 ();
 sg13g2_fill_1 FILLER_78_24 ();
 sg13g2_fill_1 FILLER_78_44 ();
 sg13g2_fill_2 FILLER_78_59 ();
 sg13g2_fill_1 FILLER_78_105 ();
 sg13g2_fill_1 FILLER_78_116 ();
 sg13g2_fill_1 FILLER_78_164 ();
 sg13g2_fill_1 FILLER_78_263 ();
 sg13g2_fill_2 FILLER_78_303 ();
 sg13g2_fill_1 FILLER_78_314 ();
 sg13g2_fill_1 FILLER_78_354 ();
 sg13g2_fill_1 FILLER_78_364 ();
 sg13g2_fill_1 FILLER_78_388 ();
 sg13g2_fill_1 FILLER_78_495 ();
 sg13g2_fill_1 FILLER_78_517 ();
 sg13g2_fill_1 FILLER_78_532 ();
 sg13g2_fill_2 FILLER_78_589 ();
 sg13g2_fill_2 FILLER_78_606 ();
 sg13g2_fill_1 FILLER_78_627 ();
 sg13g2_fill_1 FILLER_78_668 ();
 sg13g2_fill_1 FILLER_78_687 ();
 sg13g2_fill_1 FILLER_78_779 ();
 sg13g2_fill_2 FILLER_78_839 ();
 sg13g2_fill_2 FILLER_78_864 ();
 sg13g2_fill_1 FILLER_78_866 ();
 sg13g2_fill_1 FILLER_78_886 ();
 sg13g2_fill_2 FILLER_78_915 ();
 sg13g2_fill_1 FILLER_78_970 ();
 sg13g2_fill_2 FILLER_78_1023 ();
 sg13g2_fill_1 FILLER_78_1025 ();
 sg13g2_fill_1 FILLER_78_1033 ();
 sg13g2_fill_2 FILLER_78_1058 ();
 sg13g2_fill_2 FILLER_78_1068 ();
 sg13g2_fill_1 FILLER_78_1070 ();
 sg13g2_decap_8 FILLER_78_1113 ();
 sg13g2_decap_4 FILLER_78_1120 ();
 sg13g2_fill_2 FILLER_78_1158 ();
 sg13g2_fill_1 FILLER_78_1160 ();
 sg13g2_fill_2 FILLER_78_1196 ();
 sg13g2_fill_2 FILLER_78_1233 ();
 sg13g2_fill_1 FILLER_78_1235 ();
 sg13g2_fill_1 FILLER_78_1305 ();
 sg13g2_fill_1 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_36 ();
 sg13g2_fill_1 FILLER_79_202 ();
 sg13g2_fill_2 FILLER_79_234 ();
 sg13g2_fill_1 FILLER_79_279 ();
 sg13g2_fill_1 FILLER_79_345 ();
 sg13g2_fill_2 FILLER_79_372 ();
 sg13g2_fill_1 FILLER_79_427 ();
 sg13g2_fill_2 FILLER_79_454 ();
 sg13g2_fill_1 FILLER_79_605 ();
 sg13g2_fill_2 FILLER_79_668 ();
 sg13g2_fill_2 FILLER_79_675 ();
 sg13g2_fill_2 FILLER_79_691 ();
 sg13g2_fill_1 FILLER_79_754 ();
 sg13g2_fill_2 FILLER_79_808 ();
 sg13g2_fill_1 FILLER_79_810 ();
 sg13g2_fill_2 FILLER_79_837 ();
 sg13g2_fill_1 FILLER_79_910 ();
 sg13g2_fill_1 FILLER_79_921 ();
 sg13g2_fill_1 FILLER_79_927 ();
 sg13g2_fill_1 FILLER_79_984 ();
 sg13g2_fill_2 FILLER_79_1034 ();
 sg13g2_fill_1 FILLER_79_1067 ();
 sg13g2_fill_2 FILLER_79_1172 ();
 sg13g2_fill_1 FILLER_79_1174 ();
 sg13g2_fill_1 FILLER_79_1189 ();
 sg13g2_fill_2 FILLER_79_1255 ();
 sg13g2_fill_1 FILLER_79_1257 ();
 sg13g2_fill_2 FILLER_79_1275 ();
 sg13g2_fill_2 FILLER_79_1286 ();
 sg13g2_fill_1 FILLER_79_1288 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_86 ();
 sg13g2_fill_2 FILLER_80_122 ();
 sg13g2_fill_1 FILLER_80_147 ();
 sg13g2_fill_1 FILLER_80_226 ();
 sg13g2_fill_2 FILLER_80_381 ();
 sg13g2_fill_2 FILLER_80_437 ();
 sg13g2_fill_2 FILLER_80_492 ();
 sg13g2_fill_1 FILLER_80_494 ();
 sg13g2_decap_8 FILLER_80_502 ();
 sg13g2_decap_4 FILLER_80_509 ();
 sg13g2_fill_2 FILLER_80_517 ();
 sg13g2_fill_1 FILLER_80_519 ();
 sg13g2_fill_1 FILLER_80_525 ();
 sg13g2_fill_1 FILLER_80_541 ();
 sg13g2_fill_2 FILLER_80_576 ();
 sg13g2_fill_1 FILLER_80_598 ();
 sg13g2_fill_2 FILLER_80_608 ();
 sg13g2_fill_2 FILLER_80_626 ();
 sg13g2_fill_2 FILLER_80_706 ();
 sg13g2_fill_2 FILLER_80_717 ();
 sg13g2_fill_1 FILLER_80_746 ();
 sg13g2_fill_2 FILLER_80_752 ();
 sg13g2_fill_1 FILLER_80_777 ();
 sg13g2_fill_2 FILLER_80_839 ();
 sg13g2_fill_1 FILLER_80_841 ();
 sg13g2_fill_2 FILLER_80_864 ();
 sg13g2_fill_1 FILLER_80_866 ();
 sg13g2_fill_2 FILLER_80_876 ();
 sg13g2_fill_1 FILLER_80_878 ();
 sg13g2_fill_1 FILLER_80_897 ();
 sg13g2_fill_2 FILLER_80_1023 ();
 sg13g2_decap_8 FILLER_80_1055 ();
 sg13g2_fill_2 FILLER_80_1072 ();
 sg13g2_fill_2 FILLER_80_1090 ();
 sg13g2_fill_1 FILLER_80_1092 ();
 sg13g2_decap_8 FILLER_80_1096 ();
 sg13g2_decap_4 FILLER_80_1107 ();
 sg13g2_fill_1 FILLER_80_1111 ();
 sg13g2_decap_8 FILLER_80_1115 ();
 sg13g2_decap_4 FILLER_80_1126 ();
 sg13g2_decap_8 FILLER_80_1133 ();
 sg13g2_fill_2 FILLER_80_1140 ();
 sg13g2_fill_1 FILLER_80_1142 ();
 sg13g2_fill_2 FILLER_80_1147 ();
 sg13g2_fill_1 FILLER_80_1149 ();
 sg13g2_fill_2 FILLER_80_1162 ();
 sg13g2_fill_1 FILLER_80_1164 ();
 sg13g2_fill_2 FILLER_80_1229 ();
 sg13g2_fill_1 FILLER_80_1231 ();
 sg13g2_fill_2 FILLER_80_1257 ();
 sg13g2_fill_1 FILLER_80_1279 ();
 sg13g2_fill_1 FILLER_80_1284 ();
 sg13g2_fill_2 FILLER_80_1293 ();
 sg13g2_fill_1 FILLER_80_1295 ();
 sg13g2_fill_2 FILLER_80_1304 ();
endmodule

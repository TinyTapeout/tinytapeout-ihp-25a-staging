module tt_um_reemashivva_fifo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire clknet_0_clk;
 wire \clk_div_inst.r_clk ;
 wire \clk_div_inst.rd_counter[0] ;
 wire \clk_div_inst.rd_counter[1] ;
 wire \clk_div_inst.rd_counter[2] ;
 wire \clk_div_inst.w_clk ;
 wire \clk_div_inst.wr_counter[0] ;
 wire \clk_div_inst.wr_counter[1] ;
 wire \clk_div_inst.wr_counter[2] ;
 wire empty;
 wire \empty_inst.bin[0] ;
 wire \empty_inst.bin[1] ;
 wire \empty_inst.bin[2] ;
 wire \empty_inst.bin[3] ;
 wire \empty_inst.binnext[0] ;
 wire \empty_inst.binnext[1] ;
 wire \empty_inst.binnext[2] ;
 wire \empty_inst.binnext[3] ;
 wire \empty_inst.graynext[0] ;
 wire \empty_inst.graynext[1] ;
 wire \empty_inst.graynext[2] ;
 wire \empty_inst.rptr[0] ;
 wire \empty_inst.rptr[1] ;
 wire \empty_inst.rptr[2] ;
 wire \empty_inst.rsync_ptr2[0] ;
 wire \empty_inst.rsync_ptr2[1] ;
 wire \empty_inst.rsync_ptr2[2] ;
 wire \empty_inst.rsync_ptr2[3] ;
 wire \fifomem_inst.fifo[0][0] ;
 wire \fifomem_inst.fifo[0][1] ;
 wire \fifomem_inst.fifo[0][2] ;
 wire \fifomem_inst.fifo[0][3] ;
 wire \fifomem_inst.fifo[1][0] ;
 wire \fifomem_inst.fifo[1][1] ;
 wire \fifomem_inst.fifo[1][2] ;
 wire \fifomem_inst.fifo[1][3] ;
 wire \fifomem_inst.fifo[2][0] ;
 wire \fifomem_inst.fifo[2][1] ;
 wire \fifomem_inst.fifo[2][2] ;
 wire \fifomem_inst.fifo[2][3] ;
 wire \fifomem_inst.fifo[3][0] ;
 wire \fifomem_inst.fifo[3][1] ;
 wire \fifomem_inst.fifo[3][2] ;
 wire \fifomem_inst.fifo[3][3] ;
 wire \fifomem_inst.fifo[4][0] ;
 wire \fifomem_inst.fifo[4][1] ;
 wire \fifomem_inst.fifo[4][2] ;
 wire \fifomem_inst.fifo[4][3] ;
 wire \fifomem_inst.fifo[5][0] ;
 wire \fifomem_inst.fifo[5][1] ;
 wire \fifomem_inst.fifo[5][2] ;
 wire \fifomem_inst.fifo[5][3] ;
 wire \fifomem_inst.fifo[6][0] ;
 wire \fifomem_inst.fifo[6][1] ;
 wire \fifomem_inst.fifo[6][2] ;
 wire \fifomem_inst.fifo[6][3] ;
 wire \fifomem_inst.fifo[7][0] ;
 wire \fifomem_inst.fifo[7][1] ;
 wire \fifomem_inst.fifo[7][2] ;
 wire \fifomem_inst.fifo[7][3] ;
 wire \fifomem_inst.full ;
 wire \fifomem_inst.waddr[0] ;
 wire \fifomem_inst.waddr[1] ;
 wire \fifomem_inst.waddr[2] ;
 wire \full_inst.bin[3] ;
 wire \full_inst.binnext[0] ;
 wire \full_inst.binnext[1] ;
 wire \full_inst.binnext[2] ;
 wire \full_inst.binnext[3] ;
 wire \full_inst.fulln ;
 wire \full_inst.graynext[0] ;
 wire \full_inst.graynext[1] ;
 wire \full_inst.graynext[2] ;
 wire \full_inst.wptr[0] ;
 wire \full_inst.wptr[1] ;
 wire \full_inst.wptr[2] ;
 wire \full_inst.wsync_ptr2[0] ;
 wire \full_inst.wsync_ptr2[1] ;
 wire \full_inst.wsync_ptr2[2] ;
 wire \full_inst.wsync_ptr2[3] ;
 wire \sync_r2w_inst.wsync_ptr1[0] ;
 wire \sync_r2w_inst.wsync_ptr1[1] ;
 wire \sync_r2w_inst.wsync_ptr1[2] ;
 wire \sync_r2w_inst.wsync_ptr1[3] ;
 wire \sync_w2r_inst.rsync_ptr1[0] ;
 wire \sync_w2r_inst.rsync_ptr1[1] ;
 wire \sync_w2r_inst.rsync_ptr1[2] ;
 wire \sync_w2r_inst.rsync_ptr1[3] ;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;

 sg13g2_inv_1 _228_ (.Y(_003_),
    .A(net65));
 sg13g2_inv_2 _229_ (.Y(_052_),
    .A(net77));
 sg13g2_nand2b_2 _230_ (.Y(_053_),
    .B(net2),
    .A_N(empty));
 sg13g2_nor2_1 _231_ (.A(_007_),
    .B(_053_),
    .Y(_054_));
 sg13g2_nor3_1 _232_ (.A(_052_),
    .B(_007_),
    .C(_053_),
    .Y(_055_));
 sg13g2_nor4_1 _233_ (.A(_052_),
    .B(_007_),
    .C(_009_),
    .D(_053_),
    .Y(_056_));
 sg13g2_xnor2_1 _234_ (.Y(_057_),
    .A(\empty_inst.bin[3] ),
    .B(_056_));
 sg13g2_inv_1 _235_ (.Y(\empty_inst.binnext[3] ),
    .A(_057_));
 sg13g2_xnor2_1 _236_ (.Y(_058_),
    .A(net76),
    .B(_055_));
 sg13g2_inv_1 _237_ (.Y(\empty_inst.binnext[2] ),
    .A(_058_));
 sg13g2_xor2_1 _238_ (.B(_058_),
    .A(_057_),
    .X(\empty_inst.graynext[2] ));
 sg13g2_xnor2_1 _239_ (.Y(_059_),
    .A(\empty_inst.rsync_ptr2[2] ),
    .B(\empty_inst.graynext[2] ));
 sg13g2_xnor2_1 _240_ (.Y(\empty_inst.binnext[0] ),
    .A(net79),
    .B(_053_));
 sg13g2_xnor2_1 _241_ (.Y(\empty_inst.binnext[1] ),
    .A(_008_),
    .B(_054_));
 sg13g2_xor2_1 _242_ (.B(\empty_inst.binnext[1] ),
    .A(\empty_inst.binnext[0] ),
    .X(\empty_inst.graynext[0] ));
 sg13g2_xnor2_1 _243_ (.Y(_060_),
    .A(\empty_inst.rsync_ptr2[0] ),
    .B(\empty_inst.graynext[0] ));
 sg13g2_xor2_1 _244_ (.B(_057_),
    .A(\empty_inst.rsync_ptr2[3] ),
    .X(_061_));
 sg13g2_xnor2_1 _245_ (.Y(\empty_inst.graynext[1] ),
    .A(_058_),
    .B(\empty_inst.binnext[1] ));
 sg13g2_xnor2_1 _246_ (.Y(_062_),
    .A(\empty_inst.rsync_ptr2[1] ),
    .B(\empty_inst.graynext[1] ));
 sg13g2_nand4_1 _247_ (.B(_060_),
    .C(_061_),
    .A(_059_),
    .Y(_013_),
    .D(_062_));
 sg13g2_nor2b_2 _248_ (.A(\fifomem_inst.full ),
    .B_N(net1),
    .Y(_063_));
 sg13g2_nand2_1 _249_ (.Y(_064_),
    .A(\fifomem_inst.waddr[0] ),
    .B(_063_));
 sg13g2_nand3_1 _250_ (.B(net80),
    .C(_063_),
    .A(\fifomem_inst.waddr[0] ),
    .Y(_065_));
 sg13g2_a21oi_1 _251_ (.A1(\fifomem_inst.waddr[0] ),
    .A2(_063_),
    .Y(_066_),
    .B1(net80));
 sg13g2_xnor2_1 _252_ (.Y(\full_inst.binnext[1] ),
    .A(\fifomem_inst.waddr[1] ),
    .B(_064_));
 sg13g2_nand2_2 _253_ (.Y(_067_),
    .A(net80),
    .B(\fifomem_inst.waddr[2] ));
 sg13g2_nor2_1 _254_ (.A(_064_),
    .B(_067_),
    .Y(_068_));
 sg13g2_nor2b_1 _255_ (.A(\fifomem_inst.waddr[2] ),
    .B_N(_065_),
    .Y(_069_));
 sg13g2_nor2_1 _256_ (.A(_068_),
    .B(_069_),
    .Y(\full_inst.binnext[2] ));
 sg13g2_xnor2_1 _257_ (.Y(\full_inst.graynext[1] ),
    .A(\fifomem_inst.waddr[2] ),
    .B(_066_));
 sg13g2_xor2_1 _258_ (.B(_068_),
    .A(\full_inst.bin[3] ),
    .X(\full_inst.binnext[3] ));
 sg13g2_xnor2_1 _259_ (.Y(\full_inst.graynext[2] ),
    .A(\full_inst.bin[3] ),
    .B(_069_));
 sg13g2_xnor2_1 _260_ (.Y(_070_),
    .A(\full_inst.wsync_ptr2[2] ),
    .B(\full_inst.graynext[2] ));
 sg13g2_xor2_1 _261_ (.B(\full_inst.graynext[1] ),
    .A(\full_inst.wsync_ptr2[1] ),
    .X(_071_));
 sg13g2_nor2_1 _262_ (.A(\fifomem_inst.waddr[0] ),
    .B(_063_),
    .Y(_072_));
 sg13g2_xnor2_1 _263_ (.Y(\full_inst.graynext[0] ),
    .A(net80),
    .B(_072_));
 sg13g2_xor2_1 _264_ (.B(\full_inst.graynext[0] ),
    .A(\full_inst.wsync_ptr2[0] ),
    .X(_073_));
 sg13g2_xnor2_1 _265_ (.Y(_074_),
    .A(\full_inst.wsync_ptr2[3] ),
    .B(\full_inst.binnext[3] ));
 sg13g2_nor4_1 _266_ (.A(_070_),
    .B(_071_),
    .C(_073_),
    .D(_074_),
    .Y(\full_inst.fulln ));
 sg13g2_nand2_1 _267_ (.Y(_075_),
    .A(net65),
    .B(net73));
 sg13g2_nand2b_1 _268_ (.Y(_076_),
    .B(net65),
    .A_N(net66));
 sg13g2_o21ai_1 _269_ (.B1(_076_),
    .Y(_077_),
    .A1(net65),
    .A2(net73));
 sg13g2_nor2b_1 _270_ (.A(_077_),
    .B_N(_075_),
    .Y(_004_));
 sg13g2_xnor2_1 _271_ (.Y(_005_),
    .A(net66),
    .B(_075_));
 sg13g2_nor2b_1 _272_ (.A(net70),
    .B_N(net72),
    .Y(_078_));
 sg13g2_nor2_1 _273_ (.A(net68),
    .B(_078_),
    .Y(_000_));
 sg13g2_nand2_1 _274_ (.Y(_079_),
    .A(\clk_div_inst.rd_counter[1] ),
    .B(net68));
 sg13g2_xnor2_1 _275_ (.Y(_080_),
    .A(net72),
    .B(net68));
 sg13g2_nor2_1 _276_ (.A(_078_),
    .B(_080_),
    .Y(_001_));
 sg13g2_xnor2_1 _277_ (.Y(_002_),
    .A(net70),
    .B(_079_));
 sg13g2_xor2_1 _278_ (.B(_063_),
    .A(\fifomem_inst.waddr[0] ),
    .X(\full_inst.binnext[0] ));
 sg13g2_nand2b_2 _279_ (.Y(_081_),
    .B(_063_),
    .A_N(_006_));
 sg13g2_nor2_2 _280_ (.A(_067_),
    .B(_081_),
    .Y(_082_));
 sg13g2_mux2_1 _281_ (.A0(\fifomem_inst.fifo[7][0] ),
    .A1(net3),
    .S(_082_),
    .X(_014_));
 sg13g2_mux2_1 _282_ (.A0(\fifomem_inst.fifo[7][1] ),
    .A1(net4),
    .S(_082_),
    .X(_015_));
 sg13g2_mux2_1 _283_ (.A0(\fifomem_inst.fifo[7][2] ),
    .A1(net5),
    .S(_082_),
    .X(_016_));
 sg13g2_mux2_1 _284_ (.A0(\fifomem_inst.fifo[7][3] ),
    .A1(net6),
    .S(_082_),
    .X(_017_));
 sg13g2_nor2b_1 _285_ (.A(\clk_div_inst.rd_counter[0] ),
    .B_N(_078_),
    .Y(_083_));
 sg13g2_mux2_1 _286_ (.A0(net89),
    .A1(net63),
    .S(_083_),
    .X(_018_));
 sg13g2_nand2b_1 _287_ (.Y(_084_),
    .B(\fifomem_inst.waddr[2] ),
    .A_N(net80));
 sg13g2_nor2_2 _288_ (.A(_081_),
    .B(_084_),
    .Y(_085_));
 sg13g2_mux2_1 _289_ (.A0(\fifomem_inst.fifo[5][0] ),
    .A1(net3),
    .S(_085_),
    .X(_019_));
 sg13g2_mux2_1 _290_ (.A0(\fifomem_inst.fifo[5][1] ),
    .A1(net4),
    .S(_085_),
    .X(_020_));
 sg13g2_mux2_1 _291_ (.A0(\fifomem_inst.fifo[5][2] ),
    .A1(net5),
    .S(_085_),
    .X(_021_));
 sg13g2_mux2_1 _292_ (.A0(\fifomem_inst.fifo[5][3] ),
    .A1(net6),
    .S(_085_),
    .X(_022_));
 sg13g2_nand2b_1 _293_ (.Y(_086_),
    .B(net80),
    .A_N(\fifomem_inst.waddr[2] ));
 sg13g2_nor2_2 _294_ (.A(_081_),
    .B(_086_),
    .Y(_087_));
 sg13g2_mux2_1 _295_ (.A0(\fifomem_inst.fifo[3][0] ),
    .A1(net3),
    .S(_087_),
    .X(_023_));
 sg13g2_mux2_1 _296_ (.A0(\fifomem_inst.fifo[3][1] ),
    .A1(net4),
    .S(_087_),
    .X(_024_));
 sg13g2_mux2_1 _297_ (.A0(\fifomem_inst.fifo[3][2] ),
    .A1(net5),
    .S(_087_),
    .X(_025_));
 sg13g2_mux2_1 _298_ (.A0(\fifomem_inst.fifo[3][3] ),
    .A1(net6),
    .S(_087_),
    .X(_026_));
 sg13g2_nor2_1 _299_ (.A(\clk_div_inst.wr_counter[1] ),
    .B(_076_),
    .Y(_088_));
 sg13g2_mux2_1 _300_ (.A0(net88),
    .A1(net61),
    .S(_088_),
    .X(_027_));
 sg13g2_mux4_1 _301_ (.S0(net78),
    .A0(\fifomem_inst.fifo[0][0] ),
    .A1(\fifomem_inst.fifo[1][0] ),
    .A2(\fifomem_inst.fifo[2][0] ),
    .A3(\fifomem_inst.fifo[3][0] ),
    .S1(net77),
    .X(_089_));
 sg13g2_nor2_1 _302_ (.A(net76),
    .B(_089_),
    .Y(_090_));
 sg13g2_mux2_1 _303_ (.A0(\fifomem_inst.fifo[4][0] ),
    .A1(\fifomem_inst.fifo[5][0] ),
    .S(net78),
    .X(_091_));
 sg13g2_nor2b_1 _304_ (.A(\fifomem_inst.fifo[7][0] ),
    .B_N(net78),
    .Y(_092_));
 sg13g2_o21ai_1 _305_ (.B1(net77),
    .Y(_093_),
    .A1(\empty_inst.bin[0] ),
    .A2(\fifomem_inst.fifo[6][0] ));
 sg13g2_o21ai_1 _306_ (.B1(net76),
    .Y(_094_),
    .A1(_092_),
    .A2(_093_));
 sg13g2_a21oi_1 _307_ (.A1(_052_),
    .A2(_091_),
    .Y(_095_),
    .B1(_094_));
 sg13g2_nor3_1 _308_ (.A(_053_),
    .B(_090_),
    .C(_095_),
    .Y(_028_));
 sg13g2_mux4_1 _309_ (.S0(net79),
    .A0(\fifomem_inst.fifo[0][1] ),
    .A1(\fifomem_inst.fifo[1][1] ),
    .A2(\fifomem_inst.fifo[2][1] ),
    .A3(\fifomem_inst.fifo[3][1] ),
    .S1(net77),
    .X(_096_));
 sg13g2_nor2_1 _310_ (.A(\empty_inst.bin[2] ),
    .B(_096_),
    .Y(_097_));
 sg13g2_mux2_1 _311_ (.A0(\fifomem_inst.fifo[4][1] ),
    .A1(\fifomem_inst.fifo[5][1] ),
    .S(net79),
    .X(_098_));
 sg13g2_nor2b_1 _312_ (.A(\fifomem_inst.fifo[7][1] ),
    .B_N(\empty_inst.bin[0] ),
    .Y(_099_));
 sg13g2_o21ai_1 _313_ (.B1(net77),
    .Y(_100_),
    .A1(net79),
    .A2(\fifomem_inst.fifo[6][1] ));
 sg13g2_o21ai_1 _314_ (.B1(net76),
    .Y(_101_),
    .A1(_099_),
    .A2(_100_));
 sg13g2_a21oi_1 _315_ (.A1(_052_),
    .A2(_098_),
    .Y(_102_),
    .B1(_101_));
 sg13g2_nor3_1 _316_ (.A(_053_),
    .B(_097_),
    .C(_102_),
    .Y(_029_));
 sg13g2_mux4_1 _317_ (.S0(net78),
    .A0(\fifomem_inst.fifo[0][2] ),
    .A1(\fifomem_inst.fifo[1][2] ),
    .A2(\fifomem_inst.fifo[2][2] ),
    .A3(\fifomem_inst.fifo[3][2] ),
    .S1(net77),
    .X(_103_));
 sg13g2_nor2_1 _318_ (.A(net76),
    .B(_103_),
    .Y(_104_));
 sg13g2_mux2_1 _319_ (.A0(\fifomem_inst.fifo[4][2] ),
    .A1(\fifomem_inst.fifo[5][2] ),
    .S(net79),
    .X(_105_));
 sg13g2_nor2b_1 _320_ (.A(\fifomem_inst.fifo[7][2] ),
    .B_N(net78),
    .Y(_106_));
 sg13g2_o21ai_1 _321_ (.B1(net77),
    .Y(_107_),
    .A1(net79),
    .A2(\fifomem_inst.fifo[6][2] ));
 sg13g2_o21ai_1 _322_ (.B1(net76),
    .Y(_108_),
    .A1(_106_),
    .A2(_107_));
 sg13g2_a21oi_1 _323_ (.A1(_052_),
    .A2(_105_),
    .Y(_109_),
    .B1(_108_));
 sg13g2_nor3_1 _324_ (.A(_053_),
    .B(_104_),
    .C(_109_),
    .Y(_030_));
 sg13g2_mux4_1 _325_ (.S0(net78),
    .A0(\fifomem_inst.fifo[0][3] ),
    .A1(\fifomem_inst.fifo[1][3] ),
    .A2(\fifomem_inst.fifo[2][3] ),
    .A3(\fifomem_inst.fifo[3][3] ),
    .S1(net77),
    .X(_110_));
 sg13g2_nor2_1 _326_ (.A(net76),
    .B(_110_),
    .Y(_111_));
 sg13g2_mux2_1 _327_ (.A0(\fifomem_inst.fifo[4][3] ),
    .A1(\fifomem_inst.fifo[5][3] ),
    .S(net78),
    .X(_112_));
 sg13g2_nor2b_1 _328_ (.A(\fifomem_inst.fifo[7][3] ),
    .B_N(net78),
    .Y(_113_));
 sg13g2_o21ai_1 _329_ (.B1(\empty_inst.bin[1] ),
    .Y(_114_),
    .A1(net79),
    .A2(\fifomem_inst.fifo[6][3] ));
 sg13g2_o21ai_1 _330_ (.B1(net76),
    .Y(_115_),
    .A1(_113_),
    .A2(_114_));
 sg13g2_a21oi_1 _331_ (.A1(_052_),
    .A2(_112_),
    .Y(_116_),
    .B1(_115_));
 sg13g2_nor3_1 _332_ (.A(_053_),
    .B(_111_),
    .C(_116_),
    .Y(_031_));
 sg13g2_nand2b_2 _333_ (.Y(_117_),
    .B(_063_),
    .A_N(\fifomem_inst.waddr[0] ));
 sg13g2_nor2_2 _334_ (.A(_067_),
    .B(_117_),
    .Y(_118_));
 sg13g2_mux2_1 _335_ (.A0(\fifomem_inst.fifo[6][0] ),
    .A1(net3),
    .S(_118_),
    .X(_032_));
 sg13g2_mux2_1 _336_ (.A0(\fifomem_inst.fifo[6][1] ),
    .A1(net4),
    .S(_118_),
    .X(_033_));
 sg13g2_mux2_1 _337_ (.A0(\fifomem_inst.fifo[6][2] ),
    .A1(net5),
    .S(_118_),
    .X(_034_));
 sg13g2_mux2_1 _338_ (.A0(\fifomem_inst.fifo[6][3] ),
    .A1(net6),
    .S(_118_),
    .X(_035_));
 sg13g2_nor3_2 _339_ (.A(net80),
    .B(\fifomem_inst.waddr[2] ),
    .C(_117_),
    .Y(_119_));
 sg13g2_mux2_1 _340_ (.A0(\fifomem_inst.fifo[0][0] ),
    .A1(net3),
    .S(_119_),
    .X(_036_));
 sg13g2_mux2_1 _341_ (.A0(\fifomem_inst.fifo[0][1] ),
    .A1(net4),
    .S(_119_),
    .X(_037_));
 sg13g2_mux2_1 _342_ (.A0(\fifomem_inst.fifo[0][2] ),
    .A1(net5),
    .S(_119_),
    .X(_038_));
 sg13g2_mux2_1 _343_ (.A0(\fifomem_inst.fifo[0][3] ),
    .A1(net6),
    .S(_119_),
    .X(_039_));
 sg13g2_nor2_2 _344_ (.A(_086_),
    .B(_117_),
    .Y(_120_));
 sg13g2_mux2_1 _345_ (.A0(\fifomem_inst.fifo[2][0] ),
    .A1(net3),
    .S(_120_),
    .X(_040_));
 sg13g2_mux2_1 _346_ (.A0(\fifomem_inst.fifo[2][1] ),
    .A1(net4),
    .S(_120_),
    .X(_041_));
 sg13g2_mux2_1 _347_ (.A0(\fifomem_inst.fifo[2][2] ),
    .A1(net5),
    .S(_120_),
    .X(_042_));
 sg13g2_mux2_1 _348_ (.A0(\fifomem_inst.fifo[2][3] ),
    .A1(net6),
    .S(_120_),
    .X(_043_));
 sg13g2_nor3_2 _349_ (.A(net80),
    .B(\fifomem_inst.waddr[2] ),
    .C(_081_),
    .Y(_121_));
 sg13g2_mux2_1 _350_ (.A0(\fifomem_inst.fifo[1][0] ),
    .A1(net3),
    .S(_121_),
    .X(_044_));
 sg13g2_mux2_1 _351_ (.A0(\fifomem_inst.fifo[1][1] ),
    .A1(net4),
    .S(_121_),
    .X(_045_));
 sg13g2_mux2_1 _352_ (.A0(\fifomem_inst.fifo[1][2] ),
    .A1(net5),
    .S(_121_),
    .X(_046_));
 sg13g2_mux2_1 _353_ (.A0(\fifomem_inst.fifo[1][3] ),
    .A1(net6),
    .S(_121_),
    .X(_047_));
 sg13g2_nor2_2 _354_ (.A(_084_),
    .B(_117_),
    .Y(_122_));
 sg13g2_mux2_1 _355_ (.A0(\fifomem_inst.fifo[4][0] ),
    .A1(net3),
    .S(_122_),
    .X(_048_));
 sg13g2_mux2_1 _356_ (.A0(\fifomem_inst.fifo[4][1] ),
    .A1(net4),
    .S(_122_),
    .X(_049_));
 sg13g2_mux2_1 _357_ (.A0(\fifomem_inst.fifo[4][2] ),
    .A1(net5),
    .S(_122_),
    .X(_050_));
 sg13g2_mux2_1 _358_ (.A0(\fifomem_inst.fifo[4][3] ),
    .A1(net6),
    .S(_122_),
    .X(_051_));
 sg13g2_dfrbp_1 _359_ (.CLK(net82),
    .RESET_B(net27),
    .D(_014_),
    .Q_N(_173_),
    .Q(\fifomem_inst.fifo[7][0] ));
 sg13g2_dfrbp_1 _360_ (.CLK(net85),
    .RESET_B(net30),
    .D(_015_),
    .Q_N(_172_),
    .Q(\fifomem_inst.fifo[7][1] ));
 sg13g2_dfrbp_1 _361_ (.CLK(net82),
    .RESET_B(net29),
    .D(_016_),
    .Q_N(_171_),
    .Q(\fifomem_inst.fifo[7][2] ));
 sg13g2_dfrbp_1 _362_ (.CLK(net83),
    .RESET_B(net28),
    .D(_017_),
    .Q_N(_174_),
    .Q(\fifomem_inst.fifo[7][3] ));
 sg13g2_dfrbp_1 _363_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net97),
    .D(net69),
    .Q_N(_175_),
    .Q(\clk_div_inst.rd_counter[0] ));
 sg13g2_dfrbp_1 _364_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net96),
    .D(_001_),
    .Q_N(_176_),
    .Q(\clk_div_inst.rd_counter[1] ));
 sg13g2_dfrbp_1 _365_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net96),
    .D(net71),
    .Q_N(_170_),
    .Q(\clk_div_inst.rd_counter[2] ));
 sg13g2_dfrbp_1 _366_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net96),
    .D(net64),
    .Q_N(_011_),
    .Q(\clk_div_inst.r_clk ));
 sg13g2_dfrbp_1 _367_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net96),
    .D(_003_),
    .Q_N(_177_),
    .Q(\clk_div_inst.wr_counter[0] ));
 sg13g2_dfrbp_1 _368_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net96),
    .D(_004_),
    .Q_N(_178_),
    .Q(\clk_div_inst.wr_counter[1] ));
 sg13g2_dfrbp_1 _369_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net96),
    .D(net67),
    .Q_N(_179_),
    .Q(\clk_div_inst.wr_counter[2] ));
 sg13g2_dfrbp_1 _370_ (.CLK(net88),
    .RESET_B(net92),
    .D(\sync_r2w_inst.wsync_ptr1[0] ),
    .Q_N(_180_),
    .Q(\full_inst.wsync_ptr2[0] ));
 sg13g2_dfrbp_1 _371_ (.CLK(net86),
    .RESET_B(net95),
    .D(\sync_r2w_inst.wsync_ptr1[1] ),
    .Q_N(_181_),
    .Q(\full_inst.wsync_ptr2[1] ));
 sg13g2_dfrbp_1 _372_ (.CLK(net86),
    .RESET_B(net95),
    .D(\sync_r2w_inst.wsync_ptr1[2] ),
    .Q_N(_182_),
    .Q(\full_inst.wsync_ptr2[2] ));
 sg13g2_dfrbp_1 _373_ (.CLK(net86),
    .RESET_B(net94),
    .D(\sync_r2w_inst.wsync_ptr1[3] ),
    .Q_N(_183_),
    .Q(\full_inst.wsync_ptr2[3] ));
 sg13g2_dfrbp_1 _374_ (.CLK(net87),
    .RESET_B(net92),
    .D(\empty_inst.rptr[0] ),
    .Q_N(_184_),
    .Q(\sync_r2w_inst.wsync_ptr1[0] ));
 sg13g2_dfrbp_1 _375_ (.CLK(net86),
    .RESET_B(net95),
    .D(\empty_inst.rptr[1] ),
    .Q_N(_185_),
    .Q(\sync_r2w_inst.wsync_ptr1[1] ));
 sg13g2_dfrbp_1 _376_ (.CLK(net86),
    .RESET_B(net95),
    .D(\empty_inst.rptr[2] ),
    .Q_N(_186_),
    .Q(\sync_r2w_inst.wsync_ptr1[2] ));
 sg13g2_dfrbp_1 _377_ (.CLK(net87),
    .RESET_B(net93),
    .D(\empty_inst.bin[3] ),
    .Q_N(_187_),
    .Q(\sync_r2w_inst.wsync_ptr1[3] ));
 sg13g2_dfrbp_1 _378_ (.CLK(net89),
    .RESET_B(net92),
    .D(\sync_w2r_inst.rsync_ptr1[0] ),
    .Q_N(_188_),
    .Q(\empty_inst.rsync_ptr2[0] ));
 sg13g2_dfrbp_1 _379_ (.CLK(net90),
    .RESET_B(net94),
    .D(\sync_w2r_inst.rsync_ptr1[1] ),
    .Q_N(_189_),
    .Q(\empty_inst.rsync_ptr2[1] ));
 sg13g2_dfrbp_1 _380_ (.CLK(net90),
    .RESET_B(net94),
    .D(\sync_w2r_inst.rsync_ptr1[2] ),
    .Q_N(_190_),
    .Q(\empty_inst.rsync_ptr2[2] ));
 sg13g2_dfrbp_1 _381_ (.CLK(net89),
    .RESET_B(net93),
    .D(\sync_w2r_inst.rsync_ptr1[3] ),
    .Q_N(_191_),
    .Q(\empty_inst.rsync_ptr2[3] ));
 sg13g2_dfrbp_1 _382_ (.CLK(net89),
    .RESET_B(net92),
    .D(\full_inst.wptr[0] ),
    .Q_N(_123_),
    .Q(\sync_w2r_inst.rsync_ptr1[0] ));
 sg13g2_dfrbp_1 _383_ (.CLK(net90),
    .RESET_B(net94),
    .D(\full_inst.wptr[1] ),
    .Q_N(_124_),
    .Q(\sync_w2r_inst.rsync_ptr1[1] ));
 sg13g2_dfrbp_1 _384_ (.CLK(net90),
    .RESET_B(net95),
    .D(\full_inst.wptr[2] ),
    .Q_N(_125_),
    .Q(\sync_w2r_inst.rsync_ptr1[2] ));
 sg13g2_dfrbp_1 _385_ (.CLK(net89),
    .RESET_B(net93),
    .D(\full_inst.bin[3] ),
    .Q_N(_169_),
    .Q(\sync_w2r_inst.rsync_ptr1[3] ));
 sg13g2_dfrbp_1 _386_ (.CLK(net82),
    .RESET_B(net26),
    .D(_019_),
    .Q_N(_168_),
    .Q(\fifomem_inst.fifo[5][0] ));
 sg13g2_dfrbp_1 _387_ (.CLK(net85),
    .RESET_B(net25),
    .D(_020_),
    .Q_N(_167_),
    .Q(\fifomem_inst.fifo[5][1] ));
 sg13g2_dfrbp_1 _388_ (.CLK(net82),
    .RESET_B(net60),
    .D(_021_),
    .Q_N(_166_),
    .Q(\fifomem_inst.fifo[5][2] ));
 sg13g2_dfrbp_1 _389_ (.CLK(net82),
    .RESET_B(net59),
    .D(_022_),
    .Q_N(_165_),
    .Q(\fifomem_inst.fifo[5][3] ));
 sg13g2_dfrbp_1 _390_ (.CLK(net81),
    .RESET_B(net58),
    .D(_023_),
    .Q_N(_164_),
    .Q(\fifomem_inst.fifo[3][0] ));
 sg13g2_dfrbp_1 _391_ (.CLK(net84),
    .RESET_B(net57),
    .D(_024_),
    .Q_N(_163_),
    .Q(\fifomem_inst.fifo[3][1] ));
 sg13g2_dfrbp_1 _392_ (.CLK(net84),
    .RESET_B(net56),
    .D(_025_),
    .Q_N(_162_),
    .Q(\fifomem_inst.fifo[3][2] ));
 sg13g2_dfrbp_1 _393_ (.CLK(net81),
    .RESET_B(net54),
    .D(_026_),
    .Q_N(_161_),
    .Q(\fifomem_inst.fifo[3][3] ));
 sg13g2_dfrbp_1 _394_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net96),
    .D(net62),
    .Q_N(_010_),
    .Q(\clk_div_inst.w_clk ));
 sg13g2_dfrbp_1 _395_ (.CLK(net91),
    .RESET_B(net53),
    .D(_028_),
    .Q_N(_160_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _396_ (.CLK(net91),
    .RESET_B(net52),
    .D(_029_),
    .Q_N(_159_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _397_ (.CLK(net91),
    .RESET_B(net51),
    .D(_030_),
    .Q_N(_158_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _398_ (.CLK(net91),
    .RESET_B(net50),
    .D(_031_),
    .Q_N(_157_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _399_ (.CLK(net84),
    .RESET_B(net49),
    .D(_032_),
    .Q_N(_156_),
    .Q(\fifomem_inst.fifo[6][0] ));
 sg13g2_dfrbp_1 _400_ (.CLK(net84),
    .RESET_B(net48),
    .D(_033_),
    .Q_N(_155_),
    .Q(\fifomem_inst.fifo[6][1] ));
 sg13g2_dfrbp_1 _401_ (.CLK(net85),
    .RESET_B(net47),
    .D(_034_),
    .Q_N(_154_),
    .Q(\fifomem_inst.fifo[6][2] ));
 sg13g2_dfrbp_1 _402_ (.CLK(net84),
    .RESET_B(net44),
    .D(_035_),
    .Q_N(_126_),
    .Q(\fifomem_inst.fifo[6][3] ));
 sg13g2_dfrbp_1 _403_ (.CLK(net87),
    .RESET_B(net98),
    .D(\full_inst.graynext[0] ),
    .Q_N(_127_),
    .Q(\full_inst.wptr[0] ));
 sg13g2_dfrbp_1 _404_ (.CLK(net86),
    .RESET_B(net94),
    .D(\full_inst.graynext[1] ),
    .Q_N(_128_),
    .Q(\full_inst.wptr[1] ));
 sg13g2_dfrbp_1 _405_ (.CLK(net86),
    .RESET_B(net94),
    .D(\full_inst.graynext[2] ),
    .Q_N(_129_),
    .Q(\full_inst.wptr[2] ));
 sg13g2_dfrbp_1 _406_ (.CLK(net86),
    .RESET_B(net93),
    .D(\full_inst.binnext[3] ),
    .Q_N(_130_),
    .Q(\full_inst.bin[3] ));
 sg13g2_dfrbp_1 _407_ (.CLK(net87),
    .RESET_B(net96),
    .D(\full_inst.fulln ),
    .Q_N(_131_),
    .Q(\fifomem_inst.full ));
 sg13g2_dfrbp_1 _408_ (.CLK(net87),
    .RESET_B(net93),
    .D(\full_inst.binnext[0] ),
    .Q_N(_006_),
    .Q(\fifomem_inst.waddr[0] ));
 sg13g2_dfrbp_1 _409_ (.CLK(net87),
    .RESET_B(net93),
    .D(\full_inst.binnext[1] ),
    .Q_N(_132_),
    .Q(\fifomem_inst.waddr[1] ));
 sg13g2_dfrbp_1 _410_ (.CLK(net87),
    .RESET_B(net93),
    .D(\full_inst.binnext[2] ),
    .Q_N(_153_),
    .Q(\fifomem_inst.waddr[2] ));
 sg13g2_dfrbp_1 _411_ (.CLK(net81),
    .RESET_B(net46),
    .D(_036_),
    .Q_N(_152_),
    .Q(\fifomem_inst.fifo[0][0] ));
 sg13g2_dfrbp_1 _412_ (.CLK(net84),
    .RESET_B(net45),
    .D(_037_),
    .Q_N(_151_),
    .Q(\fifomem_inst.fifo[0][1] ));
 sg13g2_dfrbp_1 _413_ (.CLK(net83),
    .RESET_B(net43),
    .D(_038_),
    .Q_N(_150_),
    .Q(\fifomem_inst.fifo[0][2] ));
 sg13g2_dfrbp_1 _414_ (.CLK(net81),
    .RESET_B(net42),
    .D(_039_),
    .Q_N(_149_),
    .Q(\fifomem_inst.fifo[0][3] ));
 sg13g2_dfrbp_1 _415_ (.CLK(net81),
    .RESET_B(net41),
    .D(_040_),
    .Q_N(_148_),
    .Q(\fifomem_inst.fifo[2][0] ));
 sg13g2_dfrbp_1 _416_ (.CLK(net84),
    .RESET_B(net40),
    .D(_041_),
    .Q_N(_147_),
    .Q(\fifomem_inst.fifo[2][1] ));
 sg13g2_dfrbp_1 _417_ (.CLK(net83),
    .RESET_B(net39),
    .D(_042_),
    .Q_N(_146_),
    .Q(\fifomem_inst.fifo[2][2] ));
 sg13g2_dfrbp_1 _418_ (.CLK(net81),
    .RESET_B(net38),
    .D(_043_),
    .Q_N(_145_),
    .Q(\fifomem_inst.fifo[2][3] ));
 sg13g2_dfrbp_1 _419_ (.CLK(net81),
    .RESET_B(net37),
    .D(_044_),
    .Q_N(_144_),
    .Q(\fifomem_inst.fifo[1][0] ));
 sg13g2_dfrbp_1 _420_ (.CLK(net84),
    .RESET_B(net36),
    .D(_045_),
    .Q_N(_143_),
    .Q(\fifomem_inst.fifo[1][1] ));
 sg13g2_dfrbp_1 _421_ (.CLK(net83),
    .RESET_B(net35),
    .D(_046_),
    .Q_N(_142_),
    .Q(\fifomem_inst.fifo[1][2] ));
 sg13g2_dfrbp_1 _422_ (.CLK(net81),
    .RESET_B(net55),
    .D(_047_),
    .Q_N(_133_),
    .Q(\fifomem_inst.fifo[1][3] ));
 sg13g2_dfrbp_1 _423_ (.CLK(net89),
    .RESET_B(net92),
    .D(\empty_inst.graynext[0] ),
    .Q_N(_134_),
    .Q(\empty_inst.rptr[0] ));
 sg13g2_dfrbp_1 _424_ (.CLK(net90),
    .RESET_B(net94),
    .D(\empty_inst.graynext[1] ),
    .Q_N(_135_),
    .Q(\empty_inst.rptr[1] ));
 sg13g2_dfrbp_1 _425_ (.CLK(net90),
    .RESET_B(net94),
    .D(\empty_inst.graynext[2] ),
    .Q_N(_136_),
    .Q(\empty_inst.rptr[2] ));
 sg13g2_dfrbp_1 _426_ (.CLK(net89),
    .RESET_B(net93),
    .D(\empty_inst.binnext[3] ),
    .Q_N(_141_),
    .Q(\empty_inst.bin[3] ));
 sg13g2_dfrbp_1 _427_ (.CLK(net89),
    .RESET_B(net98),
    .D(_013_),
    .Q_N(empty),
    .Q(_012_));
 sg13g2_dfrbp_1 _428_ (.CLK(net91),
    .RESET_B(net92),
    .D(\empty_inst.binnext[0] ),
    .Q_N(_007_),
    .Q(\empty_inst.bin[0] ));
 sg13g2_dfrbp_1 _429_ (.CLK(net91),
    .RESET_B(net92),
    .D(\empty_inst.binnext[1] ),
    .Q_N(_008_),
    .Q(\empty_inst.bin[1] ));
 sg13g2_dfrbp_1 _430_ (.CLK(net91),
    .RESET_B(net92),
    .D(\empty_inst.binnext[2] ),
    .Q_N(_009_),
    .Q(\empty_inst.bin[2] ));
 sg13g2_dfrbp_1 _431_ (.CLK(net82),
    .RESET_B(net34),
    .D(_048_),
    .Q_N(_140_),
    .Q(\fifomem_inst.fifo[4][0] ));
 sg13g2_dfrbp_1 _432_ (.CLK(net85),
    .RESET_B(net33),
    .D(_049_),
    .Q_N(_139_),
    .Q(\fifomem_inst.fifo[4][1] ));
 sg13g2_dfrbp_1 _433_ (.CLK(net82),
    .RESET_B(net32),
    .D(_050_),
    .Q_N(_138_),
    .Q(\fifomem_inst.fifo[4][2] ));
 sg13g2_dfrbp_1 _434_ (.CLK(net82),
    .RESET_B(net31),
    .D(_051_),
    .Q_N(_137_),
    .Q(\fifomem_inst.fifo[4][3] ));
 sg13g2_tiehi _386__26 (.L_HI(net26));
 sg13g2_tiehi _359__27 (.L_HI(net27));
 sg13g2_tiehi _362__28 (.L_HI(net28));
 sg13g2_tiehi _361__29 (.L_HI(net29));
 sg13g2_tiehi _360__30 (.L_HI(net30));
 sg13g2_tiehi _434__31 (.L_HI(net31));
 sg13g2_tiehi _433__32 (.L_HI(net32));
 sg13g2_tiehi _432__33 (.L_HI(net33));
 sg13g2_tiehi _431__34 (.L_HI(net34));
 sg13g2_tiehi _421__35 (.L_HI(net35));
 sg13g2_tiehi _420__36 (.L_HI(net36));
 sg13g2_tiehi _419__37 (.L_HI(net37));
 sg13g2_tiehi _418__38 (.L_HI(net38));
 sg13g2_tiehi _417__39 (.L_HI(net39));
 sg13g2_tiehi _416__40 (.L_HI(net40));
 sg13g2_tiehi _415__41 (.L_HI(net41));
 sg13g2_tiehi _414__42 (.L_HI(net42));
 sg13g2_tiehi _413__43 (.L_HI(net43));
 sg13g2_tiehi _402__44 (.L_HI(net44));
 sg13g2_tiehi _412__45 (.L_HI(net45));
 sg13g2_tiehi _411__46 (.L_HI(net46));
 sg13g2_tiehi _401__47 (.L_HI(net47));
 sg13g2_tiehi _400__48 (.L_HI(net48));
 sg13g2_tiehi _399__49 (.L_HI(net49));
 sg13g2_tiehi _398__50 (.L_HI(net50));
 sg13g2_tiehi _397__51 (.L_HI(net51));
 sg13g2_tiehi _396__52 (.L_HI(net52));
 sg13g2_tiehi _395__53 (.L_HI(net53));
 sg13g2_tiehi _393__54 (.L_HI(net54));
 sg13g2_tiehi _422__55 (.L_HI(net55));
 sg13g2_tiehi _392__56 (.L_HI(net56));
 sg13g2_tiehi _391__57 (.L_HI(net57));
 sg13g2_tiehi _390__58 (.L_HI(net58));
 sg13g2_tiehi _389__59 (.L_HI(net59));
 sg13g2_tiehi _388__60 (.L_HI(net60));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_reemashivva_fifo_8 (.L_LO(net8));
 sg13g2_tielo tt_um_reemashivva_fifo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_reemashivva_fifo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_reemashivva_fifo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_reemashivva_fifo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_reemashivva_fifo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_reemashivva_fifo_14 (.L_LO(net14));
 sg13g2_tielo tt_um_reemashivva_fifo_15 (.L_LO(net15));
 sg13g2_tielo tt_um_reemashivva_fifo_16 (.L_LO(net16));
 sg13g2_tielo tt_um_reemashivva_fifo_17 (.L_LO(net17));
 sg13g2_tielo tt_um_reemashivva_fifo_18 (.L_LO(net18));
 sg13g2_tielo tt_um_reemashivva_fifo_19 (.L_LO(net19));
 sg13g2_tielo tt_um_reemashivva_fifo_20 (.L_LO(net20));
 sg13g2_tielo tt_um_reemashivva_fifo_21 (.L_LO(net21));
 sg13g2_tielo tt_um_reemashivva_fifo_22 (.L_LO(net22));
 sg13g2_tielo tt_um_reemashivva_fifo_23 (.L_LO(net23));
 sg13g2_tielo tt_um_reemashivva_fifo_24 (.L_LO(net24));
 sg13g2_tiehi _387__25 (.L_HI(net25));
 sg13g2_buf_1 _489_ (.A(\fifomem_inst.full ),
    .X(uo_out[0]));
 sg13g2_buf_1 _490_ (.A(empty),
    .X(uo_out[1]));
 sg13g2_buf_2 fanout76 (.A(\empty_inst.bin[2] ),
    .X(net76));
 sg13g2_buf_4 fanout77 (.X(net77),
    .A(\empty_inst.bin[1] ));
 sg13g2_buf_4 fanout78 (.X(net78),
    .A(net79));
 sg13g2_buf_4 fanout79 (.X(net79),
    .A(\empty_inst.bin[0] ));
 sg13g2_buf_2 fanout80 (.A(\fifomem_inst.waddr[1] ),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(net83),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(net83),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(net88),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(net88),
    .X(net84));
 sg13g2_buf_1 fanout85 (.A(net88),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(net87),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(net88),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(\clk_div_inst.w_clk ),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(\clk_div_inst.r_clk ),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(net91),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(\clk_div_inst.r_clk ),
    .X(net91));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(net98));
 sg13g2_buf_4 fanout93 (.X(net93),
    .A(net98));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(net97));
 sg13g2_buf_2 fanout95 (.A(net97),
    .X(net95));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(net97));
 sg13g2_buf_2 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(rst_n),
    .X(net98));
 sg13g2_buf_1 input1 (.A(ui_in[2]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[4]));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[5]));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[6]));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[7]));
 sg13g2_tielo tt_um_reemashivva_fifo_7 (.L_LO(net7));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_010_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold2 (.A(_027_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold3 (.A(_011_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold4 (.A(_018_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold5 (.A(\clk_div_inst.wr_counter[0] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold6 (.A(\clk_div_inst.wr_counter[2] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold7 (.A(_005_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold8 (.A(\clk_div_inst.rd_counter[0] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold9 (.A(_000_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold10 (.A(\clk_div_inst.rd_counter[2] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold11 (.A(_002_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold12 (.A(\clk_div_inst.rd_counter[1] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold13 (.A(\clk_div_inst.wr_counter[1] ),
    .X(net73));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_4 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_174 ();
 sg13g2_decap_8 FILLER_24_181 ();
 sg13g2_decap_8 FILLER_24_188 ();
 sg13g2_fill_2 FILLER_24_195 ();
 sg13g2_decap_8 FILLER_24_223 ();
 sg13g2_decap_8 FILLER_24_230 ();
 sg13g2_decap_8 FILLER_24_237 ();
 sg13g2_decap_8 FILLER_24_244 ();
 sg13g2_decap_8 FILLER_24_251 ();
 sg13g2_decap_8 FILLER_24_258 ();
 sg13g2_decap_8 FILLER_24_265 ();
 sg13g2_decap_8 FILLER_24_272 ();
 sg13g2_decap_8 FILLER_24_279 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_293 ();
 sg13g2_decap_8 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_307 ();
 sg13g2_decap_8 FILLER_24_314 ();
 sg13g2_decap_8 FILLER_24_321 ();
 sg13g2_decap_8 FILLER_24_328 ();
 sg13g2_decap_8 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_349 ();
 sg13g2_decap_8 FILLER_24_356 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_4 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_137 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_decap_8 FILLER_25_177 ();
 sg13g2_decap_8 FILLER_25_184 ();
 sg13g2_decap_8 FILLER_25_191 ();
 sg13g2_fill_1 FILLER_25_198 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_decap_8 FILLER_25_232 ();
 sg13g2_decap_8 FILLER_25_239 ();
 sg13g2_decap_8 FILLER_25_246 ();
 sg13g2_decap_8 FILLER_25_253 ();
 sg13g2_decap_8 FILLER_25_260 ();
 sg13g2_decap_8 FILLER_25_267 ();
 sg13g2_decap_8 FILLER_25_274 ();
 sg13g2_decap_8 FILLER_25_281 ();
 sg13g2_decap_8 FILLER_25_288 ();
 sg13g2_decap_8 FILLER_25_295 ();
 sg13g2_decap_8 FILLER_25_302 ();
 sg13g2_decap_8 FILLER_25_309 ();
 sg13g2_decap_8 FILLER_25_316 ();
 sg13g2_decap_8 FILLER_25_323 ();
 sg13g2_decap_8 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_25_337 ();
 sg13g2_decap_8 FILLER_25_344 ();
 sg13g2_decap_8 FILLER_25_351 ();
 sg13g2_decap_8 FILLER_25_358 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_4 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_decap_4 FILLER_26_145 ();
 sg13g2_fill_1 FILLER_26_149 ();
 sg13g2_decap_8 FILLER_26_180 ();
 sg13g2_decap_4 FILLER_26_187 ();
 sg13g2_fill_1 FILLER_26_191 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_fill_2 FILLER_26_256 ();
 sg13g2_decap_8 FILLER_26_267 ();
 sg13g2_decap_8 FILLER_26_274 ();
 sg13g2_decap_4 FILLER_26_281 ();
 sg13g2_fill_2 FILLER_26_293 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_decap_8 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_84 ();
 sg13g2_fill_1 FILLER_27_86 ();
 sg13g2_fill_1 FILLER_27_107 ();
 sg13g2_fill_2 FILLER_27_128 ();
 sg13g2_decap_4 FILLER_27_184 ();
 sg13g2_fill_2 FILLER_27_188 ();
 sg13g2_decap_8 FILLER_27_234 ();
 sg13g2_decap_4 FILLER_27_241 ();
 sg13g2_fill_2 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_fill_1 FILLER_27_280 ();
 sg13g2_decap_4 FILLER_27_333 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_decap_4 FILLER_27_370 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_131 ();
 sg13g2_decap_8 FILLER_28_138 ();
 sg13g2_decap_4 FILLER_28_145 ();
 sg13g2_decap_8 FILLER_28_180 ();
 sg13g2_decap_8 FILLER_28_187 ();
 sg13g2_decap_4 FILLER_28_194 ();
 sg13g2_decap_8 FILLER_28_229 ();
 sg13g2_fill_1 FILLER_28_236 ();
 sg13g2_fill_1 FILLER_28_280 ();
 sg13g2_decap_4 FILLER_28_320 ();
 sg13g2_fill_1 FILLER_28_324 ();
 sg13g2_decap_8 FILLER_28_341 ();
 sg13g2_decap_8 FILLER_28_348 ();
 sg13g2_decap_4 FILLER_28_355 ();
 sg13g2_fill_1 FILLER_28_359 ();
 sg13g2_decap_8 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_131 ();
 sg13g2_decap_8 FILLER_29_138 ();
 sg13g2_decap_8 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_decap_8 FILLER_29_167 ();
 sg13g2_decap_8 FILLER_29_174 ();
 sg13g2_decap_8 FILLER_29_181 ();
 sg13g2_decap_8 FILLER_29_188 ();
 sg13g2_fill_2 FILLER_29_195 ();
 sg13g2_fill_1 FILLER_29_197 ();
 sg13g2_decap_8 FILLER_29_221 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_fill_2 FILLER_29_235 ();
 sg13g2_fill_1 FILLER_29_237 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_fill_2 FILLER_29_287 ();
 sg13g2_fill_1 FILLER_29_292 ();
 sg13g2_fill_2 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_4 FILLER_30_70 ();
 sg13g2_fill_1 FILLER_30_108 ();
 sg13g2_fill_2 FILLER_30_130 ();
 sg13g2_fill_1 FILLER_30_132 ();
 sg13g2_fill_2 FILLER_30_143 ();
 sg13g2_fill_1 FILLER_30_145 ();
 sg13g2_decap_8 FILLER_30_172 ();
 sg13g2_decap_8 FILLER_30_179 ();
 sg13g2_fill_2 FILLER_30_186 ();
 sg13g2_fill_1 FILLER_30_188 ();
 sg13g2_decap_8 FILLER_30_219 ();
 sg13g2_decap_8 FILLER_30_226 ();
 sg13g2_fill_2 FILLER_30_233 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_285 ();
 sg13g2_fill_1 FILLER_30_287 ();
 sg13g2_decap_4 FILLER_30_296 ();
 sg13g2_decap_4 FILLER_30_316 ();
 sg13g2_fill_1 FILLER_30_320 ();
 sg13g2_decap_8 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_84 ();
 sg13g2_decap_4 FILLER_31_89 ();
 sg13g2_fill_2 FILLER_31_113 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_4 FILLER_31_178 ();
 sg13g2_fill_1 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_226 ();
 sg13g2_fill_2 FILLER_31_243 ();
 sg13g2_fill_1 FILLER_31_248 ();
 sg13g2_decap_8 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_31_296 ();
 sg13g2_fill_1 FILLER_31_318 ();
 sg13g2_fill_2 FILLER_31_371 ();
 sg13g2_fill_1 FILLER_31_373 ();
 sg13g2_fill_1 FILLER_31_404 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_4 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_114 ();
 sg13g2_decap_8 FILLER_32_121 ();
 sg13g2_decap_8 FILLER_32_128 ();
 sg13g2_fill_2 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_226 ();
 sg13g2_decap_8 FILLER_32_281 ();
 sg13g2_decap_4 FILLER_32_288 ();
 sg13g2_fill_2 FILLER_32_300 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_fill_2 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_353 ();
 sg13g2_fill_2 FILLER_32_392 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_4 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_124 ();
 sg13g2_decap_8 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_138 ();
 sg13g2_decap_8 FILLER_33_143 ();
 sg13g2_fill_2 FILLER_33_150 ();
 sg13g2_fill_2 FILLER_33_157 ();
 sg13g2_decap_8 FILLER_33_179 ();
 sg13g2_decap_8 FILLER_33_186 ();
 sg13g2_fill_1 FILLER_33_193 ();
 sg13g2_fill_2 FILLER_33_199 ();
 sg13g2_fill_1 FILLER_33_207 ();
 sg13g2_fill_1 FILLER_33_212 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_decap_4 FILLER_33_277 ();
 sg13g2_fill_1 FILLER_33_323 ();
 sg13g2_fill_2 FILLER_33_343 ();
 sg13g2_fill_1 FILLER_33_375 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_fill_2 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_110 ();
 sg13g2_decap_4 FILLER_34_122 ();
 sg13g2_fill_2 FILLER_34_136 ();
 sg13g2_fill_1 FILLER_34_172 ();
 sg13g2_fill_2 FILLER_34_178 ();
 sg13g2_decap_8 FILLER_34_185 ();
 sg13g2_decap_4 FILLER_34_192 ();
 sg13g2_fill_2 FILLER_34_196 ();
 sg13g2_fill_1 FILLER_34_241 ();
 sg13g2_decap_8 FILLER_34_276 ();
 sg13g2_decap_8 FILLER_34_283 ();
 sg13g2_fill_2 FILLER_34_290 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_fill_1 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_93 ();
 sg13g2_fill_2 FILLER_35_160 ();
 sg13g2_fill_2 FILLER_35_167 ();
 sg13g2_decap_8 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_191 ();
 sg13g2_fill_1 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_223 ();
 sg13g2_decap_8 FILLER_35_230 ();
 sg13g2_fill_2 FILLER_35_237 ();
 sg13g2_decap_8 FILLER_35_265 ();
 sg13g2_decap_8 FILLER_35_272 ();
 sg13g2_fill_2 FILLER_35_279 ();
 sg13g2_fill_1 FILLER_35_281 ();
 sg13g2_fill_2 FILLER_35_316 ();
 sg13g2_fill_1 FILLER_35_358 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_127 ();
 sg13g2_fill_1 FILLER_36_129 ();
 sg13g2_decap_4 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_237 ();
 sg13g2_decap_4 FILLER_36_268 ();
 sg13g2_fill_1 FILLER_36_272 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_4 FILLER_37_117 ();
 sg13g2_fill_1 FILLER_37_121 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_fill_2 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_135 ();
 sg13g2_decap_8 FILLER_37_176 ();
 sg13g2_decap_8 FILLER_37_183 ();
 sg13g2_fill_1 FILLER_37_194 ();
 sg13g2_decap_8 FILLER_37_225 ();
 sg13g2_decap_8 FILLER_37_232 ();
 sg13g2_fill_2 FILLER_37_239 ();
 sg13g2_decap_8 FILLER_37_267 ();
 sg13g2_decap_8 FILLER_37_274 ();
 sg13g2_decap_4 FILLER_37_281 ();
 sg13g2_fill_1 FILLER_37_311 ();
 sg13g2_fill_2 FILLER_37_360 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_92 ();
 sg13g2_fill_2 FILLER_38_110 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_fill_2 FILLER_38_158 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_fill_2 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_223 ();
 sg13g2_decap_8 FILLER_38_230 ();
 sg13g2_decap_8 FILLER_38_237 ();
 sg13g2_decap_4 FILLER_38_244 ();
 sg13g2_fill_2 FILLER_38_248 ();
 sg13g2_decap_8 FILLER_38_262 ();
 sg13g2_decap_8 FILLER_38_269 ();
 sg13g2_decap_8 FILLER_38_276 ();
 sg13g2_decap_8 FILLER_38_283 ();
 sg13g2_decap_8 FILLER_38_290 ();
 sg13g2_fill_2 FILLER_38_297 ();
 sg13g2_fill_1 FILLER_38_299 ();
 sg13g2_fill_2 FILLER_38_328 ();
 sg13g2_fill_1 FILLER_38_339 ();
 sg13g2_fill_2 FILLER_38_372 ();
 assign uio_oe[0] = net7;
 assign uio_oe[1] = net8;
 assign uio_oe[2] = net9;
 assign uio_oe[3] = net10;
 assign uio_oe[4] = net11;
 assign uio_oe[5] = net12;
 assign uio_oe[6] = net13;
 assign uio_oe[7] = net14;
 assign uio_out[0] = net15;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
 assign uio_out[3] = net18;
 assign uio_out[4] = net19;
 assign uio_out[5] = net20;
 assign uio_out[6] = net21;
 assign uio_out[7] = net22;
 assign uo_out[6] = net23;
 assign uo_out[7] = net24;
endmodule

module tt_um_MichaelBell_canon (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire \crotchet[0] ;
 wire \crotchet[1] ;
 wire \crotchet[2] ;
 wire \crotchet[3] ;
 wire \crotchet[4] ;
 wire \crotchet[5] ;
 wire \crotchet[6] ;
 wire \i_display.colour[0] ;
 wire \i_display.colour[1] ;
 wire \i_display.colour[2] ;
 wire \i_display.colour[3] ;
 wire \i_display.colour[4] ;
 wire \i_display.colour[5] ;
 wire \i_display.frame[0] ;
 wire \i_display.frame[1] ;
 wire \i_display.frame[2] ;
 wire \i_display.frame[3] ;
 wire \i_display.frame[4] ;
 wire \i_display.frame[5] ;
 wire \i_display.frame[6] ;
 wire \i_display.frame[7] ;
 wire \i_display.frame[8] ;
 wire \i_display.frame[9] ;
 wire \i_display.frame_crotchet[0] ;
 wire \i_display.frame_crotchet[1] ;
 wire \i_display.frame_crotchet[2] ;
 wire \i_display.frame_crotchet[3] ;
 wire \i_display.frame_crotchet[4] ;
 wire \i_display.frame_crotchet[5] ;
 wire \i_display.frame_crotchet[6] ;
 wire \i_display.hsync ;
 wire \i_display.i_vga.hblank ;
 wire \i_display.i_vga.hblank_tmp ;
 wire \i_display.i_vga.hsync_tmp ;
 wire \i_display.i_vga.low_count[0] ;
 wire \i_display.i_vga.low_count[1] ;
 wire \i_display.i_vga.low_count[2] ;
 wire \i_display.i_vga.low_count[3] ;
 wire \i_display.i_vga.low_count[4] ;
 wire \i_display.i_vga.low_count[5] ;
 wire \i_display.i_vga.low_count[6] ;
 wire \i_display.i_vga.low_count[7] ;
 wire \i_display.i_vga.low_count[8] ;
 wire \i_display.i_vga.low_count[9] ;
 wire \i_display.i_vga.timing_ver.blank ;
 wire \i_display.i_vga.timing_ver.counter[0] ;
 wire \i_display.i_vga.timing_ver.counter[10] ;
 wire \i_display.i_vga.timing_ver.counter[1] ;
 wire \i_display.i_vga.timing_ver.counter[2] ;
 wire \i_display.i_vga.timing_ver.counter[3] ;
 wire \i_display.i_vga.timing_ver.counter[4] ;
 wire \i_display.i_vga.timing_ver.counter[5] ;
 wire \i_display.i_vga.timing_ver.counter[6] ;
 wire \i_display.i_vga.timing_ver.counter[7] ;
 wire \i_display.i_vga.timing_ver.counter[8] ;
 wire \i_display.i_vga.timing_ver.counter[9] ;
 wire \i_display.i_vga.timing_ver.sync ;
 wire \i_display.i_vga.timing_ver.sync_tmp ;
 wire \i_display.i_vga.vblank ;
 wire \i_display.in_line ;
 wire \i_display.x_idx[0] ;
 wire \i_display.x_idx[1] ;
 wire \i_display.x_idx[2] ;
 wire \i_display.x_idx[3] ;
 wire \i_display.x_idx[4] ;
 wire \i_display.x_idx[5] ;
 wire \i_display.x_idx[6] ;
 wire \i_display.x_idx[7] ;
 wire \i_display.x_idx[8] ;
 wire \i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[-1] ;
 wire \i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[-2] ;
 wire \i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[-3] ;
 wire \i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[-4] ;
 wire \i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[-5] ;
 wire \i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[0] ;
 wire \i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[1] ;
 wire \i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[2] ;
 wire \i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[0] ;
 wire \i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[1] ;
 wire \i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[2] ;
 wire \i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[3] ;
 wire \i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[4] ;
 wire \i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[5] ;
 wire \i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[6] ;
 wire \i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[7] ;
 wire \i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[8] ;
 wire \i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[9] ;
 wire \i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[0] ;
 wire \i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[10] ;
 wire \i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[1] ;
 wire \i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[2] ;
 wire \i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[3] ;
 wire \i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[4] ;
 wire \i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[5] ;
 wire \i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[6] ;
 wire \i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[7] ;
 wire \i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[8] ;
 wire \i_music.count[10] ;
 wire \i_music.count[11] ;
 wire \i_music.count[12] ;
 wire \i_music.count[13] ;
 wire \i_music.count[14] ;
 wire \i_music.count[15] ;
 wire \i_music.count[16] ;
 wire \i_music.count[17] ;
 wire \i_music.count[18] ;
 wire \i_music.count[19] ;
 wire \i_music.count[20] ;
 wire \i_music.count[21] ;
 wire \i_music.count[22] ;
 wire \i_music.count[23] ;
 wire \i_music.count[24] ;
 wire \i_music.i_pwm.count[0] ;
 wire \i_music.i_pwm.count[1] ;
 wire \i_music.i_pwm.count[2] ;
 wire \i_music.i_pwm.count[3] ;
 wire \i_music.i_pwm.count[4] ;
 wire \i_music.i_pwm.count[5] ;
 wire \i_music.i_pwm.count[6] ;
 wire \i_music.i_pwm.count[7] ;
 wire \i_music.i_pwm.pwm ;
 wire \i_music.i_pwm.sample[0] ;
 wire \i_music.i_pwm.sample[1] ;
 wire \i_music.i_pwm.sample[2] ;
 wire \i_music.i_pwm.sample[3] ;
 wire \i_music.i_pwm.sample[4] ;
 wire \i_music.i_pwm.sample[5] ;
 wire \i_music.i_pwm.sample[6] ;
 wire \i_music.i_pwm.sample[7] ;
 wire \i_music.i_sample.sample_acc[0] ;
 wire \i_music.i_sample.sample_acc[1] ;
 wire \i_music.i_sample.sample_acc[2] ;
 wire \i_music.i_sample.sample_acc[3] ;
 wire \i_music.i_sample.sample_acc[4] ;
 wire \i_music.i_sample.sample_acc[5] ;
 wire \i_music.i_sample.sample_acc[6] ;
 wire \i_music.i_sample.sample_acc[7] ;
 wire \i_music.i_sample.sample_acc[8] ;
 wire \i_music.i_sample.sample_idx[0] ;
 wire \i_music.i_sample.sample_idx[1] ;
 wire \i_music.i_sample.sample_idx[2] ;
 wire \i_music.i_sample.sample_idx[3] ;
 wire \i_music.i_sample.sample_idx[4] ;
 wire \i_music.i_sample.sample_idx[5] ;
 wire \i_music.i_sample.sample_idx[6] ;
 wire \i_music.i_sample.sample_idx[7] ;
 wire \i_music.i_sample.t1.CG.GCLK ;
 wire \i_music.i_sample.t1.genblk1[0].state.D ;
 wire \i_music.i_sample.t1.genblk1[0].state.Q ;
 wire \i_music.i_sample.t1.genblk1[10].state.D ;
 wire \i_music.i_sample.t1.genblk1[10].state.Q ;
 wire \i_music.i_sample.t1.genblk1[11].state.D ;
 wire \i_music.i_sample.t1.genblk1[11].state.Q ;
 wire \i_music.i_sample.t1.genblk1[12].state.D ;
 wire \i_music.i_sample.t1.genblk1[12].state.Q ;
 wire \i_music.i_sample.t1.genblk1[13].state.D ;
 wire \i_music.i_sample.t1.genblk1[13].state.Q ;
 wire \i_music.i_sample.t1.genblk1[14].state.D ;
 wire \i_music.i_sample.t1.genblk1[14].state.Q ;
 wire \i_music.i_sample.t1.genblk1[15].state.D ;
 wire \i_music.i_sample.t1.genblk1[15].state.Q ;
 wire \i_music.i_sample.t1.genblk1[16].state.D ;
 wire \i_music.i_sample.t1.genblk1[16].state.Q ;
 wire \i_music.i_sample.t1.genblk1[17].state.D ;
 wire \i_music.i_sample.t1.genblk1[17].state.Q ;
 wire \i_music.i_sample.t1.genblk1[18].state.D ;
 wire \i_music.i_sample.t1.genblk1[18].state.Q ;
 wire \i_music.i_sample.t1.genblk1[1].state.D ;
 wire \i_music.i_sample.t1.genblk1[1].state.Q ;
 wire \i_music.i_sample.t1.genblk1[2].state.D ;
 wire \i_music.i_sample.t1.genblk1[2].state.Q ;
 wire \i_music.i_sample.t1.genblk1[3].state.D ;
 wire \i_music.i_sample.t1.genblk1[3].state.Q ;
 wire \i_music.i_sample.t1.genblk1[4].state.D ;
 wire \i_music.i_sample.t1.genblk1[4].state.Q ;
 wire \i_music.i_sample.t1.genblk1[5].state.D ;
 wire \i_music.i_sample.t1.genblk1[5].state.Q ;
 wire \i_music.i_sample.t1.genblk1[6].state.D ;
 wire \i_music.i_sample.t1.genblk1[6].state.Q ;
 wire \i_music.i_sample.t1.genblk1[7].state.D ;
 wire \i_music.i_sample.t1.genblk1[7].state.Q ;
 wire \i_music.i_sample.t1.genblk1[8].state.D ;
 wire \i_music.i_sample.t1.genblk1[8].state.Q ;
 wire \i_music.i_sample.t1.genblk1[9].state.D ;
 wire \i_music.i_sample.t1.genblk1[9].state.Q ;
 wire \i_music.i_sample.t2.CG.GCLK ;
 wire \i_music.i_sample.t2.genblk1[0].state.Q ;
 wire \i_music.i_sample.t2.genblk1[10].state.Q ;
 wire \i_music.i_sample.t2.genblk1[11].state.Q ;
 wire \i_music.i_sample.t2.genblk1[12].state.Q ;
 wire \i_music.i_sample.t2.genblk1[13].state.Q ;
 wire \i_music.i_sample.t2.genblk1[14].state.Q ;
 wire \i_music.i_sample.t2.genblk1[15].state.Q ;
 wire \i_music.i_sample.t2.genblk1[16].state.Q ;
 wire \i_music.i_sample.t2.genblk1[17].state.Q ;
 wire \i_music.i_sample.t2.genblk1[1].state.Q ;
 wire \i_music.i_sample.t2.genblk1[2].state.Q ;
 wire \i_music.i_sample.t2.genblk1[3].state.Q ;
 wire \i_music.i_sample.t2.genblk1[4].state.Q ;
 wire \i_music.i_sample.t2.genblk1[5].state.Q ;
 wire \i_music.i_sample.t2.genblk1[6].state.Q ;
 wire \i_music.i_sample.t2.genblk1[7].state.Q ;
 wire \i_music.i_sample.t2.genblk1[8].state.Q ;
 wire \i_music.i_sample.t2.genblk1[9].state.Q ;
 wire \i_music.i_sample.t3.CG.GCLK ;
 wire \i_music.i_sample.t3.genblk1[0].state.Q ;
 wire \i_music.i_sample.t3.genblk1[10].state.Q ;
 wire \i_music.i_sample.t3.genblk1[11].state.Q ;
 wire \i_music.i_sample.t3.genblk1[12].state.Q ;
 wire \i_music.i_sample.t3.genblk1[13].state.Q ;
 wire \i_music.i_sample.t3.genblk1[14].state.Q ;
 wire \i_music.i_sample.t3.genblk1[15].state.Q ;
 wire \i_music.i_sample.t3.genblk1[16].state.Q ;
 wire \i_music.i_sample.t3.genblk1[17].state.Q ;
 wire \i_music.i_sample.t3.genblk1[1].state.Q ;
 wire \i_music.i_sample.t3.genblk1[2].state.Q ;
 wire \i_music.i_sample.t3.genblk1[3].state.Q ;
 wire \i_music.i_sample.t3.genblk1[4].state.Q ;
 wire \i_music.i_sample.t3.genblk1[5].state.Q ;
 wire \i_music.i_sample.t3.genblk1[6].state.Q ;
 wire \i_music.i_sample.t3.genblk1[7].state.Q ;
 wire \i_music.i_sample.t3.genblk1[8].state.Q ;
 wire \i_music.i_sample.t3.genblk1[9].state.Q ;
 wire \i_music.i_sample.t4.CG.GCLK ;
 wire \i_music.i_sample.t4.genblk1[0].state.Q ;
 wire \i_music.i_sample.t4.genblk1[10].state.Q ;
 wire \i_music.i_sample.t4.genblk1[11].state.Q ;
 wire \i_music.i_sample.t4.genblk1[12].state.Q ;
 wire \i_music.i_sample.t4.genblk1[13].state.Q ;
 wire \i_music.i_sample.t4.genblk1[14].state.Q ;
 wire \i_music.i_sample.t4.genblk1[15].state.Q ;
 wire \i_music.i_sample.t4.genblk1[16].state.Q ;
 wire \i_music.i_sample.t4.genblk1[17].state.Q ;
 wire \i_music.i_sample.t4.genblk1[1].state.Q ;
 wire \i_music.i_sample.t4.genblk1[2].state.Q ;
 wire \i_music.i_sample.t4.genblk1[3].state.Q ;
 wire \i_music.i_sample.t4.genblk1[4].state.Q ;
 wire \i_music.i_sample.t4.genblk1[5].state.Q ;
 wire \i_music.i_sample.t4.genblk1[6].state.Q ;
 wire \i_music.i_sample.t4.genblk1[7].state.Q ;
 wire \i_music.i_sample.t4.genblk1[8].state.Q ;
 wire \i_music.i_sample.t4.genblk1[9].state.Q ;
 wire \i_music.i_sample.thresh[0] ;
 wire \i_music.i_sample.thresh[10] ;
 wire \i_music.i_sample.thresh[1] ;
 wire \i_music.i_sample.thresh[2] ;
 wire \i_music.i_sample.thresh[3] ;
 wire \i_music.i_sample.thresh[4] ;
 wire \i_music.i_sample.thresh[5] ;
 wire \i_music.i_sample.thresh[6] ;
 wire \i_music.i_sample.thresh[7] ;
 wire \i_music.i_sample.thresh[8] ;
 wire \i_music.i_sample.thresh[9] ;
 wire \i_music.violin_note_idx[1][0] ;
 wire \i_music.violin_note_idx[1][1] ;
 wire \i_music.violin_note_idx[1][2] ;
 wire \i_music.violin_note_idx[1][3] ;
 wire \i_music.violin_note_idx[1][4] ;
 wire \i_music.violin_note_idx[1][5] ;
 wire \i_music.violin_note_idx[1][6] ;
 wire \i_music.violin_note_idx[1][7] ;
 wire \i_music.violin_note_idx[1][8] ;
 wire \i_music.violin_note_idx[2][0] ;
 wire \i_music.violin_note_idx[2][1] ;
 wire \i_music.violin_note_idx[2][2] ;
 wire \i_music.violin_note_idx[2][3] ;
 wire \i_music.violin_note_idx[2][4] ;
 wire \i_music.violin_note_idx[2][5] ;
 wire \i_music.violin_note_idx[2][6] ;
 wire \i_music.violin_note_idx[2][7] ;
 wire \i_music.violin_note_idx[2][8] ;
 wire \i_music.violin_note_idx[3][0] ;
 wire \i_music.violin_note_idx[3][1] ;
 wire \i_music.violin_note_idx[3][2] ;
 wire \i_music.violin_note_idx[3][3] ;
 wire \i_music.violin_note_idx[3][4] ;
 wire \i_music.violin_note_idx[3][5] ;
 wire \i_music.violin_note_idx[3][6] ;
 wire \i_music.violin_note_idx[3][7] ;
 wire \i_music.violin_note_idx[3][8] ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clk_regs;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire clknet_0__1501_;
 wire clknet_1_0__leaf__1501_;
 wire clknet_1_1__leaf__1501_;
 wire \clknet_0_i_music.i_sample.t4.CG.GCLK ;
 wire \clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ;
 wire \clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ;
 wire \clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ;
 wire \clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ;
 wire \clknet_0_i_music.i_sample.t3.CG.GCLK ;
 wire \clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ;
 wire \clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ;
 wire \clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ;
 wire \clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ;
 wire \clknet_0_i_music.i_sample.t2.CG.GCLK ;
 wire \clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ;
 wire \clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ;
 wire \clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ;
 wire \clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ;
 wire \clknet_0_i_music.i_sample.t1.CG.GCLK ;
 wire \clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ;
 wire \clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ;
 wire \clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ;
 wire \clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ;
 wire delaynet_0_clk;
 wire delaynet_1_clk;
 wire delaynet_2_clk;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;

 sg13g2_inv_1 _3606_ (.Y(_2908_),
    .A(net326));
 sg13g2_inv_1 _3607_ (.Y(_2909_),
    .A(\i_display.in_line ));
 sg13g2_inv_1 _3608_ (.Y(_2910_),
    .A(_0096_));
 sg13g2_inv_2 _3609_ (.Y(_2911_),
    .A(net1104));
 sg13g2_inv_1 _3610_ (.Y(_2912_),
    .A(net1111));
 sg13g2_inv_2 _3611_ (.Y(_2913_),
    .A(net1113));
 sg13g2_inv_2 _3612_ (.Y(_2914_),
    .A(net1114));
 sg13g2_inv_1 _3613_ (.Y(_2915_),
    .A(net1119));
 sg13g2_inv_2 _3614_ (.Y(_2916_),
    .A(net1122));
 sg13g2_inv_2 _3615_ (.Y(_2917_),
    .A(net1123));
 sg13g2_inv_1 _3616_ (.Y(_2918_),
    .A(net1126));
 sg13g2_inv_1 _3617_ (.Y(_2919_),
    .A(net1127));
 sg13g2_inv_1 _3618_ (.Y(_2920_),
    .A(net368));
 sg13g2_inv_1 _3619_ (.Y(_2921_),
    .A(net375));
 sg13g2_inv_1 _3620_ (.Y(_2922_),
    .A(net1130));
 sg13g2_inv_1 _3621_ (.Y(_2923_),
    .A(net1167));
 sg13g2_inv_1 _3622_ (.Y(_2924_),
    .A(\crotchet[2] ));
 sg13g2_inv_1 _3623_ (.Y(_2925_),
    .A(\i_music.violin_note_idx[2][0] ));
 sg13g2_inv_1 _3624_ (.Y(_2926_),
    .A(net301));
 sg13g2_inv_1 _3625_ (.Y(_2927_),
    .A(\i_display.i_vga.low_count[6] ));
 sg13g2_inv_1 _3626_ (.Y(_2928_),
    .A(\i_display.i_vga.low_count[8] ));
 sg13g2_inv_2 _3627_ (.Y(_2929_),
    .A(net330));
 sg13g2_inv_1 _3628_ (.Y(_2930_),
    .A(net1149));
 sg13g2_inv_1 _3629_ (.Y(_2931_),
    .A(\i_display.i_vga.low_count[4] ));
 sg13g2_inv_2 _3630_ (.Y(_2932_),
    .A(_0069_));
 sg13g2_inv_2 _3631_ (.Y(_2933_),
    .A(_0075_));
 sg13g2_inv_2 _3632_ (.Y(_2934_),
    .A(_0077_));
 sg13g2_inv_2 _3633_ (.Y(_2935_),
    .A(_0081_));
 sg13g2_inv_1 _3634_ (.Y(_2936_),
    .A(_0085_));
 sg13g2_inv_1 _3635_ (.Y(_2937_),
    .A(_0087_));
 sg13g2_inv_2 _3636_ (.Y(_2938_),
    .A(_0089_));
 sg13g2_inv_1 _3637_ (.Y(_2939_),
    .A(_0092_));
 sg13g2_inv_1 _3638_ (.Y(_2940_),
    .A(_0094_));
 sg13g2_inv_1 _3639_ (.Y(_2941_),
    .A(_0095_));
 sg13g2_inv_1 _3640_ (.Y(_2942_),
    .A(_0028_));
 sg13g2_inv_1 _3641_ (.Y(_2943_),
    .A(_0083_));
 sg13g2_inv_1 _3642_ (.Y(_2944_),
    .A(net262));
 sg13g2_inv_1 _3643_ (.Y(_2945_),
    .A(net344));
 sg13g2_inv_1 _3644_ (.Y(_2946_),
    .A(\i_music.count[22] ));
 sg13g2_inv_1 _3645_ (.Y(_2947_),
    .A(\i_music.violin_note_idx[3][5] ));
 sg13g2_inv_1 _3646_ (.Y(_2948_),
    .A(\i_music.violin_note_idx[2][5] ));
 sg13g2_inv_2 _3647_ (.Y(_2949_),
    .A(net333));
 sg13g2_inv_1 _3648_ (.Y(_2950_),
    .A(net222));
 sg13g2_inv_1 _3649_ (.Y(_2951_),
    .A(\i_music.violin_note_idx[3][4] ));
 sg13g2_inv_1 _3650_ (.Y(_2952_),
    .A(net311));
 sg13g2_inv_1 _3651_ (.Y(_2953_),
    .A(\i_music.violin_note_idx[2][6] ));
 sg13g2_inv_1 _3652_ (.Y(_2954_),
    .A(\i_music.violin_note_idx[3][1] ));
 sg13g2_inv_1 _3653_ (.Y(_2955_),
    .A(net250));
 sg13g2_inv_1 _3654_ (.Y(_2956_),
    .A(\i_music.violin_note_idx[3][0] ));
 sg13g2_inv_1 _3655_ (.Y(_2957_),
    .A(net306));
 sg13g2_inv_1 _3656_ (.Y(_2958_),
    .A(\i_music.violin_note_idx[2][2] ));
 sg13g2_inv_1 _3657_ (.Y(_2959_),
    .A(\i_music.violin_note_idx[2][8] ));
 sg13g2_inv_1 _3658_ (.Y(_2960_),
    .A(\i_music.i_pwm.count[1] ));
 sg13g2_inv_1 _3659_ (.Y(_2961_),
    .A(\i_music.i_pwm.count[4] ));
 sg13g2_inv_1 _3660_ (.Y(_2962_),
    .A(\i_music.i_pwm.count[7] ));
 sg13g2_inv_1 _3661_ (.Y(_2963_),
    .A(_0047_));
 sg13g2_inv_2 _3662_ (.Y(_2964_),
    .A(net351));
 sg13g2_inv_1 _3663_ (.Y(_2965_),
    .A(net280));
 sg13g2_inv_1 _3664_ (.Y(_2966_),
    .A(net968));
 sg13g2_inv_1 _3665_ (.Y(_2967_),
    .A(net959));
 sg13g2_inv_1 _3666_ (.Y(_2968_),
    .A(net953));
 sg13g2_inv_2 _3667_ (.Y(_2969_),
    .A(net975));
 sg13g2_inv_1 _3668_ (.Y(_2970_),
    .A(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[4] ));
 sg13g2_inv_1 _3669_ (.Y(_2971_),
    .A(\i_music.i_sample.t1.genblk1[8].state.Q ));
 sg13g2_inv_1 _3670_ (.Y(_2972_),
    .A(\i_music.i_sample.t1.genblk1[9].state.Q ));
 sg13g2_inv_1 _3671_ (.Y(_2973_),
    .A(\i_music.i_sample.t1.genblk1[10].state.Q ));
 sg13g2_inv_1 _3672_ (.Y(_2974_),
    .A(\i_music.i_sample.t1.genblk1[11].state.Q ));
 sg13g2_inv_1 _3673_ (.Y(_2975_),
    .A(\i_music.i_sample.t1.genblk1[12].state.Q ));
 sg13g2_inv_1 _3674_ (.Y(_2976_),
    .A(\i_music.i_sample.t1.genblk1[13].state.Q ));
 sg13g2_inv_1 _3675_ (.Y(_2977_),
    .A(\i_music.i_sample.t1.genblk1[14].state.Q ));
 sg13g2_inv_1 _3676_ (.Y(_2978_),
    .A(\i_music.i_sample.t1.genblk1[15].state.Q ));
 sg13g2_inv_1 _3677_ (.Y(_2979_),
    .A(\i_music.i_sample.t1.genblk1[16].state.Q ));
 sg13g2_inv_1 _3678_ (.Y(_2980_),
    .A(\i_music.i_sample.t1.genblk1[17].state.Q ));
 sg13g2_inv_1 _3679_ (.Y(_2981_),
    .A(\i_music.i_sample.thresh[8] ));
 sg13g2_inv_1 _3680_ (.Y(_2982_),
    .A(net376));
 sg13g2_inv_1 _3681_ (.Y(_2983_),
    .A(\i_music.i_sample.sample_idx[4] ));
 sg13g2_inv_1 _3682_ (.Y(_2984_),
    .A(net372));
 sg13g2_inv_1 _3683_ (.Y(_2985_),
    .A(net1));
 sg13g2_inv_1 _3684_ (.Y(_2986_),
    .A(net271));
 sg13g2_inv_2 _3685_ (.Y(_2987_),
    .A(net240));
 sg13g2_inv_1 _3686_ (.Y(_2988_),
    .A(\i_music.i_pwm.sample[4] ));
 sg13g2_inv_1 _3687_ (.Y(_2989_),
    .A(net254));
 sg13g2_inv_1 _3688_ (.Y(_2990_),
    .A(\i_music.i_pwm.sample[1] ));
 sg13g2_inv_1 _3689_ (.Y(_2991_),
    .A(net206));
 sg13g2_or2_1 _3690_ (.X(_2992_),
    .B(\i_display.i_vga.low_count[5] ),
    .A(\i_display.i_vga.low_count[6] ));
 sg13g2_nor3_2 _3691_ (.A(_2928_),
    .B(net1142),
    .C(_2992_),
    .Y(_2993_));
 sg13g2_nor3_1 _3692_ (.A(_2929_),
    .B(net210),
    .C(_2993_),
    .Y(_2994_));
 sg13g2_and2_1 _3693_ (.A(net1154),
    .B(net1148),
    .X(_2995_));
 sg13g2_nand2_2 _3694_ (.Y(_2996_),
    .A(net1153),
    .B(net1147));
 sg13g2_and3_1 _3695_ (.X(_2997_),
    .A(\i_display.i_vga.low_count[2] ),
    .B(\i_display.i_vga.low_count[3] ),
    .C(net1088));
 sg13g2_nand4_1 _3696_ (.B(\i_display.i_vga.low_count[2] ),
    .C(net1148),
    .A(net1153),
    .Y(_2998_),
    .D(\i_display.i_vga.low_count[3] ));
 sg13g2_nand3b_1 _3697_ (.B(\i_display.i_vga.low_count[9] ),
    .C(\i_display.i_vga.low_count[8] ),
    .Y(_2999_),
    .A_N(net1141));
 sg13g2_nor4_2 _3698_ (.A(_2931_),
    .B(_2992_),
    .C(_2998_),
    .Y(_3000_),
    .D(_2999_));
 sg13g2_nor3_2 _3699_ (.A(_2929_),
    .B(_2931_),
    .C(_2998_),
    .Y(_3001_));
 sg13g2_or2_1 _3700_ (.X(\i_display.i_vga.hblank_tmp ),
    .B(_3000_),
    .A(_2994_));
 sg13g2_nand4_1 _3701_ (.B(\i_display.i_vga.low_count[5] ),
    .C(\i_display.i_vga.low_count[4] ),
    .A(_2927_),
    .Y(_3002_),
    .D(\i_display.i_vga.low_count[3] ));
 sg13g2_a21oi_1 _3702_ (.A1(net245),
    .A2(_3002_),
    .Y(\i_display.i_vga.hsync_tmp ),
    .B1(_2999_));
 sg13g2_nand3b_1 _3703_ (.B(net212),
    .C(\i_display.i_vga.timing_ver.counter[7] ),
    .Y(_3003_),
    .A_N(\i_display.i_vga.timing_ver.counter[4] ));
 sg13g2_nand4_1 _3704_ (.B(\i_display.i_vga.timing_ver.counter[8] ),
    .C(\i_display.i_vga.timing_ver.counter[6] ),
    .A(\i_display.i_vga.timing_ver.counter[9] ),
    .Y(_3004_),
    .D(\i_display.i_vga.timing_ver.counter[5] ));
 sg13g2_or3_1 _3705_ (.A(\i_display.i_vga.timing_ver.counter[2] ),
    .B(net1130),
    .C(_3004_),
    .X(_3005_));
 sg13g2_nor3_2 _3706_ (.A(net207),
    .B(net213),
    .C(_3005_),
    .Y(\i_display.i_vga.timing_ver.sync_tmp ));
 sg13g2_mux2_1 _3707_ (.A0(\i_music.i_sample.t2.genblk1[0].state.Q ),
    .A1(\i_music.i_sample.t4.genblk1[0].state.Q ),
    .S(net1143),
    .X(_3006_));
 sg13g2_inv_1 _3708_ (.Y(_3007_),
    .A(_3006_));
 sg13g2_nor2b_2 _3709_ (.A(net1144),
    .B_N(net1150),
    .Y(_3008_));
 sg13g2_inv_1 _3710_ (.Y(_3009_),
    .A(_3008_));
 sg13g2_a22oi_1 _3711_ (.Y(_3010_),
    .B1(net1082),
    .B2(\i_music.i_sample.t3.genblk1[0].state.Q ),
    .A2(net1084),
    .A1(net943));
 sg13g2_o21ai_1 _3712_ (.B1(_3010_),
    .Y(_0237_),
    .A1(net1150),
    .A2(_3007_));
 sg13g2_mux2_1 _3713_ (.A0(\i_music.i_sample.t2.genblk1[1].state.Q ),
    .A1(\i_music.i_sample.t4.genblk1[1].state.Q ),
    .S(net1143),
    .X(_3011_));
 sg13g2_inv_1 _3714_ (.Y(_3012_),
    .A(_3011_));
 sg13g2_a22oi_1 _3715_ (.Y(_3013_),
    .B1(net1082),
    .B2(\i_music.i_sample.t3.genblk1[1].state.Q ),
    .A2(net1084),
    .A1(net948));
 sg13g2_o21ai_1 _3716_ (.B1(_3013_),
    .Y(_0238_),
    .A1(net1150),
    .A2(_3012_));
 sg13g2_mux2_1 _3717_ (.A0(\i_music.i_sample.t2.genblk1[2].state.Q ),
    .A1(\i_music.i_sample.t4.genblk1[2].state.Q ),
    .S(net1143),
    .X(_3014_));
 sg13g2_inv_1 _3718_ (.Y(_3015_),
    .A(_3014_));
 sg13g2_a22oi_1 _3719_ (.Y(_3016_),
    .B1(net1082),
    .B2(\i_music.i_sample.t3.genblk1[2].state.Q ),
    .A2(net1084),
    .A1(net952));
 sg13g2_o21ai_1 _3720_ (.B1(_3016_),
    .Y(_0239_),
    .A1(net1150),
    .A2(_3015_));
 sg13g2_mux2_1 _3721_ (.A0(\i_music.i_sample.t2.genblk1[3].state.Q ),
    .A1(\i_music.i_sample.t4.genblk1[3].state.Q ),
    .S(net1143),
    .X(_3017_));
 sg13g2_inv_1 _3722_ (.Y(_3018_),
    .A(_3017_));
 sg13g2_a22oi_1 _3723_ (.Y(_3019_),
    .B1(net1082),
    .B2(\i_music.i_sample.t3.genblk1[3].state.Q ),
    .A2(net1084),
    .A1(net958));
 sg13g2_o21ai_1 _3724_ (.B1(_3019_),
    .Y(_0240_),
    .A1(net1150),
    .A2(_3018_));
 sg13g2_mux2_1 _3725_ (.A0(\i_music.i_sample.t2.genblk1[4].state.Q ),
    .A1(\i_music.i_sample.t4.genblk1[4].state.Q ),
    .S(net1144),
    .X(_3020_));
 sg13g2_inv_1 _3726_ (.Y(_3021_),
    .A(_3020_));
 sg13g2_a22oi_1 _3727_ (.Y(_3022_),
    .B1(net1082),
    .B2(\i_music.i_sample.t3.genblk1[4].state.Q ),
    .A2(net1085),
    .A1(net965));
 sg13g2_o21ai_1 _3728_ (.B1(_3022_),
    .Y(_0241_),
    .A1(net1152),
    .A2(_3021_));
 sg13g2_mux2_1 _3729_ (.A0(\i_music.i_sample.t2.genblk1[5].state.Q ),
    .A1(\i_music.i_sample.t4.genblk1[5].state.Q ),
    .S(net1145),
    .X(_3023_));
 sg13g2_inv_1 _3730_ (.Y(_3024_),
    .A(_3023_));
 sg13g2_a22oi_1 _3731_ (.Y(_3025_),
    .B1(_3008_),
    .B2(\i_music.i_sample.t3.genblk1[5].state.Q ),
    .A2(net1085),
    .A1(\i_music.i_sample.t1.genblk1[5].state.Q ));
 sg13g2_o21ai_1 _3732_ (.B1(_3025_),
    .Y(_0242_),
    .A1(net1152),
    .A2(_3024_));
 sg13g2_mux2_1 _3733_ (.A0(\i_music.i_sample.t2.genblk1[6].state.Q ),
    .A1(\i_music.i_sample.t4.genblk1[6].state.Q ),
    .S(net1145),
    .X(_3026_));
 sg13g2_inv_1 _3734_ (.Y(_3027_),
    .A(_3026_));
 sg13g2_a22oi_1 _3735_ (.Y(_3028_),
    .B1(net1083),
    .B2(\i_music.i_sample.t3.genblk1[6].state.Q ),
    .A2(net1088),
    .A1(net974));
 sg13g2_o21ai_1 _3736_ (.B1(_3028_),
    .Y(_0243_),
    .A1(net1153),
    .A2(_3027_));
 sg13g2_mux2_1 _3737_ (.A0(\i_music.i_sample.t2.genblk1[7].state.Q ),
    .A1(\i_music.i_sample.t4.genblk1[7].state.Q ),
    .S(net1145),
    .X(_3029_));
 sg13g2_inv_1 _3738_ (.Y(_3030_),
    .A(_3029_));
 sg13g2_a22oi_1 _3739_ (.Y(_3031_),
    .B1(net1083),
    .B2(\i_music.i_sample.t3.genblk1[7].state.Q ),
    .A2(net1088),
    .A1(net976));
 sg13g2_o21ai_1 _3740_ (.B1(_3031_),
    .Y(_0244_),
    .A1(net1153),
    .A2(_3030_));
 sg13g2_nor2b_1 _3741_ (.A(net1154),
    .B_N(net1148),
    .Y(_3032_));
 sg13g2_nand2b_1 _3742_ (.Y(_3033_),
    .B(net1143),
    .A_N(net1152));
 sg13g2_o21ai_1 _3743_ (.B1(net1146),
    .Y(_3034_),
    .A1(net1151),
    .A2(\i_music.i_sample.t4.genblk1[8].state.Q ));
 sg13g2_nor2_1 _3744_ (.A(net1153),
    .B(net1145),
    .Y(_3035_));
 sg13g2_or2_1 _3745_ (.X(_3036_),
    .B(net1148),
    .A(net1153));
 sg13g2_a22oi_1 _3746_ (.Y(_3037_),
    .B1(net1070),
    .B2(\i_music.i_sample.t2.genblk1[8].state.Q ),
    .A2(net1083),
    .A1(\i_music.i_sample.t3.genblk1[8].state.Q ));
 sg13g2_a22oi_1 _3747_ (.Y(_0245_),
    .B1(_3034_),
    .B2(_3037_),
    .A2(net1086),
    .A1(_2971_));
 sg13g2_nand2_1 _3748_ (.Y(_3038_),
    .A(\i_music.i_sample.t2.genblk1[9].state.Q ),
    .B(net1070));
 sg13g2_a221oi_1 _3749_ (.B2(net1083),
    .C1(net1086),
    .B1(\i_music.i_sample.t3.genblk1[9].state.Q ),
    .A1(net1146),
    .Y(_3039_),
    .A2(\i_music.i_sample.t4.genblk1[9].state.Q ));
 sg13g2_a22oi_1 _3750_ (.Y(_0246_),
    .B1(_3038_),
    .B2(_3039_),
    .A2(net1086),
    .A1(_2972_));
 sg13g2_nand2_1 _3751_ (.Y(_3040_),
    .A(\i_music.i_sample.t2.genblk1[10].state.Q ),
    .B(net1070));
 sg13g2_a221oi_1 _3752_ (.B2(net1083),
    .C1(net1086),
    .B1(\i_music.i_sample.t3.genblk1[10].state.Q ),
    .A1(net1146),
    .Y(_3041_),
    .A2(\i_music.i_sample.t4.genblk1[10].state.Q ));
 sg13g2_a22oi_1 _3753_ (.Y(_0247_),
    .B1(_3040_),
    .B2(_3041_),
    .A2(net1086),
    .A1(_2973_));
 sg13g2_o21ai_1 _3754_ (.B1(net1146),
    .Y(_3042_),
    .A1(net1150),
    .A2(\i_music.i_sample.t4.genblk1[11].state.Q ));
 sg13g2_a22oi_1 _3755_ (.Y(_3043_),
    .B1(\i_music.i_sample.t2.genblk1[11].state.Q ),
    .B2(net1070),
    .A2(\i_music.i_sample.t3.genblk1[11].state.Q ),
    .A1(net1150));
 sg13g2_a22oi_1 _3756_ (.Y(_0248_),
    .B1(_3042_),
    .B2(_3043_),
    .A2(net1085),
    .A1(_2974_));
 sg13g2_o21ai_1 _3757_ (.B1(net1144),
    .Y(_3044_),
    .A1(net1151),
    .A2(\i_music.i_sample.t4.genblk1[12].state.Q ));
 sg13g2_a22oi_1 _3758_ (.Y(_3045_),
    .B1(\i_music.i_sample.t2.genblk1[12].state.Q ),
    .B2(net1070),
    .A2(\i_music.i_sample.t3.genblk1[12].state.Q ),
    .A1(net1151));
 sg13g2_a22oi_1 _3759_ (.Y(_0249_),
    .B1(_3044_),
    .B2(_3045_),
    .A2(net1085),
    .A1(_2975_));
 sg13g2_o21ai_1 _3760_ (.B1(net1144),
    .Y(_3046_),
    .A1(net1151),
    .A2(\i_music.i_sample.t4.genblk1[13].state.Q ));
 sg13g2_a22oi_1 _3761_ (.Y(_3047_),
    .B1(net1070),
    .B2(\i_music.i_sample.t2.genblk1[13].state.Q ),
    .A2(net1082),
    .A1(\i_music.i_sample.t3.genblk1[13].state.Q ));
 sg13g2_a22oi_1 _3762_ (.Y(_0250_),
    .B1(_3046_),
    .B2(_3047_),
    .A2(net1084),
    .A1(_2976_));
 sg13g2_nand2_1 _3763_ (.Y(_3048_),
    .A(\i_music.i_sample.t2.genblk1[14].state.Q ),
    .B(net1070));
 sg13g2_a221oi_1 _3764_ (.B2(net1082),
    .C1(net1084),
    .B1(\i_music.i_sample.t3.genblk1[14].state.Q ),
    .A1(net1143),
    .Y(_3049_),
    .A2(\i_music.i_sample.t4.genblk1[14].state.Q ));
 sg13g2_a22oi_1 _3765_ (.Y(_0251_),
    .B1(_3048_),
    .B2(_3049_),
    .A2(net1084),
    .A1(_2977_));
 sg13g2_o21ai_1 _3766_ (.B1(net1143),
    .Y(_3050_),
    .A1(net1150),
    .A2(\i_music.i_sample.t4.genblk1[15].state.Q ));
 sg13g2_a22oi_1 _3767_ (.Y(_3051_),
    .B1(\i_music.i_sample.t2.genblk1[15].state.Q ),
    .B2(net1070),
    .A2(\i_music.i_sample.t3.genblk1[15].state.Q ),
    .A1(net1151));
 sg13g2_a22oi_1 _3768_ (.Y(_0252_),
    .B1(_3050_),
    .B2(_3051_),
    .A2(net1084),
    .A1(_2978_));
 sg13g2_o21ai_1 _3769_ (.B1(net1143),
    .Y(_3052_),
    .A1(net1152),
    .A2(\i_music.i_sample.t4.genblk1[16].state.Q ));
 sg13g2_a22oi_1 _3770_ (.Y(_3053_),
    .B1(net1072),
    .B2(\i_music.i_sample.t2.genblk1[16].state.Q ),
    .A2(net1082),
    .A1(\i_music.i_sample.t3.genblk1[16].state.Q ));
 sg13g2_a22oi_1 _3771_ (.Y(_0253_),
    .B1(_3052_),
    .B2(_3053_),
    .A2(net1085),
    .A1(_2979_));
 sg13g2_nand2_1 _3772_ (.Y(_3054_),
    .A(\i_music.i_sample.t2.genblk1[17].state.Q ),
    .B(net1074));
 sg13g2_a221oi_1 _3773_ (.B2(net1083),
    .C1(net1088),
    .B1(\i_music.i_sample.t3.genblk1[17].state.Q ),
    .A1(net1145),
    .Y(_3055_),
    .A2(\i_music.i_sample.t4.genblk1[17].state.Q ));
 sg13g2_a22oi_1 _3774_ (.Y(_0254_),
    .B1(_3054_),
    .B2(_3055_),
    .A2(net1088),
    .A1(_2980_));
 sg13g2_nor2_1 _3775_ (.A(net1132),
    .B(\i_display.i_vga.hblank ),
    .Y(_3056_));
 sg13g2_and2_1 _3776_ (.A(\i_display.colour[5] ),
    .B(net1066),
    .X(uo_out[0]));
 sg13g2_and2_2 _3777_ (.A(\i_display.colour[3] ),
    .B(net1066),
    .X(uo_out[1]));
 sg13g2_and2_1 _3778_ (.A(\i_display.colour[1] ),
    .B(net1066),
    .X(uo_out[2]));
 sg13g2_and2_1 _3779_ (.A(\i_display.colour[4] ),
    .B(net1066),
    .X(uo_out[4]));
 sg13g2_and2_1 _3780_ (.A(\i_display.colour[2] ),
    .B(net1066),
    .X(uo_out[5]));
 sg13g2_and2_1 _3781_ (.A(\i_display.colour[0] ),
    .B(net1066),
    .X(uo_out[6]));
 sg13g2_and3_1 _3782_ (.X(_3057_),
    .A(\i_display.i_vga.low_count[5] ),
    .B(\i_display.i_vga.low_count[4] ),
    .C(_2997_));
 sg13g2_nand3_1 _3783_ (.B(net1141),
    .C(_3057_),
    .A(\i_display.i_vga.low_count[6] ),
    .Y(_3058_));
 sg13g2_or3_1 _3784_ (.A(_2928_),
    .B(_2929_),
    .C(_3058_),
    .X(_3059_));
 sg13g2_nor2_1 _3785_ (.A(_2945_),
    .B(_3059_),
    .Y(_3060_));
 sg13g2_and2_1 _3786_ (.A(net287),
    .B(_3060_),
    .X(_3061_));
 sg13g2_and2_1 _3787_ (.A(net260),
    .B(_3061_),
    .X(_3062_));
 sg13g2_and2_1 _3788_ (.A(net273),
    .B(_3062_),
    .X(_3063_));
 sg13g2_and2_1 _3789_ (.A(net293),
    .B(_3063_),
    .X(_3064_));
 sg13g2_and2_1 _3790_ (.A(net296),
    .B(_3064_),
    .X(_3065_));
 sg13g2_and2_1 _3791_ (.A(net288),
    .B(_3065_),
    .X(_3066_));
 sg13g2_and2_1 _3792_ (.A(net300),
    .B(_3066_),
    .X(_3067_));
 sg13g2_and2_1 _3793_ (.A(net274),
    .B(_3067_),
    .X(_3068_));
 sg13g2_and2_1 _3794_ (.A(net353),
    .B(_3068_),
    .X(_3069_));
 sg13g2_and2_1 _3795_ (.A(net360),
    .B(_3069_),
    .X(_3070_));
 sg13g2_and2_1 _3796_ (.A(\i_music.count[21] ),
    .B(_3070_),
    .X(_3071_));
 sg13g2_and2_1 _3797_ (.A(net347),
    .B(_3071_),
    .X(_3072_));
 sg13g2_and3_1 _3798_ (.X(_3073_),
    .A(net382),
    .B(net225),
    .C(_3072_));
 sg13g2_nand3_1 _3799_ (.B(\crotchet[0] ),
    .C(_3073_),
    .A(\crotchet[1] ),
    .Y(_3074_));
 sg13g2_nand2_1 _3800_ (.Y(_3075_),
    .A(_2924_),
    .B(_3074_));
 sg13g2_nor2_2 _3801_ (.A(_2924_),
    .B(_3074_),
    .Y(_3076_));
 sg13g2_nand3b_1 _3802_ (.B(net1168),
    .C(_3075_),
    .Y(_3077_),
    .A_N(_3076_));
 sg13g2_inv_1 _3803_ (.Y(_0162_),
    .A(_3077_));
 sg13g2_a21oi_1 _3804_ (.A1(_2963_),
    .A2(_3073_),
    .Y(_3078_),
    .B1(net1157));
 sg13g2_o21ai_1 _3805_ (.B1(_3078_),
    .Y(_3079_),
    .A1(_2963_),
    .A2(_3073_));
 sg13g2_inv_1 _3806_ (.Y(_0160_),
    .A(_3079_));
 sg13g2_a21o_1 _3807_ (.A2(_3073_),
    .A1(\crotchet[0] ),
    .B1(\crotchet[1] ),
    .X(_3080_));
 sg13g2_and2_1 _3808_ (.A(_3074_),
    .B(_3080_),
    .X(_3081_));
 sg13g2_nand2_1 _3809_ (.Y(_3082_),
    .A(net1168),
    .B(_3081_));
 sg13g2_inv_1 _3810_ (.Y(_0161_),
    .A(_3082_));
 sg13g2_o21ai_1 _3811_ (.B1(_3077_),
    .Y(_3083_),
    .A1(_0160_),
    .A2(_0161_));
 sg13g2_o21ai_1 _3812_ (.B1(_0162_),
    .Y(_3084_),
    .A1(_3079_),
    .A2(_3081_));
 sg13g2_nand2_1 _3813_ (.Y(_3085_),
    .A(_3083_),
    .B(_3084_));
 sg13g2_inv_1 _3814_ (.Y(_0019_),
    .A(_3085_));
 sg13g2_nand2_1 _3815_ (.Y(_3086_),
    .A(_3077_),
    .B(_3082_));
 sg13g2_nand2_1 _3816_ (.Y(_3087_),
    .A(_0160_),
    .B(_3081_));
 sg13g2_o21ai_1 _3817_ (.B1(_3086_),
    .Y(_0020_),
    .A1(_3077_),
    .A2(_3087_));
 sg13g2_nand2_1 _3818_ (.Y(_0185_),
    .A(_2924_),
    .B(_0161_));
 sg13g2_inv_1 _3819_ (.Y(_0184_),
    .A(_0185_));
 sg13g2_nand2_1 _3820_ (.Y(_0021_),
    .A(_3079_),
    .B(_0185_));
 sg13g2_nand2_1 _3821_ (.Y(_0181_),
    .A(_0162_),
    .B(_3079_));
 sg13g2_nand3_1 _3822_ (.B(_3087_),
    .C(_0181_),
    .A(_3086_),
    .Y(_0022_));
 sg13g2_mux2_1 _3823_ (.A0(_3077_),
    .A1(_3083_),
    .S(_3087_),
    .X(_0023_));
 sg13g2_and2_2 _3824_ (.A(\i_display.i_vga.timing_ver.counter[0] ),
    .B(_3000_),
    .X(_3088_));
 sg13g2_and2_2 _3825_ (.A(\i_display.i_vga.timing_ver.sync_tmp ),
    .B(_3088_),
    .X(_3089_));
 sg13g2_nand2_2 _3826_ (.Y(_3090_),
    .A(\i_display.i_vga.timing_ver.sync_tmp ),
    .B(_3088_));
 sg13g2_nand2_2 _3827_ (.Y(_3091_),
    .A(net1174),
    .B(net1005));
 sg13g2_and3_2 _3828_ (.X(_3092_),
    .A(\i_display.i_vga.timing_ver.counter[0] ),
    .B(_2993_),
    .C(_3001_));
 sg13g2_and2_2 _3829_ (.A(\i_display.i_vga.timing_ver.sync_tmp ),
    .B(_3092_),
    .X(_3093_));
 sg13g2_inv_1 _3830_ (.Y(_3094_),
    .A(_3093_));
 sg13g2_nand2b_1 _3831_ (.Y(_3095_),
    .B(net1001),
    .A_N(net341));
 sg13g2_xnor2_1 _3832_ (.Y(_3096_),
    .A(net6),
    .B(\crotchet[4] ));
 sg13g2_xor2_1 _3833_ (.B(\crotchet[4] ),
    .A(net6),
    .X(_3097_));
 sg13g2_o21ai_1 _3834_ (.B1(_3095_),
    .Y(_0018_),
    .A1(net1001),
    .A2(_3096_));
 sg13g2_inv_1 _3835_ (.Y(_0017_),
    .A(_0018_));
 sg13g2_nor2_1 _3836_ (.A(\i_display.hsync ),
    .B(_3000_),
    .Y(_3098_));
 sg13g2_or2_1 _3837_ (.X(_3099_),
    .B(_3000_),
    .A(\i_display.hsync ));
 sg13g2_nand2b_2 _3838_ (.Y(_3100_),
    .B(net1099),
    .A_N(net1097));
 sg13g2_nor2_2 _3839_ (.A(net1093),
    .B(\i_display.x_idx[0] ),
    .Y(_3101_));
 sg13g2_or2_2 _3840_ (.X(_3102_),
    .B(net1096),
    .A(net1092));
 sg13g2_nor2_2 _3841_ (.A(_0088_),
    .B(_3102_),
    .Y(_3103_));
 sg13g2_nand2b_2 _3842_ (.Y(_3104_),
    .B(_3101_),
    .A_N(_0088_));
 sg13g2_a21oi_1 _3843_ (.A1(_2937_),
    .A2(_3103_),
    .Y(_3105_),
    .B1(net1090));
 sg13g2_nor2_1 _3844_ (.A(net1113),
    .B(_3104_),
    .Y(_3106_));
 sg13g2_nor2_2 _3845_ (.A(net1109),
    .B(_3106_),
    .Y(_3107_));
 sg13g2_o21ai_1 _3846_ (.B1(net1090),
    .Y(_3108_),
    .A1(net1112),
    .A2(_3104_));
 sg13g2_nand2b_2 _3847_ (.Y(_3109_),
    .B(net1096),
    .A_N(net1093));
 sg13g2_nor2_1 _3848_ (.A(_0088_),
    .B(_3109_),
    .Y(_3110_));
 sg13g2_nand2_1 _3849_ (.Y(_3111_),
    .A(net1113),
    .B(_3110_));
 sg13g2_nand2b_1 _3850_ (.Y(_3112_),
    .B(_3111_),
    .A_N(_3106_));
 sg13g2_a21oi_1 _3851_ (.A1(_3107_),
    .A2(_3111_),
    .Y(_3113_),
    .B1(_3105_));
 sg13g2_nor2_1 _3852_ (.A(net1105),
    .B(net1090),
    .Y(_3114_));
 sg13g2_nor2_1 _3853_ (.A(net1093),
    .B(_2913_),
    .Y(_3115_));
 sg13g2_nor2_2 _3854_ (.A(_3101_),
    .B(_3115_),
    .Y(_3116_));
 sg13g2_nor2_2 _3855_ (.A(_2913_),
    .B(_2914_),
    .Y(_3117_));
 sg13g2_nand2_2 _3856_ (.Y(_3118_),
    .A(net1113),
    .B(net1115));
 sg13g2_nor2_2 _3857_ (.A(net1094),
    .B(_2914_),
    .Y(_3119_));
 sg13g2_nor2_2 _3858_ (.A(net1113),
    .B(net1114),
    .Y(_3120_));
 sg13g2_or2_2 _3859_ (.X(_3121_),
    .B(net1115),
    .A(net1113));
 sg13g2_nor3_1 _3860_ (.A(net1094),
    .B(_3117_),
    .C(_3120_),
    .Y(_3122_));
 sg13g2_nor2_1 _3861_ (.A(net1104),
    .B(net1109),
    .Y(_3123_));
 sg13g2_nor4_1 _3862_ (.A(net1105),
    .B(net1110),
    .C(net1062),
    .D(_3122_),
    .Y(_3124_));
 sg13g2_a21oi_1 _3863_ (.A1(_3114_),
    .A2(_3116_),
    .Y(_3125_),
    .B1(_3124_));
 sg13g2_o21ai_1 _3864_ (.B1(_3125_),
    .Y(_3126_),
    .A1(_2911_),
    .A2(_3113_));
 sg13g2_nand2b_1 _3865_ (.Y(_3127_),
    .B(_3126_),
    .A_N(_3100_));
 sg13g2_or2_1 _3866_ (.X(_3128_),
    .B(net1099),
    .A(net1097));
 sg13g2_a21oi_1 _3867_ (.A1(_2936_),
    .A2(_3113_),
    .Y(_3129_),
    .B1(_3128_));
 sg13g2_nor2b_2 _3868_ (.A(net1099),
    .B_N(net1097),
    .Y(_3130_));
 sg13g2_nand2b_2 _3869_ (.Y(_3131_),
    .B(net1097),
    .A_N(net1099));
 sg13g2_nor2_1 _3870_ (.A(net1112),
    .B(_2914_),
    .Y(_3132_));
 sg13g2_nand2b_2 _3871_ (.Y(_3133_),
    .B(net1114),
    .A_N(net1112));
 sg13g2_nor2_1 _3872_ (.A(net1092),
    .B(_3133_),
    .Y(_3134_));
 sg13g2_nand2_2 _3873_ (.Y(_3135_),
    .A(_2913_),
    .B(_3119_));
 sg13g2_o21ai_1 _3874_ (.B1(_3130_),
    .Y(_3136_),
    .A1(net1101),
    .A2(_3135_));
 sg13g2_nor2_1 _3875_ (.A(_2911_),
    .B(net1109),
    .Y(_3137_));
 sg13g2_a21oi_1 _3876_ (.A1(_3112_),
    .A2(_3137_),
    .Y(_3138_),
    .B1(_3136_));
 sg13g2_nand2_1 _3877_ (.Y(_3139_),
    .A(_0071_),
    .B(net1027));
 sg13g2_and2_1 _3878_ (.A(net1097),
    .B(net1099),
    .X(_3140_));
 sg13g2_nand2_1 _3879_ (.Y(_3141_),
    .A(net1097),
    .B(net1099));
 sg13g2_nor2_2 _3880_ (.A(net1104),
    .B(net1062),
    .Y(_3142_));
 sg13g2_a21oi_1 _3881_ (.A1(_3114_),
    .A2(_3121_),
    .Y(_3143_),
    .B1(_3142_));
 sg13g2_nor2_2 _3882_ (.A(net1094),
    .B(net1114),
    .Y(_3144_));
 sg13g2_or2_1 _3883_ (.X(_3145_),
    .B(net1114),
    .A(net1093));
 sg13g2_nand2_1 _3884_ (.Y(_3146_),
    .A(_2937_),
    .B(_3144_));
 sg13g2_o21ai_1 _3885_ (.B1(net1104),
    .Y(_3147_),
    .A1(_0086_),
    .A2(_3146_));
 sg13g2_a21oi_1 _3886_ (.A1(_3143_),
    .A2(_3147_),
    .Y(_3148_),
    .B1(_3141_));
 sg13g2_nor4_1 _3887_ (.A(_3129_),
    .B(_3138_),
    .C(net1002),
    .D(_3148_),
    .Y(_3149_));
 sg13g2_a22oi_1 _3888_ (.Y(_3150_),
    .B1(_3127_),
    .B2(_3149_),
    .A2(net1024),
    .A1(_0032_));
 sg13g2_and2_1 _3889_ (.A(_0072_),
    .B(net1021),
    .X(_3151_));
 sg13g2_nand2_2 _3890_ (.Y(_3152_),
    .A(_0072_),
    .B(net1021));
 sg13g2_a21o_2 _3891_ (.A2(net1114),
    .A1(net1093),
    .B1(net1112),
    .X(_3153_));
 sg13g2_nand2b_2 _3892_ (.Y(_3154_),
    .B(_0071_),
    .A_N(net1101));
 sg13g2_nand2_1 _3893_ (.Y(_3155_),
    .A(net1096),
    .B(net1107));
 sg13g2_nor4_1 _3894_ (.A(net1061),
    .B(_3144_),
    .C(_3153_),
    .D(_3154_),
    .Y(_3156_));
 sg13g2_nor3_2 _3895_ (.A(net1090),
    .B(net1061),
    .C(_3154_),
    .Y(_3157_));
 sg13g2_nand2b_2 _3896_ (.Y(_3158_),
    .B(_3156_),
    .A_N(_3155_));
 sg13g2_nand2_1 _3897_ (.Y(_3159_),
    .A(net1096),
    .B(net1113));
 sg13g2_nor2_1 _3898_ (.A(_3145_),
    .B(_3159_),
    .Y(_3160_));
 sg13g2_nor3_2 _3899_ (.A(net1107),
    .B(net1061),
    .C(_3154_),
    .Y(_3161_));
 sg13g2_nor2_1 _3900_ (.A(_3109_),
    .B(_3121_),
    .Y(_3162_));
 sg13g2_a22oi_1 _3901_ (.Y(_3163_),
    .B1(_3162_),
    .B2(_3157_),
    .A2(_3161_),
    .A1(_3160_));
 sg13g2_nand4_1 _3902_ (.B(net1100),
    .C(net1106),
    .A(net1098),
    .Y(_3164_),
    .D(net1111));
 sg13g2_nor4_2 _3903_ (.A(\i_display.x_idx[8] ),
    .B(_3145_),
    .C(_3159_),
    .Y(_3165_),
    .D(_3164_));
 sg13g2_inv_1 _3904_ (.Y(_3166_),
    .A(_3165_));
 sg13g2_nand3b_1 _3905_ (.B(_0071_),
    .C(net1102),
    .Y(_3167_),
    .A_N(net1108));
 sg13g2_nor4_2 _3906_ (.A(net1092),
    .B(_3133_),
    .C(net1060),
    .Y(_3168_),
    .D(_3167_));
 sg13g2_nor4_2 _3907_ (.A(\i_display.hsync ),
    .B(_3000_),
    .C(_3165_),
    .Y(_3169_),
    .D(_3168_));
 sg13g2_nand2_1 _3908_ (.Y(_3170_),
    .A(_3134_),
    .B(_3161_));
 sg13g2_nor4_2 _3909_ (.A(_3109_),
    .B(_3118_),
    .C(net1061),
    .Y(_3171_),
    .D(_3154_));
 sg13g2_nor2_1 _3910_ (.A(_2913_),
    .B(_3102_),
    .Y(_3172_));
 sg13g2_nor2_1 _3911_ (.A(_3102_),
    .B(_3118_),
    .Y(_3173_));
 sg13g2_nor2_1 _3912_ (.A(_3109_),
    .B(_3133_),
    .Y(_3174_));
 sg13g2_a221oi_1 _3913_ (.B2(_3161_),
    .C1(_3171_),
    .B1(_3174_),
    .A1(_3157_),
    .Y(_3175_),
    .A2(_3173_));
 sg13g2_and4_1 _3914_ (.A(_3158_),
    .B(_3163_),
    .C(_3169_),
    .D(_3175_),
    .X(_3176_));
 sg13g2_nand4_1 _3915_ (.B(_3163_),
    .C(_3169_),
    .A(_3158_),
    .Y(_3177_),
    .D(_3175_));
 sg13g2_nor2_2 _3916_ (.A(_3151_),
    .B(_3176_),
    .Y(_3178_));
 sg13g2_inv_1 _3917_ (.Y(_3179_),
    .A(net1000));
 sg13g2_nand3_1 _3918_ (.B(_3152_),
    .C(_3177_),
    .A(net1116),
    .Y(_3180_));
 sg13g2_nor2_1 _3919_ (.A(_3102_),
    .B(_3121_),
    .Y(_3181_));
 sg13g2_nand3_1 _3920_ (.B(net1107),
    .C(_0071_),
    .A(net1101),
    .Y(_3182_));
 sg13g2_nor4_2 _3921_ (.A(_3102_),
    .B(_3121_),
    .C(net1060),
    .Y(_3183_),
    .D(_3182_));
 sg13g2_nor3_1 _3922_ (.A(\i_display.hsync ),
    .B(_3000_),
    .C(_3183_),
    .Y(_3184_));
 sg13g2_or2_1 _3923_ (.X(_3185_),
    .B(_3154_),
    .A(_3131_));
 sg13g2_nand3b_1 _3924_ (.B(net1107),
    .C(_0071_),
    .Y(_3186_),
    .A_N(net1101));
 sg13g2_nor2_1 _3925_ (.A(_3131_),
    .B(_3186_),
    .Y(_3187_));
 sg13g2_nand2b_2 _3926_ (.Y(_3188_),
    .B(net1092),
    .A_N(net1096));
 sg13g2_nor4_1 _3927_ (.A(_3131_),
    .B(_3133_),
    .C(_3186_),
    .D(_3188_),
    .Y(_3189_));
 sg13g2_nand2_1 _3928_ (.Y(_3190_),
    .A(net1094),
    .B(net1096));
 sg13g2_nand4_1 _3929_ (.B(net1096),
    .C(_3132_),
    .A(net1092),
    .Y(_3191_),
    .D(_3187_));
 sg13g2_nand3_1 _3930_ (.B(_3132_),
    .C(_3187_),
    .A(net1092),
    .Y(_3192_));
 sg13g2_and3_2 _3931_ (.X(_3193_),
    .A(_3170_),
    .B(_3184_),
    .C(_3192_));
 sg13g2_a22oi_1 _3932_ (.Y(_3194_),
    .B1(_3181_),
    .B2(_3157_),
    .A2(_3172_),
    .A1(_3161_));
 sg13g2_and2_1 _3933_ (.A(_3163_),
    .B(_3194_),
    .X(_3195_));
 sg13g2_nor2_1 _3934_ (.A(_3153_),
    .B(_3182_),
    .Y(_3196_));
 sg13g2_nor3_1 _3935_ (.A(net1092),
    .B(_3120_),
    .C(_3167_),
    .Y(_3197_));
 sg13g2_o21ai_1 _3936_ (.B1(_3130_),
    .Y(_3198_),
    .A1(_3196_),
    .A2(_3197_));
 sg13g2_and4_2 _3937_ (.A(_3163_),
    .B(_3166_),
    .C(_3194_),
    .D(_3198_),
    .X(_3199_));
 sg13g2_a22oi_1 _3938_ (.Y(_3200_),
    .B1(_3193_),
    .B2(_3199_),
    .A2(net1021),
    .A1(_0070_));
 sg13g2_inv_1 _3939_ (.Y(_3201_),
    .A(_3200_));
 sg13g2_a221oi_1 _3940_ (.B2(_3199_),
    .C1(_0095_),
    .B1(_3193_),
    .A1(_0070_),
    .Y(_3202_),
    .A2(net1021));
 sg13g2_nand2b_1 _3941_ (.Y(_3203_),
    .B(_3202_),
    .A_N(_3180_));
 sg13g2_nor4_2 _3942_ (.A(_3100_),
    .B(_3102_),
    .C(_3118_),
    .Y(_3204_),
    .D(_3182_));
 sg13g2_nor2_1 _3943_ (.A(_3171_),
    .B(_3204_),
    .Y(_3205_));
 sg13g2_nand2b_1 _3944_ (.Y(_3206_),
    .B(net1114),
    .A_N(net1107));
 sg13g2_or4_1 _3945_ (.A(_3109_),
    .B(net1060),
    .C(_3154_),
    .D(_3206_),
    .X(_3207_));
 sg13g2_nor4_1 _3946_ (.A(net1060),
    .B(_3154_),
    .C(_3188_),
    .D(_3206_),
    .Y(_3208_));
 sg13g2_nor3_1 _3947_ (.A(_3165_),
    .B(_3168_),
    .C(_3208_),
    .Y(_3209_));
 sg13g2_nor3_1 _3948_ (.A(_3171_),
    .B(_3189_),
    .C(_3204_),
    .Y(_3210_));
 sg13g2_and3_1 _3949_ (.X(_3211_),
    .A(_3198_),
    .B(_3207_),
    .C(_3210_));
 sg13g2_a221oi_1 _3950_ (.B2(_3187_),
    .C1(\i_display.hsync ),
    .B1(_3174_),
    .A1(_2993_),
    .Y(_3212_),
    .A2(_3001_));
 sg13g2_and4_1 _3951_ (.A(_3158_),
    .B(_3163_),
    .C(_3209_),
    .D(_3212_),
    .X(_3213_));
 sg13g2_a22oi_1 _3952_ (.Y(_3214_),
    .B1(_3211_),
    .B2(_3213_),
    .A2(net1023),
    .A1(_0073_));
 sg13g2_nand2_1 _3953_ (.Y(_3215_),
    .A(net1120),
    .B(net999));
 sg13g2_a21oi_1 _3954_ (.A1(\i_display.frame[7] ),
    .A2(_3178_),
    .Y(_3216_),
    .B1(_3202_));
 sg13g2_xnor2_1 _3955_ (.Y(_3217_),
    .A(_3180_),
    .B(_3202_));
 sg13g2_o21ai_1 _3956_ (.B1(_3203_),
    .Y(_3218_),
    .A1(_3215_),
    .A2(_3216_));
 sg13g2_nand2_1 _3957_ (.Y(_3219_),
    .A(net1118),
    .B(_3214_));
 sg13g2_a221oi_1 _3958_ (.B2(_3199_),
    .C1(_0028_),
    .B1(_3193_),
    .A1(_0070_),
    .Y(_3220_),
    .A2(net1022));
 sg13g2_nand3_1 _3959_ (.B(_3152_),
    .C(_3177_),
    .A(\i_display.frame[8] ),
    .Y(_3221_));
 sg13g2_nand3_1 _3960_ (.B(_3178_),
    .C(_3220_),
    .A(\i_display.frame[8] ),
    .Y(_3222_));
 sg13g2_xor2_1 _3961_ (.B(_3221_),
    .A(_3220_),
    .X(_3223_));
 sg13g2_xor2_1 _3962_ (.B(_3223_),
    .A(_3219_),
    .X(_3224_));
 sg13g2_nand2_1 _3963_ (.Y(_3225_),
    .A(_3218_),
    .B(_3224_));
 sg13g2_nor2_1 _3964_ (.A(_3102_),
    .B(_3133_),
    .Y(_3226_));
 sg13g2_a22oi_1 _3965_ (.Y(_3227_),
    .B1(_3226_),
    .B2(_3161_),
    .A2(_3173_),
    .A1(_3157_));
 sg13g2_nand3_1 _3966_ (.B(_3194_),
    .C(_3227_),
    .A(_3163_),
    .Y(_3228_));
 sg13g2_nand2_1 _3967_ (.Y(_3229_),
    .A(_3166_),
    .B(_3207_));
 sg13g2_nor4_1 _3968_ (.A(net1023),
    .B(_3204_),
    .C(_3228_),
    .D(_3229_),
    .Y(_3230_));
 sg13g2_a21oi_2 _3969_ (.B1(_3230_),
    .Y(_3231_),
    .A2(net1023),
    .A1(_0080_));
 sg13g2_inv_1 _3970_ (.Y(_3232_),
    .A(_3231_));
 sg13g2_nand2_1 _3971_ (.Y(_3233_),
    .A(net1121),
    .B(net993));
 sg13g2_nor2_1 _3972_ (.A(_3121_),
    .B(_3188_),
    .Y(_3234_));
 sg13g2_nand2_1 _3973_ (.Y(_3235_),
    .A(net1107),
    .B(_3171_));
 sg13g2_o21ai_1 _3974_ (.B1(_3157_),
    .Y(_3236_),
    .A1(_3226_),
    .A2(_3234_));
 sg13g2_and3_1 _3975_ (.X(_3237_),
    .A(_3158_),
    .B(_3235_),
    .C(_3236_));
 sg13g2_a22oi_1 _3976_ (.Y(_3238_),
    .B1(_3193_),
    .B2(_3237_),
    .A2(net1023),
    .A1(_0076_));
 sg13g2_nand2_1 _3977_ (.Y(_3239_),
    .A(net1116),
    .B(net998));
 sg13g2_and4_1 _3978_ (.A(net1027),
    .B(_3191_),
    .C(_3205_),
    .D(_3209_),
    .X(_3240_));
 sg13g2_a22oi_1 _3979_ (.Y(_3241_),
    .B1(_3195_),
    .B2(_3240_),
    .A2(net1023),
    .A1(_0078_));
 sg13g2_nand2_1 _3980_ (.Y(_3242_),
    .A(net1120),
    .B(net996));
 sg13g2_xor2_1 _3981_ (.B(_3242_),
    .A(_3239_),
    .X(_3243_));
 sg13g2_nand2b_1 _3982_ (.Y(_3244_),
    .B(_3243_),
    .A_N(_3233_));
 sg13g2_xor2_1 _3983_ (.B(_3243_),
    .A(_3233_),
    .X(_3245_));
 sg13g2_xnor2_1 _3984_ (.Y(_3246_),
    .A(_3218_),
    .B(_3224_));
 sg13g2_o21ai_1 _3985_ (.B1(_3225_),
    .Y(_3247_),
    .A1(_3245_),
    .A2(_3246_));
 sg13g2_nand2_1 _3986_ (.Y(_3248_),
    .A(net1120),
    .B(net993));
 sg13g2_nand2_1 _3987_ (.Y(_3249_),
    .A(\i_display.frame[8] ),
    .B(net998));
 sg13g2_nand2_1 _3988_ (.Y(_3250_),
    .A(net1118),
    .B(net996));
 sg13g2_xor2_1 _3989_ (.B(_3250_),
    .A(_3249_),
    .X(_3251_));
 sg13g2_nand2b_1 _3990_ (.Y(_3252_),
    .B(_3251_),
    .A_N(_3248_));
 sg13g2_xnor2_1 _3991_ (.Y(_3253_),
    .A(_3248_),
    .B(_3251_));
 sg13g2_nand2_2 _3992_ (.Y(_3254_),
    .A(\i_display.frame[9] ),
    .B(net999));
 sg13g2_nor2_1 _3993_ (.A(_3180_),
    .B(_3254_),
    .Y(_3255_));
 sg13g2_a22oi_1 _3994_ (.Y(_3256_),
    .B1(net999),
    .B2(net1116),
    .A2(_3178_),
    .A1(\i_display.frame[9] ));
 sg13g2_nor2_1 _3995_ (.A(_3255_),
    .B(_3256_),
    .Y(_3257_));
 sg13g2_o21ai_1 _3996_ (.B1(_3222_),
    .Y(_3258_),
    .A1(_3219_),
    .A2(_3223_));
 sg13g2_and2_1 _3997_ (.A(_3257_),
    .B(_3258_),
    .X(_3259_));
 sg13g2_xor2_1 _3998_ (.B(_3258_),
    .A(_3257_),
    .X(_3260_));
 sg13g2_xnor2_1 _3999_ (.Y(_3261_),
    .A(_3253_),
    .B(_3260_));
 sg13g2_nand2b_1 _4000_ (.Y(_3262_),
    .B(_3247_),
    .A_N(_3261_));
 sg13g2_nand3_1 _4001_ (.B(_3198_),
    .C(_3207_),
    .A(_3192_),
    .Y(_3263_));
 sg13g2_o21ai_1 _4002_ (.B1(_3169_),
    .Y(_3264_),
    .A1(_3135_),
    .A2(_3185_));
 sg13g2_nor4_1 _4003_ (.A(_3204_),
    .B(_3228_),
    .C(_3263_),
    .D(_3264_),
    .Y(_3265_));
 sg13g2_a21o_2 _4004_ (.A2(net1023),
    .A1(_0090_),
    .B1(_3265_),
    .X(_3266_));
 sg13g2_inv_1 _4005_ (.Y(_3267_),
    .A(_3266_));
 sg13g2_nor2_1 _4006_ (.A(_0075_),
    .B(net992),
    .Y(_3268_));
 sg13g2_nor4_1 _4007_ (.A(net1023),
    .B(_3183_),
    .C(_3228_),
    .D(_3263_),
    .Y(_3269_));
 sg13g2_a21o_2 _4008_ (.A2(net1023),
    .A1(_0093_),
    .B1(_3269_),
    .X(_3270_));
 sg13g2_inv_2 _4009_ (.Y(_3271_),
    .A(_3270_));
 sg13g2_nor2_1 _4010_ (.A(net1125),
    .B(_3270_),
    .Y(_3272_));
 sg13g2_and2_1 _4011_ (.A(_3268_),
    .B(_3272_),
    .X(_3273_));
 sg13g2_o21ai_1 _4012_ (.B1(_3244_),
    .Y(_3274_),
    .A1(_3239_),
    .A2(_3242_));
 sg13g2_nor2_1 _4013_ (.A(_0074_),
    .B(net992),
    .Y(_3275_));
 sg13g2_nor2_1 _4014_ (.A(net1124),
    .B(_3270_),
    .Y(_3276_));
 sg13g2_and2_1 _4015_ (.A(_3275_),
    .B(_3276_),
    .X(_3277_));
 sg13g2_xor2_1 _4016_ (.B(_3276_),
    .A(_3275_),
    .X(_3278_));
 sg13g2_and2_1 _4017_ (.A(_3274_),
    .B(_3278_),
    .X(_3279_));
 sg13g2_xor2_1 _4018_ (.B(_3278_),
    .A(_3274_),
    .X(_3280_));
 sg13g2_xnor2_1 _4019_ (.Y(_3281_),
    .A(_3273_),
    .B(_3280_));
 sg13g2_xor2_1 _4020_ (.B(_3261_),
    .A(_3247_),
    .X(_3282_));
 sg13g2_o21ai_1 _4021_ (.B1(_3262_),
    .Y(_3283_),
    .A1(_3281_),
    .A2(_3282_));
 sg13g2_o21ai_1 _4022_ (.B1(_3252_),
    .Y(_3284_),
    .A1(_3249_),
    .A2(_3250_));
 sg13g2_nor2_1 _4023_ (.A(_0069_),
    .B(net992),
    .Y(_3285_));
 sg13g2_nor2_1 _4024_ (.A(net1122),
    .B(_3270_),
    .Y(_3286_));
 sg13g2_and2_1 _4025_ (.A(_3285_),
    .B(_3286_),
    .X(_3287_));
 sg13g2_inv_1 _4026_ (.Y(_3288_),
    .A(_3287_));
 sg13g2_xor2_1 _4027_ (.B(_3286_),
    .A(_3285_),
    .X(_3289_));
 sg13g2_xor2_1 _4028_ (.B(_3289_),
    .A(_3284_),
    .X(_3290_));
 sg13g2_and2_1 _4029_ (.A(_3277_),
    .B(_3290_),
    .X(_3291_));
 sg13g2_xnor2_1 _4030_ (.Y(_3292_),
    .A(_3277_),
    .B(_3290_));
 sg13g2_a21o_1 _4031_ (.A2(_3260_),
    .A1(_3253_),
    .B1(_3259_),
    .X(_3293_));
 sg13g2_a21oi_1 _4032_ (.A1(_2941_),
    .A2(net999),
    .Y(_3294_),
    .B1(_3255_));
 sg13g2_a21oi_1 _4033_ (.A1(_2941_),
    .A2(_3255_),
    .Y(_3295_),
    .B1(_3294_));
 sg13g2_nand2_1 _4034_ (.Y(_3296_),
    .A(net1118),
    .B(_3231_));
 sg13g2_nand2_1 _4035_ (.Y(_3297_),
    .A(\i_display.frame[9] ),
    .B(net996));
 sg13g2_nand2_1 _4036_ (.Y(_3298_),
    .A(\i_display.frame[9] ),
    .B(net998));
 sg13g2_nand2_1 _4037_ (.Y(_3299_),
    .A(net1116),
    .B(net996));
 sg13g2_xor2_1 _4038_ (.B(_3299_),
    .A(_3298_),
    .X(_3300_));
 sg13g2_nand2b_1 _4039_ (.Y(_3301_),
    .B(_3300_),
    .A_N(_3296_));
 sg13g2_xnor2_1 _4040_ (.Y(_3302_),
    .A(_3296_),
    .B(_3300_));
 sg13g2_xor2_1 _4041_ (.B(_3302_),
    .A(_3295_),
    .X(_3303_));
 sg13g2_nand2_1 _4042_ (.Y(_3304_),
    .A(_3293_),
    .B(_3303_));
 sg13g2_xnor2_1 _4043_ (.Y(_3305_),
    .A(_3293_),
    .B(_3303_));
 sg13g2_xor2_1 _4044_ (.B(_3305_),
    .A(_3292_),
    .X(_3306_));
 sg13g2_a21o_1 _4045_ (.A2(_3280_),
    .A1(_3273_),
    .B1(_3279_),
    .X(_3307_));
 sg13g2_xnor2_1 _4046_ (.Y(_3308_),
    .A(_3283_),
    .B(_3306_));
 sg13g2_nor2b_1 _4047_ (.A(_3308_),
    .B_N(_3307_),
    .Y(_3309_));
 sg13g2_a21o_1 _4048_ (.A2(_3306_),
    .A1(_3283_),
    .B1(_3309_),
    .X(_3310_));
 sg13g2_a21o_1 _4049_ (.A2(_3289_),
    .A1(_3284_),
    .B1(_3291_),
    .X(_3311_));
 sg13g2_o21ai_1 _4050_ (.B1(_3304_),
    .Y(_3312_),
    .A1(_3292_),
    .A2(_3305_));
 sg13g2_nand2_1 _4051_ (.Y(_3313_),
    .A(_2941_),
    .B(net996));
 sg13g2_nor2_1 _4052_ (.A(_0092_),
    .B(_3232_),
    .Y(_3314_));
 sg13g2_nor3_1 _4053_ (.A(_0092_),
    .B(_3232_),
    .C(_3313_),
    .Y(_3315_));
 sg13g2_xnor2_1 _4054_ (.Y(_3316_),
    .A(_3313_),
    .B(_3314_));
 sg13g2_nor2b_1 _4055_ (.A(_3254_),
    .B_N(_3316_),
    .Y(_0255_));
 sg13g2_xnor2_1 _4056_ (.Y(_0256_),
    .A(_3254_),
    .B(_3316_));
 sg13g2_a22oi_1 _4057_ (.Y(_0257_),
    .B1(_3295_),
    .B2(_3302_),
    .A2(_3255_),
    .A1(_2941_));
 sg13g2_nor2b_1 _4058_ (.A(_0257_),
    .B_N(_0256_),
    .Y(_0258_));
 sg13g2_xnor2_1 _4059_ (.Y(_0259_),
    .A(_0256_),
    .B(_0257_));
 sg13g2_o21ai_1 _4060_ (.B1(_3301_),
    .Y(_0260_),
    .A1(_3298_),
    .A2(_3299_));
 sg13g2_nor2_1 _4061_ (.A(_0089_),
    .B(net992),
    .Y(_0261_));
 sg13g2_nor2_1 _4062_ (.A(net1120),
    .B(_3270_),
    .Y(_0262_));
 sg13g2_and2_1 _4063_ (.A(_0261_),
    .B(_0262_),
    .X(_0263_));
 sg13g2_xor2_1 _4064_ (.B(_0262_),
    .A(_0261_),
    .X(_0264_));
 sg13g2_nand2_1 _4065_ (.Y(_0265_),
    .A(_0260_),
    .B(_0264_));
 sg13g2_xnor2_1 _4066_ (.Y(_0266_),
    .A(_0260_),
    .B(_0264_));
 sg13g2_xnor2_1 _4067_ (.Y(_0267_),
    .A(_3287_),
    .B(_0266_));
 sg13g2_xnor2_1 _4068_ (.Y(_0268_),
    .A(_0259_),
    .B(_0267_));
 sg13g2_inv_1 _4069_ (.Y(_0269_),
    .A(_0268_));
 sg13g2_xor2_1 _4070_ (.B(_0268_),
    .A(_3312_),
    .X(_0270_));
 sg13g2_nor2b_1 _4071_ (.A(_0270_),
    .B_N(_3311_),
    .Y(_0271_));
 sg13g2_xor2_1 _4072_ (.B(_0270_),
    .A(_3311_),
    .X(_0272_));
 sg13g2_nor2b_1 _4073_ (.A(_0272_),
    .B_N(_3310_),
    .Y(_0273_));
 sg13g2_a221oi_1 _4074_ (.B2(_3199_),
    .C1(_0092_),
    .B1(_3193_),
    .A1(_0070_),
    .Y(_0274_),
    .A2(net1021));
 sg13g2_nand3_1 _4075_ (.B(_3152_),
    .C(_3177_),
    .A(net1118),
    .Y(_0275_));
 sg13g2_nand3_1 _4076_ (.B(net1000),
    .C(_0274_),
    .A(net1117),
    .Y(_0276_));
 sg13g2_nand2_1 _4077_ (.Y(_0277_),
    .A(net1121),
    .B(_3214_));
 sg13g2_nor2b_1 _4078_ (.A(_0274_),
    .B_N(_0275_),
    .Y(_0278_));
 sg13g2_xnor2_1 _4079_ (.Y(_0279_),
    .A(_0274_),
    .B(_0275_));
 sg13g2_o21ai_1 _4080_ (.B1(_0276_),
    .Y(_0280_),
    .A1(_0277_),
    .A2(_0278_));
 sg13g2_xnor2_1 _4081_ (.Y(_0281_),
    .A(_3215_),
    .B(_3217_));
 sg13g2_nand2_1 _4082_ (.Y(_0282_),
    .A(_0280_),
    .B(_0281_));
 sg13g2_nand2_1 _4083_ (.Y(_0283_),
    .A(net1124),
    .B(net993));
 sg13g2_and4_1 _4084_ (.A(net1121),
    .B(_2938_),
    .C(net998),
    .D(net996),
    .X(_0284_));
 sg13g2_nand4_1 _4085_ (.B(_2938_),
    .C(net998),
    .A(net1121),
    .Y(_0285_),
    .D(net995));
 sg13g2_a22oi_1 _4086_ (.Y(_0286_),
    .B1(net995),
    .B2(net1121),
    .A2(net998),
    .A1(_2938_));
 sg13g2_nor2_1 _4087_ (.A(_0284_),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_xor2_1 _4088_ (.B(_0287_),
    .A(_0283_),
    .X(_0288_));
 sg13g2_xnor2_1 _4089_ (.Y(_0289_),
    .A(_0280_),
    .B(_0281_));
 sg13g2_o21ai_1 _4090_ (.B1(_0282_),
    .Y(_0290_),
    .A1(_0288_),
    .A2(_0289_));
 sg13g2_xnor2_1 _4091_ (.Y(_0291_),
    .A(_3245_),
    .B(_3246_));
 sg13g2_nand2b_1 _4092_ (.Y(_0292_),
    .B(_0290_),
    .A_N(_0291_));
 sg13g2_nor2_1 _4093_ (.A(_0081_),
    .B(net992),
    .Y(_0293_));
 sg13g2_nor2_1 _4094_ (.A(net1127),
    .B(_3270_),
    .Y(_0294_));
 sg13g2_and2_1 _4095_ (.A(_0293_),
    .B(_0294_),
    .X(_0295_));
 sg13g2_o21ai_1 _4096_ (.B1(_0285_),
    .Y(_0296_),
    .A1(_0283_),
    .A2(_0286_));
 sg13g2_xor2_1 _4097_ (.B(_3272_),
    .A(_3268_),
    .X(_0297_));
 sg13g2_and2_1 _4098_ (.A(_0296_),
    .B(_0297_),
    .X(_0298_));
 sg13g2_xor2_1 _4099_ (.B(_0297_),
    .A(_0296_),
    .X(_0299_));
 sg13g2_xnor2_1 _4100_ (.Y(_0300_),
    .A(_0295_),
    .B(_0299_));
 sg13g2_xor2_1 _4101_ (.B(_0291_),
    .A(_0290_),
    .X(_0301_));
 sg13g2_o21ai_1 _4102_ (.B1(_0292_),
    .Y(_0302_),
    .A1(_0300_),
    .A2(_0301_));
 sg13g2_xor2_1 _4103_ (.B(_3282_),
    .A(_3281_),
    .X(_0303_));
 sg13g2_a21o_1 _4104_ (.A2(_0299_),
    .A1(_0295_),
    .B1(_0298_),
    .X(_0304_));
 sg13g2_xnor2_1 _4105_ (.Y(_0305_),
    .A(_0302_),
    .B(_0303_));
 sg13g2_nor2b_1 _4106_ (.A(_0305_),
    .B_N(_0304_),
    .Y(_0306_));
 sg13g2_a21o_1 _4107_ (.A2(_0303_),
    .A1(_0302_),
    .B1(_0306_),
    .X(_0307_));
 sg13g2_xor2_1 _4108_ (.B(_3308_),
    .A(_3307_),
    .X(_0308_));
 sg13g2_nand2b_1 _4109_ (.Y(_0309_),
    .B(_0307_),
    .A_N(_0308_));
 sg13g2_a221oi_1 _4110_ (.B2(_3199_),
    .C1(_0089_),
    .B1(_3193_),
    .A1(_0070_),
    .Y(_0310_),
    .A2(net1021));
 sg13g2_nand3_1 _4111_ (.B(_3152_),
    .C(_3177_),
    .A(net1120),
    .Y(_0311_));
 sg13g2_nand3_1 _4112_ (.B(net1000),
    .C(_0310_),
    .A(net1119),
    .Y(_0312_));
 sg13g2_nand2_1 _4113_ (.Y(_0313_),
    .A(net1124),
    .B(net999));
 sg13g2_nor2b_1 _4114_ (.A(_0310_),
    .B_N(_0311_),
    .Y(_0314_));
 sg13g2_xnor2_1 _4115_ (.Y(_0315_),
    .A(_0310_),
    .B(_0311_));
 sg13g2_o21ai_1 _4116_ (.B1(_0312_),
    .Y(_0316_),
    .A1(_0313_),
    .A2(_0314_));
 sg13g2_xnor2_1 _4117_ (.Y(_0317_),
    .A(_0277_),
    .B(_0279_));
 sg13g2_nand2_1 _4118_ (.Y(_0318_),
    .A(_0316_),
    .B(_0317_));
 sg13g2_nand2_1 _4119_ (.Y(_0319_),
    .A(net1125),
    .B(net993));
 sg13g2_and4_1 _4120_ (.A(net1123),
    .B(_2932_),
    .C(net997),
    .D(net995),
    .X(_0320_));
 sg13g2_nand4_1 _4121_ (.B(_2932_),
    .C(net997),
    .A(net1123),
    .Y(_0321_),
    .D(net995));
 sg13g2_a22oi_1 _4122_ (.Y(_0322_),
    .B1(net995),
    .B2(net1123),
    .A2(net997),
    .A1(_2932_));
 sg13g2_nor2_1 _4123_ (.A(_0320_),
    .B(_0322_),
    .Y(_0323_));
 sg13g2_xor2_1 _4124_ (.B(_0323_),
    .A(_0319_),
    .X(_0324_));
 sg13g2_xnor2_1 _4125_ (.Y(_0325_),
    .A(_0316_),
    .B(_0317_));
 sg13g2_o21ai_1 _4126_ (.B1(_0318_),
    .Y(_0326_),
    .A1(_0324_),
    .A2(_0325_));
 sg13g2_xnor2_1 _4127_ (.Y(_0327_),
    .A(_0288_),
    .B(_0289_));
 sg13g2_nand2b_1 _4128_ (.Y(_0328_),
    .B(_0326_),
    .A_N(_0327_));
 sg13g2_nor2_1 _4129_ (.A(_0077_),
    .B(net992),
    .Y(_0329_));
 sg13g2_o21ai_1 _4130_ (.B1(_3271_),
    .Y(_0330_),
    .A1(_0079_),
    .A2(_0329_));
 sg13g2_o21ai_1 _4131_ (.B1(_0321_),
    .Y(_0331_),
    .A1(_0319_),
    .A2(_0322_));
 sg13g2_xor2_1 _4132_ (.B(_0294_),
    .A(_0293_),
    .X(_0332_));
 sg13g2_nand2_1 _4133_ (.Y(_0333_),
    .A(_0331_),
    .B(_0332_));
 sg13g2_xnor2_1 _4134_ (.Y(_0334_),
    .A(_0331_),
    .B(_0332_));
 sg13g2_xnor2_1 _4135_ (.Y(_0335_),
    .A(_0330_),
    .B(_0334_));
 sg13g2_xor2_1 _4136_ (.B(_0327_),
    .A(_0326_),
    .X(_0336_));
 sg13g2_o21ai_1 _4137_ (.B1(_0328_),
    .Y(_0337_),
    .A1(_0335_),
    .A2(_0336_));
 sg13g2_xor2_1 _4138_ (.B(_0301_),
    .A(_0300_),
    .X(_0338_));
 sg13g2_nand2_1 _4139_ (.Y(_0339_),
    .A(_0337_),
    .B(_0338_));
 sg13g2_o21ai_1 _4140_ (.B1(_0333_),
    .Y(_0340_),
    .A1(_0330_),
    .A2(_0334_));
 sg13g2_inv_1 _4141_ (.Y(_0341_),
    .A(_0340_));
 sg13g2_xnor2_1 _4142_ (.Y(_0342_),
    .A(_0337_),
    .B(_0338_));
 sg13g2_o21ai_1 _4143_ (.B1(_0339_),
    .Y(_0343_),
    .A1(_0341_),
    .A2(_0342_));
 sg13g2_xor2_1 _4144_ (.B(_0305_),
    .A(_0304_),
    .X(_0344_));
 sg13g2_nor2b_1 _4145_ (.A(_0344_),
    .B_N(_0343_),
    .Y(_0345_));
 sg13g2_inv_1 _4146_ (.Y(_0346_),
    .A(_0345_));
 sg13g2_a221oi_1 _4147_ (.B2(_3199_),
    .C1(_0069_),
    .B1(_3193_),
    .A1(_0070_),
    .Y(_0347_),
    .A2(net1021));
 sg13g2_nand3_1 _4148_ (.B(_3152_),
    .C(_3177_),
    .A(net1121),
    .Y(_0348_));
 sg13g2_nand3_1 _4149_ (.B(net1000),
    .C(_0347_),
    .A(net1121),
    .Y(_0349_));
 sg13g2_nand2_1 _4150_ (.Y(_0350_),
    .A(net1125),
    .B(net999));
 sg13g2_nor2b_1 _4151_ (.A(_0347_),
    .B_N(_0348_),
    .Y(_0351_));
 sg13g2_xnor2_1 _4152_ (.Y(_0352_),
    .A(_0347_),
    .B(_0348_));
 sg13g2_o21ai_1 _4153_ (.B1(_0349_),
    .Y(_0353_),
    .A1(_0350_),
    .A2(_0351_));
 sg13g2_xnor2_1 _4154_ (.Y(_0354_),
    .A(_0313_),
    .B(_0315_));
 sg13g2_nand2_1 _4155_ (.Y(_0355_),
    .A(_0353_),
    .B(_0354_));
 sg13g2_nand2_1 _4156_ (.Y(_0356_),
    .A(net1128),
    .B(net993));
 sg13g2_nand2_1 _4157_ (.Y(_0357_),
    .A(net1125),
    .B(net997));
 sg13g2_nand2_1 _4158_ (.Y(_0358_),
    .A(net1125),
    .B(net995));
 sg13g2_nand2_1 _4159_ (.Y(_0359_),
    .A(net1121),
    .B(net998));
 sg13g2_xor2_1 _4160_ (.B(_0359_),
    .A(_0358_),
    .X(_0360_));
 sg13g2_nand2b_1 _4161_ (.Y(_0361_),
    .B(_0360_),
    .A_N(_0356_));
 sg13g2_xor2_1 _4162_ (.B(_0360_),
    .A(_0356_),
    .X(_0362_));
 sg13g2_xnor2_1 _4163_ (.Y(_0363_),
    .A(_0353_),
    .B(_0354_));
 sg13g2_o21ai_1 _4164_ (.B1(_0355_),
    .Y(_0364_),
    .A1(_0362_),
    .A2(_0363_));
 sg13g2_xnor2_1 _4165_ (.Y(_0365_),
    .A(_0324_),
    .B(_0325_));
 sg13g2_nand2b_1 _4166_ (.Y(_0366_),
    .B(_0364_),
    .A_N(_0365_));
 sg13g2_o21ai_1 _4167_ (.B1(_0361_),
    .Y(_0367_),
    .A1(_0358_),
    .A2(_0359_));
 sg13g2_nor2_1 _4168_ (.A(_0079_),
    .B(_3270_),
    .Y(_0368_));
 sg13g2_xor2_1 _4169_ (.B(_0368_),
    .A(_0329_),
    .X(_0369_));
 sg13g2_nand2_1 _4170_ (.Y(_0370_),
    .A(_0367_),
    .B(_0369_));
 sg13g2_xnor2_1 _4171_ (.Y(_0371_),
    .A(_0367_),
    .B(_0369_));
 sg13g2_xor2_1 _4172_ (.B(_0365_),
    .A(_0364_),
    .X(_0372_));
 sg13g2_o21ai_1 _4173_ (.B1(_0366_),
    .Y(_0373_),
    .A1(_0371_),
    .A2(_0372_));
 sg13g2_xnor2_1 _4174_ (.Y(_0374_),
    .A(_0335_),
    .B(_0336_));
 sg13g2_nor2b_1 _4175_ (.A(_0374_),
    .B_N(_0373_),
    .Y(_0375_));
 sg13g2_xor2_1 _4176_ (.B(_0374_),
    .A(_0373_),
    .X(_0376_));
 sg13g2_nor2_1 _4177_ (.A(_0370_),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_xnor2_1 _4178_ (.Y(_0378_),
    .A(_0340_),
    .B(_0342_));
 sg13g2_nor3_1 _4179_ (.A(_0375_),
    .B(_0377_),
    .C(_0378_),
    .Y(_0379_));
 sg13g2_and4_1 _4180_ (.A(net1126),
    .B(_2933_),
    .C(net1000),
    .D(_3200_),
    .X(_0380_));
 sg13g2_nand4_1 _4181_ (.B(_2933_),
    .C(net1000),
    .A(net1125),
    .Y(_0381_),
    .D(_3200_));
 sg13g2_nand2_1 _4182_ (.Y(_0382_),
    .A(net1129),
    .B(net999));
 sg13g2_a22oi_1 _4183_ (.Y(_0383_),
    .B1(_3200_),
    .B2(_2933_),
    .A2(net1000),
    .A1(net1125));
 sg13g2_nor3_1 _4184_ (.A(_0380_),
    .B(_0382_),
    .C(_0383_),
    .Y(_0384_));
 sg13g2_o21ai_1 _4185_ (.B1(_0381_),
    .Y(_0385_),
    .A1(_0382_),
    .A2(_0383_));
 sg13g2_nand2_1 _4186_ (.Y(_0386_),
    .A(net1127),
    .B(net999));
 sg13g2_a221oi_1 _4187_ (.B2(_3199_),
    .C1(_0074_),
    .B1(_3193_),
    .A1(_0070_),
    .Y(_0387_),
    .A2(net1021));
 sg13g2_nor3_1 _4188_ (.A(_2917_),
    .B(_3151_),
    .C(_3176_),
    .Y(_0388_));
 sg13g2_nand2_1 _4189_ (.Y(_0389_),
    .A(_0387_),
    .B(_0388_));
 sg13g2_xnor2_1 _4190_ (.Y(_0390_),
    .A(_0387_),
    .B(_0388_));
 sg13g2_xor2_1 _4191_ (.B(_0390_),
    .A(_0386_),
    .X(_0391_));
 sg13g2_nand2_1 _4192_ (.Y(_0392_),
    .A(_0385_),
    .B(_0391_));
 sg13g2_nand2_1 _4193_ (.Y(_0393_),
    .A(net1129),
    .B(net995));
 sg13g2_or2_1 _4194_ (.X(_0394_),
    .B(_0393_),
    .A(_0357_));
 sg13g2_xnor2_1 _4195_ (.Y(_0395_),
    .A(_0357_),
    .B(_0393_));
 sg13g2_xnor2_1 _4196_ (.Y(_0396_),
    .A(_0385_),
    .B(_0391_));
 sg13g2_o21ai_1 _4197_ (.B1(_0392_),
    .Y(_0397_),
    .A1(_0395_),
    .A2(_0396_));
 sg13g2_nand2b_1 _4198_ (.Y(_0398_),
    .B(net993),
    .A_N(_0079_));
 sg13g2_and2_1 _4199_ (.A(_2933_),
    .B(net997),
    .X(_0399_));
 sg13g2_and2_1 _4200_ (.A(_2934_),
    .B(net995),
    .X(_0400_));
 sg13g2_xor2_1 _4201_ (.B(_0400_),
    .A(_0399_),
    .X(_0401_));
 sg13g2_nor2b_1 _4202_ (.A(_0398_),
    .B_N(_0401_),
    .Y(_0402_));
 sg13g2_xor2_1 _4203_ (.B(_0401_),
    .A(_0398_),
    .X(_0403_));
 sg13g2_o21ai_1 _4204_ (.B1(_0389_),
    .Y(_0404_),
    .A1(_0386_),
    .A2(_0390_));
 sg13g2_xnor2_1 _4205_ (.Y(_0405_),
    .A(_0350_),
    .B(_0352_));
 sg13g2_nand2_1 _4206_ (.Y(_0406_),
    .A(_0404_),
    .B(_0405_));
 sg13g2_xnor2_1 _4207_ (.Y(_0407_),
    .A(_0404_),
    .B(_0405_));
 sg13g2_xor2_1 _4208_ (.B(_0407_),
    .A(_0403_),
    .X(_0408_));
 sg13g2_nand2_1 _4209_ (.Y(_0409_),
    .A(_0397_),
    .B(_0408_));
 sg13g2_xnor2_1 _4210_ (.Y(_0410_),
    .A(_0397_),
    .B(_0408_));
 sg13g2_o21ai_1 _4211_ (.B1(_0409_),
    .Y(_0411_),
    .A1(_0394_),
    .A2(_0410_));
 sg13g2_a21oi_2 _4212_ (.B1(_0402_),
    .Y(_0412_),
    .A2(_0400_),
    .A1(_0399_));
 sg13g2_nor2_1 _4213_ (.A(_0079_),
    .B(net992),
    .Y(_0413_));
 sg13g2_nand2b_1 _4214_ (.Y(_0414_),
    .B(_0413_),
    .A_N(_0412_));
 sg13g2_xor2_1 _4215_ (.B(_0413_),
    .A(_0412_),
    .X(_0415_));
 sg13g2_o21ai_1 _4216_ (.B1(_0406_),
    .Y(_0416_),
    .A1(_0403_),
    .A2(_0407_));
 sg13g2_xnor2_1 _4217_ (.Y(_0417_),
    .A(_0362_),
    .B(_0363_));
 sg13g2_nand2b_1 _4218_ (.Y(_0418_),
    .B(_0416_),
    .A_N(_0417_));
 sg13g2_xor2_1 _4219_ (.B(_0417_),
    .A(_0416_),
    .X(_0419_));
 sg13g2_xor2_1 _4220_ (.B(_0419_),
    .A(_0415_),
    .X(_0420_));
 sg13g2_nand2_1 _4221_ (.Y(_0421_),
    .A(_0411_),
    .B(_0420_));
 sg13g2_o21ai_1 _4222_ (.B1(_0418_),
    .Y(_0422_),
    .A1(_0415_),
    .A2(_0419_));
 sg13g2_xnor2_1 _4223_ (.Y(_0423_),
    .A(_0371_),
    .B(_0372_));
 sg13g2_nand2b_1 _4224_ (.Y(_0424_),
    .B(_0422_),
    .A_N(_0423_));
 sg13g2_xor2_1 _4225_ (.B(_0423_),
    .A(_0422_),
    .X(_0425_));
 sg13g2_xor2_1 _4226_ (.B(_0425_),
    .A(_0414_),
    .X(_0426_));
 sg13g2_nor2b_1 _4227_ (.A(_0421_),
    .B_N(_0426_),
    .Y(_0427_));
 sg13g2_o21ai_1 _4228_ (.B1(_0382_),
    .Y(_0428_),
    .A1(_0380_),
    .A2(_0383_));
 sg13g2_nor2b_1 _4229_ (.A(_0384_),
    .B_N(_0428_),
    .Y(_0429_));
 sg13g2_nor4_2 _4230_ (.A(_0077_),
    .B(_0081_),
    .C(_3179_),
    .Y(_0430_),
    .D(_3201_));
 sg13g2_nand2_1 _4231_ (.Y(_0431_),
    .A(_0429_),
    .B(_0430_));
 sg13g2_nand2_1 _4232_ (.Y(_0432_),
    .A(net1127),
    .B(net997));
 sg13g2_xnor2_1 _4233_ (.Y(_0433_),
    .A(_0429_),
    .B(_0430_));
 sg13g2_or2_1 _4234_ (.X(_0434_),
    .B(_0433_),
    .A(_0432_));
 sg13g2_xnor2_1 _4235_ (.Y(_0435_),
    .A(_0395_),
    .B(_0396_));
 sg13g2_a21oi_2 _4236_ (.B1(_0435_),
    .Y(_0436_),
    .A2(_0434_),
    .A1(_0431_));
 sg13g2_xor2_1 _4237_ (.B(_0410_),
    .A(_0394_),
    .X(_0437_));
 sg13g2_nand2_1 _4238_ (.Y(_0438_),
    .A(_0436_),
    .B(_0437_));
 sg13g2_xnor2_1 _4239_ (.Y(_0439_),
    .A(_0411_),
    .B(_0420_));
 sg13g2_or2_1 _4240_ (.X(_0440_),
    .B(_0439_),
    .A(_0438_));
 sg13g2_and3_1 _4241_ (.X(_0441_),
    .A(_0431_),
    .B(_0434_),
    .C(_0435_));
 sg13g2_nor4_1 _4242_ (.A(_2919_),
    .B(_0079_),
    .C(_3179_),
    .D(_3201_),
    .Y(_0442_));
 sg13g2_a22oi_1 _4243_ (.Y(_0443_),
    .B1(_3200_),
    .B2(_2935_),
    .A2(net1000),
    .A1(_2934_));
 sg13g2_or2_1 _4244_ (.X(_0444_),
    .B(_0443_),
    .A(_0430_));
 sg13g2_nand3_1 _4245_ (.B(net997),
    .C(_0442_),
    .A(net1129),
    .Y(_0445_));
 sg13g2_a21oi_1 _4246_ (.A1(net1129),
    .A2(net997),
    .Y(_0446_),
    .B1(_0442_));
 sg13g2_a221oi_1 _4247_ (.B2(_0445_),
    .C1(_0446_),
    .B1(_0444_),
    .A1(_0432_),
    .Y(_0447_),
    .A2(_0433_));
 sg13g2_nand2_1 _4248_ (.Y(_0448_),
    .A(_0434_),
    .B(_0447_));
 sg13g2_nor3_1 _4249_ (.A(_0436_),
    .B(_0441_),
    .C(_0448_),
    .Y(_0449_));
 sg13g2_nand2_1 _4250_ (.Y(_0450_),
    .A(_0437_),
    .B(_0449_));
 sg13g2_xnor2_1 _4251_ (.Y(_0451_),
    .A(_0438_),
    .B(_0439_));
 sg13g2_o21ai_1 _4252_ (.B1(_0440_),
    .Y(_0452_),
    .A1(_0450_),
    .A2(_0451_));
 sg13g2_xnor2_1 _4253_ (.Y(_0453_),
    .A(_0421_),
    .B(_0426_));
 sg13g2_a21oi_2 _4254_ (.B1(_0427_),
    .Y(_0454_),
    .A2(_0453_),
    .A1(_0452_));
 sg13g2_xor2_1 _4255_ (.B(_0376_),
    .A(_0370_),
    .X(_0455_));
 sg13g2_o21ai_1 _4256_ (.B1(_0424_),
    .Y(_0456_),
    .A1(_0414_),
    .A2(_0425_));
 sg13g2_nand2_1 _4257_ (.Y(_0457_),
    .A(_0455_),
    .B(_0456_));
 sg13g2_xor2_1 _4258_ (.B(_0456_),
    .A(_0455_),
    .X(_0458_));
 sg13g2_inv_1 _4259_ (.Y(_0459_),
    .A(_0458_));
 sg13g2_o21ai_1 _4260_ (.B1(_0378_),
    .Y(_0460_),
    .A1(_0375_),
    .A2(_0377_));
 sg13g2_and2_1 _4261_ (.A(_0457_),
    .B(_0460_),
    .X(_0461_));
 sg13g2_o21ai_1 _4262_ (.B1(_0461_),
    .Y(_0462_),
    .A1(_0454_),
    .A2(_0459_));
 sg13g2_nor2b_1 _4263_ (.A(_0379_),
    .B_N(_0462_),
    .Y(_0463_));
 sg13g2_xor2_1 _4264_ (.B(_0344_),
    .A(_0343_),
    .X(_0464_));
 sg13g2_inv_1 _4265_ (.Y(_0465_),
    .A(_0464_));
 sg13g2_nand3b_1 _4266_ (.B(_0462_),
    .C(_0465_),
    .Y(_0466_),
    .A_N(_0379_));
 sg13g2_xor2_1 _4267_ (.B(_0308_),
    .A(_0307_),
    .X(_0467_));
 sg13g2_a21o_1 _4268_ (.A2(_0466_),
    .A1(_0346_),
    .B1(_0467_),
    .X(_0468_));
 sg13g2_xor2_1 _4269_ (.B(_0272_),
    .A(_3310_),
    .X(_0469_));
 sg13g2_a21oi_2 _4270_ (.B1(_0469_),
    .Y(_0470_),
    .A2(_0468_),
    .A1(_0309_));
 sg13g2_a21oi_1 _4271_ (.A1(_3312_),
    .A2(_0269_),
    .Y(_0471_),
    .B1(_0271_));
 sg13g2_o21ai_1 _4272_ (.B1(_0265_),
    .Y(_0472_),
    .A1(_3288_),
    .A2(_0266_));
 sg13g2_a21o_1 _4273_ (.A2(_0267_),
    .A1(_0259_),
    .B1(_0258_),
    .X(_0473_));
 sg13g2_nand2_1 _4274_ (.Y(_0474_),
    .A(\i_display.frame[8] ),
    .B(net993));
 sg13g2_or2_1 _4275_ (.X(_0475_),
    .B(_0474_),
    .A(_3297_));
 sg13g2_xor2_1 _4276_ (.B(_0474_),
    .A(_3297_),
    .X(_0476_));
 sg13g2_xnor2_1 _4277_ (.Y(_0477_),
    .A(_0255_),
    .B(_0476_));
 sg13g2_nor2_1 _4278_ (.A(_0092_),
    .B(net992),
    .Y(_0478_));
 sg13g2_nor2_1 _4279_ (.A(net1117),
    .B(_3270_),
    .Y(_0479_));
 sg13g2_and2_1 _4280_ (.A(_0478_),
    .B(_0479_),
    .X(_0480_));
 sg13g2_xnor2_1 _4281_ (.Y(_0481_),
    .A(_0478_),
    .B(_0479_));
 sg13g2_nor4_1 _4282_ (.A(_0092_),
    .B(_3232_),
    .C(_3313_),
    .D(_0481_),
    .Y(_0482_));
 sg13g2_xnor2_1 _4283_ (.Y(_0483_),
    .A(_3315_),
    .B(_0481_));
 sg13g2_xnor2_1 _4284_ (.Y(_0484_),
    .A(_0263_),
    .B(_0483_));
 sg13g2_nor2_1 _4285_ (.A(_0477_),
    .B(_0484_),
    .Y(_0485_));
 sg13g2_xor2_1 _4286_ (.B(_0484_),
    .A(_0477_),
    .X(_0486_));
 sg13g2_and2_1 _4287_ (.A(_0473_),
    .B(_0486_),
    .X(_0487_));
 sg13g2_xor2_1 _4288_ (.B(_0486_),
    .A(_0473_),
    .X(_0488_));
 sg13g2_xnor2_1 _4289_ (.Y(_0489_),
    .A(_0472_),
    .B(_0488_));
 sg13g2_xor2_1 _4290_ (.B(_0489_),
    .A(_0471_),
    .X(_0490_));
 sg13g2_o21ai_1 _4291_ (.B1(_0490_),
    .Y(_0491_),
    .A1(_0273_),
    .A2(_0470_));
 sg13g2_or3_1 _4292_ (.A(_0273_),
    .B(_0470_),
    .C(_0490_),
    .X(_0492_));
 sg13g2_and2_1 _4293_ (.A(_0491_),
    .B(_0492_),
    .X(_0493_));
 sg13g2_nand2_1 _4294_ (.Y(_0494_),
    .A(_3150_),
    .B(_0493_));
 sg13g2_nand2_1 _4295_ (.Y(_0495_),
    .A(_0031_),
    .B(net1025));
 sg13g2_nor2_2 _4296_ (.A(net1110),
    .B(_3115_),
    .Y(_0496_));
 sg13g2_o21ai_1 _4297_ (.B1(net1108),
    .Y(_0497_),
    .A1(net1092),
    .A2(_3121_));
 sg13g2_a21oi_1 _4298_ (.A1(net1112),
    .A2(_3103_),
    .Y(_0498_),
    .B1(_0497_));
 sg13g2_nor2_1 _4299_ (.A(_0496_),
    .B(_0498_),
    .Y(_0499_));
 sg13g2_o21ai_1 _4300_ (.B1(net1103),
    .Y(_0500_),
    .A1(_0496_),
    .A2(_0498_));
 sg13g2_nor2_1 _4301_ (.A(_3101_),
    .B(_3144_),
    .Y(_0501_));
 sg13g2_a21oi_2 _4302_ (.B1(net1062),
    .Y(_0502_),
    .A2(_3144_),
    .A1(net1112));
 sg13g2_nor2b_2 _4303_ (.A(_3119_),
    .B_N(_3142_),
    .Y(_0503_));
 sg13g2_inv_1 _4304_ (.Y(_0504_),
    .A(_0503_));
 sg13g2_a22oi_1 _4305_ (.Y(_0505_),
    .B1(_0503_),
    .B2(net1109),
    .A2(_0502_),
    .A1(_3123_));
 sg13g2_a21oi_1 _4306_ (.A1(_0500_),
    .A2(_0505_),
    .Y(_0506_),
    .B1(_3100_));
 sg13g2_nor2_1 _4307_ (.A(net1115),
    .B(_3116_),
    .Y(_0507_));
 sg13g2_nor3_1 _4308_ (.A(net1115),
    .B(_0086_),
    .C(_3116_),
    .Y(_0508_));
 sg13g2_o21ai_1 _4309_ (.B1(_3143_),
    .Y(_0509_),
    .A1(_2911_),
    .A2(_0508_));
 sg13g2_a21oi_1 _4310_ (.A1(_2936_),
    .A2(_0499_),
    .Y(_0510_),
    .B1(net1061));
 sg13g2_a21oi_1 _4311_ (.A1(net1095),
    .A2(net1090),
    .Y(_0511_),
    .B1(_3133_));
 sg13g2_a21oi_1 _4312_ (.A1(_2911_),
    .A2(_0511_),
    .Y(_0512_),
    .B1(_3131_));
 sg13g2_nand3b_1 _4313_ (.B(_0497_),
    .C(net1103),
    .Y(_0513_),
    .A_N(_0496_));
 sg13g2_a221oi_1 _4314_ (.B2(_0513_),
    .C1(net1002),
    .B1(_0512_),
    .A1(_3140_),
    .Y(_0514_),
    .A2(_0509_));
 sg13g2_nand2b_1 _4315_ (.Y(_0515_),
    .B(_0514_),
    .A_N(_0510_));
 sg13g2_o21ai_1 _4316_ (.B1(_0495_),
    .Y(_0516_),
    .A1(_0506_),
    .A2(_0515_));
 sg13g2_nand3_1 _4317_ (.B(_0468_),
    .C(_0469_),
    .A(_0309_),
    .Y(_0517_));
 sg13g2_nand2b_1 _4318_ (.Y(_0518_),
    .B(_0517_),
    .A_N(_0470_));
 sg13g2_nor2_1 _4319_ (.A(_0516_),
    .B(_0518_),
    .Y(_0519_));
 sg13g2_o21ai_1 _4320_ (.B1(net1112),
    .Y(_0520_),
    .A1(net1062),
    .A2(_3119_));
 sg13g2_o21ai_1 _4321_ (.B1(net1090),
    .Y(_0521_),
    .A1(_0088_),
    .A2(_3109_));
 sg13g2_a21oi_1 _4322_ (.A1(_2913_),
    .A2(_3110_),
    .Y(_0522_),
    .B1(net1109));
 sg13g2_and2_1 _4323_ (.A(_0520_),
    .B(_0522_),
    .X(_0523_));
 sg13g2_nand2_1 _4324_ (.Y(_0524_),
    .A(net1108),
    .B(_3153_));
 sg13g2_o21ai_1 _4325_ (.B1(_3155_),
    .Y(_0525_),
    .A1(_3103_),
    .A2(_0524_));
 sg13g2_o21ai_1 _4326_ (.B1(net1102),
    .Y(_0526_),
    .A1(_0523_),
    .A2(_0525_));
 sg13g2_a21oi_1 _4327_ (.A1(net1110),
    .A2(_3121_),
    .Y(_0527_),
    .B1(_0496_));
 sg13g2_nor4_2 _4328_ (.A(net1100),
    .B(net1105),
    .C(_3119_),
    .Y(_0528_),
    .D(_0527_));
 sg13g2_nor2b_1 _4329_ (.A(net1106),
    .B_N(net1100),
    .Y(_0529_));
 sg13g2_nand2_1 _4330_ (.Y(_0530_),
    .A(net1090),
    .B(_3162_));
 sg13g2_nand3b_1 _4331_ (.B(_3159_),
    .C(_0530_),
    .Y(_0531_),
    .A_N(net1093));
 sg13g2_a21oi_1 _4332_ (.A1(_0529_),
    .A2(_0531_),
    .Y(_0532_),
    .B1(_0528_));
 sg13g2_a21oi_1 _4333_ (.A1(_0526_),
    .A2(_0532_),
    .Y(_0533_),
    .B1(net1097));
 sg13g2_nor2b_1 _4334_ (.A(_3181_),
    .B_N(_3114_),
    .Y(_0534_));
 sg13g2_o21ai_1 _4335_ (.B1(_3190_),
    .Y(_0535_),
    .A1(net1114),
    .A2(net1062));
 sg13g2_a21oi_1 _4336_ (.A1(_2911_),
    .A2(_0535_),
    .Y(_0536_),
    .B1(_0534_));
 sg13g2_nor2_1 _4337_ (.A(net1090),
    .B(_0507_),
    .Y(_0537_));
 sg13g2_o21ai_1 _4338_ (.B1(net1104),
    .Y(_0538_),
    .A1(_3107_),
    .A2(_0537_));
 sg13g2_a21oi_1 _4339_ (.A1(_0536_),
    .A2(_0538_),
    .Y(_0539_),
    .B1(net1060));
 sg13g2_nand3_1 _4340_ (.B(_3155_),
    .C(_0524_),
    .A(net1101),
    .Y(_0540_));
 sg13g2_o21ai_1 _4341_ (.B1(_0512_),
    .Y(_0541_),
    .A1(_0523_),
    .A2(_0540_));
 sg13g2_nor3_1 _4342_ (.A(net1002),
    .B(_0533_),
    .C(_0539_),
    .Y(_0542_));
 sg13g2_a22oi_1 _4343_ (.Y(_0543_),
    .B1(_0541_),
    .B2(_0542_),
    .A2(net1024),
    .A1(_0030_));
 sg13g2_nand3_1 _4344_ (.B(_0466_),
    .C(_0467_),
    .A(_0346_),
    .Y(_0544_));
 sg13g2_and3_1 _4345_ (.X(_0545_),
    .A(_0468_),
    .B(_0543_),
    .C(_0544_));
 sg13g2_o21ai_1 _4346_ (.B1(net1104),
    .Y(_0546_),
    .A1(_0522_),
    .A2(_0537_));
 sg13g2_a21oi_1 _4347_ (.A1(_0536_),
    .A2(_0546_),
    .Y(_0547_),
    .B1(net1060));
 sg13g2_o21ai_1 _4348_ (.B1(net1104),
    .Y(_0548_),
    .A1(_3105_),
    .A2(_3107_));
 sg13g2_o21ai_1 _4349_ (.B1(net1110),
    .Y(_0549_),
    .A1(net1062),
    .A2(_3144_));
 sg13g2_nand3_1 _4350_ (.B(_0502_),
    .C(_0549_),
    .A(net1100),
    .Y(_0550_));
 sg13g2_nor2b_1 _4351_ (.A(_0528_),
    .B_N(_0550_),
    .Y(_0551_));
 sg13g2_a21oi_2 _4352_ (.B1(net1098),
    .Y(_0552_),
    .A2(_0551_),
    .A1(_0548_));
 sg13g2_o21ai_1 _4353_ (.B1(net1107),
    .Y(_0553_),
    .A1(net1101),
    .A2(_3133_));
 sg13g2_a21oi_1 _4354_ (.A1(_3108_),
    .A2(_0553_),
    .Y(_0554_),
    .B1(_3131_));
 sg13g2_nor4_2 _4355_ (.A(net1002),
    .B(_0547_),
    .C(_0552_),
    .Y(_0555_),
    .D(_0554_));
 sg13g2_a21oi_2 _4356_ (.B1(_0555_),
    .Y(_0556_),
    .A2(net1024),
    .A1(_0029_));
 sg13g2_xnor2_1 _4357_ (.Y(_0557_),
    .A(_0463_),
    .B(_0464_));
 sg13g2_nor2_1 _4358_ (.A(_0556_),
    .B(_0557_),
    .Y(_0558_));
 sg13g2_nand2_1 _4359_ (.Y(_0559_),
    .A(net1109),
    .B(_3146_));
 sg13g2_o21ai_1 _4360_ (.B1(_0559_),
    .Y(_0560_),
    .A1(net1108),
    .A2(_3134_));
 sg13g2_nand2_1 _4361_ (.Y(_0561_),
    .A(net1102),
    .B(_0560_));
 sg13g2_a21oi_1 _4362_ (.A1(net1095),
    .A2(_2914_),
    .Y(_0562_),
    .B1(net1096));
 sg13g2_a21oi_1 _4363_ (.A1(_0497_),
    .A2(_0562_),
    .Y(_0563_),
    .B1(net1102));
 sg13g2_a21o_1 _4364_ (.A2(_0560_),
    .A1(net1101),
    .B1(_0563_),
    .X(_0564_));
 sg13g2_nand2_1 _4365_ (.Y(_0565_),
    .A(_3140_),
    .B(_0564_));
 sg13g2_nor3_2 _4366_ (.A(_0087_),
    .B(_0086_),
    .C(_3104_),
    .Y(_0566_));
 sg13g2_a21oi_1 _4367_ (.A1(_2936_),
    .A2(_0566_),
    .Y(_0567_),
    .B1(net1061));
 sg13g2_nor2_1 _4368_ (.A(net1104),
    .B(_3116_),
    .Y(_0568_));
 sg13g2_a21oi_1 _4369_ (.A1(net1103),
    .A2(_0566_),
    .Y(_0569_),
    .B1(_3100_));
 sg13g2_nor2b_1 _4370_ (.A(_0568_),
    .B_N(_0569_),
    .Y(_0570_));
 sg13g2_nor3_1 _4371_ (.A(net1002),
    .B(_0567_),
    .C(_0570_),
    .Y(_0571_));
 sg13g2_nand3_1 _4372_ (.B(_0565_),
    .C(_0571_),
    .A(_3136_),
    .Y(_0572_));
 sg13g2_o21ai_1 _4373_ (.B1(_0572_),
    .Y(_0573_),
    .A1(_2940_),
    .A2(net1027));
 sg13g2_inv_1 _4374_ (.Y(_0574_),
    .A(_0573_));
 sg13g2_xnor2_1 _4375_ (.Y(_0575_),
    .A(_0454_),
    .B(_0458_));
 sg13g2_nand2_1 _4376_ (.Y(_0576_),
    .A(_0574_),
    .B(_0575_));
 sg13g2_nand3_1 _4377_ (.B(_3103_),
    .C(_0521_),
    .A(net1112),
    .Y(_0577_));
 sg13g2_o21ai_1 _4378_ (.B1(net1109),
    .Y(_0578_),
    .A1(_3144_),
    .A2(_3153_));
 sg13g2_nand2_1 _4379_ (.Y(_0579_),
    .A(_0521_),
    .B(_0578_));
 sg13g2_nand3_1 _4380_ (.B(_0577_),
    .C(_0579_),
    .A(net1103),
    .Y(_0580_));
 sg13g2_a21oi_1 _4381_ (.A1(_0504_),
    .A2(_0580_),
    .Y(_0581_),
    .B1(_3100_));
 sg13g2_a21oi_1 _4382_ (.A1(_3108_),
    .A2(_0559_),
    .Y(_0582_),
    .B1(_2911_));
 sg13g2_o21ai_1 _4383_ (.B1(_3140_),
    .Y(_0583_),
    .A1(_0563_),
    .A2(_0582_));
 sg13g2_a21oi_1 _4384_ (.A1(_0577_),
    .A2(_0579_),
    .Y(_0584_),
    .B1(_0085_));
 sg13g2_a21oi_1 _4385_ (.A1(net1107),
    .A2(_3135_),
    .Y(_0585_),
    .B1(_3107_));
 sg13g2_nor2_1 _4386_ (.A(net1101),
    .B(_0585_),
    .Y(_0586_));
 sg13g2_a21oi_1 _4387_ (.A1(net1103),
    .A2(_0579_),
    .Y(_0587_),
    .B1(_0586_));
 sg13g2_nor2_1 _4388_ (.A(_3131_),
    .B(_0587_),
    .Y(_0588_));
 sg13g2_o21ai_1 _4389_ (.B1(_0583_),
    .Y(_0589_),
    .A1(net1061),
    .A2(_0584_));
 sg13g2_nor4_1 _4390_ (.A(net1002),
    .B(_0581_),
    .C(_0588_),
    .D(_0589_),
    .Y(_0590_));
 sg13g2_a21o_1 _4391_ (.A2(net1024),
    .A1(_0091_),
    .B1(_0590_),
    .X(_0591_));
 sg13g2_xnor2_1 _4392_ (.Y(_0592_),
    .A(_0452_),
    .B(_0453_));
 sg13g2_nor2_1 _4393_ (.A(_0591_),
    .B(_0592_),
    .Y(_0593_));
 sg13g2_a21o_1 _4394_ (.A2(_0520_),
    .A1(_3107_),
    .B1(_0525_),
    .X(_0594_));
 sg13g2_a21oi_1 _4395_ (.A1(net1103),
    .A2(_0594_),
    .Y(_0595_),
    .B1(_3142_));
 sg13g2_nor2_1 _4396_ (.A(_3100_),
    .B(_0595_),
    .Y(_0596_));
 sg13g2_a221oi_1 _4397_ (.B2(net1099),
    .C1(_0540_),
    .B1(_0564_),
    .A1(_3107_),
    .Y(_0597_),
    .A2(_0520_));
 sg13g2_a21oi_1 _4398_ (.A1(_3136_),
    .A2(_0565_),
    .Y(_0598_),
    .B1(_0597_));
 sg13g2_nor2_1 _4399_ (.A(_0085_),
    .B(_0594_),
    .Y(_0599_));
 sg13g2_nor2_1 _4400_ (.A(net1061),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_nor4_1 _4401_ (.A(net1002),
    .B(_0596_),
    .C(_0598_),
    .D(_0600_),
    .Y(_0601_));
 sg13g2_a21o_1 _4402_ (.A2(net1024),
    .A1(_0082_),
    .B1(_0601_),
    .X(_0602_));
 sg13g2_xor2_1 _4403_ (.B(_0451_),
    .A(_0450_),
    .X(_0603_));
 sg13g2_nand2b_1 _4404_ (.Y(_0604_),
    .B(_0603_),
    .A_N(_0602_));
 sg13g2_nor2_1 _4405_ (.A(_0096_),
    .B(net1020),
    .Y(_0605_));
 sg13g2_nor2_1 _4406_ (.A(_0436_),
    .B(_0449_),
    .Y(_0606_));
 sg13g2_xnor2_1 _4407_ (.Y(_0607_),
    .A(_0437_),
    .B(_0606_));
 sg13g2_nand2_1 _4408_ (.Y(_0608_),
    .A(_0605_),
    .B(_0607_));
 sg13g2_xor2_1 _4409_ (.B(_0603_),
    .A(_0602_),
    .X(_0609_));
 sg13g2_o21ai_1 _4410_ (.B1(_0604_),
    .Y(_0610_),
    .A1(_0608_),
    .A2(_0609_));
 sg13g2_xor2_1 _4411_ (.B(_0592_),
    .A(_0591_),
    .X(_0611_));
 sg13g2_a21oi_1 _4412_ (.A1(_0610_),
    .A2(_0611_),
    .Y(_0612_),
    .B1(_0593_));
 sg13g2_nor2_1 _4413_ (.A(_0574_),
    .B(_0575_),
    .Y(_0613_));
 sg13g2_xnor2_1 _4414_ (.Y(_0614_),
    .A(_0573_),
    .B(_0575_));
 sg13g2_o21ai_1 _4415_ (.B1(_0576_),
    .Y(_0615_),
    .A1(_0612_),
    .A2(_0613_));
 sg13g2_nand2_1 _4416_ (.Y(_0616_),
    .A(_0027_),
    .B(net1025));
 sg13g2_o21ai_1 _4417_ (.B1(_3137_),
    .Y(_0617_),
    .A1(_0087_),
    .A2(_0501_));
 sg13g2_nand4_1 _4418_ (.B(net1110),
    .C(_3104_),
    .A(net1105),
    .Y(_0618_),
    .D(_3153_));
 sg13g2_o21ai_1 _4419_ (.B1(_0529_),
    .Y(_0619_),
    .A1(net1093),
    .A2(_2912_));
 sg13g2_nor2_1 _4420_ (.A(net1062),
    .B(_0619_),
    .Y(_0620_));
 sg13g2_nor2_1 _4421_ (.A(net1098),
    .B(_0620_),
    .Y(_0621_));
 sg13g2_nand3b_1 _4422_ (.B(_0618_),
    .C(_0621_),
    .Y(_0622_),
    .A_N(_0528_));
 sg13g2_o21ai_1 _4423_ (.B1(_3130_),
    .Y(_0623_),
    .A1(_2911_),
    .A2(_0524_));
 sg13g2_o21ai_1 _4424_ (.B1(_0622_),
    .Y(_0624_),
    .A1(_0586_),
    .A2(_0623_));
 sg13g2_nor4_1 _4425_ (.A(net1060),
    .B(_0503_),
    .C(_0534_),
    .D(_0582_),
    .Y(_0625_));
 sg13g2_a21oi_1 _4426_ (.A1(_0617_),
    .A2(_0624_),
    .Y(_0626_),
    .B1(_0625_));
 sg13g2_o21ai_1 _4427_ (.B1(_0616_),
    .Y(_0627_),
    .A1(_3139_),
    .A2(_0626_));
 sg13g2_nor2b_1 _4428_ (.A(_0379_),
    .B_N(_0460_),
    .Y(_0628_));
 sg13g2_o21ai_1 _4429_ (.B1(_0457_),
    .Y(_0629_),
    .A1(_0454_),
    .A2(_0459_));
 sg13g2_xnor2_1 _4430_ (.Y(_0630_),
    .A(_0628_),
    .B(_0629_));
 sg13g2_nor2_1 _4431_ (.A(_0627_),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_xor2_1 _4432_ (.B(_0630_),
    .A(_0627_),
    .X(_0632_));
 sg13g2_a221oi_1 _4433_ (.B2(_0632_),
    .C1(_0631_),
    .B1(_0615_),
    .A1(_0556_),
    .Y(_0633_),
    .A2(_0557_));
 sg13g2_xnor2_1 _4434_ (.Y(_0634_),
    .A(_0556_),
    .B(_0557_));
 sg13g2_nor2_1 _4435_ (.A(_0558_),
    .B(_0633_),
    .Y(_0635_));
 sg13g2_a21oi_1 _4436_ (.A1(_0468_),
    .A2(_0544_),
    .Y(_0636_),
    .B1(_0543_));
 sg13g2_nor2_1 _4437_ (.A(_0545_),
    .B(_0636_),
    .Y(_0637_));
 sg13g2_a21o_1 _4438_ (.A2(_0637_),
    .A1(_0635_),
    .B1(_0545_),
    .X(_0638_));
 sg13g2_xor2_1 _4439_ (.B(_0518_),
    .A(_0516_),
    .X(_0639_));
 sg13g2_a21oi_2 _4440_ (.B1(_0519_),
    .Y(_0640_),
    .A2(_0639_),
    .A1(_0638_));
 sg13g2_xnor2_1 _4441_ (.Y(_0641_),
    .A(_3150_),
    .B(_0493_));
 sg13g2_o21ai_1 _4442_ (.B1(_0494_),
    .Y(_0642_),
    .A1(_0640_),
    .A2(_0641_));
 sg13g2_a21o_1 _4443_ (.A2(_3119_),
    .A1(net1113),
    .B1(net1062),
    .X(_0643_));
 sg13g2_a21oi_1 _4444_ (.A1(_2912_),
    .A2(_0643_),
    .Y(_0644_),
    .B1(_0619_));
 sg13g2_nor4_1 _4445_ (.A(_2911_),
    .B(net1111),
    .C(_3122_),
    .D(_3172_),
    .Y(_0645_));
 sg13g2_nor3_1 _4446_ (.A(_0528_),
    .B(_0644_),
    .C(_0645_),
    .Y(_0646_));
 sg13g2_a21oi_1 _4447_ (.A1(_0618_),
    .A2(_0646_),
    .Y(_0647_),
    .B1(net1097));
 sg13g2_a21oi_1 _4448_ (.A1(_0536_),
    .A2(_0561_),
    .Y(_0648_),
    .B1(net1060));
 sg13g2_nor4_2 _4449_ (.A(net1110),
    .B(_0088_),
    .C(_0087_),
    .Y(_0649_),
    .D(_3109_));
 sg13g2_a21oi_1 _4450_ (.A1(net1106),
    .A2(_0649_),
    .Y(_0650_),
    .B1(_3136_));
 sg13g2_nor4_1 _4451_ (.A(net1002),
    .B(_0647_),
    .C(_0648_),
    .D(_0650_),
    .Y(_0651_));
 sg13g2_a21o_1 _4452_ (.A2(net1024),
    .A1(_0033_),
    .B1(_0651_),
    .X(_0652_));
 sg13g2_o21ai_1 _4453_ (.B1(_0491_),
    .Y(_0653_),
    .A1(_0471_),
    .A2(_0489_));
 sg13g2_a21oi_1 _4454_ (.A1(_0472_),
    .A2(_0488_),
    .Y(_0654_),
    .B1(_0487_));
 sg13g2_a21oi_1 _4455_ (.A1(_0263_),
    .A2(_0483_),
    .Y(_0655_),
    .B1(_0482_));
 sg13g2_nand2_1 _4456_ (.Y(_0656_),
    .A(\i_display.frame[9] ),
    .B(net993));
 sg13g2_nand2_1 _4457_ (.Y(_0657_),
    .A(\i_display.frame[8] ),
    .B(_3267_));
 sg13g2_nand2_1 _4458_ (.Y(_0658_),
    .A(_0092_),
    .B(_3271_));
 sg13g2_nor2_1 _4459_ (.A(_0657_),
    .B(_0658_),
    .Y(_0659_));
 sg13g2_xor2_1 _4460_ (.B(_0658_),
    .A(_0657_),
    .X(_0660_));
 sg13g2_nor2b_1 _4461_ (.A(_0475_),
    .B_N(_0660_),
    .Y(_0661_));
 sg13g2_xnor2_1 _4462_ (.Y(_0662_),
    .A(_0475_),
    .B(_0660_));
 sg13g2_xnor2_1 _4463_ (.Y(_0663_),
    .A(_0480_),
    .B(_0662_));
 sg13g2_nor2_1 _4464_ (.A(_0656_),
    .B(_0663_),
    .Y(_0664_));
 sg13g2_xor2_1 _4465_ (.B(_0663_),
    .A(_0656_),
    .X(_0665_));
 sg13g2_a21oi_1 _4466_ (.A1(_0255_),
    .A2(_0476_),
    .Y(_0666_),
    .B1(_0485_));
 sg13g2_nand2b_1 _4467_ (.Y(_0667_),
    .B(_0665_),
    .A_N(_0666_));
 sg13g2_xnor2_1 _4468_ (.Y(_0668_),
    .A(_0665_),
    .B(_0666_));
 sg13g2_nor2b_1 _4469_ (.A(_0655_),
    .B_N(_0668_),
    .Y(_0669_));
 sg13g2_xor2_1 _4470_ (.B(_0668_),
    .A(_0655_),
    .X(_0670_));
 sg13g2_nor2_1 _4471_ (.A(_0654_),
    .B(_0670_),
    .Y(_0671_));
 sg13g2_xor2_1 _4472_ (.B(_0670_),
    .A(_0654_),
    .X(_0672_));
 sg13g2_xnor2_1 _4473_ (.Y(_0673_),
    .A(_0653_),
    .B(_0672_));
 sg13g2_nor2_1 _4474_ (.A(_0652_),
    .B(_0673_),
    .Y(_0674_));
 sg13g2_nand2_1 _4475_ (.Y(_0675_),
    .A(_0652_),
    .B(_0673_));
 sg13g2_xnor2_1 _4476_ (.Y(_0676_),
    .A(_0652_),
    .B(_0673_));
 sg13g2_xnor2_1 _4477_ (.Y(_0677_),
    .A(_0642_),
    .B(_0676_));
 sg13g2_nor2_1 _4478_ (.A(_2920_),
    .B(net1132),
    .Y(_0678_));
 sg13g2_nand2_1 _4479_ (.Y(_0679_),
    .A(\i_display.i_vga.low_count[9] ),
    .B(net1064));
 sg13g2_nand2_1 _4480_ (.Y(_0680_),
    .A(net1027),
    .B(_0679_));
 sg13g2_o21ai_1 _4481_ (.B1(_0680_),
    .Y(_0681_),
    .A1(net1026),
    .A2(_0678_));
 sg13g2_xnor2_1 _4482_ (.Y(_0682_),
    .A(_0677_),
    .B(_0681_));
 sg13g2_xnor2_1 _4483_ (.Y(_0683_),
    .A(_0640_),
    .B(_0641_));
 sg13g2_nand2b_2 _4484_ (.Y(_0684_),
    .B(\i_display.i_vga.timing_ver.counter[8] ),
    .A_N(net1132));
 sg13g2_and2_1 _4485_ (.A(\i_display.i_vga.low_count[8] ),
    .B(net1064),
    .X(_0685_));
 sg13g2_nor2_1 _4486_ (.A(net1019),
    .B(_0685_),
    .Y(_0686_));
 sg13g2_a21oi_2 _4487_ (.B1(_0686_),
    .Y(_0687_),
    .A2(_0684_),
    .A1(net1019));
 sg13g2_nor2_1 _4488_ (.A(_0683_),
    .B(_0687_),
    .Y(_0688_));
 sg13g2_nand2_1 _4489_ (.Y(_0689_),
    .A(_0683_),
    .B(_0687_));
 sg13g2_xor2_1 _4490_ (.B(_0639_),
    .A(_0638_),
    .X(_0690_));
 sg13g2_nand2b_1 _4491_ (.Y(_0691_),
    .B(\i_display.i_vga.timing_ver.counter[7] ),
    .A_N(net1132));
 sg13g2_a21oi_1 _4492_ (.A1(net1142),
    .A2(net1063),
    .Y(_0692_),
    .B1(net1019));
 sg13g2_a21o_1 _4493_ (.A2(_0691_),
    .A1(net1019),
    .B1(_0692_),
    .X(_0693_));
 sg13g2_or2_1 _4494_ (.X(_0694_),
    .B(_0693_),
    .A(_0690_));
 sg13g2_nand2_1 _4495_ (.Y(_0695_),
    .A(_0690_),
    .B(_0693_));
 sg13g2_xnor2_1 _4496_ (.Y(_0696_),
    .A(_0635_),
    .B(_0637_));
 sg13g2_nand2b_2 _4497_ (.Y(_0697_),
    .B(\i_display.i_vga.timing_ver.counter[6] ),
    .A_N(net1131));
 sg13g2_a21oi_1 _4498_ (.A1(\i_display.i_vga.low_count[6] ),
    .A2(net1064),
    .Y(_0698_),
    .B1(net1020));
 sg13g2_a21oi_1 _4499_ (.A1(net1020),
    .A2(_0697_),
    .Y(_0699_),
    .B1(_0698_));
 sg13g2_nor2_1 _4500_ (.A(_0696_),
    .B(_0699_),
    .Y(_0700_));
 sg13g2_nand2_1 _4501_ (.Y(_0701_),
    .A(_0696_),
    .B(_0699_));
 sg13g2_xnor2_1 _4502_ (.Y(_0702_),
    .A(_0615_),
    .B(_0632_));
 sg13g2_nand2b_2 _4503_ (.Y(_0703_),
    .B(\i_display.i_vga.timing_ver.counter[4] ),
    .A_N(net1131));
 sg13g2_nand2_2 _4504_ (.Y(_0704_),
    .A(\i_display.i_vga.low_count[4] ),
    .B(net1063));
 sg13g2_and2_1 _4505_ (.A(net1026),
    .B(_0704_),
    .X(_0705_));
 sg13g2_a21oi_2 _4506_ (.B1(_0705_),
    .Y(_0706_),
    .A2(_0703_),
    .A1(net1019));
 sg13g2_nand2_1 _4507_ (.Y(_0707_),
    .A(_0702_),
    .B(_0706_));
 sg13g2_xnor2_1 _4508_ (.Y(_0708_),
    .A(_0612_),
    .B(_0614_));
 sg13g2_nor2b_2 _4509_ (.A(net1131),
    .B_N(\i_display.i_vga.timing_ver.counter[3] ),
    .Y(_0709_));
 sg13g2_nand2_2 _4510_ (.Y(_0710_),
    .A(\i_display.i_vga.low_count[3] ),
    .B(net1063));
 sg13g2_inv_2 _4511_ (.Y(_0711_),
    .A(_0710_));
 sg13g2_nor2_1 _4512_ (.A(net1019),
    .B(_0710_),
    .Y(_0712_));
 sg13g2_a21oi_1 _4513_ (.A1(net1019),
    .A2(_0709_),
    .Y(_0713_),
    .B1(_0712_));
 sg13g2_nor2_1 _4514_ (.A(_0708_),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_xor2_1 _4515_ (.B(_0611_),
    .A(_0610_),
    .X(_0715_));
 sg13g2_nand2_2 _4516_ (.Y(_0716_),
    .A(\i_display.i_vga.low_count[2] ),
    .B(net1063));
 sg13g2_nand2b_2 _4517_ (.Y(_0717_),
    .B(\i_display.i_vga.timing_ver.counter[2] ),
    .A_N(net1131));
 sg13g2_mux2_1 _4518_ (.A0(_0716_),
    .A1(_0717_),
    .S(net1019),
    .X(_0718_));
 sg13g2_xor2_1 _4519_ (.B(_0609_),
    .A(_0608_),
    .X(_0719_));
 sg13g2_nand2_2 _4520_ (.Y(_0720_),
    .A(net1148),
    .B(net1065));
 sg13g2_nor2_2 _4521_ (.A(_2922_),
    .B(net1131),
    .Y(_0721_));
 sg13g2_nand2b_1 _4522_ (.Y(_0722_),
    .B(net1130),
    .A_N(net1131));
 sg13g2_nor2_1 _4523_ (.A(net1026),
    .B(_0721_),
    .Y(_0723_));
 sg13g2_a21oi_2 _4524_ (.B1(_0723_),
    .Y(_0724_),
    .A2(_0720_),
    .A1(net1026));
 sg13g2_xnor2_1 _4525_ (.Y(_0725_),
    .A(_0719_),
    .B(_0724_));
 sg13g2_xor2_1 _4526_ (.B(_0607_),
    .A(_0605_),
    .X(_0726_));
 sg13g2_nor2b_2 _4527_ (.A(net1132),
    .B_N(\i_display.i_vga.timing_ver.counter[0] ),
    .Y(_0727_));
 sg13g2_nand2b_1 _4528_ (.Y(_0728_),
    .B(\i_display.i_vga.timing_ver.counter[0] ),
    .A_N(net1131));
 sg13g2_nor2_1 _4529_ (.A(net1026),
    .B(_0728_),
    .Y(_0729_));
 sg13g2_and2_2 _4530_ (.A(net1153),
    .B(net1063),
    .X(_0730_));
 sg13g2_a21oi_1 _4531_ (.A1(net1026),
    .A2(_0730_),
    .Y(_0731_),
    .B1(_0729_));
 sg13g2_xnor2_1 _4532_ (.Y(_0732_),
    .A(_0726_),
    .B(_0731_));
 sg13g2_o21ai_1 _4533_ (.B1(_0725_),
    .Y(_0733_),
    .A1(_0715_),
    .A2(_0718_));
 sg13g2_nor2_1 _4534_ (.A(_0714_),
    .B(_0733_),
    .Y(_0734_));
 sg13g2_o21ai_1 _4535_ (.B1(_0734_),
    .Y(_0735_),
    .A1(_0702_),
    .A2(_0706_));
 sg13g2_a221oi_1 _4536_ (.B2(_0718_),
    .C1(_0732_),
    .B1(_0715_),
    .A1(_0708_),
    .Y(_0736_),
    .A2(_0713_));
 sg13g2_nand2_1 _4537_ (.Y(_0737_),
    .A(_0707_),
    .B(_0736_));
 sg13g2_a21oi_1 _4538_ (.A1(_0615_),
    .A2(_0632_),
    .Y(_0738_),
    .B1(_0631_));
 sg13g2_nand2_1 _4539_ (.Y(_0739_),
    .A(\i_display.i_vga.low_count[5] ),
    .B(net1063));
 sg13g2_nor2b_2 _4540_ (.A(net1131),
    .B_N(\i_display.i_vga.timing_ver.counter[5] ),
    .Y(_0740_));
 sg13g2_nor2_1 _4541_ (.A(net1026),
    .B(_0740_),
    .Y(_0741_));
 sg13g2_a21oi_1 _4542_ (.A1(net1026),
    .A2(_0739_),
    .Y(_0742_),
    .B1(_0741_));
 sg13g2_xnor2_1 _4543_ (.Y(_0743_),
    .A(_0634_),
    .B(_0742_));
 sg13g2_xnor2_1 _4544_ (.Y(_0744_),
    .A(_0738_),
    .B(_0743_));
 sg13g2_nor4_1 _4545_ (.A(_0700_),
    .B(_0735_),
    .C(_0737_),
    .D(_0744_),
    .Y(_0745_));
 sg13g2_and4_1 _4546_ (.A(_0694_),
    .B(_0695_),
    .C(_0701_),
    .D(_0745_),
    .X(_0746_));
 sg13g2_nand3b_1 _4547_ (.B(_0689_),
    .C(_0746_),
    .Y(_0747_),
    .A_N(_0688_));
 sg13g2_a21oi_1 _4548_ (.A1(_0642_),
    .A2(_0675_),
    .Y(_0748_),
    .B1(_0674_));
 sg13g2_a21oi_1 _4549_ (.A1(_0653_),
    .A2(_0672_),
    .Y(_0749_),
    .B1(_0671_));
 sg13g2_xnor2_1 _4550_ (.Y(_0750_),
    .A(_0664_),
    .B(_0669_));
 sg13g2_nand2_1 _4551_ (.Y(_0751_),
    .A(_0667_),
    .B(_0750_));
 sg13g2_a21oi_1 _4552_ (.A1(_0480_),
    .A2(_0662_),
    .Y(_0752_),
    .B1(_0661_));
 sg13g2_nor2_1 _4553_ (.A(net1100),
    .B(_0085_),
    .Y(_0753_));
 sg13g2_nand4_1 _4554_ (.B(_2943_),
    .C(_0649_),
    .A(_0071_),
    .Y(_0754_),
    .D(_0753_));
 sg13g2_nand2_1 _4555_ (.Y(_0755_),
    .A(\i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[9] ),
    .B(net1024));
 sg13g2_o21ai_1 _4556_ (.B1(_0755_),
    .Y(_0756_),
    .A1(net1025),
    .A2(_0754_));
 sg13g2_xor2_1 _4557_ (.B(_0756_),
    .A(_0659_),
    .X(_0757_));
 sg13g2_nand2_1 _4558_ (.Y(_0758_),
    .A(\i_display.frame[9] ),
    .B(_3267_));
 sg13g2_nand2_1 _4559_ (.Y(_0759_),
    .A(_0095_),
    .B(_3271_));
 sg13g2_xnor2_1 _4560_ (.Y(_0760_),
    .A(_0758_),
    .B(_0759_));
 sg13g2_xnor2_1 _4561_ (.Y(_0761_),
    .A(_0757_),
    .B(_0760_));
 sg13g2_xnor2_1 _4562_ (.Y(_0762_),
    .A(_0752_),
    .B(_0761_));
 sg13g2_xnor2_1 _4563_ (.Y(_0763_),
    .A(_0751_),
    .B(_0762_));
 sg13g2_xor2_1 _4564_ (.B(_0763_),
    .A(_0749_),
    .X(_0764_));
 sg13g2_xnor2_1 _4565_ (.Y(_0765_),
    .A(_0748_),
    .B(_0764_));
 sg13g2_nor3_2 _4566_ (.A(_0682_),
    .B(_0747_),
    .C(_0765_),
    .Y(_0766_));
 sg13g2_nor4_2 _4567_ (.A(net1027),
    .B(_0682_),
    .C(_0747_),
    .Y(_0767_),
    .D(_0765_));
 sg13g2_or4_2 _4568_ (.A(net1027),
    .B(_0682_),
    .C(_0747_),
    .D(_0765_),
    .X(_0768_));
 sg13g2_nor2_2 _4569_ (.A(_3093_),
    .B(_0767_),
    .Y(_0769_));
 sg13g2_nand3b_1 _4570_ (.B(net1003),
    .C(_0768_),
    .Y(_0770_),
    .A_N(_0086_));
 sg13g2_nand2_1 _4571_ (.Y(_0771_),
    .A(net1110),
    .B(_3117_));
 sg13g2_nand2_1 _4572_ (.Y(_0772_),
    .A(_2912_),
    .B(_3118_));
 sg13g2_nand3_1 _4573_ (.B(_0771_),
    .C(_0772_),
    .A(net1004),
    .Y(_0773_));
 sg13g2_xnor2_1 _4574_ (.Y(_0774_),
    .A(net8),
    .B(\crotchet[6] ));
 sg13g2_xor2_1 _4575_ (.B(\crotchet[6] ),
    .A(net8),
    .X(_0775_));
 sg13g2_xnor2_1 _4576_ (.Y(_0776_),
    .A(\crotchet[5] ),
    .B(net7));
 sg13g2_xor2_1 _4577_ (.B(net7),
    .A(\crotchet[5] ),
    .X(_0777_));
 sg13g2_xnor2_1 _4578_ (.Y(_0778_),
    .A(net5),
    .B(\crotchet[3] ));
 sg13g2_xor2_1 _4579_ (.B(\crotchet[3] ),
    .A(net5),
    .X(_0779_));
 sg13g2_nor2_1 _4580_ (.A(_3097_),
    .B(_0779_),
    .Y(_0780_));
 sg13g2_xnor2_1 _4581_ (.Y(_0781_),
    .A(net4),
    .B(\crotchet[2] ));
 sg13g2_xor2_1 _4582_ (.B(\crotchet[2] ),
    .A(net4),
    .X(_0782_));
 sg13g2_nand3_1 _4583_ (.B(_0779_),
    .C(_0782_),
    .A(_3097_),
    .Y(_0783_));
 sg13g2_nand2b_1 _4584_ (.Y(_0784_),
    .B(_0783_),
    .A_N(_0780_));
 sg13g2_a21oi_1 _4585_ (.A1(net1058),
    .A2(_0784_),
    .Y(_0785_),
    .B1(_0774_));
 sg13g2_nor2_1 _4586_ (.A(net1057),
    .B(_0781_),
    .Y(_0786_));
 sg13g2_nand2_1 _4587_ (.Y(_0787_),
    .A(_0778_),
    .B(_0782_));
 sg13g2_nand2_1 _4588_ (.Y(_0788_),
    .A(net1057),
    .B(_0781_));
 sg13g2_nand3_1 _4589_ (.B(_0776_),
    .C(_0788_),
    .A(_3096_),
    .Y(_0789_));
 sg13g2_nand2_1 _4590_ (.Y(_0790_),
    .A(_3097_),
    .B(_0776_));
 sg13g2_nand2_1 _4591_ (.Y(_0791_),
    .A(_3096_),
    .B(net1059));
 sg13g2_nand3_1 _4592_ (.B(_0790_),
    .C(_0791_),
    .A(_0774_),
    .Y(_0792_));
 sg13g2_xor2_1 _4593_ (.B(\crotchet[1] ),
    .A(net3),
    .X(_0793_));
 sg13g2_nor2_1 _4594_ (.A(\crotchet[0] ),
    .B(_0793_),
    .Y(_0794_));
 sg13g2_nor3_1 _4595_ (.A(\crotchet[0] ),
    .B(_0782_),
    .C(_0793_),
    .Y(_0795_));
 sg13g2_nand3_1 _4596_ (.B(_0778_),
    .C(_0795_),
    .A(_0776_),
    .Y(_0796_));
 sg13g2_nand2b_1 _4597_ (.Y(_0797_),
    .B(_0796_),
    .A_N(_0792_));
 sg13g2_o21ai_1 _4598_ (.B1(_0785_),
    .Y(_0798_),
    .A1(_0786_),
    .A2(_0789_));
 sg13g2_a21oi_1 _4599_ (.A1(_0785_),
    .A2(_0790_),
    .Y(_0799_),
    .B1(_0788_));
 sg13g2_a21oi_1 _4600_ (.A1(_0797_),
    .A2(_0798_),
    .Y(_0800_),
    .B1(_0799_));
 sg13g2_o21ai_1 _4601_ (.B1(_0773_),
    .Y(_0801_),
    .A1(net1004),
    .A2(_0800_));
 sg13g2_o21ai_1 _4602_ (.B1(_0801_),
    .Y(_0802_),
    .A1(_3093_),
    .A2(_0767_));
 sg13g2_and2_1 _4603_ (.A(_0770_),
    .B(_0802_),
    .X(_0803_));
 sg13g2_nand2_2 _4604_ (.Y(_0804_),
    .A(_0770_),
    .B(_0802_));
 sg13g2_nand3_1 _4605_ (.B(net1003),
    .C(_0768_),
    .A(_2943_),
    .Y(_0805_));
 sg13g2_nand3_1 _4606_ (.B(net1111),
    .C(_3117_),
    .A(net1106),
    .Y(_0806_));
 sg13g2_nor2_1 _4607_ (.A(_0084_),
    .B(_0806_),
    .Y(_0807_));
 sg13g2_xnor2_1 _4608_ (.Y(_0808_),
    .A(_2943_),
    .B(_0807_));
 sg13g2_a21oi_1 _4609_ (.A1(net1058),
    .A2(_0783_),
    .Y(_0809_),
    .B1(_0774_));
 sg13g2_nand2_1 _4610_ (.Y(_0810_),
    .A(_0780_),
    .B(_0781_));
 sg13g2_nand2_1 _4611_ (.Y(_0811_),
    .A(_0809_),
    .B(_0810_));
 sg13g2_nand2_1 _4612_ (.Y(_0812_),
    .A(_0780_),
    .B(_0795_));
 sg13g2_nor3_1 _4613_ (.A(_0775_),
    .B(net1058),
    .C(_0812_),
    .Y(_0813_));
 sg13g2_nor2_1 _4614_ (.A(net1003),
    .B(_0813_),
    .Y(_0814_));
 sg13g2_a22oi_1 _4615_ (.Y(_0815_),
    .B1(_0811_),
    .B2(_0814_),
    .A2(_0808_),
    .A1(net1004));
 sg13g2_o21ai_1 _4616_ (.B1(_0815_),
    .Y(_0816_),
    .A1(_3089_),
    .A2(_0767_));
 sg13g2_and2_2 _4617_ (.A(_0805_),
    .B(_0816_),
    .X(_0817_));
 sg13g2_nand3b_1 _4618_ (.B(net1003),
    .C(_0768_),
    .Y(_0818_),
    .A_N(_0084_));
 sg13g2_a21o_1 _4619_ (.A2(_0806_),
    .A1(_0084_),
    .B1(_3093_),
    .X(_0819_));
 sg13g2_nor2_1 _4620_ (.A(net1057),
    .B(_0795_),
    .Y(_0820_));
 sg13g2_o21ai_1 _4621_ (.B1(_0809_),
    .Y(_0821_),
    .A1(_3097_),
    .A2(_0781_));
 sg13g2_o21ai_1 _4622_ (.B1(_0821_),
    .Y(_0822_),
    .A1(_0792_),
    .A2(_0820_));
 sg13g2_nand2_1 _4623_ (.Y(_0823_),
    .A(_3097_),
    .B(_0778_));
 sg13g2_nand3_1 _4624_ (.B(_0822_),
    .C(_0823_),
    .A(_3089_),
    .Y(_0824_));
 sg13g2_o21ai_1 _4625_ (.B1(_0824_),
    .Y(_0825_),
    .A1(_0807_),
    .A2(_0819_));
 sg13g2_o21ai_1 _4626_ (.B1(_0825_),
    .Y(_0826_),
    .A1(net1005),
    .A2(_0767_));
 sg13g2_and2_1 _4627_ (.A(_0818_),
    .B(_0826_),
    .X(_0827_));
 sg13g2_a21oi_1 _4628_ (.A1(_0818_),
    .A2(_0826_),
    .Y(_0828_),
    .B1(net1160));
 sg13g2_a21oi_2 _4629_ (.B1(net1160),
    .Y(_0829_),
    .A2(_0816_),
    .A1(_0805_));
 sg13g2_nand2b_2 _4630_ (.Y(_0830_),
    .B(net1172),
    .A_N(_0817_));
 sg13g2_nor2b_2 _4631_ (.A(_0817_),
    .B_N(net896),
    .Y(_0831_));
 sg13g2_nand2b_2 _4632_ (.Y(_0832_),
    .B(net896),
    .A_N(_0817_));
 sg13g2_nand3_1 _4633_ (.B(net1003),
    .C(_0768_),
    .A(_2936_),
    .Y(_0833_));
 sg13g2_xnor2_1 _4634_ (.Y(_0834_),
    .A(_0085_),
    .B(_0771_));
 sg13g2_a21oi_1 _4635_ (.A1(_3097_),
    .A2(net1057),
    .Y(_0835_),
    .B1(net1058));
 sg13g2_a22oi_1 _4636_ (.Y(_0836_),
    .B1(_0812_),
    .B2(_0835_),
    .A2(_0787_),
    .A1(net1058));
 sg13g2_o21ai_1 _4637_ (.B1(_0776_),
    .Y(_0837_),
    .A1(_0787_),
    .A2(_0794_));
 sg13g2_and2_1 _4638_ (.A(_3096_),
    .B(_0837_),
    .X(_0838_));
 sg13g2_o21ai_1 _4639_ (.B1(_0774_),
    .Y(_0839_),
    .A1(_0836_),
    .A2(_0838_));
 sg13g2_nand3_1 _4640_ (.B(_0782_),
    .C(_0823_),
    .A(_0776_),
    .Y(_0840_));
 sg13g2_nor2_1 _4641_ (.A(_0788_),
    .B(_0791_),
    .Y(_0841_));
 sg13g2_nor2_1 _4642_ (.A(_0774_),
    .B(_0841_),
    .Y(_0842_));
 sg13g2_a21oi_1 _4643_ (.A1(_0840_),
    .A2(_0842_),
    .Y(_0843_),
    .B1(net1004));
 sg13g2_a22oi_1 _4644_ (.Y(_0844_),
    .B1(_0839_),
    .B2(_0843_),
    .A2(_0834_),
    .A1(net1004));
 sg13g2_o21ai_1 _4645_ (.B1(_0844_),
    .Y(_0845_),
    .A1(net1005),
    .A2(_0767_));
 sg13g2_and2_1 _4646_ (.A(_0833_),
    .B(_0845_),
    .X(_0846_));
 sg13g2_nand2_2 _4647_ (.Y(_0847_),
    .A(_0833_),
    .B(_0845_));
 sg13g2_a21oi_1 _4648_ (.A1(_0833_),
    .A2(_0845_),
    .Y(_0848_),
    .B1(net1162));
 sg13g2_nand2_1 _4649_ (.Y(_0849_),
    .A(net1172),
    .B(_0847_));
 sg13g2_nor3_1 _4650_ (.A(_0804_),
    .B(_0832_),
    .C(net893),
    .Y(_0850_));
 sg13g2_nand3_1 _4651_ (.B(net1003),
    .C(_0768_),
    .A(_2937_),
    .Y(_0851_));
 sg13g2_nand3_1 _4652_ (.B(_3118_),
    .C(_3121_),
    .A(net1003),
    .Y(_0852_));
 sg13g2_nor2_1 _4653_ (.A(_0778_),
    .B(_0793_),
    .Y(_0853_));
 sg13g2_a21oi_1 _4654_ (.A1(_0785_),
    .A2(_0810_),
    .Y(_0854_),
    .B1(_3094_));
 sg13g2_o21ai_1 _4655_ (.B1(_0854_),
    .Y(_0855_),
    .A1(_0797_),
    .A2(_0853_));
 sg13g2_nand2_1 _4656_ (.Y(_0856_),
    .A(_0852_),
    .B(_0855_));
 sg13g2_inv_1 _4657_ (.Y(_0857_),
    .A(_0856_));
 sg13g2_o21ai_1 _4658_ (.B1(_0856_),
    .Y(_0858_),
    .A1(_3089_),
    .A2(_0767_));
 sg13g2_and2_1 _4659_ (.A(_0851_),
    .B(_0858_),
    .X(_0859_));
 sg13g2_nand2_1 _4660_ (.Y(_0860_),
    .A(_0851_),
    .B(_0858_));
 sg13g2_nand2_2 _4661_ (.Y(_0861_),
    .A(net1172),
    .B(net891));
 sg13g2_or2_1 _4662_ (.X(_0862_),
    .B(net894),
    .A(net898));
 sg13g2_nor3_2 _4663_ (.A(net896),
    .B(_0829_),
    .C(net893),
    .Y(_0863_));
 sg13g2_a21oi_1 _4664_ (.A1(_0770_),
    .A2(_0802_),
    .Y(_0864_),
    .B1(net1162));
 sg13g2_nand2_2 _4665_ (.Y(_0865_),
    .A(net1173),
    .B(_0804_));
 sg13g2_a21oi_1 _4666_ (.A1(net1172),
    .A2(net890),
    .Y(_0866_),
    .B1(net889));
 sg13g2_a21o_1 _4667_ (.A2(_0866_),
    .A1(_0863_),
    .B1(_0850_),
    .X(_0009_));
 sg13g2_nand3b_1 _4668_ (.B(net1003),
    .C(_0768_),
    .Y(_0867_),
    .A_N(_0088_));
 sg13g2_a21oi_1 _4669_ (.A1(_0047_),
    .A2(net1057),
    .Y(_0868_),
    .B1(_0797_));
 sg13g2_nand2b_1 _4670_ (.Y(_0869_),
    .B(_0854_),
    .A_N(_0868_));
 sg13g2_o21ai_1 _4671_ (.B1(_0869_),
    .Y(_0870_),
    .A1(net1115),
    .A2(net1005));
 sg13g2_o21ai_1 _4672_ (.B1(_0870_),
    .Y(_0871_),
    .A1(_3093_),
    .A2(_0767_));
 sg13g2_and2_2 _4673_ (.A(_0867_),
    .B(_0871_),
    .X(_0872_));
 sg13g2_a21oi_1 _4674_ (.A1(_0867_),
    .A2(_0871_),
    .Y(_0873_),
    .B1(net1162));
 sg13g2_nand2_1 _4675_ (.Y(_0874_),
    .A(net895),
    .B(net887));
 sg13g2_nand2_2 _4676_ (.Y(_0875_),
    .A(_0804_),
    .B(net887));
 sg13g2_nor2_1 _4677_ (.A(net899),
    .B(_0861_),
    .Y(_0876_));
 sg13g2_nand2_2 _4678_ (.Y(_0877_),
    .A(net890),
    .B(net888));
 sg13g2_nor2_1 _4679_ (.A(_0803_),
    .B(_0877_),
    .Y(_0878_));
 sg13g2_o21ai_1 _4680_ (.B1(net893),
    .Y(_0879_),
    .A1(net899),
    .A2(_0877_));
 sg13g2_and2_1 _4681_ (.A(_0817_),
    .B(net896),
    .X(_0880_));
 sg13g2_nand2_2 _4682_ (.Y(_0881_),
    .A(_0817_),
    .B(net898));
 sg13g2_a21oi_1 _4683_ (.A1(_0874_),
    .A2(_0879_),
    .Y(_0882_),
    .B1(_0881_));
 sg13g2_nand3_1 _4684_ (.B(net893),
    .C(net892),
    .A(_0804_),
    .Y(_0883_));
 sg13g2_nand3_1 _4685_ (.B(net895),
    .C(net887),
    .A(net899),
    .Y(_0884_));
 sg13g2_a21oi_1 _4686_ (.A1(_0883_),
    .A2(_0884_),
    .Y(_0885_),
    .B1(_0832_));
 sg13g2_or2_2 _4687_ (.X(_0886_),
    .B(net887),
    .A(net889));
 sg13g2_nor3_1 _4688_ (.A(_0829_),
    .B(_0862_),
    .C(_0886_),
    .Y(_0887_));
 sg13g2_or3_1 _4689_ (.A(_0882_),
    .B(_0885_),
    .C(_0887_),
    .X(_0010_));
 sg13g2_and2_1 _4690_ (.A(net896),
    .B(_0847_),
    .X(_0888_));
 sg13g2_and4_1 _4691_ (.A(_0831_),
    .B(_0847_),
    .C(_0861_),
    .D(_0875_),
    .X(_0889_));
 sg13g2_a21o_1 _4692_ (.A2(net887),
    .A1(_0850_),
    .B1(_0889_),
    .X(_0890_));
 sg13g2_nand3_1 _4693_ (.B(net895),
    .C(net890),
    .A(net1172),
    .Y(_0891_));
 sg13g2_a21oi_1 _4694_ (.A1(_0879_),
    .A2(_0891_),
    .Y(_0892_),
    .B1(_0881_));
 sg13g2_nand2_2 _4695_ (.Y(_0893_),
    .A(net892),
    .B(_0872_));
 sg13g2_a21oi_2 _4696_ (.B1(net1162),
    .Y(_0894_),
    .A2(_0872_),
    .A1(net892));
 sg13g2_a21oi_2 _4697_ (.B1(net889),
    .Y(_0895_),
    .A2(_0894_),
    .A1(_0877_));
 sg13g2_and2_1 _4698_ (.A(net892),
    .B(net887),
    .X(_0896_));
 sg13g2_nand2_2 _4699_ (.Y(_0897_),
    .A(net892),
    .B(net887));
 sg13g2_o21ai_1 _4700_ (.B1(_0863_),
    .Y(_0898_),
    .A1(net884),
    .A2(_0896_));
 sg13g2_and2_1 _4701_ (.A(_0827_),
    .B(_0829_),
    .X(_0899_));
 sg13g2_nand3_1 _4702_ (.B(_0861_),
    .C(_0899_),
    .A(_0846_),
    .Y(_0900_));
 sg13g2_o21ai_1 _4703_ (.B1(_0900_),
    .Y(_0901_),
    .A1(_0895_),
    .A2(_0898_));
 sg13g2_or3_1 _4704_ (.A(_0890_),
    .B(_0892_),
    .C(_0901_),
    .X(_0011_));
 sg13g2_nand3_1 _4705_ (.B(_0875_),
    .C(_0886_),
    .A(net885),
    .Y(_0902_));
 sg13g2_nand2_1 _4706_ (.Y(_0903_),
    .A(_0847_),
    .B(net890));
 sg13g2_o21ai_1 _4707_ (.B1(_0880_),
    .Y(_0904_),
    .A1(_0875_),
    .A2(_0903_));
 sg13g2_nand2b_1 _4708_ (.Y(_0905_),
    .B(_0902_),
    .A_N(_0904_));
 sg13g2_o21ai_1 _4709_ (.B1(net892),
    .Y(_0906_),
    .A1(net889),
    .A2(net888));
 sg13g2_nand3_1 _4710_ (.B(_0863_),
    .C(_0886_),
    .A(net892),
    .Y(_0907_));
 sg13g2_nand3b_1 _4711_ (.B(_0905_),
    .C(_0907_),
    .Y(_0012_),
    .A_N(_0890_));
 sg13g2_nor3_1 _4712_ (.A(_0832_),
    .B(net893),
    .C(_0886_),
    .Y(_0908_));
 sg13g2_nand3_1 _4713_ (.B(net899),
    .C(net890),
    .A(net1172),
    .Y(_0909_));
 sg13g2_a221oi_1 _4714_ (.B2(_0897_),
    .C1(_0832_),
    .B1(net889),
    .A1(_0833_),
    .Y(_0910_),
    .A2(_0845_));
 sg13g2_a21oi_1 _4715_ (.A1(_0909_),
    .A2(_0910_),
    .Y(_0911_),
    .B1(_0908_));
 sg13g2_a21o_1 _4716_ (.A2(_0894_),
    .A1(_0877_),
    .B1(net884),
    .X(_0912_));
 sg13g2_and2_2 _4717_ (.A(net896),
    .B(net895),
    .X(_0913_));
 sg13g2_nand2_1 _4718_ (.Y(_0914_),
    .A(net897),
    .B(net895));
 sg13g2_and3_1 _4719_ (.X(_0915_),
    .A(net886),
    .B(_0909_),
    .C(_0913_));
 sg13g2_nand3_1 _4720_ (.B(net890),
    .C(_0872_),
    .A(net1172),
    .Y(_0916_));
 sg13g2_nand4_1 _4721_ (.B(net899),
    .C(net890),
    .A(net1172),
    .Y(_0917_),
    .D(_0872_));
 sg13g2_o21ai_1 _4722_ (.B1(_0917_),
    .Y(_0918_),
    .A1(net884),
    .A2(_0897_));
 sg13g2_a22oi_1 _4723_ (.Y(_0919_),
    .B1(_0918_),
    .B2(_0863_),
    .A2(_0915_),
    .A1(_0912_));
 sg13g2_nand2_1 _4724_ (.Y(_0013_),
    .A(_0911_),
    .B(_0919_));
 sg13g2_nand3_1 _4725_ (.B(net884),
    .C(_0877_),
    .A(_0863_),
    .Y(_0920_));
 sg13g2_and2_1 _4726_ (.A(_0900_),
    .B(_0920_),
    .X(_0921_));
 sg13g2_o21ai_1 _4727_ (.B1(net893),
    .Y(_0922_),
    .A1(net884),
    .A2(_0893_));
 sg13g2_a21oi_1 _4728_ (.A1(net885),
    .A2(_0886_),
    .Y(_0923_),
    .B1(_0832_));
 sg13g2_nand2_1 _4729_ (.Y(_0924_),
    .A(_0922_),
    .B(_0923_));
 sg13g2_nand2_1 _4730_ (.Y(_0925_),
    .A(net889),
    .B(_0893_));
 sg13g2_nand3_1 _4731_ (.B(_0913_),
    .C(_0925_),
    .A(_0817_),
    .Y(_0926_));
 sg13g2_nand3_1 _4732_ (.B(_0924_),
    .C(_0926_),
    .A(_0921_),
    .Y(_0014_));
 sg13g2_nand3_1 _4733_ (.B(_0911_),
    .C(_0920_),
    .A(_0904_),
    .Y(_0015_));
 sg13g2_nor4_1 _4734_ (.A(_0832_),
    .B(net895),
    .C(net884),
    .D(_0897_),
    .Y(_0927_));
 sg13g2_nor2_1 _4735_ (.A(_0908_),
    .B(_0927_),
    .Y(_0928_));
 sg13g2_nand2_1 _4736_ (.Y(_0016_),
    .A(_0921_),
    .B(_0928_));
 sg13g2_nand3_1 _4737_ (.B(_0875_),
    .C(_0916_),
    .A(net893),
    .Y(_0929_));
 sg13g2_and3_1 _4738_ (.X(_0930_),
    .A(_0827_),
    .B(net891),
    .C(net889));
 sg13g2_nand3_1 _4739_ (.B(net891),
    .C(_0864_),
    .A(_0827_),
    .Y(_0931_));
 sg13g2_nand3_1 _4740_ (.B(net885),
    .C(_0931_),
    .A(_0830_),
    .Y(_0932_));
 sg13g2_a21oi_1 _4741_ (.A1(_0929_),
    .A2(_0932_),
    .Y(_0933_),
    .B1(_0831_));
 sg13g2_nor3_1 _4742_ (.A(_0889_),
    .B(_0908_),
    .C(_0933_),
    .Y(_0000_));
 sg13g2_nand2_1 _4743_ (.Y(_0934_),
    .A(net899),
    .B(net887));
 sg13g2_a221oi_1 _4744_ (.B2(_0871_),
    .C1(net1162),
    .B1(_0867_),
    .A1(_0804_),
    .Y(_0935_),
    .A2(net891));
 sg13g2_o21ai_1 _4745_ (.B1(net886),
    .Y(_0936_),
    .A1(net894),
    .A2(_0931_));
 sg13g2_a221oi_1 _4746_ (.B2(_0913_),
    .C1(_0829_),
    .B1(_0935_),
    .A1(_0849_),
    .Y(_0937_),
    .A2(_0930_));
 sg13g2_a221oi_1 _4747_ (.B2(_0913_),
    .C1(_0830_),
    .B1(_0909_),
    .A1(_0888_),
    .Y(_0938_),
    .A2(_0893_));
 sg13g2_a21oi_1 _4748_ (.A1(_0859_),
    .A2(net888),
    .Y(_0939_),
    .B1(net894));
 sg13g2_nand2_1 _4749_ (.Y(_0940_),
    .A(net885),
    .B(_0897_));
 sg13g2_a21o_1 _4750_ (.A2(_0940_),
    .A1(_0938_),
    .B1(_0937_),
    .X(_0941_));
 sg13g2_nand2b_1 _4751_ (.Y(_0942_),
    .B(net893),
    .A_N(_0895_));
 sg13g2_a22oi_1 _4752_ (.Y(_0001_),
    .B1(_0941_),
    .B2(_0942_),
    .A2(_0938_),
    .A1(net896));
 sg13g2_nor2b_1 _4753_ (.A(net897),
    .B_N(_0891_),
    .Y(_0943_));
 sg13g2_nand2_1 _4754_ (.Y(_0944_),
    .A(net894),
    .B(_0917_));
 sg13g2_a21o_1 _4755_ (.A2(_0934_),
    .A1(_0861_),
    .B1(net885),
    .X(_0945_));
 sg13g2_nor2_1 _4756_ (.A(_0847_),
    .B(_0865_),
    .Y(_0946_));
 sg13g2_nand2_1 _4757_ (.Y(_0947_),
    .A(net895),
    .B(net889));
 sg13g2_and2_1 _4758_ (.A(net897),
    .B(_0947_),
    .X(_0948_));
 sg13g2_a221oi_1 _4759_ (.B2(_0948_),
    .C1(net886),
    .B1(_0945_),
    .A1(_0943_),
    .Y(_0949_),
    .A2(_0944_));
 sg13g2_o21ai_1 _4760_ (.B1(_0913_),
    .Y(_0950_),
    .A1(net884),
    .A2(_0893_));
 sg13g2_or2_1 _4761_ (.X(_0951_),
    .B(_0950_),
    .A(_0895_));
 sg13g2_o21ai_1 _4762_ (.B1(net886),
    .Y(_0952_),
    .A1(net885),
    .A2(_0917_));
 sg13g2_inv_1 _4763_ (.Y(_0953_),
    .A(_0952_));
 sg13g2_a21o_1 _4764_ (.A2(_0953_),
    .A1(_0951_),
    .B1(_0949_),
    .X(_0002_));
 sg13g2_a21oi_1 _4765_ (.A1(net899),
    .A2(net894),
    .Y(_0954_),
    .B1(net896));
 sg13g2_a21o_1 _4766_ (.A2(_0848_),
    .A1(_0803_),
    .B1(net898),
    .X(_0955_));
 sg13g2_xnor2_1 _4767_ (.Y(_0956_),
    .A(_0865_),
    .B(_0939_));
 sg13g2_a21oi_1 _4768_ (.A1(_0862_),
    .A2(_0956_),
    .Y(_0957_),
    .B1(_0936_));
 sg13g2_a21oi_1 _4769_ (.A1(_0938_),
    .A2(_0955_),
    .Y(_0003_),
    .B1(_0957_));
 sg13g2_a221oi_1 _4770_ (.B2(_0861_),
    .C1(net886),
    .B1(_0954_),
    .A1(_0945_),
    .Y(_0958_),
    .A2(_0948_));
 sg13g2_a21o_1 _4771_ (.A2(_0934_),
    .A1(_0861_),
    .B1(_0914_),
    .X(_0959_));
 sg13g2_nand3_1 _4772_ (.B(_0883_),
    .C(_0959_),
    .A(net886),
    .Y(_0960_));
 sg13g2_nand2b_1 _4773_ (.Y(_0004_),
    .B(_0960_),
    .A_N(_0958_));
 sg13g2_nand2_1 _4774_ (.Y(_0961_),
    .A(net894),
    .B(_0934_));
 sg13g2_nand2b_1 _4775_ (.Y(_0962_),
    .B(_0899_),
    .A_N(_0939_));
 sg13g2_a21oi_1 _4776_ (.A1(_0906_),
    .A2(_0909_),
    .Y(_0963_),
    .B1(_0914_));
 sg13g2_o21ai_1 _4777_ (.B1(_0962_),
    .Y(_0964_),
    .A1(_0936_),
    .A2(_0963_));
 sg13g2_nand3_1 _4778_ (.B(_0891_),
    .C(_0947_),
    .A(net897),
    .Y(_0965_));
 sg13g2_a21oi_1 _4779_ (.A1(net892),
    .A2(_0875_),
    .Y(_0966_),
    .B1(_0849_));
 sg13g2_nor3_1 _4780_ (.A(_0817_),
    .B(_0965_),
    .C(_0966_),
    .Y(_0967_));
 sg13g2_a21oi_1 _4781_ (.A1(_0961_),
    .A2(_0964_),
    .Y(_0005_),
    .B1(_0967_));
 sg13g2_nor3_1 _4782_ (.A(_0831_),
    .B(_0895_),
    .C(_0922_),
    .Y(_0968_));
 sg13g2_and2_1 _4783_ (.A(_0886_),
    .B(_0913_),
    .X(_0969_));
 sg13g2_a21o_1 _4784_ (.A2(_0969_),
    .A1(_0912_),
    .B1(_0936_),
    .X(_0970_));
 sg13g2_o21ai_1 _4785_ (.B1(net897),
    .Y(_0971_),
    .A1(net885),
    .A2(net890));
 sg13g2_a21oi_1 _4786_ (.A1(net895),
    .A2(_0893_),
    .Y(_0972_),
    .B1(net886));
 sg13g2_nand2_1 _4787_ (.Y(_0973_),
    .A(_0971_),
    .B(_0972_));
 sg13g2_a21o_1 _4788_ (.A2(_0973_),
    .A1(_0970_),
    .B1(_0968_),
    .X(_0006_));
 sg13g2_a21o_1 _4789_ (.A2(_0877_),
    .A1(net884),
    .B1(net885),
    .X(_0974_));
 sg13g2_nor2b_1 _4790_ (.A(_0965_),
    .B_N(_0903_),
    .Y(_0975_));
 sg13g2_a21o_1 _4791_ (.A2(_0974_),
    .A1(_0943_),
    .B1(net886),
    .X(_0976_));
 sg13g2_nand3_1 _4792_ (.B(_0913_),
    .C(_0916_),
    .A(_0909_),
    .Y(_0977_));
 sg13g2_nand3_1 _4793_ (.B(net894),
    .C(_0877_),
    .A(net899),
    .Y(_0978_));
 sg13g2_nand3_1 _4794_ (.B(_0977_),
    .C(_0978_),
    .A(_0830_),
    .Y(_0979_));
 sg13g2_o21ai_1 _4795_ (.B1(_0979_),
    .Y(_0007_),
    .A1(_0975_),
    .A2(_0976_));
 sg13g2_o21ai_1 _4796_ (.B1(_0831_),
    .Y(_0980_),
    .A1(_0946_),
    .A2(_0966_));
 sg13g2_nor2b_1 _4797_ (.A(_0947_),
    .B_N(_0877_),
    .Y(_0981_));
 sg13g2_a221oi_1 _4798_ (.B2(net898),
    .C1(_0829_),
    .B1(_0981_),
    .A1(_0876_),
    .Y(_0982_),
    .A2(_0914_));
 sg13g2_and3_1 _4799_ (.X(_0983_),
    .A(_0829_),
    .B(_0862_),
    .C(_0931_));
 sg13g2_o21ai_1 _4800_ (.B1(_0980_),
    .Y(_0008_),
    .A1(_0982_),
    .A2(_0983_));
 sg13g2_nor2_1 _4801_ (.A(\i_music.violin_note_idx[3][6] ),
    .B(_2996_),
    .Y(_0984_));
 sg13g2_a22oi_1 _4802_ (.Y(_0985_),
    .B1(net1081),
    .B2(_2953_),
    .A2(_0039_),
    .A1(_2930_));
 sg13g2_nor2b_2 _4803_ (.A(_0984_),
    .B_N(_0985_),
    .Y(_0986_));
 sg13g2_nand2b_2 _4804_ (.Y(_0987_),
    .B(_0985_),
    .A_N(_0984_));
 sg13g2_nor2b_1 _4805_ (.A(net1149),
    .B_N(_0036_),
    .Y(_0988_));
 sg13g2_a21oi_1 _4806_ (.A1(_2947_),
    .A2(net1087),
    .Y(_0989_),
    .B1(_0988_));
 sg13g2_a221oi_1 _4807_ (.B2(_2948_),
    .C1(_0988_),
    .B1(net1080),
    .A1(_2947_),
    .Y(_0990_),
    .A2(net1087));
 sg13g2_o21ai_1 _4808_ (.B1(_0989_),
    .Y(_0991_),
    .A1(\i_music.violin_note_idx[2][5] ),
    .A2(net1079));
 sg13g2_nor2_2 _4809_ (.A(_0986_),
    .B(net1056),
    .Y(_0992_));
 sg13g2_nand2_2 _4810_ (.Y(_0993_),
    .A(_0987_),
    .B(net1017));
 sg13g2_nor2_1 _4811_ (.A(\i_music.violin_note_idx[3][1] ),
    .B(_2996_),
    .Y(_0994_));
 sg13g2_nor2b_1 _4812_ (.A(net1146),
    .B_N(_0040_),
    .Y(_0995_));
 sg13g2_a21o_1 _4813_ (.A2(net1080),
    .A1(_2955_),
    .B1(_0995_),
    .X(_0996_));
 sg13g2_a221oi_1 _4814_ (.B2(_2955_),
    .C1(_0995_),
    .B1(net1080),
    .A1(_2954_),
    .Y(_0997_),
    .A2(net1087));
 sg13g2_nor2b_1 _4815_ (.A(net1146),
    .B_N(_0038_),
    .Y(_0998_));
 sg13g2_a21oi_1 _4816_ (.A1(_2951_),
    .A2(net1087),
    .Y(_0999_),
    .B1(_0998_));
 sg13g2_a221oi_1 _4817_ (.B2(_2952_),
    .C1(_0998_),
    .B1(net1080),
    .A1(_2951_),
    .Y(_1000_),
    .A2(net1087));
 sg13g2_o21ai_1 _4818_ (.B1(_0999_),
    .Y(_1001_),
    .A1(\i_music.violin_note_idx[2][4] ),
    .A2(net1079));
 sg13g2_nor4_2 _4819_ (.A(_0993_),
    .B(_0994_),
    .C(_0996_),
    .Y(_1002_),
    .D(net1051));
 sg13g2_a22oi_1 _4820_ (.Y(_1003_),
    .B1(net1081),
    .B2(_2959_),
    .A2(_0044_),
    .A1(_2930_));
 sg13g2_o21ai_1 _4821_ (.B1(_1003_),
    .Y(_1004_),
    .A1(\i_music.violin_note_idx[3][8] ),
    .A2(_2996_));
 sg13g2_a22oi_1 _4822_ (.Y(_1005_),
    .B1(net1089),
    .B2(_0043_),
    .A2(_0042_),
    .A1(_2930_));
 sg13g2_o21ai_1 _4823_ (.B1(_1005_),
    .Y(_1006_),
    .A1(\i_music.violin_note_idx[2][7] ),
    .A2(net1079));
 sg13g2_nor2b_1 _4824_ (.A(_1006_),
    .B_N(_1004_),
    .Y(_1007_));
 sg13g2_nand2b_2 _4825_ (.Y(_1008_),
    .B(_1004_),
    .A_N(_1006_));
 sg13g2_nor2b_1 _4826_ (.A(net1147),
    .B_N(_0037_),
    .Y(_1009_));
 sg13g2_a21oi_1 _4827_ (.A1(_2950_),
    .A2(net1080),
    .Y(_1010_),
    .B1(_1009_));
 sg13g2_a221oi_1 _4828_ (.B2(_2950_),
    .C1(_1009_),
    .B1(net1080),
    .A1(_2949_),
    .Y(_1011_),
    .A2(net1087));
 sg13g2_o21ai_1 _4829_ (.B1(_1010_),
    .Y(_1012_),
    .A1(\i_music.violin_note_idx[3][3] ),
    .A2(_2996_));
 sg13g2_nor2b_1 _4830_ (.A(net1146),
    .B_N(_0041_),
    .Y(_1013_));
 sg13g2_a221oi_1 _4831_ (.B2(_2958_),
    .C1(_1013_),
    .B1(net1080),
    .A1(_2957_),
    .Y(_1014_),
    .A2(net1087));
 sg13g2_inv_2 _4832_ (.Y(_1015_),
    .A(net1039));
 sg13g2_nor2_2 _4833_ (.A(net1047),
    .B(net1040),
    .Y(_1016_));
 sg13g2_and3_2 _4834_ (.X(_1017_),
    .A(_1002_),
    .B(_1007_),
    .C(_1016_));
 sg13g2_nor2_2 _4835_ (.A(net1053),
    .B(net1038),
    .Y(_1018_));
 sg13g2_or2_2 _4836_ (.X(_1019_),
    .B(net1037),
    .A(net1052));
 sg13g2_nor2b_1 _4837_ (.A(net1146),
    .B_N(_0100_),
    .Y(_1020_));
 sg13g2_a221oi_1 _4838_ (.B2(_2925_),
    .C1(_1020_),
    .B1(net1080),
    .A1(_2956_),
    .Y(_1021_),
    .A2(net1087));
 sg13g2_inv_2 _4839_ (.Y(_1022_),
    .A(net1033));
 sg13g2_and2_2 _4840_ (.A(net1042),
    .B(net1033),
    .X(_1023_));
 sg13g2_nand2_2 _4841_ (.Y(_1024_),
    .A(net1043),
    .B(net1032));
 sg13g2_nand2_1 _4842_ (.Y(_1025_),
    .A(net1042),
    .B(net1038));
 sg13g2_nor2_2 _4843_ (.A(net1039),
    .B(net1034),
    .Y(_1026_));
 sg13g2_or2_1 _4844_ (.X(_1027_),
    .B(net1035),
    .A(net1040));
 sg13g2_o21ai_1 _4845_ (.B1(net1047),
    .Y(_1028_),
    .A1(net1041),
    .A2(net1036));
 sg13g2_nor2_1 _4846_ (.A(_1018_),
    .B(_1028_),
    .Y(_1029_));
 sg13g2_nand2b_2 _4847_ (.Y(_1030_),
    .B(net1054),
    .A_N(net1035));
 sg13g2_nor2_1 _4848_ (.A(net1039),
    .B(_1030_),
    .Y(_1031_));
 sg13g2_or4_2 _4849_ (.A(_0994_),
    .B(_0996_),
    .C(net1040),
    .D(net1035),
    .X(_1032_));
 sg13g2_a21oi_1 _4850_ (.A1(net1010),
    .A2(_1031_),
    .Y(_1033_),
    .B1(_1029_));
 sg13g2_nand3_1 _4851_ (.B(net1014),
    .C(_1033_),
    .A(net1056),
    .Y(_1034_));
 sg13g2_nor2_1 _4852_ (.A(net1052),
    .B(net1033),
    .Y(_1035_));
 sg13g2_or2_1 _4853_ (.X(_1036_),
    .B(net1034),
    .A(net1053));
 sg13g2_nor2_1 _4854_ (.A(net1008),
    .B(_1035_),
    .Y(_1037_));
 sg13g2_nor2_2 _4855_ (.A(net1042),
    .B(net1032),
    .Y(_1038_));
 sg13g2_or2_1 _4856_ (.X(_1039_),
    .B(net1032),
    .A(net1042));
 sg13g2_nor2b_2 _4857_ (.A(net1035),
    .B_N(net1040),
    .Y(_1040_));
 sg13g2_nand2b_2 _4858_ (.Y(_1041_),
    .B(net1038),
    .A_N(net1034));
 sg13g2_nor2_1 _4859_ (.A(net1043),
    .B(_1041_),
    .Y(_1042_));
 sg13g2_nand2_1 _4860_ (.Y(_1043_),
    .A(_0990_),
    .B(net1051));
 sg13g2_a21oi_1 _4861_ (.A1(net1010),
    .A2(_1040_),
    .Y(_1044_),
    .B1(net1015));
 sg13g2_a221oi_1 _4862_ (.B2(net1010),
    .C1(_1043_),
    .B1(_1040_),
    .A1(_1019_),
    .Y(_1045_),
    .A2(_1037_));
 sg13g2_nor2_1 _4863_ (.A(net1048),
    .B(_1018_),
    .Y(_1046_));
 sg13g2_a21oi_1 _4864_ (.A1(net1008),
    .A2(_1018_),
    .Y(_1047_),
    .B1(net1049));
 sg13g2_nor2b_1 _4865_ (.A(net1044),
    .B_N(net1048),
    .Y(_1048_));
 sg13g2_nand2b_1 _4866_ (.Y(_1049_),
    .B(net1051),
    .A_N(net1047));
 sg13g2_nand2b_1 _4867_ (.Y(_1050_),
    .B(net1048),
    .A_N(net1052));
 sg13g2_o21ai_1 _4868_ (.B1(net1017),
    .Y(_1051_),
    .A1(_1019_),
    .A2(_1049_));
 sg13g2_nor2_1 _4869_ (.A(_1047_),
    .B(_1051_),
    .Y(_1052_));
 sg13g2_nor2_1 _4870_ (.A(_1045_),
    .B(_1052_),
    .Y(_1053_));
 sg13g2_a21oi_1 _4871_ (.A1(_1034_),
    .A2(_1053_),
    .Y(_1054_),
    .B1(_0987_));
 sg13g2_or3_2 _4872_ (.A(net1055),
    .B(net1040),
    .C(net1036),
    .X(_1055_));
 sg13g2_and2_2 _4873_ (.A(net1052),
    .B(net1037),
    .X(_1056_));
 sg13g2_nand2_2 _4874_ (.Y(_1057_),
    .A(net1052),
    .B(net1037));
 sg13g2_nand2_2 _4875_ (.Y(_1058_),
    .A(net1040),
    .B(net1035));
 sg13g2_o21ai_1 _4876_ (.B1(net1039),
    .Y(_1059_),
    .A1(net1054),
    .A2(net1036));
 sg13g2_nand3_1 _4877_ (.B(_1055_),
    .C(_1059_),
    .A(net1008),
    .Y(_1060_));
 sg13g2_nand2_1 _4878_ (.Y(_1061_),
    .A(net1049),
    .B(_1025_));
 sg13g2_nor2b_1 _4879_ (.A(_1061_),
    .B_N(_1060_),
    .Y(_1062_));
 sg13g2_nor2b_2 _4880_ (.A(net1053),
    .B_N(net1034),
    .Y(_1063_));
 sg13g2_a21oi_1 _4881_ (.A1(net1045),
    .A2(_1058_),
    .Y(_1064_),
    .B1(_1063_));
 sg13g2_nor4_1 _4882_ (.A(net1049),
    .B(_1018_),
    .C(_1026_),
    .D(_1064_),
    .Y(_1065_));
 sg13g2_nor2_2 _4883_ (.A(_0986_),
    .B(net1016),
    .Y(_1066_));
 sg13g2_nand2_2 _4884_ (.Y(_1067_),
    .A(net1018),
    .B(net1056));
 sg13g2_nor3_1 _4885_ (.A(_1062_),
    .B(_1065_),
    .C(_1067_),
    .Y(_1068_));
 sg13g2_and2_1 _4886_ (.A(_1004_),
    .B(_1006_),
    .X(_1069_));
 sg13g2_nand2_1 _4887_ (.Y(_1070_),
    .A(_1004_),
    .B(_1006_));
 sg13g2_nand2_1 _4888_ (.Y(_1071_),
    .A(net1052),
    .B(net1033));
 sg13g2_a21oi_1 _4889_ (.A1(_1016_),
    .A2(net1007),
    .Y(_1072_),
    .B1(net1014));
 sg13g2_nand3b_1 _4890_ (.B(net1041),
    .C(net1035),
    .Y(_1073_),
    .A_N(net1055));
 sg13g2_nor2_2 _4891_ (.A(net1051),
    .B(_1073_),
    .Y(_1074_));
 sg13g2_nor2_2 _4892_ (.A(_1000_),
    .B(net1047),
    .Y(_1075_));
 sg13g2_nor3_1 _4893_ (.A(_1072_),
    .B(_1074_),
    .C(_1075_),
    .Y(_1076_));
 sg13g2_o21ai_1 _4894_ (.B1(_1069_),
    .Y(_1077_),
    .A1(_0993_),
    .A2(_1076_));
 sg13g2_nor3_2 _4895_ (.A(_1054_),
    .B(_1068_),
    .C(_1077_),
    .Y(_1078_));
 sg13g2_nand3b_1 _4896_ (.B(_1006_),
    .C(net1018),
    .Y(_1079_),
    .A_N(_1004_));
 sg13g2_xor2_1 _4897_ (.B(net1035),
    .A(net1054),
    .X(_1080_));
 sg13g2_xnor2_1 _4898_ (.Y(_1081_),
    .A(net1053),
    .B(net1034));
 sg13g2_nand4_1 _4899_ (.B(net1014),
    .C(_1016_),
    .A(net1056),
    .Y(_1082_),
    .D(_1080_));
 sg13g2_nor2_1 _4900_ (.A(_0990_),
    .B(net1051),
    .Y(_1083_));
 sg13g2_inv_1 _4901_ (.Y(_1084_),
    .A(net1006));
 sg13g2_nand2_1 _4902_ (.Y(_1085_),
    .A(net1034),
    .B(_1056_));
 sg13g2_nor2_1 _4903_ (.A(_1024_),
    .B(_1057_),
    .Y(_1086_));
 sg13g2_nor2b_2 _4904_ (.A(net1056),
    .B_N(net1049),
    .Y(_1087_));
 sg13g2_nand2_1 _4905_ (.Y(_1088_),
    .A(net1016),
    .B(net1050));
 sg13g2_a22oi_1 _4906_ (.Y(_1089_),
    .B1(_1086_),
    .B2(_1087_),
    .A2(net1006),
    .A1(_1038_));
 sg13g2_a21oi_1 _4907_ (.A1(_1082_),
    .A2(_1089_),
    .Y(_1090_),
    .B1(_1079_));
 sg13g2_nor2_1 _4908_ (.A(net1013),
    .B(_1026_),
    .Y(_1091_));
 sg13g2_a21oi_1 _4909_ (.A1(_1037_),
    .A2(_1091_),
    .Y(_1092_),
    .B1(_1074_));
 sg13g2_or4_1 _4910_ (.A(net1052),
    .B(net1048),
    .C(net1044),
    .D(net1037),
    .X(_1093_));
 sg13g2_nand3_1 _4911_ (.B(_1092_),
    .C(_1093_),
    .A(net1056),
    .Y(_1094_));
 sg13g2_nand4_1 _4912_ (.B(_1028_),
    .C(_1058_),
    .A(net1054),
    .Y(_1095_),
    .D(_1083_));
 sg13g2_a21oi_1 _4913_ (.A1(_1094_),
    .A2(_1095_),
    .Y(_1096_),
    .B1(_0986_));
 sg13g2_nor2_1 _4914_ (.A(net1018),
    .B(_0990_),
    .Y(_1097_));
 sg13g2_a221oi_1 _4915_ (.B2(_1023_),
    .C1(net1048),
    .B1(_1056_),
    .A1(net1008),
    .Y(_1098_),
    .A2(_1055_));
 sg13g2_o21ai_1 _4916_ (.B1(_0986_),
    .Y(_1099_),
    .A1(net1016),
    .A2(_1098_));
 sg13g2_nor2_1 _4917_ (.A(net1033),
    .B(_1093_),
    .Y(_1100_));
 sg13g2_nor2_1 _4918_ (.A(net1013),
    .B(net1008),
    .Y(_1101_));
 sg13g2_nand2_1 _4919_ (.Y(_1102_),
    .A(net1048),
    .B(net1044));
 sg13g2_a21oi_1 _4920_ (.A1(_1019_),
    .A2(_1101_),
    .Y(_1103_),
    .B1(_1100_));
 sg13g2_a21oi_1 _4921_ (.A1(net1016),
    .A2(_1103_),
    .Y(_1104_),
    .B1(_1099_));
 sg13g2_nor3_1 _4922_ (.A(_0993_),
    .B(_1049_),
    .C(_1085_),
    .Y(_1105_));
 sg13g2_nor4_2 _4923_ (.A(_1008_),
    .B(_1096_),
    .C(_1104_),
    .Y(_1106_),
    .D(_1105_));
 sg13g2_nor3_2 _4924_ (.A(_1078_),
    .B(_1090_),
    .C(_1106_),
    .Y(_1107_));
 sg13g2_or3_1 _4925_ (.A(_1078_),
    .B(_1090_),
    .C(_1106_),
    .X(_1108_));
 sg13g2_nand3b_1 _4926_ (.B(net1045),
    .C(_1058_),
    .Y(_1109_),
    .A_N(_1063_));
 sg13g2_nand2_1 _4927_ (.Y(_1110_),
    .A(net1037),
    .B(net1007));
 sg13g2_nand3_1 _4928_ (.B(net1038),
    .C(net1007),
    .A(net1009),
    .Y(_1111_));
 sg13g2_nand3_1 _4929_ (.B(_1109_),
    .C(_1111_),
    .A(_1091_),
    .Y(_1112_));
 sg13g2_nand2_2 _4930_ (.Y(_1113_),
    .A(_1022_),
    .B(_1056_));
 sg13g2_nand3_1 _4931_ (.B(_1055_),
    .C(_1113_),
    .A(net1009),
    .Y(_1114_));
 sg13g2_nand3_1 _4932_ (.B(_1024_),
    .C(_1114_),
    .A(net1012),
    .Y(_1115_));
 sg13g2_nand3_1 _4933_ (.B(_1112_),
    .C(_1115_),
    .A(net1017),
    .Y(_1116_));
 sg13g2_a21oi_1 _4934_ (.A1(_1031_),
    .A2(_1075_),
    .Y(_1117_),
    .B1(net1017));
 sg13g2_nand2b_2 _4935_ (.Y(_1118_),
    .B(net1016),
    .A_N(_1079_));
 sg13g2_nor2_1 _4936_ (.A(_1079_),
    .B(_1117_),
    .Y(_1119_));
 sg13g2_nand2_1 _4937_ (.Y(_1120_),
    .A(_1063_),
    .B(_1075_));
 sg13g2_nor2_1 _4938_ (.A(net1010),
    .B(_1040_),
    .Y(_1121_));
 sg13g2_nor2_1 _4939_ (.A(net1039),
    .B(_1080_),
    .Y(_1122_));
 sg13g2_a221oi_1 _4940_ (.B2(net1053),
    .C1(net1012),
    .B1(_1121_),
    .A1(_1015_),
    .Y(_1123_),
    .A2(_1081_));
 sg13g2_nand4_1 _4941_ (.B(net1050),
    .C(_1015_),
    .A(net1052),
    .Y(_1124_),
    .D(_1023_));
 sg13g2_nor2_1 _4942_ (.A(_1019_),
    .B(_1022_),
    .Y(_1125_));
 sg13g2_nand3_1 _4943_ (.B(_1041_),
    .C(_1057_),
    .A(net1043),
    .Y(_1126_));
 sg13g2_o21ai_1 _4944_ (.B1(net1013),
    .Y(_1127_),
    .A1(_1125_),
    .A2(_1126_));
 sg13g2_nand3b_1 _4945_ (.B(_1124_),
    .C(_1127_),
    .Y(_1128_),
    .A_N(_1123_));
 sg13g2_a21oi_1 _4946_ (.A1(_1120_),
    .A2(_1128_),
    .Y(_1129_),
    .B1(_1067_));
 sg13g2_nand2_2 _4947_ (.Y(_1130_),
    .A(_0986_),
    .B(net1056));
 sg13g2_nor2_1 _4948_ (.A(_1022_),
    .B(_1093_),
    .Y(_1131_));
 sg13g2_nand2_1 _4949_ (.Y(_1132_),
    .A(_1032_),
    .B(_1058_));
 sg13g2_nand3_1 _4950_ (.B(_1032_),
    .C(_1058_),
    .A(net1009),
    .Y(_1133_));
 sg13g2_nor2_1 _4951_ (.A(net1050),
    .B(_1063_),
    .Y(_1134_));
 sg13g2_a21oi_1 _4952_ (.A1(_1133_),
    .A2(_1134_),
    .Y(_1135_),
    .B1(_1131_));
 sg13g2_o21ai_1 _4953_ (.B1(net1032),
    .Y(_1136_),
    .A1(net1043),
    .A2(net1038));
 sg13g2_a21oi_1 _4954_ (.A1(_1018_),
    .A2(_1024_),
    .Y(_1137_),
    .B1(net1012));
 sg13g2_o21ai_1 _4955_ (.B1(_1137_),
    .Y(_1138_),
    .A1(_1018_),
    .A2(_1136_));
 sg13g2_a21o_1 _4956_ (.A2(_1138_),
    .A1(_1135_),
    .B1(_1130_),
    .X(_1139_));
 sg13g2_o21ai_1 _4957_ (.B1(net1054),
    .Y(_1140_),
    .A1(net1040),
    .A2(net1035));
 sg13g2_nand2_1 _4958_ (.Y(_1141_),
    .A(_1055_),
    .B(_1140_));
 sg13g2_a21o_1 _4959_ (.A2(_1030_),
    .A1(net1040),
    .B1(net1046),
    .X(_1142_));
 sg13g2_a221oi_1 _4960_ (.B2(_1142_),
    .C1(net1051),
    .B1(_1141_),
    .A1(_1016_),
    .Y(_1143_),
    .A2(_1080_));
 sg13g2_a21oi_1 _4961_ (.A1(net1054),
    .A2(_1058_),
    .Y(_1144_),
    .B1(_1028_));
 sg13g2_and3_1 _4962_ (.X(_1145_),
    .A(net1054),
    .B(net1011),
    .C(_1058_));
 sg13g2_nor3_1 _4963_ (.A(net1014),
    .B(_1144_),
    .C(_1145_),
    .Y(_1146_));
 sg13g2_o21ai_1 _4964_ (.B1(_1097_),
    .Y(_1147_),
    .A1(_1143_),
    .A2(_1146_));
 sg13g2_a21oi_1 _4965_ (.A1(_1015_),
    .A2(_1081_),
    .Y(_1148_),
    .B1(_1040_));
 sg13g2_nand3_1 _4966_ (.B(_1019_),
    .C(_1071_),
    .A(net1046),
    .Y(_1149_));
 sg13g2_nand2b_2 _4967_ (.Y(_1150_),
    .B(net1046),
    .A_N(net1034));
 sg13g2_a221oi_1 _4968_ (.B2(_1149_),
    .C1(net1014),
    .B1(_1148_),
    .A1(net1046),
    .Y(_1151_),
    .A2(_1040_));
 sg13g2_nand3_1 _4969_ (.B(_1041_),
    .C(_1080_),
    .A(net1045),
    .Y(_1152_));
 sg13g2_nand2b_1 _4970_ (.Y(_1153_),
    .B(net1014),
    .A_N(_1152_));
 sg13g2_nand3b_1 _4971_ (.B(_1153_),
    .C(_0992_),
    .Y(_1154_),
    .A_N(_1151_));
 sg13g2_nand4_1 _4972_ (.B(_1139_),
    .C(_1147_),
    .A(_1006_),
    .Y(_1155_),
    .D(_1154_));
 sg13g2_a21oi_1 _4973_ (.A1(_1133_),
    .A2(_1152_),
    .Y(_1156_),
    .B1(_1088_));
 sg13g2_a21oi_1 _4974_ (.A1(_1036_),
    .A2(_1041_),
    .Y(_1157_),
    .B1(net1012));
 sg13g2_nor2_1 _4975_ (.A(_1015_),
    .B(_1080_),
    .Y(_1158_));
 sg13g2_nor4_1 _4976_ (.A(net1016),
    .B(_1038_),
    .C(_1157_),
    .D(_1158_),
    .Y(_1159_));
 sg13g2_o21ai_1 _4977_ (.B1(net1006),
    .Y(_1160_),
    .A1(net1046),
    .A2(_1081_));
 sg13g2_a21oi_1 _4978_ (.A1(_1081_),
    .A2(_1121_),
    .Y(_1161_),
    .B1(_1160_));
 sg13g2_or4_1 _4979_ (.A(net1018),
    .B(_1156_),
    .C(_1159_),
    .D(_1161_),
    .X(_1162_));
 sg13g2_a221oi_1 _4980_ (.B2(net1010),
    .C1(net1015),
    .B1(_1141_),
    .A1(net1054),
    .Y(_1163_),
    .A2(_1121_));
 sg13g2_o21ai_1 _4981_ (.B1(_0992_),
    .Y(_1164_),
    .A1(_1074_),
    .A2(_1163_));
 sg13g2_a221oi_1 _4982_ (.B2(net1039),
    .C1(_1067_),
    .B1(_1081_),
    .A1(net1046),
    .Y(_1165_),
    .A2(_1026_));
 sg13g2_o21ai_1 _4983_ (.B1(_1165_),
    .Y(_1166_),
    .A1(net1050),
    .A2(_1148_));
 sg13g2_a21oi_1 _4984_ (.A1(_1002_),
    .A2(_1028_),
    .Y(_1167_),
    .B1(_1006_));
 sg13g2_nand4_1 _4985_ (.B(_1164_),
    .C(_1166_),
    .A(_1162_),
    .Y(_1168_),
    .D(_1167_));
 sg13g2_o21ai_1 _4986_ (.B1(_1168_),
    .Y(_1169_),
    .A1(_1129_),
    .A2(_1155_));
 sg13g2_a22oi_1 _4987_ (.Y(_1170_),
    .B1(_1169_),
    .B2(_1004_),
    .A2(_1119_),
    .A1(_1116_));
 sg13g2_nand4_1 _4988_ (.B(_1019_),
    .C(_1027_),
    .A(net1046),
    .Y(_1171_),
    .D(_1057_));
 sg13g2_and2_1 _4989_ (.A(_1028_),
    .B(_1032_),
    .X(_1172_));
 sg13g2_a221oi_1 _4990_ (.B2(net1014),
    .C1(net1017),
    .B1(_1172_),
    .A1(_1044_),
    .Y(_1173_),
    .A2(_1171_));
 sg13g2_a22oi_1 _4991_ (.Y(_1174_),
    .B1(_1055_),
    .B2(net1010),
    .A2(_1027_),
    .A1(net1055));
 sg13g2_nor2_1 _4992_ (.A(net1043),
    .B(_1057_),
    .Y(_1175_));
 sg13g2_o21ai_1 _4993_ (.B1(net1006),
    .Y(_1176_),
    .A1(net1046),
    .A2(_1057_));
 sg13g2_nand2_1 _4994_ (.Y(_1177_),
    .A(_1087_),
    .B(_1150_));
 sg13g2_nand3_1 _4995_ (.B(_1087_),
    .C(_1150_),
    .A(_1018_),
    .Y(_1178_));
 sg13g2_o21ai_1 _4996_ (.B1(_1178_),
    .Y(_1179_),
    .A1(_1174_),
    .A2(_1176_));
 sg13g2_o21ai_1 _4997_ (.B1(_0986_),
    .Y(_1180_),
    .A1(_1173_),
    .A2(_1179_));
 sg13g2_a21o_1 _4998_ (.A2(_1073_),
    .A1(_1055_),
    .B1(net1010),
    .X(_1181_));
 sg13g2_a21oi_1 _4999_ (.A1(_1072_),
    .A2(_1181_),
    .Y(_1182_),
    .B1(_0993_));
 sg13g2_o21ai_1 _5000_ (.B1(_1182_),
    .Y(_1183_),
    .A1(net1051),
    .A2(_1181_));
 sg13g2_o21ai_1 _5001_ (.B1(net1009),
    .Y(_1184_),
    .A1(_1026_),
    .A2(_1063_));
 sg13g2_nand2b_1 _5002_ (.Y(_1185_),
    .B(_1059_),
    .A_N(_1028_));
 sg13g2_a21oi_1 _5003_ (.A1(_1184_),
    .A2(_1185_),
    .Y(_1186_),
    .B1(net1049));
 sg13g2_a22oi_1 _5004_ (.Y(_1187_),
    .B1(_1050_),
    .B2(_1061_),
    .A2(_1036_),
    .A1(_1016_));
 sg13g2_o21ai_1 _5005_ (.B1(_1066_),
    .Y(_1188_),
    .A1(_1186_),
    .A2(_1187_));
 sg13g2_nand4_1 _5006_ (.B(_1180_),
    .C(_1183_),
    .A(_1069_),
    .Y(_1189_),
    .D(_1188_));
 sg13g2_a21oi_1 _5007_ (.A1(_1050_),
    .A2(_1061_),
    .Y(_1190_),
    .B1(_1022_));
 sg13g2_nor2b_1 _5008_ (.A(net1042),
    .B_N(net1032),
    .Y(_1191_));
 sg13g2_nand2b_2 _5009_ (.Y(_1192_),
    .B(net1032),
    .A_N(net1042));
 sg13g2_nor3_1 _5010_ (.A(net1016),
    .B(_1019_),
    .C(_1192_),
    .Y(_1193_));
 sg13g2_a21oi_1 _5011_ (.A1(net1056),
    .A2(_1190_),
    .Y(_1194_),
    .B1(_1079_));
 sg13g2_o21ai_1 _5012_ (.B1(_1194_),
    .Y(_1195_),
    .A1(_1190_),
    .A2(_1193_));
 sg13g2_o21ai_1 _5013_ (.B1(_1060_),
    .Y(_1196_),
    .A1(net1008),
    .A2(_1122_));
 sg13g2_a221oi_1 _5014_ (.B2(net1006),
    .C1(_1099_),
    .B1(_1196_),
    .A1(_1033_),
    .Y(_1197_),
    .A2(_1087_));
 sg13g2_and3_1 _5015_ (.X(_1198_),
    .A(net1042),
    .B(net1037),
    .C(net1032));
 sg13g2_nand2_1 _5016_ (.Y(_1199_),
    .A(net1037),
    .B(_1023_));
 sg13g2_nand2_1 _5017_ (.Y(_1200_),
    .A(_0992_),
    .B(_1102_));
 sg13g2_a221oi_1 _5018_ (.B2(_1047_),
    .C1(_0993_),
    .B1(_1199_),
    .A1(_1101_),
    .Y(_1201_),
    .A2(_1110_));
 sg13g2_nor4_1 _5019_ (.A(net1013),
    .B(net1044),
    .C(_1026_),
    .D(_1036_),
    .Y(_1202_));
 sg13g2_nor3_1 _5020_ (.A(_1067_),
    .B(_1100_),
    .C(_1202_),
    .Y(_1203_));
 sg13g2_a21o_1 _5021_ (.A2(_1203_),
    .A1(_1092_),
    .B1(_1201_),
    .X(_1204_));
 sg13g2_o21ai_1 _5022_ (.B1(_1007_),
    .Y(_1205_),
    .A1(_1197_),
    .A2(_1204_));
 sg13g2_nand3_1 _5023_ (.B(_1195_),
    .C(_1205_),
    .A(_1189_),
    .Y(_1206_));
 sg13g2_inv_1 _5024_ (.Y(_1207_),
    .A(_1206_));
 sg13g2_nand2_1 _5025_ (.Y(_1208_),
    .A(net985),
    .B(_1207_));
 sg13g2_nand4_1 _5026_ (.B(_1032_),
    .C(_1041_),
    .A(net1043),
    .Y(_1209_),
    .D(_1057_));
 sg13g2_a21oi_1 _5027_ (.A1(_1192_),
    .A2(_1209_),
    .Y(_1210_),
    .B1(_1084_));
 sg13g2_nand2_1 _5028_ (.Y(_1211_),
    .A(net1032),
    .B(_1057_));
 sg13g2_nor2_1 _5029_ (.A(_1056_),
    .B(_1192_),
    .Y(_1212_));
 sg13g2_nor2_1 _5030_ (.A(_1177_),
    .B(_1212_),
    .Y(_1213_));
 sg13g2_o21ai_1 _5031_ (.B1(_0986_),
    .Y(_1214_),
    .A1(_1210_),
    .A2(_1213_));
 sg13g2_nor2_1 _5032_ (.A(_1025_),
    .B(_1081_),
    .Y(_1215_));
 sg13g2_o21ai_1 _5033_ (.B1(net1012),
    .Y(_1216_),
    .A1(_1212_),
    .A2(_1215_));
 sg13g2_o21ai_1 _5034_ (.B1(net1044),
    .Y(_1217_),
    .A1(_1022_),
    .A2(_1056_));
 sg13g2_nand3_1 _5035_ (.B(_1133_),
    .C(_1217_),
    .A(net1050),
    .Y(_1218_));
 sg13g2_nand3_1 _5036_ (.B(_1216_),
    .C(_1218_),
    .A(_0992_),
    .Y(_1219_));
 sg13g2_a221oi_1 _5037_ (.B2(_1192_),
    .C1(_1035_),
    .B1(_1102_),
    .A1(net1037),
    .Y(_1220_),
    .A2(_1022_));
 sg13g2_a21oi_1 _5038_ (.A1(_1015_),
    .A2(_1030_),
    .Y(_1221_),
    .B1(net1050));
 sg13g2_and3_1 _5039_ (.X(_1222_),
    .A(net1044),
    .B(_1113_),
    .C(_1221_));
 sg13g2_o21ai_1 _5040_ (.B1(_1066_),
    .Y(_1223_),
    .A1(_1220_),
    .A2(_1222_));
 sg13g2_nand3_1 _5041_ (.B(_1113_),
    .C(_1211_),
    .A(_1101_),
    .Y(_1224_));
 sg13g2_nand3_1 _5042_ (.B(_1030_),
    .C(_1150_),
    .A(_1027_),
    .Y(_1225_));
 sg13g2_a221oi_1 _5043_ (.B2(net1013),
    .C1(_1130_),
    .B1(_1225_),
    .A1(net1009),
    .Y(_1226_),
    .A2(_1157_));
 sg13g2_a21oi_1 _5044_ (.A1(_1224_),
    .A2(_1226_),
    .Y(_1227_),
    .B1(_1008_));
 sg13g2_nand4_1 _5045_ (.B(_1219_),
    .C(_1223_),
    .A(_1214_),
    .Y(_1228_),
    .D(_1227_));
 sg13g2_nand3_1 _5046_ (.B(_1135_),
    .C(_1192_),
    .A(net1007),
    .Y(_1229_));
 sg13g2_a21oi_1 _5047_ (.A1(net1007),
    .A2(_1192_),
    .Y(_1230_),
    .B1(net1048));
 sg13g2_nor2_1 _5048_ (.A(_1118_),
    .B(_1230_),
    .Y(_1231_));
 sg13g2_nand2_1 _5049_ (.Y(_1232_),
    .A(_1229_),
    .B(_1231_));
 sg13g2_nand3_1 _5050_ (.B(_1113_),
    .C(_1211_),
    .A(net1008),
    .Y(_1233_));
 sg13g2_nor2_1 _5051_ (.A(_1023_),
    .B(_1088_),
    .Y(_1234_));
 sg13g2_nand3_1 _5052_ (.B(net1007),
    .C(_1192_),
    .A(net1038),
    .Y(_1235_));
 sg13g2_nand3_1 _5053_ (.B(_1015_),
    .C(_1081_),
    .A(net1043),
    .Y(_1236_));
 sg13g2_nor3_1 _5054_ (.A(net1050),
    .B(_1038_),
    .C(_1198_),
    .Y(_1237_));
 sg13g2_a21oi_1 _5055_ (.A1(_1039_),
    .A2(_1136_),
    .Y(_1238_),
    .B1(net1012));
 sg13g2_a221oi_1 _5056_ (.B2(_1235_),
    .C1(net1016),
    .B1(_1238_),
    .A1(_1236_),
    .Y(_1239_),
    .A2(_1237_));
 sg13g2_a21o_1 _5057_ (.A2(_1132_),
    .A1(_1111_),
    .B1(_1042_),
    .X(_1240_));
 sg13g2_a221oi_1 _5058_ (.B2(net1006),
    .C1(_1239_),
    .B1(_1240_),
    .A1(_1233_),
    .Y(_1241_),
    .A2(_1234_));
 sg13g2_a221oi_1 _5059_ (.B2(_1057_),
    .C1(net1012),
    .B1(_1191_),
    .A1(net1042),
    .Y(_1242_),
    .A2(net1007));
 sg13g2_a21o_1 _5060_ (.A2(_1024_),
    .A1(net1012),
    .B1(_1242_),
    .X(_1243_));
 sg13g2_nand2b_1 _5061_ (.Y(_1244_),
    .B(_1048_),
    .A_N(_1059_));
 sg13g2_a22oi_1 _5062_ (.Y(_1245_),
    .B1(_1048_),
    .B2(_1018_),
    .A2(_1023_),
    .A1(net1048));
 sg13g2_nand4_1 _5063_ (.B(net1044),
    .C(_1019_),
    .A(net1013),
    .Y(_1246_),
    .D(net1007));
 sg13g2_nand3_1 _5064_ (.B(_1030_),
    .C(_1075_),
    .A(net1041),
    .Y(_1247_));
 sg13g2_nand4_1 _5065_ (.B(_1245_),
    .C(_1246_),
    .A(_1244_),
    .Y(_1248_),
    .D(_1247_));
 sg13g2_a221oi_1 _5066_ (.B2(_1066_),
    .C1(_1070_),
    .B1(_1248_),
    .A1(_0992_),
    .Y(_1249_),
    .A2(_1243_));
 sg13g2_o21ai_1 _5067_ (.B1(_1249_),
    .Y(_1250_),
    .A1(net1018),
    .A2(_1241_));
 sg13g2_and3_2 _5068_ (.X(_1251_),
    .A(_1228_),
    .B(_1232_),
    .C(_1250_));
 sg13g2_nand3_1 _5069_ (.B(_1232_),
    .C(_1250_),
    .A(_1228_),
    .Y(_1252_));
 sg13g2_nand2_1 _5070_ (.Y(_1253_),
    .A(_1206_),
    .B(_1252_));
 sg13g2_or2_1 _5071_ (.X(_1254_),
    .B(_1253_),
    .A(net986));
 sg13g2_nand2_1 _5072_ (.Y(_1255_),
    .A(_1207_),
    .B(_1251_));
 sg13g2_o21ai_1 _5073_ (.B1(_1207_),
    .Y(_1256_),
    .A1(net985),
    .A2(_1251_));
 sg13g2_a21o_1 _5074_ (.A2(_1256_),
    .A1(_1254_),
    .B1(net987),
    .X(_1257_));
 sg13g2_a221oi_1 _5075_ (.B2(_1004_),
    .C1(_1252_),
    .B1(_1169_),
    .A1(_1116_),
    .Y(_1258_),
    .A2(_1119_));
 sg13g2_nand2_1 _5076_ (.Y(_1259_),
    .A(net986),
    .B(_1251_));
 sg13g2_nand3_1 _5077_ (.B(_1254_),
    .C(_1259_),
    .A(net987),
    .Y(_1260_));
 sg13g2_a21oi_1 _5078_ (.A1(_1257_),
    .A2(_1260_),
    .Y(_1261_),
    .B1(_1017_));
 sg13g2_nor2_1 _5079_ (.A(net1071),
    .B(_1017_),
    .Y(_1262_));
 sg13g2_or2_1 _5080_ (.X(_1263_),
    .B(_1017_),
    .A(net1073));
 sg13g2_a21oi_1 _5081_ (.A1(net1068),
    .A2(_1251_),
    .Y(_1264_),
    .B1(_1262_));
 sg13g2_xor2_1 _5082_ (.B(\i_music.count[20] ),
    .A(\i_music.count[21] ),
    .X(_1265_));
 sg13g2_xnor2_1 _5083_ (.Y(_1266_),
    .A(\i_music.count[21] ),
    .B(\i_music.count[20] ));
 sg13g2_xnor2_1 _5084_ (.Y(_1267_),
    .A(\i_music.count[19] ),
    .B(\i_music.count[21] ));
 sg13g2_xor2_1 _5085_ (.B(\i_music.count[21] ),
    .A(\i_music.count[19] ),
    .X(_1268_));
 sg13g2_nor3_1 _5086_ (.A(_2946_),
    .B(_1266_),
    .C(_1268_),
    .Y(_1269_));
 sg13g2_a21oi_1 _5087_ (.A1(_1265_),
    .A2(_1267_),
    .Y(_1270_),
    .B1(\i_music.count[22] ));
 sg13g2_or2_1 _5088_ (.X(_1271_),
    .B(_1270_),
    .A(_1269_));
 sg13g2_and2_1 _5089_ (.A(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[0] ),
    .B(_1271_),
    .X(_1272_));
 sg13g2_o21ai_1 _5090_ (.B1(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[0] ),
    .Y(_1273_),
    .A1(_1269_),
    .A2(_1270_));
 sg13g2_nand2_1 _5091_ (.Y(_1274_),
    .A(\i_music.violin_note_idx[1][7] ),
    .B(\i_music.violin_note_idx[1][8] ));
 sg13g2_and2_1 _5092_ (.A(net1072),
    .B(_1274_),
    .X(_1275_));
 sg13g2_nand2_2 _5093_ (.Y(_1276_),
    .A(net1072),
    .B(_1274_));
 sg13g2_o21ai_1 _5094_ (.B1(_1275_),
    .Y(_1277_),
    .A1(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[0] ),
    .A2(_1271_));
 sg13g2_nand2b_1 _5095_ (.Y(_1278_),
    .B(_1273_),
    .A_N(_1277_));
 sg13g2_o21ai_1 _5096_ (.B1(_1278_),
    .Y(_1279_),
    .A1(_1261_),
    .A2(_1264_));
 sg13g2_or2_1 _5097_ (.X(_1280_),
    .B(_1279_),
    .A(\i_music.i_sample.thresh[0] ));
 sg13g2_nand2_1 _5098_ (.Y(_1281_),
    .A(\i_music.i_sample.thresh[0] ),
    .B(_1279_));
 sg13g2_and3_1 _5099_ (.X(\i_music.i_sample.t1.genblk1[8].state.D ),
    .A(net1171),
    .B(_1280_),
    .C(_1281_));
 sg13g2_o21ai_1 _5100_ (.B1(_1206_),
    .Y(_1282_),
    .A1(_1107_),
    .A2(net985));
 sg13g2_nor2b_1 _5101_ (.A(_1017_),
    .B_N(_1282_),
    .Y(_1283_));
 sg13g2_a21o_1 _5102_ (.A2(net985),
    .A1(_1107_),
    .B1(_1252_),
    .X(_1284_));
 sg13g2_nor2_1 _5103_ (.A(_1252_),
    .B(_1283_),
    .Y(_1285_));
 sg13g2_a21o_1 _5104_ (.A2(_1284_),
    .A1(_1283_),
    .B1(net1071),
    .X(_1286_));
 sg13g2_o21ai_1 _5105_ (.B1(\i_music.count[22] ),
    .Y(_1287_),
    .A1(_1265_),
    .A2(_1268_));
 sg13g2_nand3_1 _5106_ (.B(_1266_),
    .C(_1267_),
    .A(_2946_),
    .Y(_1288_));
 sg13g2_and2_1 _5107_ (.A(_1287_),
    .B(_1288_),
    .X(_1289_));
 sg13g2_nand3_1 _5108_ (.B(_1287_),
    .C(_1288_),
    .A(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[1] ),
    .Y(_1290_));
 sg13g2_a21oi_1 _5109_ (.A1(_1287_),
    .A2(_1288_),
    .Y(_1291_),
    .B1(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[1] ));
 sg13g2_xor2_1 _5110_ (.B(_1289_),
    .A(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[1] ),
    .X(_1292_));
 sg13g2_and2_1 _5111_ (.A(_1272_),
    .B(_1292_),
    .X(_1293_));
 sg13g2_nor2_1 _5112_ (.A(_1276_),
    .B(_1293_),
    .Y(_1294_));
 sg13g2_o21ai_1 _5113_ (.B1(_1294_),
    .Y(_1295_),
    .A1(_1272_),
    .A2(_1292_));
 sg13g2_o21ai_1 _5114_ (.B1(_1295_),
    .Y(_1296_),
    .A1(_1285_),
    .A2(_1286_));
 sg13g2_xor2_1 _5115_ (.B(_1296_),
    .A(_0056_),
    .X(_1297_));
 sg13g2_nor2_1 _5116_ (.A(_1281_),
    .B(_1297_),
    .Y(_1298_));
 sg13g2_a21oi_1 _5117_ (.A1(_1281_),
    .A2(_1297_),
    .Y(_1299_),
    .B1(net1158));
 sg13g2_nor2b_1 _5118_ (.A(_1298_),
    .B_N(_1299_),
    .Y(\i_music.i_sample.t1.genblk1[9].state.D ));
 sg13g2_a21o_1 _5119_ (.A2(_1296_),
    .A1(\i_music.i_sample.thresh[1] ),
    .B1(_1298_),
    .X(_1300_));
 sg13g2_and3_1 _5120_ (.X(_1301_),
    .A(_1108_),
    .B(_1253_),
    .C(_1255_));
 sg13g2_nor2_1 _5121_ (.A(net987),
    .B(_1255_),
    .Y(_1302_));
 sg13g2_o21ai_1 _5122_ (.B1(_1262_),
    .Y(_1303_),
    .A1(net986),
    .A2(_1302_));
 sg13g2_xnor2_1 _5123_ (.Y(_1304_),
    .A(_0035_),
    .B(_1265_));
 sg13g2_nand2_1 _5124_ (.Y(_1305_),
    .A(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[2] ),
    .B(_1304_));
 sg13g2_xnor2_1 _5125_ (.Y(_1306_),
    .A(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[2] ),
    .B(_1304_));
 sg13g2_a21oi_1 _5126_ (.A1(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[1] ),
    .A2(_1289_),
    .Y(_1307_),
    .B1(_1293_));
 sg13g2_o21ai_1 _5127_ (.B1(_1290_),
    .Y(_1308_),
    .A1(_1273_),
    .A2(_1291_));
 sg13g2_nand2b_1 _5128_ (.Y(_1309_),
    .B(_1308_),
    .A_N(_1306_));
 sg13g2_a22oi_1 _5129_ (.Y(_1310_),
    .B1(_1306_),
    .B2(_1307_),
    .A2(\i_music.violin_note_idx[1][8] ),
    .A1(\i_music.violin_note_idx[1][7] ));
 sg13g2_a21o_1 _5130_ (.A2(_1310_),
    .A1(_1309_),
    .B1(net1068),
    .X(_1311_));
 sg13g2_o21ai_1 _5131_ (.B1(_1311_),
    .Y(_1312_),
    .A1(_1301_),
    .A2(_1303_));
 sg13g2_nor2_1 _5132_ (.A(_1206_),
    .B(_1258_),
    .Y(_1313_));
 sg13g2_o21ai_1 _5133_ (.B1(_1251_),
    .Y(_1314_),
    .A1(net985),
    .A2(_1206_));
 sg13g2_and2_1 _5134_ (.A(_1107_),
    .B(_1314_),
    .X(_1315_));
 sg13g2_nand2_1 _5135_ (.Y(_1316_),
    .A(net987),
    .B(net986));
 sg13g2_nand2b_1 _5136_ (.Y(_1317_),
    .B(_1316_),
    .A_N(_1017_));
 sg13g2_nor3_1 _5137_ (.A(_1301_),
    .B(_1315_),
    .C(_1317_),
    .Y(_1318_));
 sg13g2_nand2_1 _5138_ (.Y(_1319_),
    .A(_2946_),
    .B(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[3] ));
 sg13g2_xor2_1 _5139_ (.B(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[3] ),
    .A(\i_music.count[22] ),
    .X(_1320_));
 sg13g2_a21o_1 _5140_ (.A2(_1309_),
    .A1(_1305_),
    .B1(_1320_),
    .X(_1321_));
 sg13g2_nand3_1 _5141_ (.B(_1319_),
    .C(_1321_),
    .A(_2970_),
    .Y(_1322_));
 sg13g2_a21oi_2 _5142_ (.B1(_2970_),
    .Y(_1323_),
    .A2(_1321_),
    .A1(_1319_));
 sg13g2_nand3b_1 _5143_ (.B(_1275_),
    .C(_1322_),
    .Y(_1324_),
    .A_N(_1323_));
 sg13g2_o21ai_1 _5144_ (.B1(_1324_),
    .Y(_1325_),
    .A1(net1071),
    .A2(_1318_));
 sg13g2_nand2_1 _5145_ (.Y(_1326_),
    .A(_1107_),
    .B(_1208_));
 sg13g2_xnor2_1 _5146_ (.Y(_1327_),
    .A(net985),
    .B(_1251_));
 sg13g2_a21o_1 _5147_ (.A2(_1327_),
    .A1(_1206_),
    .B1(_1326_),
    .X(_1328_));
 sg13g2_a21oi_1 _5148_ (.A1(net987),
    .A2(_1313_),
    .Y(_1329_),
    .B1(_1017_));
 sg13g2_a21oi_1 _5149_ (.A1(_1328_),
    .A2(_1329_),
    .Y(_1330_),
    .B1(net1071));
 sg13g2_a21oi_1 _5150_ (.A1(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[5] ),
    .A2(_1323_),
    .Y(_1331_),
    .B1(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[6] ));
 sg13g2_and3_1 _5151_ (.X(_1332_),
    .A(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[5] ),
    .B(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[6] ),
    .C(_1323_));
 sg13g2_nor3_1 _5152_ (.A(_1276_),
    .B(_1331_),
    .C(_1332_),
    .Y(_1333_));
 sg13g2_nor2_1 _5153_ (.A(_1330_),
    .B(_1333_),
    .Y(_1334_));
 sg13g2_nor4_1 _5154_ (.A(_1296_),
    .B(_1325_),
    .C(_1330_),
    .D(_1333_),
    .Y(_1335_));
 sg13g2_a21o_1 _5155_ (.A2(_1252_),
    .A1(net985),
    .B1(_1207_),
    .X(_1336_));
 sg13g2_nand3_1 _5156_ (.B(_1256_),
    .C(_1336_),
    .A(net987),
    .Y(_1337_));
 sg13g2_o21ai_1 _5157_ (.B1(_1206_),
    .Y(_1338_),
    .A1(net985),
    .A2(_1252_));
 sg13g2_nand3b_1 _5158_ (.B(_1338_),
    .C(_1107_),
    .Y(_1339_),
    .A_N(_1313_));
 sg13g2_a21oi_1 _5159_ (.A1(_1337_),
    .A2(_1339_),
    .Y(_1340_),
    .B1(_1017_));
 sg13g2_nand3_1 _5160_ (.B(_1309_),
    .C(_1320_),
    .A(_1305_),
    .Y(_1341_));
 sg13g2_nand3_1 _5161_ (.B(_1321_),
    .C(_1341_),
    .A(_1275_),
    .Y(_1342_));
 sg13g2_o21ai_1 _5162_ (.B1(_1342_),
    .Y(_1343_),
    .A1(_1264_),
    .A2(_1340_));
 sg13g2_o21ai_1 _5163_ (.B1(_1326_),
    .Y(_1344_),
    .A1(_1255_),
    .A2(_1316_));
 sg13g2_and2_1 _5164_ (.A(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[7] ),
    .B(_1332_),
    .X(_1345_));
 sg13g2_o21ai_1 _5165_ (.B1(_1275_),
    .Y(_1346_),
    .A1(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[8] ),
    .A2(_1345_));
 sg13g2_a21oi_1 _5166_ (.A1(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[8] ),
    .A2(_1345_),
    .Y(_1347_),
    .B1(_1346_));
 sg13g2_a21oi_2 _5167_ (.B1(_1347_),
    .Y(_1348_),
    .A2(_1344_),
    .A1(_1262_));
 sg13g2_a21oi_1 _5168_ (.A1(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[8] ),
    .A2(_1345_),
    .Y(_1349_),
    .B1(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[0] ));
 sg13g2_nand3_1 _5169_ (.B(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[8] ),
    .C(_1345_),
    .A(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[0] ),
    .Y(_1350_));
 sg13g2_nor2_1 _5170_ (.A(_1276_),
    .B(_1349_),
    .Y(_1351_));
 sg13g2_nor4_1 _5171_ (.A(net987),
    .B(_1208_),
    .C(_1251_),
    .D(_1263_),
    .Y(_1352_));
 sg13g2_a21o_1 _5172_ (.A2(_1351_),
    .A1(_1350_),
    .B1(_1352_),
    .X(_1353_));
 sg13g2_xor2_1 _5173_ (.B(_1350_),
    .A(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[10] ),
    .X(_1354_));
 sg13g2_nor2_1 _5174_ (.A(_1276_),
    .B(_1354_),
    .Y(_1355_));
 sg13g2_nor2_1 _5175_ (.A(_1206_),
    .B(_1327_),
    .Y(_1356_));
 sg13g2_nor2b_1 _5176_ (.A(_1356_),
    .B_N(_1283_),
    .Y(_1357_));
 sg13g2_a21oi_1 _5177_ (.A1(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[5] ),
    .A2(_1323_),
    .Y(_1358_),
    .B1(_1276_));
 sg13g2_o21ai_1 _5178_ (.B1(_1358_),
    .Y(_1359_),
    .A1(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[5] ),
    .A2(_1323_));
 sg13g2_o21ai_1 _5179_ (.B1(_1359_),
    .Y(_1360_),
    .A1(net1073),
    .A2(_1357_));
 sg13g2_or2_1 _5180_ (.X(_1361_),
    .B(_1258_),
    .A(_1207_));
 sg13g2_a22oi_1 _5181_ (.Y(_1362_),
    .B1(_1361_),
    .B2(_1208_),
    .A2(_1259_),
    .A1(net987));
 sg13g2_nor2_1 _5182_ (.A(_1276_),
    .B(_1345_),
    .Y(_1363_));
 sg13g2_o21ai_1 _5183_ (.B1(_1363_),
    .Y(_1364_),
    .A1(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[7] ),
    .A2(_1332_));
 sg13g2_o21ai_1 _5184_ (.B1(_1364_),
    .Y(_1365_),
    .A1(_1263_),
    .A2(_1362_));
 sg13g2_or3_1 _5185_ (.A(_1353_),
    .B(_1355_),
    .C(_1365_),
    .X(_1366_));
 sg13g2_nor4_1 _5186_ (.A(_1279_),
    .B(_1343_),
    .C(_1360_),
    .D(_1366_),
    .Y(_1367_));
 sg13g2_nand4_1 _5187_ (.B(_1335_),
    .C(_1348_),
    .A(_1312_),
    .Y(_1368_),
    .D(_1367_));
 sg13g2_inv_2 _5188_ (.Y(_1369_),
    .A(net983));
 sg13g2_and2_1 _5189_ (.A(_1312_),
    .B(net983),
    .X(_1370_));
 sg13g2_nor2_1 _5190_ (.A(_0057_),
    .B(_1370_),
    .Y(_1371_));
 sg13g2_xnor2_1 _5191_ (.Y(_1372_),
    .A(_0057_),
    .B(_1370_));
 sg13g2_nand2b_1 _5192_ (.Y(_1373_),
    .B(_1372_),
    .A_N(_1300_));
 sg13g2_nand2b_1 _5193_ (.Y(_1374_),
    .B(_1300_),
    .A_N(_1372_));
 sg13g2_and3_1 _5194_ (.X(\i_music.i_sample.t1.genblk1[10].state.D ),
    .A(net1171),
    .B(_1373_),
    .C(_1374_));
 sg13g2_nor2b_1 _5195_ (.A(_1371_),
    .B_N(_1374_),
    .Y(_1375_));
 sg13g2_inv_1 _5196_ (.Y(_1376_),
    .A(_1375_));
 sg13g2_xor2_1 _5197_ (.B(_1343_),
    .A(\i_music.i_sample.thresh[3] ),
    .X(_1377_));
 sg13g2_nor2b_1 _5198_ (.A(_1375_),
    .B_N(_1377_),
    .Y(_1378_));
 sg13g2_o21ai_1 _5199_ (.B1(net1171),
    .Y(_1379_),
    .A1(_1376_),
    .A2(_1377_));
 sg13g2_nor2_2 _5200_ (.A(_1378_),
    .B(_1379_),
    .Y(\i_music.i_sample.t1.genblk1[11].state.D ));
 sg13g2_nor2b_1 _5201_ (.A(_0058_),
    .B_N(_1343_),
    .Y(_1380_));
 sg13g2_xor2_1 _5202_ (.B(_1325_),
    .A(\i_music.i_sample.thresh[4] ),
    .X(_1381_));
 sg13g2_nor3_1 _5203_ (.A(_1378_),
    .B(_1380_),
    .C(_1381_),
    .Y(_1382_));
 sg13g2_o21ai_1 _5204_ (.B1(_1381_),
    .Y(_1383_),
    .A1(_1378_),
    .A2(_1380_));
 sg13g2_inv_1 _5205_ (.Y(_1384_),
    .A(_1383_));
 sg13g2_nor3_2 _5206_ (.A(net1158),
    .B(_1382_),
    .C(_1384_),
    .Y(\i_music.i_sample.t1.genblk1[12].state.D ));
 sg13g2_a21oi_2 _5207_ (.B1(_1384_),
    .Y(_1385_),
    .A2(_1325_),
    .A1(\i_music.i_sample.thresh[4] ));
 sg13g2_xnor2_1 _5208_ (.Y(_1386_),
    .A(\i_music.i_sample.thresh[5] ),
    .B(_1360_));
 sg13g2_o21ai_1 _5209_ (.B1(net1171),
    .Y(_1387_),
    .A1(_1385_),
    .A2(_1386_));
 sg13g2_a21oi_2 _5210_ (.B1(_1387_),
    .Y(\i_music.i_sample.t1.genblk1[13].state.D ),
    .A2(_1386_),
    .A1(_1385_));
 sg13g2_nand2b_1 _5211_ (.Y(_1388_),
    .B(_1360_),
    .A_N(_0059_));
 sg13g2_o21ai_1 _5212_ (.B1(_1388_),
    .Y(_1389_),
    .A1(_1385_),
    .A2(_1386_));
 sg13g2_nor2b_1 _5213_ (.A(_1334_),
    .B_N(\i_music.i_sample.thresh[6] ),
    .Y(_1390_));
 sg13g2_xnor2_1 _5214_ (.Y(_1391_),
    .A(\i_music.i_sample.thresh[6] ),
    .B(_1334_));
 sg13g2_nor2_1 _5215_ (.A(_1389_),
    .B(_1391_),
    .Y(_1392_));
 sg13g2_and2_1 _5216_ (.A(_1389_),
    .B(_1391_),
    .X(_1393_));
 sg13g2_nor3_2 _5217_ (.A(net1155),
    .B(_1392_),
    .C(_1393_),
    .Y(\i_music.i_sample.t1.genblk1[14].state.D ));
 sg13g2_a21oi_1 _5218_ (.A1(_1389_),
    .A2(_1391_),
    .Y(_1394_),
    .B1(_1390_));
 sg13g2_xor2_1 _5219_ (.B(_1365_),
    .A(\i_music.i_sample.thresh[7] ),
    .X(_1395_));
 sg13g2_nor2b_1 _5220_ (.A(_1395_),
    .B_N(_1394_),
    .Y(_1396_));
 sg13g2_nor2b_1 _5221_ (.A(_1394_),
    .B_N(_1395_),
    .Y(_1397_));
 sg13g2_nor3_2 _5222_ (.A(net1155),
    .B(_1396_),
    .C(_1397_),
    .Y(\i_music.i_sample.t1.genblk1[15].state.D ));
 sg13g2_a21oi_1 _5223_ (.A1(\i_music.i_sample.thresh[7] ),
    .A2(_1365_),
    .Y(_1398_),
    .B1(_1397_));
 sg13g2_xnor2_1 _5224_ (.Y(_1399_),
    .A(\i_music.i_sample.thresh[8] ),
    .B(_1348_));
 sg13g2_nand2b_1 _5225_ (.Y(_1400_),
    .B(_1398_),
    .A_N(_1399_));
 sg13g2_nand2b_1 _5226_ (.Y(_1401_),
    .B(_1399_),
    .A_N(_1398_));
 sg13g2_and3_1 _5227_ (.X(\i_music.i_sample.t1.genblk1[16].state.D ),
    .A(net1166),
    .B(_1400_),
    .C(_1401_));
 sg13g2_and2_1 _5228_ (.A(\i_music.i_sample.thresh[9] ),
    .B(_1353_),
    .X(_1402_));
 sg13g2_or2_1 _5229_ (.X(_1403_),
    .B(_1353_),
    .A(\i_music.i_sample.thresh[9] ));
 sg13g2_nor2b_1 _5230_ (.A(_1402_),
    .B_N(_1403_),
    .Y(_1404_));
 sg13g2_o21ai_1 _5231_ (.B1(_1401_),
    .Y(_1405_),
    .A1(_2981_),
    .A2(_1348_));
 sg13g2_o21ai_1 _5232_ (.B1(net1171),
    .Y(_1406_),
    .A1(_1404_),
    .A2(_1405_));
 sg13g2_a21oi_2 _5233_ (.B1(_1406_),
    .Y(\i_music.i_sample.t1.genblk1[17].state.D ),
    .A2(_1405_),
    .A1(_1404_));
 sg13g2_xnor2_1 _5234_ (.Y(_1407_),
    .A(\i_music.i_sample.thresh[10] ),
    .B(_1355_));
 sg13g2_a21oi_1 _5235_ (.A1(_1403_),
    .A2(_1405_),
    .Y(_1408_),
    .B1(_1402_));
 sg13g2_o21ai_1 _5236_ (.B1(net1171),
    .Y(_1409_),
    .A1(_1407_),
    .A2(_1408_));
 sg13g2_a21oi_1 _5237_ (.A1(_1407_),
    .A2(_1408_),
    .Y(\i_music.i_sample.t1.genblk1[18].state.D ),
    .B1(_1409_));
 sg13g2_nor2_1 _5238_ (.A(net1155),
    .B(net374),
    .Y(\i_music.i_sample.t1.genblk1[0].state.D ));
 sg13g2_o21ai_1 _5239_ (.B1(net1166),
    .Y(_1410_),
    .A1(\i_music.i_sample.sample_idx[0] ),
    .A2(\i_music.i_sample.sample_idx[1] ));
 sg13g2_a21oi_2 _5240_ (.B1(_1410_),
    .Y(\i_music.i_sample.t1.genblk1[1].state.D ),
    .A2(net377),
    .A1(net374));
 sg13g2_a21oi_1 _5241_ (.A1(\i_music.i_sample.sample_idx[0] ),
    .A2(\i_music.i_sample.sample_idx[1] ),
    .Y(_1411_),
    .B1(net373));
 sg13g2_nand3_1 _5242_ (.B(\i_music.i_sample.sample_idx[1] ),
    .C(\i_music.i_sample.sample_idx[2] ),
    .A(\i_music.i_sample.sample_idx[0] ),
    .Y(_1412_));
 sg13g2_nand2_1 _5243_ (.Y(_1413_),
    .A(net1166),
    .B(_1412_));
 sg13g2_nor2_1 _5244_ (.A(_1411_),
    .B(_1413_),
    .Y(\i_music.i_sample.t1.genblk1[2].state.D ));
 sg13g2_or2_1 _5245_ (.X(_1414_),
    .B(_1412_),
    .A(_2982_));
 sg13g2_nand2_1 _5246_ (.Y(_1415_),
    .A(net1166),
    .B(_1414_));
 sg13g2_a21oi_2 _5247_ (.B1(_1415_),
    .Y(\i_music.i_sample.t1.genblk1[3].state.D ),
    .A2(_1412_),
    .A1(_2982_));
 sg13g2_and2_1 _5248_ (.A(_2983_),
    .B(_1414_),
    .X(_1416_));
 sg13g2_nor2_2 _5249_ (.A(_2983_),
    .B(_1414_),
    .Y(_1417_));
 sg13g2_nor3_2 _5250_ (.A(net1155),
    .B(_1416_),
    .C(_1417_),
    .Y(\i_music.i_sample.t1.genblk1[4].state.D ));
 sg13g2_xnor2_1 _5251_ (.Y(_1418_),
    .A(\i_music.i_sample.sample_idx[5] ),
    .B(_1417_));
 sg13g2_nor2_1 _5252_ (.A(net1155),
    .B(_1418_),
    .Y(\i_music.i_sample.t1.genblk1[5].state.D ));
 sg13g2_a21oi_1 _5253_ (.A1(\i_music.i_sample.sample_idx[5] ),
    .A2(_1417_),
    .Y(_1419_),
    .B1(net370));
 sg13g2_nand3_1 _5254_ (.B(\i_music.i_sample.sample_idx[6] ),
    .C(_1417_),
    .A(\i_music.i_sample.sample_idx[5] ),
    .Y(_1420_));
 sg13g2_nand2_1 _5255_ (.Y(_1421_),
    .A(net1164),
    .B(_1420_));
 sg13g2_nor2_1 _5256_ (.A(_1419_),
    .B(_1421_),
    .Y(\i_music.i_sample.t1.genblk1[6].state.D ));
 sg13g2_o21ai_1 _5257_ (.B1(net1164),
    .Y(_1422_),
    .A1(_2984_),
    .A2(_1420_));
 sg13g2_a21oi_2 _5258_ (.B1(_1422_),
    .Y(\i_music.i_sample.t1.genblk1[7].state.D ),
    .A2(_1420_),
    .A1(_2984_));
 sg13g2_nor4_1 _5259_ (.A(\i_display.i_vga.timing_ver.counter[9] ),
    .B(\i_display.i_vga.timing_ver.counter[8] ),
    .C(\i_display.i_vga.timing_ver.counter[4] ),
    .D(\i_display.i_vga.timing_ver.counter[2] ),
    .Y(_1423_));
 sg13g2_nor2_1 _5260_ (.A(\i_display.i_vga.timing_ver.counter[7] ),
    .B(\i_display.i_vga.timing_ver.counter[6] ),
    .Y(_1424_));
 sg13g2_nor2_1 _5261_ (.A(net1130),
    .B(\i_display.i_vga.timing_ver.counter[0] ),
    .Y(_1425_));
 sg13g2_nor2_1 _5262_ (.A(\i_display.i_vga.timing_ver.counter[5] ),
    .B(\i_display.i_vga.timing_ver.counter[3] ),
    .Y(_1426_));
 sg13g2_nand4_1 _5263_ (.B(_1424_),
    .C(_1425_),
    .A(_1423_),
    .Y(_1427_),
    .D(_1426_));
 sg13g2_nand2_1 _5264_ (.Y(_1428_),
    .A(\i_display.i_vga.timing_ver.counter[10] ),
    .B(_1427_));
 sg13g2_o21ai_1 _5265_ (.B1(_1428_),
    .Y(\i_display.i_vga.timing_ver.blank ),
    .A1(net207),
    .A2(_1427_));
 sg13g2_nor2_1 _5266_ (.A(\i_display.i_vga.low_count[8] ),
    .B(net1074),
    .Y(_1429_));
 sg13g2_a21oi_1 _5267_ (.A1(_2929_),
    .A2(net1074),
    .Y(_1430_),
    .B1(_1429_));
 sg13g2_nor2_1 _5268_ (.A(\i_music.i_sample.thresh[9] ),
    .B(net1069),
    .Y(_1431_));
 sg13g2_a21oi_1 _5269_ (.A1(_2981_),
    .A2(net1069),
    .Y(_1432_),
    .B1(_1431_));
 sg13g2_nand2b_1 _5270_ (.Y(_1433_),
    .B(_1432_),
    .A_N(_1430_));
 sg13g2_mux2_1 _5271_ (.A0(_0046_),
    .A1(_0063_),
    .S(net1074),
    .X(_1434_));
 sg13g2_mux2_2 _5272_ (.A0(\i_music.i_sample.thresh[6] ),
    .A1(\i_music.i_sample.thresh[7] ),
    .S(net1072),
    .X(_1435_));
 sg13g2_nand2_1 _5273_ (.Y(_1436_),
    .A(_1434_),
    .B(_1435_));
 sg13g2_mux2_1 _5274_ (.A0(_0046_),
    .A1(_0064_),
    .S(net1067),
    .X(_1437_));
 sg13g2_mux2_2 _5275_ (.A0(\i_music.i_sample.thresh[5] ),
    .A1(\i_music.i_sample.thresh[6] ),
    .S(net1072),
    .X(_1438_));
 sg13g2_nand2_1 _5276_ (.Y(_1439_),
    .A(_1437_),
    .B(_1438_));
 sg13g2_xnor2_1 _5277_ (.Y(_1440_),
    .A(_1437_),
    .B(_1438_));
 sg13g2_mux2_1 _5278_ (.A0(_0062_),
    .A1(_0064_),
    .S(net1074),
    .X(_1441_));
 sg13g2_inv_1 _5279_ (.Y(_1442_),
    .A(_1441_));
 sg13g2_mux2_2 _5280_ (.A0(_0059_),
    .A1(_0065_),
    .S(net1068),
    .X(_1443_));
 sg13g2_nor2_1 _5281_ (.A(_1442_),
    .B(_1443_),
    .Y(_1444_));
 sg13g2_mux2_1 _5282_ (.A0(_0062_),
    .A1(_0066_),
    .S(net1069),
    .X(_1445_));
 sg13g2_mux2_1 _5283_ (.A0(_0058_),
    .A1(_0065_),
    .S(net1072),
    .X(_1446_));
 sg13g2_inv_1 _5284_ (.Y(_1447_),
    .A(_1446_));
 sg13g2_nor2_1 _5285_ (.A(_1445_),
    .B(_1447_),
    .Y(_1448_));
 sg13g2_nand2_1 _5286_ (.Y(_1449_),
    .A(_1445_),
    .B(_1447_));
 sg13g2_nor2b_1 _5287_ (.A(_1448_),
    .B_N(_1449_),
    .Y(_1450_));
 sg13g2_mux2_1 _5288_ (.A0(_0061_),
    .A1(_0066_),
    .S(net1074),
    .X(_1451_));
 sg13g2_mux2_2 _5289_ (.A0(_0057_),
    .A1(_0058_),
    .S(net1072),
    .X(_1452_));
 sg13g2_nor2b_1 _5290_ (.A(_1451_),
    .B_N(_1452_),
    .Y(_1453_));
 sg13g2_xnor2_1 _5291_ (.Y(_1454_),
    .A(_1451_),
    .B(_1452_));
 sg13g2_nand2b_1 _5292_ (.Y(_1455_),
    .B(net1068),
    .A_N(_0067_));
 sg13g2_o21ai_1 _5293_ (.B1(_1455_),
    .Y(_1456_),
    .A1(_0061_),
    .A2(net1068));
 sg13g2_mux2_1 _5294_ (.A0(_0056_),
    .A1(_0057_),
    .S(net1072),
    .X(_1457_));
 sg13g2_nor2_1 _5295_ (.A(_1456_),
    .B(_1457_),
    .Y(_1458_));
 sg13g2_nand2_1 _5296_ (.Y(_1459_),
    .A(_1456_),
    .B(_1457_));
 sg13g2_nor2_1 _5297_ (.A(_0056_),
    .B(net1068),
    .Y(_1460_));
 sg13g2_nor2b_1 _5298_ (.A(_0068_),
    .B_N(_0097_),
    .Y(_1461_));
 sg13g2_nor2b_1 _5299_ (.A(net1153),
    .B_N(_0067_),
    .Y(_1462_));
 sg13g2_o21ai_1 _5300_ (.B1(_1462_),
    .Y(_1463_),
    .A1(_1460_),
    .A2(_1461_));
 sg13g2_a21oi_1 _5301_ (.A1(_0097_),
    .A2(_1460_),
    .Y(_1464_),
    .B1(net1081));
 sg13g2_o21ai_1 _5302_ (.B1(_1463_),
    .Y(_1465_),
    .A1(_0068_),
    .A2(_1464_));
 sg13g2_a21oi_1 _5303_ (.A1(_1459_),
    .A2(_1465_),
    .Y(_1466_),
    .B1(_1458_));
 sg13g2_a21o_1 _5304_ (.A2(_1466_),
    .A1(_1454_),
    .B1(_1453_),
    .X(_1467_));
 sg13g2_a221oi_1 _5305_ (.B2(_1467_),
    .C1(_1448_),
    .B1(_1449_),
    .A1(_1442_),
    .Y(_1468_),
    .A2(_1443_));
 sg13g2_or2_1 _5306_ (.X(_1469_),
    .B(_1468_),
    .A(_1444_));
 sg13g2_nor2_1 _5307_ (.A(_1440_),
    .B(_1469_),
    .Y(_1470_));
 sg13g2_or2_1 _5308_ (.X(_1471_),
    .B(_1435_),
    .A(_1434_));
 sg13g2_o21ai_1 _5309_ (.B1(_1471_),
    .Y(_1472_),
    .A1(_1437_),
    .A2(_1438_));
 sg13g2_o21ai_1 _5310_ (.B1(_1436_),
    .Y(_1473_),
    .A1(_1470_),
    .A2(_1472_));
 sg13g2_mux2_1 _5311_ (.A0(_0045_),
    .A1(_0063_),
    .S(net1067),
    .X(_1474_));
 sg13g2_nand2_1 _5312_ (.Y(_1475_),
    .A(\i_music.i_sample.thresh[7] ),
    .B(net1068));
 sg13g2_o21ai_1 _5313_ (.B1(_1475_),
    .Y(_1476_),
    .A1(_2981_),
    .A2(net1067));
 sg13g2_nand2_1 _5314_ (.Y(_1477_),
    .A(_1474_),
    .B(_1476_));
 sg13g2_xnor2_1 _5315_ (.Y(_1478_),
    .A(_1474_),
    .B(_1476_));
 sg13g2_nor2_1 _5316_ (.A(_1473_),
    .B(_1478_),
    .Y(_1479_));
 sg13g2_nand2b_1 _5317_ (.Y(_1480_),
    .B(_1430_),
    .A_N(_1432_));
 sg13g2_o21ai_1 _5318_ (.B1(_1480_),
    .Y(_1481_),
    .A1(_1474_),
    .A2(_1476_));
 sg13g2_o21ai_1 _5319_ (.B1(_1433_),
    .Y(_1482_),
    .A1(_1479_),
    .A2(_1481_));
 sg13g2_a21oi_1 _5320_ (.A1(\i_music.count[10] ),
    .A2(\i_music.i_sample.thresh[10] ),
    .Y(_1483_),
    .B1(net1067));
 sg13g2_o21ai_1 _5321_ (.B1(_1483_),
    .Y(_1484_),
    .A1(\i_music.count[10] ),
    .A2(\i_music.i_sample.thresh[10] ));
 sg13g2_xnor2_1 _5322_ (.Y(_1485_),
    .A(\i_display.i_vga.low_count[9] ),
    .B(\i_music.i_sample.thresh[9] ));
 sg13g2_o21ai_1 _5323_ (.B1(_1484_),
    .Y(_1486_),
    .A1(net1074),
    .A2(_1485_));
 sg13g2_xnor2_1 _5324_ (.Y(_1487_),
    .A(_1482_),
    .B(_1486_));
 sg13g2_xnor2_1 _5325_ (.Y(_1488_),
    .A(_1440_),
    .B(_1469_));
 sg13g2_xor2_1 _5326_ (.B(_1467_),
    .A(_1450_),
    .X(_1489_));
 sg13g2_xnor2_1 _5327_ (.Y(_1490_),
    .A(_1454_),
    .B(_1466_));
 sg13g2_xnor2_1 _5328_ (.Y(_1491_),
    .A(_1441_),
    .B(_1443_));
 sg13g2_xnor2_1 _5329_ (.Y(_1492_),
    .A(_1449_),
    .B(_1491_));
 sg13g2_nand2_1 _5330_ (.Y(_1493_),
    .A(_1433_),
    .B(_1480_));
 sg13g2_xnor2_1 _5331_ (.Y(_1494_),
    .A(_1477_),
    .B(_1493_));
 sg13g2_and2_1 _5332_ (.A(_1436_),
    .B(_1471_),
    .X(_1495_));
 sg13g2_xnor2_1 _5333_ (.Y(_1496_),
    .A(_1439_),
    .B(_1495_));
 sg13g2_nand3_1 _5334_ (.B(_1492_),
    .C(_1496_),
    .A(_1490_),
    .Y(_1497_));
 sg13g2_nor3_1 _5335_ (.A(_1489_),
    .B(_1494_),
    .C(_1497_),
    .Y(_1498_));
 sg13g2_xnor2_1 _5336_ (.Y(_1499_),
    .A(_1473_),
    .B(_1478_));
 sg13g2_nand4_1 _5337_ (.B(_1488_),
    .C(_1498_),
    .A(_1487_),
    .Y(_1500_),
    .D(_1499_));
 sg13g2_a21o_1 _5338_ (.A2(_1500_),
    .A1(net1168),
    .B1(clknet_1_0__leaf_clk),
    .X(_1501_));
 sg13g2_a21oi_1 _5339_ (.A1(net1164),
    .A2(net1068),
    .Y(\i_music.i_sample.t1.CG.GCLK ),
    .B1(clknet_1_1__leaf__1501_));
 sg13g2_a21oi_1 _5340_ (.A1(net1164),
    .A2(_3009_),
    .Y(\i_music.i_sample.t2.CG.GCLK ),
    .B1(clknet_1_0__leaf__1501_));
 sg13g2_a21oi_1 _5341_ (.A1(net1164),
    .A2(net1078),
    .Y(\i_music.i_sample.t3.CG.GCLK ),
    .B1(clknet_1_0__leaf__1501_));
 sg13g2_a21oi_1 _5342_ (.A1(net1168),
    .A2(_2996_),
    .Y(\i_music.i_sample.t4.CG.GCLK ),
    .B1(clknet_1_1__leaf__1501_));
 sg13g2_a21oi_1 _5343_ (.A1(_1032_),
    .A2(_1073_),
    .Y(_1502_),
    .B1(net1015));
 sg13g2_a21o_1 _5344_ (.A2(_1158_),
    .A1(net1014),
    .B1(_1502_),
    .X(_1503_));
 sg13g2_a21oi_1 _5345_ (.A1(net1044),
    .A2(_1503_),
    .Y(_1504_),
    .B1(_1131_));
 sg13g2_nand2_1 _5346_ (.Y(_1505_),
    .A(_1066_),
    .B(_1504_));
 sg13g2_o21ai_1 _5347_ (.B1(_0992_),
    .Y(_1506_),
    .A1(_1102_),
    .A2(_1113_));
 sg13g2_a221oi_1 _5348_ (.B2(_1046_),
    .C1(_1506_),
    .B1(_1184_),
    .A1(_1048_),
    .Y(_1507_),
    .A2(_1122_));
 sg13g2_o21ai_1 _5349_ (.B1(_1192_),
    .Y(_1508_),
    .A1(_1125_),
    .A2(_1175_));
 sg13g2_a22oi_1 _5350_ (.Y(_1509_),
    .B1(_1508_),
    .B2(_1087_),
    .A2(_1236_),
    .A1(net1006));
 sg13g2_a21oi_1 _5351_ (.A1(net1008),
    .A2(_1503_),
    .Y(_1510_),
    .B1(_1130_));
 sg13g2_o21ai_1 _5352_ (.B1(_1505_),
    .Y(_1511_),
    .A1(net1018),
    .A2(_1509_));
 sg13g2_nor4_1 _5353_ (.A(_1008_),
    .B(_1507_),
    .C(_1510_),
    .D(_1511_),
    .Y(_1512_));
 sg13g2_nor3_1 _5354_ (.A(_1102_),
    .B(_1130_),
    .C(_1140_),
    .Y(_1513_));
 sg13g2_nor2_1 _5355_ (.A(_1070_),
    .B(_1513_),
    .Y(_1514_));
 sg13g2_a21oi_2 _5356_ (.B1(_1512_),
    .Y(_1515_),
    .A2(_1514_),
    .A1(_1200_));
 sg13g2_nor2_1 _5357_ (.A(_0035_),
    .B(_1515_),
    .Y(_1516_));
 sg13g2_a21oi_1 _5358_ (.A1(net1010),
    .A2(_1085_),
    .Y(_1517_),
    .B1(_1043_));
 sg13g2_nor2_1 _5359_ (.A(net1018),
    .B(_1172_),
    .Y(_1518_));
 sg13g2_nor2b_1 _5360_ (.A(_1518_),
    .B_N(_1517_),
    .Y(_1519_));
 sg13g2_or2_1 _5361_ (.X(_1520_),
    .B(net1006),
    .A(_1006_));
 sg13g2_o21ai_1 _5362_ (.B1(_1520_),
    .Y(_1521_),
    .A1(net1018),
    .A2(_1517_));
 sg13g2_o21ai_1 _5363_ (.B1(_1004_),
    .Y(_1522_),
    .A1(_1519_),
    .A2(_1521_));
 sg13g2_nor2_1 _5364_ (.A(_1516_),
    .B(_1522_),
    .Y(_1523_));
 sg13g2_nand3_1 _5365_ (.B(_1118_),
    .C(_1515_),
    .A(\i_music.count[24] ),
    .Y(_1524_));
 sg13g2_nor2b_1 _5366_ (.A(\i_music.count[23] ),
    .B_N(_0035_),
    .Y(_1525_));
 sg13g2_a21oi_2 _5367_ (.B1(_1523_),
    .Y(_1526_),
    .A2(_1525_),
    .A1(_1524_));
 sg13g2_or3_2 _5368_ (.A(\i_display.i_vga.low_count[6] ),
    .B(\i_display.i_vga.low_count[5] ),
    .C(\i_display.i_vga.low_count[4] ),
    .X(_1527_));
 sg13g2_nor4_1 _5369_ (.A(\i_display.i_vga.low_count[2] ),
    .B(\i_display.i_vga.low_count[3] ),
    .C(net287),
    .D(\i_music.count[10] ),
    .Y(_1528_));
 sg13g2_nor4_1 _5370_ (.A(\i_display.i_vga.low_count[8] ),
    .B(\i_display.i_vga.low_count[9] ),
    .C(\i_music.count[21] ),
    .D(\i_music.count[20] ),
    .Y(_1529_));
 sg13g2_nor4_1 _5371_ (.A(net300),
    .B(net288),
    .C(\i_music.count[19] ),
    .D(net274),
    .Y(_1530_));
 sg13g2_nor4_1 _5372_ (.A(net273),
    .B(net260),
    .C(net296),
    .D(net293),
    .Y(_1531_));
 sg13g2_nand4_1 _5373_ (.B(_1529_),
    .C(_1530_),
    .A(_1528_),
    .Y(_1532_),
    .D(_1531_));
 sg13g2_nor4_2 _5374_ (.A(net1142),
    .B(_1526_),
    .C(_1527_),
    .Y(_1533_),
    .D(_1532_));
 sg13g2_nand2_1 _5375_ (.Y(_1534_),
    .A(net1081),
    .B(_1533_));
 sg13g2_nand2_1 _5376_ (.Y(_1535_),
    .A(net1170),
    .B(_1534_));
 sg13g2_nor2_1 _5377_ (.A(net1169),
    .B(_2985_),
    .Y(_1536_));
 sg13g2_nor2_1 _5378_ (.A(\i_music.violin_note_idx[1][2] ),
    .B(\i_music.violin_note_idx[1][4] ),
    .Y(_1537_));
 sg13g2_nand3_1 _5379_ (.B(\i_music.violin_note_idx[1][8] ),
    .C(_1537_),
    .A(\i_music.violin_note_idx[1][5] ),
    .Y(_1538_));
 sg13g2_nand2_1 _5380_ (.Y(_1539_),
    .A(\i_music.violin_note_idx[1][7] ),
    .B(\i_music.violin_note_idx[1][6] ));
 sg13g2_nand2_1 _5381_ (.Y(_1540_),
    .A(\i_music.violin_note_idx[1][0] ),
    .B(\i_music.violin_note_idx[1][3] ));
 sg13g2_nor4_2 _5382_ (.A(\i_music.violin_note_idx[1][1] ),
    .B(_1538_),
    .C(_1539_),
    .Y(_1541_),
    .D(_1540_));
 sg13g2_or2_1 _5383_ (.X(_1542_),
    .B(\i_music.violin_note_idx[1][0] ),
    .A(net328));
 sg13g2_nor4_1 _5384_ (.A(\i_music.violin_note_idx[1][3] ),
    .B(\i_music.violin_note_idx[1][7] ),
    .C(\i_music.violin_note_idx[1][6] ),
    .D(_1542_),
    .Y(_1543_));
 sg13g2_nand2b_2 _5385_ (.Y(_1544_),
    .B(_1543_),
    .A_N(_1538_));
 sg13g2_inv_1 _5386_ (.Y(_1545_),
    .A(_1544_));
 sg13g2_nor2_2 _5387_ (.A(net1157),
    .B(_1545_),
    .Y(_1546_));
 sg13g2_nand2_2 _5388_ (.Y(_1547_),
    .A(net1169),
    .B(_1544_));
 sg13g2_nor2_1 _5389_ (.A(net1156),
    .B(_1541_),
    .Y(_1548_));
 sg13g2_nand2_2 _5390_ (.Y(_1549_),
    .A(\i_music.violin_note_idx[2][0] ),
    .B(net250));
 sg13g2_nor3_2 _5391_ (.A(_2950_),
    .B(_2958_),
    .C(_1549_),
    .Y(_1550_));
 sg13g2_xnor2_1 _5392_ (.Y(_1551_),
    .A(net311),
    .B(_1550_));
 sg13g2_nor3_1 _5393_ (.A(_1541_),
    .B(_1547_),
    .C(_1551_),
    .Y(_1552_));
 sg13g2_a21oi_1 _5394_ (.A1(net979),
    .A2(_1552_),
    .Y(_1553_),
    .B1(_1536_));
 sg13g2_o21ai_1 _5395_ (.B1(_1553_),
    .Y(_0101_),
    .A1(_2952_),
    .A2(net978));
 sg13g2_nor2_2 _5396_ (.A(net1170),
    .B(net2),
    .Y(_1554_));
 sg13g2_and3_1 _5397_ (.X(_1555_),
    .A(\i_music.violin_note_idx[2][5] ),
    .B(\i_music.violin_note_idx[2][4] ),
    .C(_1550_));
 sg13g2_a21oi_1 _5398_ (.A1(\i_music.violin_note_idx[2][4] ),
    .A2(_1550_),
    .Y(_1556_),
    .B1(\i_music.violin_note_idx[2][5] ));
 sg13g2_nor2_2 _5399_ (.A(_1541_),
    .B(_1545_),
    .Y(_1557_));
 sg13g2_o21ai_1 _5400_ (.B1(_1557_),
    .Y(_1558_),
    .A1(_1555_),
    .A2(_1556_));
 sg13g2_a21oi_1 _5401_ (.A1(net1170),
    .A2(_1558_),
    .Y(_1559_),
    .B1(_1554_));
 sg13g2_nor2_1 _5402_ (.A(net303),
    .B(net978),
    .Y(_1560_));
 sg13g2_a21oi_1 _5403_ (.A1(net978),
    .A2(_1559_),
    .Y(_0102_),
    .B1(_1560_));
 sg13g2_a21oi_2 _5404_ (.B1(_1554_),
    .Y(_1561_),
    .A2(_1541_),
    .A1(net1169));
 sg13g2_and2_1 _5405_ (.A(\i_music.violin_note_idx[2][6] ),
    .B(_1555_),
    .X(_1562_));
 sg13g2_o21ai_1 _5406_ (.B1(_1546_),
    .Y(_1563_),
    .A1(\i_music.violin_note_idx[2][6] ),
    .A2(_1555_));
 sg13g2_o21ai_1 _5407_ (.B1(_1561_),
    .Y(_1564_),
    .A1(_1562_),
    .A2(_1563_));
 sg13g2_mux2_1 _5408_ (.A0(net249),
    .A1(_1564_),
    .S(net979),
    .X(_0103_));
 sg13g2_nand2_1 _5409_ (.Y(_1565_),
    .A(\i_music.violin_note_idx[2][7] ),
    .B(_1562_));
 sg13g2_nor2_1 _5410_ (.A(\i_music.violin_note_idx[2][7] ),
    .B(_1562_),
    .Y(_1566_));
 sg13g2_nand2_1 _5411_ (.Y(_1567_),
    .A(_1546_),
    .B(_1565_));
 sg13g2_o21ai_1 _5412_ (.B1(_1561_),
    .Y(_1568_),
    .A1(_1566_),
    .A2(_1567_));
 sg13g2_mux2_1 _5413_ (.A0(net276),
    .A1(_1568_),
    .S(net979),
    .X(_0104_));
 sg13g2_o21ai_1 _5414_ (.B1(_1557_),
    .Y(_1569_),
    .A1(\i_music.violin_note_idx[2][8] ),
    .A2(_1565_));
 sg13g2_a21o_1 _5415_ (.A2(_1565_),
    .A1(net236),
    .B1(_1569_),
    .X(_1570_));
 sg13g2_a21oi_1 _5416_ (.A1(net1169),
    .A2(_1570_),
    .Y(_1571_),
    .B1(_1554_));
 sg13g2_nor2_1 _5417_ (.A(net236),
    .B(net979),
    .Y(_1572_));
 sg13g2_a21oi_1 _5418_ (.A1(net979),
    .A2(_1571_),
    .Y(_0105_),
    .B1(_1572_));
 sg13g2_nand3_1 _5419_ (.B(_2996_),
    .C(net1067),
    .A(net1164),
    .Y(_1573_));
 sg13g2_inv_2 _5420_ (.Y(_0136_),
    .A(_1573_));
 sg13g2_nor2_1 _5421_ (.A(\i_music.i_sample.t3.genblk1[6].state.Q ),
    .B(net1078),
    .Y(_1574_));
 sg13g2_a21oi_1 _5422_ (.A1(_3027_),
    .A2(net1078),
    .Y(_1575_),
    .B1(_1574_));
 sg13g2_a21o_2 _5423_ (.A2(net1078),
    .A1(_3027_),
    .B1(_1574_),
    .X(_1576_));
 sg13g2_nor2_1 _5424_ (.A(\i_music.i_sample.t3.genblk1[5].state.Q ),
    .B(net1077),
    .Y(_1577_));
 sg13g2_a21oi_1 _5425_ (.A1(_3024_),
    .A2(net1077),
    .Y(_1578_),
    .B1(_1577_));
 sg13g2_a21o_1 _5426_ (.A2(net1077),
    .A1(_3024_),
    .B1(_1577_),
    .X(_1579_));
 sg13g2_nor2_2 _5427_ (.A(_1576_),
    .B(net928),
    .Y(_1580_));
 sg13g2_nand2_2 _5428_ (.Y(_1581_),
    .A(net931),
    .B(net930));
 sg13g2_nor2_1 _5429_ (.A(\i_music.i_sample.t3.genblk1[1].state.Q ),
    .B(net1076),
    .Y(_1582_));
 sg13g2_a21oi_2 _5430_ (.B1(_1582_),
    .Y(_1583_),
    .A2(net1075),
    .A1(_3012_));
 sg13g2_a21o_1 _5431_ (.A2(net1075),
    .A1(_3012_),
    .B1(_1582_),
    .X(_1584_));
 sg13g2_nor2_1 _5432_ (.A(\i_music.i_sample.t3.genblk1[2].state.Q ),
    .B(net1076),
    .Y(_1585_));
 sg13g2_a21oi_1 _5433_ (.A1(_3015_),
    .A2(net1075),
    .Y(_1586_),
    .B1(_1585_));
 sg13g2_a21o_1 _5434_ (.A2(net1075),
    .A1(_3015_),
    .B1(_1585_),
    .X(_1587_));
 sg13g2_nor2_2 _5435_ (.A(net925),
    .B(net921),
    .Y(_1588_));
 sg13g2_nand2_2 _5436_ (.Y(_1589_),
    .A(net926),
    .B(net923));
 sg13g2_nor2_1 _5437_ (.A(\i_music.i_sample.t3.genblk1[3].state.Q ),
    .B(net1076),
    .Y(_1590_));
 sg13g2_a21oi_2 _5438_ (.B1(_1590_),
    .Y(_1591_),
    .A2(net1075),
    .A1(_3018_));
 sg13g2_a21o_1 _5439_ (.A2(net1075),
    .A1(_3018_),
    .B1(_1590_),
    .X(_1592_));
 sg13g2_nor2_2 _5440_ (.A(_1588_),
    .B(net920),
    .Y(_1593_));
 sg13g2_nor2_1 _5441_ (.A(\i_music.i_sample.t3.genblk1[4].state.Q ),
    .B(net1076),
    .Y(_1594_));
 sg13g2_a21oi_1 _5442_ (.A1(_3021_),
    .A2(net1076),
    .Y(_1595_),
    .B1(_1594_));
 sg13g2_a21o_1 _5443_ (.A2(net1075),
    .A1(_3021_),
    .B1(_1594_),
    .X(_1596_));
 sg13g2_xnor2_1 _5444_ (.Y(_1597_),
    .A(_1593_),
    .B(net906));
 sg13g2_nand2_1 _5445_ (.Y(_1598_),
    .A(_3030_),
    .B(net1078));
 sg13g2_o21ai_1 _5446_ (.B1(_1598_),
    .Y(_1599_),
    .A1(\i_music.i_sample.t3.genblk1[7].state.Q ),
    .A2(net1078));
 sg13g2_inv_2 _5447_ (.Y(_1600_),
    .A(_1599_));
 sg13g2_o21ai_1 _5448_ (.B1(_1600_),
    .Y(_1601_),
    .A1(_1581_),
    .A2(_1597_));
 sg13g2_nor2_1 _5449_ (.A(net920),
    .B(net912),
    .Y(_1602_));
 sg13g2_nand2_1 _5450_ (.Y(_1603_),
    .A(net922),
    .B(net906));
 sg13g2_nand2_2 _5451_ (.Y(_1604_),
    .A(net924),
    .B(net919));
 sg13g2_nand2_1 _5452_ (.Y(_1605_),
    .A(net907),
    .B(_1604_));
 sg13g2_nor2_1 _5453_ (.A(\i_music.i_sample.t3.genblk1[0].state.Q ),
    .B(net1076),
    .Y(_1606_));
 sg13g2_a21oi_1 _5454_ (.A1(_3007_),
    .A2(net1075),
    .Y(_1607_),
    .B1(_1606_));
 sg13g2_a21o_1 _5455_ (.A2(net1076),
    .A1(_3007_),
    .B1(_1606_),
    .X(_1608_));
 sg13g2_nor2_2 _5456_ (.A(net926),
    .B(net903),
    .Y(_1609_));
 sg13g2_nand2_1 _5457_ (.Y(_1610_),
    .A(net925),
    .B(net902));
 sg13g2_nor2_2 _5458_ (.A(net914),
    .B(_1609_),
    .Y(_1611_));
 sg13g2_nor2_2 _5459_ (.A(net926),
    .B(net923),
    .Y(_1612_));
 sg13g2_nand2_2 _5460_ (.Y(_1613_),
    .A(net925),
    .B(net921));
 sg13g2_o21ai_1 _5461_ (.B1(net920),
    .Y(_1614_),
    .A1(net924),
    .A2(_1610_));
 sg13g2_nand3_1 _5462_ (.B(net906),
    .C(_1614_),
    .A(net931),
    .Y(_1615_));
 sg13g2_nand2_2 _5463_ (.Y(_1616_),
    .A(_1576_),
    .B(net927));
 sg13g2_nor2_2 _5464_ (.A(_1576_),
    .B(net929),
    .Y(_1617_));
 sg13g2_nand2_2 _5465_ (.Y(_1618_),
    .A(net931),
    .B(net928));
 sg13g2_nand2_1 _5466_ (.Y(_1619_),
    .A(_1615_),
    .B(_1618_));
 sg13g2_nor2_2 _5467_ (.A(net931),
    .B(net928),
    .Y(_1620_));
 sg13g2_nor2_1 _5468_ (.A(_1600_),
    .B(_1620_),
    .Y(_1621_));
 sg13g2_o21ai_1 _5469_ (.B1(_1621_),
    .Y(_1622_),
    .A1(net931),
    .A2(_1602_));
 sg13g2_o21ai_1 _5470_ (.B1(_1601_),
    .Y(_1623_),
    .A1(_1619_),
    .A2(_1622_));
 sg13g2_nand2_1 _5471_ (.Y(_1624_),
    .A(net983),
    .B(_1623_));
 sg13g2_nor2_2 _5472_ (.A(net923),
    .B(net903),
    .Y(_1625_));
 sg13g2_nand2_1 _5473_ (.Y(_1626_),
    .A(net926),
    .B(net916));
 sg13g2_nand2_1 _5474_ (.Y(_1627_),
    .A(_1591_),
    .B(_1613_));
 sg13g2_nor2_2 _5475_ (.A(net925),
    .B(net902),
    .Y(_1628_));
 sg13g2_nand2_1 _5476_ (.Y(_1629_),
    .A(net926),
    .B(net903));
 sg13g2_nor2_2 _5477_ (.A(net924),
    .B(net900),
    .Y(_1630_));
 sg13g2_o21ai_1 _5478_ (.B1(net920),
    .Y(_1631_),
    .A1(net924),
    .A2(_1628_));
 sg13g2_or2_1 _5479_ (.X(_1632_),
    .B(_1631_),
    .A(net906));
 sg13g2_nand3_1 _5480_ (.B(_1597_),
    .C(_1632_),
    .A(_1580_),
    .Y(_1633_));
 sg13g2_nand2_1 _5481_ (.Y(_1634_),
    .A(net922),
    .B(net913));
 sg13g2_a21oi_2 _5482_ (.B1(net906),
    .Y(_1635_),
    .A2(_1612_),
    .A1(net913));
 sg13g2_a21oi_1 _5483_ (.A1(_1588_),
    .A2(net920),
    .Y(_1636_),
    .B1(net912));
 sg13g2_o21ai_1 _5484_ (.B1(_1617_),
    .Y(_1637_),
    .A1(_1635_),
    .A2(_1636_));
 sg13g2_nand3_1 _5485_ (.B(net908),
    .C(_1627_),
    .A(net930),
    .Y(_1638_));
 sg13g2_nor2_1 _5486_ (.A(net908),
    .B(_1604_),
    .Y(_1639_));
 sg13g2_nor2_1 _5487_ (.A(net931),
    .B(_1639_),
    .Y(_1640_));
 sg13g2_nand2_1 _5488_ (.Y(_1641_),
    .A(_1638_),
    .B(_1640_));
 sg13g2_a21oi_1 _5489_ (.A1(_1620_),
    .A2(_1638_),
    .Y(_1642_),
    .B1(net901));
 sg13g2_nand4_1 _5490_ (.B(_1637_),
    .C(_1641_),
    .A(_1633_),
    .Y(_1643_),
    .D(_1642_));
 sg13g2_nand2_1 _5491_ (.Y(_1644_),
    .A(net907),
    .B(_1631_));
 sg13g2_nand3_1 _5492_ (.B(_1632_),
    .C(_1644_),
    .A(net928),
    .Y(_1645_));
 sg13g2_nand3_1 _5493_ (.B(_1632_),
    .C(_1638_),
    .A(_1603_),
    .Y(_1646_));
 sg13g2_a22oi_1 _5494_ (.Y(_1647_),
    .B1(_1646_),
    .B2(_1576_),
    .A2(_1645_),
    .A1(_1619_));
 sg13g2_o21ai_1 _5495_ (.B1(_1643_),
    .Y(_1648_),
    .A1(_1600_),
    .A2(_1647_));
 sg13g2_nand2b_1 _5496_ (.Y(_1649_),
    .B(net982),
    .A_N(_1648_));
 sg13g2_nor2_1 _5497_ (.A(_0055_),
    .B(_1649_),
    .Y(_1650_));
 sg13g2_xor2_1 _5498_ (.B(_1649_),
    .A(_0055_),
    .X(_1651_));
 sg13g2_nor2_2 _5499_ (.A(_1584_),
    .B(_1607_),
    .Y(_1652_));
 sg13g2_nand2_2 _5500_ (.Y(_1653_),
    .A(_1583_),
    .B(net902));
 sg13g2_nor2_2 _5501_ (.A(net921),
    .B(net902),
    .Y(_1654_));
 sg13g2_nand2_2 _5502_ (.Y(_1655_),
    .A(net923),
    .B(net903));
 sg13g2_nand2_1 _5503_ (.Y(_1656_),
    .A(_1653_),
    .B(_1655_));
 sg13g2_nor2_1 _5504_ (.A(_1612_),
    .B(_1656_),
    .Y(_1657_));
 sg13g2_o21ai_1 _5505_ (.B1(net905),
    .Y(_1658_),
    .A1(net913),
    .A2(_1657_));
 sg13g2_nor2_2 _5506_ (.A(_1583_),
    .B(net921),
    .Y(_1659_));
 sg13g2_nor2_2 _5507_ (.A(net921),
    .B(net903),
    .Y(_1660_));
 sg13g2_nor2_1 _5508_ (.A(net914),
    .B(_1660_),
    .Y(_1661_));
 sg13g2_nand3b_1 _5509_ (.B(_1661_),
    .C(net910),
    .Y(_1662_),
    .A_N(_1659_));
 sg13g2_o21ai_1 _5510_ (.B1(net927),
    .Y(_1663_),
    .A1(_1657_),
    .A2(_1662_));
 sg13g2_nand2b_1 _5511_ (.Y(_1664_),
    .B(_1658_),
    .A_N(_1663_));
 sg13g2_nand2_2 _5512_ (.Y(_1665_),
    .A(net926),
    .B(net921));
 sg13g2_nor2_2 _5513_ (.A(_1584_),
    .B(net917),
    .Y(_1666_));
 sg13g2_nor2_1 _5514_ (.A(net911),
    .B(_1666_),
    .Y(_1667_));
 sg13g2_a22oi_1 _5515_ (.Y(_1668_),
    .B1(_1665_),
    .B2(_1667_),
    .A2(_1635_),
    .A1(_1631_));
 sg13g2_nor2_2 _5516_ (.A(net919),
    .B(_1652_),
    .Y(_1669_));
 sg13g2_nor2_2 _5517_ (.A(_1588_),
    .B(_1612_),
    .Y(_1670_));
 sg13g2_o21ai_1 _5518_ (.B1(_1669_),
    .Y(_1671_),
    .A1(_1588_),
    .A2(_1612_));
 sg13g2_a21oi_2 _5519_ (.B1(net908),
    .Y(_1672_),
    .A2(_1630_),
    .A1(net919));
 sg13g2_and2_1 _5520_ (.A(_1671_),
    .B(_1672_),
    .X(_1673_));
 sg13g2_o21ai_1 _5521_ (.B1(_1673_),
    .Y(_1674_),
    .A1(_1589_),
    .A2(net915));
 sg13g2_nand3_1 _5522_ (.B(_1620_),
    .C(_1674_),
    .A(_1605_),
    .Y(_1675_));
 sg13g2_o21ai_1 _5523_ (.B1(_1675_),
    .Y(_1676_),
    .A1(_1616_),
    .A2(_1668_));
 sg13g2_a21oi_1 _5524_ (.A1(_1619_),
    .A2(_1664_),
    .Y(_1677_),
    .B1(_1676_));
 sg13g2_nand2_1 _5525_ (.Y(_1678_),
    .A(_1593_),
    .B(_1655_));
 sg13g2_nand3_1 _5526_ (.B(net912),
    .C(_1655_),
    .A(_1593_),
    .Y(_1679_));
 sg13g2_o21ai_1 _5527_ (.B1(_1679_),
    .Y(_1680_),
    .A1(net920),
    .A2(_1613_));
 sg13g2_a21oi_1 _5528_ (.A1(_1602_),
    .A2(_1612_),
    .Y(_1681_),
    .B1(net930));
 sg13g2_a21oi_1 _5529_ (.A1(net928),
    .A2(_1680_),
    .Y(_1682_),
    .B1(_1641_));
 sg13g2_nand2_2 _5530_ (.Y(_1683_),
    .A(_1589_),
    .B(net917));
 sg13g2_nor2_2 _5531_ (.A(net921),
    .B(net916),
    .Y(_1684_));
 sg13g2_nand2_1 _5532_ (.Y(_1685_),
    .A(net923),
    .B(net914));
 sg13g2_o21ai_1 _5533_ (.B1(_1683_),
    .Y(_1686_),
    .A1(_1629_),
    .A2(_1685_));
 sg13g2_a22oi_1 _5534_ (.Y(_1687_),
    .B1(_1686_),
    .B2(net907),
    .A2(_1635_),
    .A1(_1627_));
 sg13g2_nor2_1 _5535_ (.A(_1618_),
    .B(_1687_),
    .Y(_1688_));
 sg13g2_nand2_1 _5536_ (.Y(_1689_),
    .A(net922),
    .B(net900));
 sg13g2_nand3_1 _5537_ (.B(_1611_),
    .C(_1689_),
    .A(_1580_),
    .Y(_1690_));
 sg13g2_nor3_1 _5538_ (.A(_1601_),
    .B(_1682_),
    .C(_1688_),
    .Y(_1691_));
 sg13g2_a22oi_1 _5539_ (.Y(_1692_),
    .B1(_1690_),
    .B2(_1691_),
    .A2(_1677_),
    .A1(net901));
 sg13g2_nor2_1 _5540_ (.A(_1369_),
    .B(_1692_),
    .Y(_1693_));
 sg13g2_nand2_1 _5541_ (.Y(_1694_),
    .A(\i_music.i_sample.sample_acc[4] ),
    .B(_1693_));
 sg13g2_nor2_1 _5542_ (.A(net926),
    .B(net902),
    .Y(_1695_));
 sg13g2_nand2_1 _5543_ (.Y(_1696_),
    .A(net925),
    .B(net903));
 sg13g2_nand2_1 _5544_ (.Y(_1697_),
    .A(net919),
    .B(_1696_));
 sg13g2_inv_1 _5545_ (.Y(_1698_),
    .A(_1697_));
 sg13g2_o21ai_1 _5546_ (.B1(_1635_),
    .Y(_1699_),
    .A1(_1669_),
    .A2(_1698_));
 sg13g2_o21ai_1 _5547_ (.B1(_1699_),
    .Y(_1700_),
    .A1(_1593_),
    .A2(_1644_));
 sg13g2_o21ai_1 _5548_ (.B1(net906),
    .Y(_1701_),
    .A1(_1593_),
    .A2(_1670_));
 sg13g2_nand2_2 _5549_ (.Y(_1702_),
    .A(net918),
    .B(_1654_));
 sg13g2_nor3_2 _5550_ (.A(net917),
    .B(net909),
    .C(net903),
    .Y(_1703_));
 sg13g2_a21oi_1 _5551_ (.A1(_1670_),
    .A2(_1702_),
    .Y(_1704_),
    .B1(_1703_));
 sg13g2_a21oi_1 _5552_ (.A1(_1701_),
    .A2(_1704_),
    .Y(_1705_),
    .B1(_1618_));
 sg13g2_nor2_1 _5553_ (.A(net924),
    .B(_1609_),
    .Y(_1706_));
 sg13g2_a21oi_1 _5554_ (.A1(net913),
    .A2(_1609_),
    .Y(_1707_),
    .B1(_1706_));
 sg13g2_o21ai_1 _5555_ (.B1(_1681_),
    .Y(_1708_),
    .A1(net906),
    .A2(_1707_));
 sg13g2_nor2_1 _5556_ (.A(net928),
    .B(_1639_),
    .Y(_1709_));
 sg13g2_a21oi_1 _5557_ (.A1(_1701_),
    .A2(_1709_),
    .Y(_1710_),
    .B1(net931));
 sg13g2_a221oi_1 _5558_ (.B2(_1710_),
    .C1(_1705_),
    .B1(_1708_),
    .A1(_1580_),
    .Y(_1711_),
    .A2(_1700_));
 sg13g2_nor2_1 _5559_ (.A(net901),
    .B(_1711_),
    .Y(_1712_));
 sg13g2_nor2_2 _5560_ (.A(_1609_),
    .B(net900),
    .Y(_1713_));
 sg13g2_inv_1 _5561_ (.Y(_1714_),
    .A(_1713_));
 sg13g2_nor2_1 _5562_ (.A(net923),
    .B(_1713_),
    .Y(_1715_));
 sg13g2_a21oi_2 _5563_ (.B1(_1630_),
    .Y(_1716_),
    .A2(_1714_),
    .A1(net924));
 sg13g2_a21oi_1 _5564_ (.A1(net922),
    .A2(_1609_),
    .Y(_1717_),
    .B1(_1716_));
 sg13g2_inv_1 _5565_ (.Y(_1718_),
    .A(_1717_));
 sg13g2_o21ai_1 _5566_ (.B1(_1678_),
    .Y(_1719_),
    .A1(net913),
    .A2(_1717_));
 sg13g2_o21ai_1 _5567_ (.B1(net912),
    .Y(_1720_),
    .A1(net913),
    .A2(_1713_));
 sg13g2_o21ai_1 _5568_ (.B1(_1617_),
    .Y(_1721_),
    .A1(_1593_),
    .A2(_1720_));
 sg13g2_a21oi_1 _5569_ (.A1(net906),
    .A2(_1719_),
    .Y(_1722_),
    .B1(_1721_));
 sg13g2_nand2_1 _5570_ (.Y(_1723_),
    .A(net923),
    .B(net900));
 sg13g2_nor2_1 _5571_ (.A(net916),
    .B(_1612_),
    .Y(_1724_));
 sg13g2_a21oi_1 _5572_ (.A1(_1723_),
    .A2(_1724_),
    .Y(_1725_),
    .B1(net904));
 sg13g2_o21ai_1 _5573_ (.B1(_1725_),
    .Y(_1726_),
    .A1(_1683_),
    .A2(_1715_));
 sg13g2_nor2_1 _5574_ (.A(net909),
    .B(_1626_),
    .Y(_1727_));
 sg13g2_nand2_1 _5575_ (.Y(_1728_),
    .A(net903),
    .B(_1727_));
 sg13g2_a21oi_1 _5576_ (.A1(net915),
    .A2(_1630_),
    .Y(_1729_),
    .B1(net912));
 sg13g2_a221oi_1 _5577_ (.B2(_1614_),
    .C1(_1581_),
    .B1(_1729_),
    .A1(net900),
    .Y(_1730_),
    .A2(_1639_));
 sg13g2_nor3_1 _5578_ (.A(net929),
    .B(_1625_),
    .C(_1659_),
    .Y(_1731_));
 sg13g2_a21oi_1 _5579_ (.A1(net913),
    .A2(_1608_),
    .Y(_1732_),
    .B1(net911));
 sg13g2_a21oi_1 _5580_ (.A1(_1726_),
    .A2(_1728_),
    .Y(_1733_),
    .B1(net927));
 sg13g2_a221oi_1 _5581_ (.B2(_1732_),
    .C1(_1733_),
    .B1(_1731_),
    .A1(net927),
    .Y(_1734_),
    .A2(_1673_));
 sg13g2_nor2_1 _5582_ (.A(net932),
    .B(_1734_),
    .Y(_1735_));
 sg13g2_nor4_1 _5583_ (.A(_1600_),
    .B(_1722_),
    .C(_1730_),
    .D(_1735_),
    .Y(_1736_));
 sg13g2_nor3_1 _5584_ (.A(_1369_),
    .B(_1712_),
    .C(_1736_),
    .Y(_1737_));
 sg13g2_nand2_1 _5585_ (.Y(_1738_),
    .A(_1604_),
    .B(_1697_));
 sg13g2_o21ai_1 _5586_ (.B1(_1738_),
    .Y(_1739_),
    .A1(net922),
    .A2(_1653_));
 sg13g2_nor2_1 _5587_ (.A(net916),
    .B(_1655_),
    .Y(_1740_));
 sg13g2_nand2_2 _5588_ (.Y(_1741_),
    .A(net914),
    .B(_1654_));
 sg13g2_nand3_1 _5589_ (.B(_1739_),
    .C(_1741_),
    .A(_1729_),
    .Y(_1742_));
 sg13g2_nor3_1 _5590_ (.A(net919),
    .B(_1628_),
    .C(_1670_),
    .Y(_1743_));
 sg13g2_a21oi_1 _5591_ (.A1(_1589_),
    .A2(_1653_),
    .Y(_1744_),
    .B1(net915));
 sg13g2_o21ai_1 _5592_ (.B1(net911),
    .Y(_1745_),
    .A1(_1743_),
    .A2(_1744_));
 sg13g2_nand3_1 _5593_ (.B(_1742_),
    .C(_1745_),
    .A(net927),
    .Y(_1746_));
 sg13g2_o21ai_1 _5594_ (.B1(_1661_),
    .Y(_1747_),
    .A1(net902),
    .A2(_1613_));
 sg13g2_and2_1 _5595_ (.A(_1725_),
    .B(_1747_),
    .X(_1748_));
 sg13g2_nor2_1 _5596_ (.A(_1627_),
    .B(_1652_),
    .Y(_1749_));
 sg13g2_nor3_1 _5597_ (.A(net911),
    .B(_1684_),
    .C(_1749_),
    .Y(_1750_));
 sg13g2_o21ai_1 _5598_ (.B1(net929),
    .Y(_1751_),
    .A1(_1748_),
    .A2(_1750_));
 sg13g2_nand3_1 _5599_ (.B(_1746_),
    .C(_1751_),
    .A(_1576_),
    .Y(_1752_));
 sg13g2_a21oi_1 _5600_ (.A1(_1684_),
    .A2(_1713_),
    .Y(_1753_),
    .B1(net910));
 sg13g2_nand2_1 _5601_ (.Y(_1754_),
    .A(net921),
    .B(_1666_));
 sg13g2_nand3_1 _5602_ (.B(_1753_),
    .C(_1754_),
    .A(_1702_),
    .Y(_1755_));
 sg13g2_a21oi_1 _5603_ (.A1(net916),
    .A2(_1660_),
    .Y(_1756_),
    .B1(net904));
 sg13g2_a21oi_1 _5604_ (.A1(_1741_),
    .A2(_1756_),
    .Y(_1757_),
    .B1(_1618_));
 sg13g2_a21oi_2 _5605_ (.B1(net910),
    .Y(_1758_),
    .A2(_1609_),
    .A1(net914));
 sg13g2_o21ai_1 _5606_ (.B1(net904),
    .Y(_1759_),
    .A1(net916),
    .A2(_1610_));
 sg13g2_o21ai_1 _5607_ (.B1(_1706_),
    .Y(_1760_),
    .A1(net920),
    .A2(net900));
 sg13g2_a21oi_1 _5608_ (.A1(_1604_),
    .A2(_1634_),
    .Y(_1761_),
    .B1(_1720_));
 sg13g2_a21o_1 _5609_ (.A2(_1760_),
    .A1(_1758_),
    .B1(_1761_),
    .X(_1762_));
 sg13g2_a22oi_1 _5610_ (.Y(_1763_),
    .B1(_1762_),
    .B2(_1580_),
    .A2(_1757_),
    .A1(_1755_));
 sg13g2_nand3_1 _5611_ (.B(_1752_),
    .C(_1763_),
    .A(net901),
    .Y(_1764_));
 sg13g2_nor3_1 _5612_ (.A(net907),
    .B(_1659_),
    .C(_1697_),
    .Y(_1765_));
 sg13g2_nor2b_1 _5613_ (.A(_1605_),
    .B_N(_1754_),
    .Y(_1766_));
 sg13g2_nor3_1 _5614_ (.A(net930),
    .B(_1765_),
    .C(_1766_),
    .Y(_1767_));
 sg13g2_nand3_1 _5615_ (.B(net904),
    .C(_1626_),
    .A(_1589_),
    .Y(_1768_));
 sg13g2_nand2_1 _5616_ (.Y(_1769_),
    .A(_1662_),
    .B(_1768_));
 sg13g2_a221oi_1 _5617_ (.B2(net929),
    .C1(net932),
    .B1(_1769_),
    .A1(_1679_),
    .Y(_1770_),
    .A2(_1767_));
 sg13g2_nor2_1 _5618_ (.A(net919),
    .B(_1696_),
    .Y(_1771_));
 sg13g2_and2_1 _5619_ (.A(_1669_),
    .B(_1670_),
    .X(_1772_));
 sg13g2_nor2_1 _5620_ (.A(_1656_),
    .B(_1772_),
    .Y(_1773_));
 sg13g2_a21oi_1 _5621_ (.A1(_1684_),
    .A2(_1695_),
    .Y(_1774_),
    .B1(_1773_));
 sg13g2_o21ai_1 _5622_ (.B1(_1753_),
    .Y(_1775_),
    .A1(_1625_),
    .A2(_1683_));
 sg13g2_o21ai_1 _5623_ (.B1(_1775_),
    .Y(_1776_),
    .A1(net904),
    .A2(_1774_));
 sg13g2_a21oi_1 _5624_ (.A1(net923),
    .A2(_1666_),
    .Y(_1777_),
    .B1(net910));
 sg13g2_nand3_1 _5625_ (.B(net916),
    .C(_1653_),
    .A(_1589_),
    .Y(_1778_));
 sg13g2_nand2_1 _5626_ (.Y(_1779_),
    .A(_1713_),
    .B(_1724_));
 sg13g2_a221oi_1 _5627_ (.B2(_1672_),
    .C1(_1581_),
    .B1(_1779_),
    .A1(_1777_),
    .Y(_1780_),
    .A2(_1778_));
 sg13g2_nor3_1 _5628_ (.A(net901),
    .B(_1770_),
    .C(_1780_),
    .Y(_1781_));
 sg13g2_o21ai_1 _5629_ (.B1(_1781_),
    .Y(_1782_),
    .A1(_1618_),
    .A2(_1776_));
 sg13g2_a21oi_1 _5630_ (.A1(_1764_),
    .A2(_1782_),
    .Y(_1783_),
    .B1(_1369_));
 sg13g2_nor3_1 _5631_ (.A(_1625_),
    .B(_1683_),
    .C(_1716_),
    .Y(_1784_));
 sg13g2_a21oi_1 _5632_ (.A1(net914),
    .A2(_1716_),
    .Y(_1785_),
    .B1(_1784_));
 sg13g2_nor3_1 _5633_ (.A(net929),
    .B(_1625_),
    .C(_1666_),
    .Y(_1786_));
 sg13g2_a221oi_1 _5634_ (.B2(_1702_),
    .C1(net909),
    .B1(_1786_),
    .A1(net929),
    .Y(_1787_),
    .A2(_1785_));
 sg13g2_o21ai_1 _5635_ (.B1(net917),
    .Y(_1788_),
    .A1(net927),
    .A2(_1660_));
 sg13g2_nor2_1 _5636_ (.A(_1731_),
    .B(_1788_),
    .Y(_1789_));
 sg13g2_o21ai_1 _5637_ (.B1(net909),
    .Y(_1790_),
    .A1(_1583_),
    .A2(_1685_));
 sg13g2_nor3_1 _5638_ (.A(net924),
    .B(net917),
    .C(_1610_),
    .Y(_1791_));
 sg13g2_nor3_1 _5639_ (.A(_1789_),
    .B(_1790_),
    .C(_1791_),
    .Y(_1792_));
 sg13g2_nor3_1 _5640_ (.A(_1576_),
    .B(_1787_),
    .C(_1792_),
    .Y(_1793_));
 sg13g2_nor2_1 _5641_ (.A(_1625_),
    .B(_1654_),
    .Y(_1794_));
 sg13g2_nor3_2 _5642_ (.A(net925),
    .B(_1625_),
    .C(_1654_),
    .Y(_1795_));
 sg13g2_a22oi_1 _5643_ (.Y(_1796_),
    .B1(_1666_),
    .B2(_1794_),
    .A2(_1665_),
    .A1(net917));
 sg13g2_o21ai_1 _5644_ (.B1(net917),
    .Y(_1797_),
    .A1(_1625_),
    .A2(_1654_));
 sg13g2_inv_1 _5645_ (.Y(_1798_),
    .A(_1797_));
 sg13g2_nand2_1 _5646_ (.Y(_1799_),
    .A(net914),
    .B(_1660_));
 sg13g2_nand4_1 _5647_ (.B(net909),
    .C(_1797_),
    .A(net926),
    .Y(_1800_),
    .D(_1799_));
 sg13g2_o21ai_1 _5648_ (.B1(_1665_),
    .Y(_1801_),
    .A1(_1703_),
    .A2(_1727_));
 sg13g2_nor4_1 _5649_ (.A(net914),
    .B(_1609_),
    .C(net900),
    .D(_1660_),
    .Y(_1802_));
 sg13g2_o21ai_1 _5650_ (.B1(net904),
    .Y(_1803_),
    .A1(_1772_),
    .A2(_1802_));
 sg13g2_o21ai_1 _5651_ (.B1(_1635_),
    .Y(_1804_),
    .A1(_1614_),
    .A2(_1795_));
 sg13g2_o21ai_1 _5652_ (.B1(_1803_),
    .Y(_1805_),
    .A1(_1740_),
    .A2(_1804_));
 sg13g2_nand2_1 _5653_ (.Y(_1806_),
    .A(_1580_),
    .B(_1805_));
 sg13g2_o21ai_1 _5654_ (.B1(_1777_),
    .Y(_1807_),
    .A1(net916),
    .A2(_1713_));
 sg13g2_a21oi_1 _5655_ (.A1(_1629_),
    .A2(_1661_),
    .Y(_1808_),
    .B1(_1807_));
 sg13g2_a221oi_1 _5656_ (.B2(net925),
    .C1(net904),
    .B1(_1798_),
    .A1(_1713_),
    .Y(_1809_),
    .A2(_1724_));
 sg13g2_o21ai_1 _5657_ (.B1(_1617_),
    .Y(_1810_),
    .A1(_1808_),
    .A2(_1809_));
 sg13g2_a21oi_1 _5658_ (.A1(_1589_),
    .A2(_1611_),
    .Y(_1811_),
    .B1(_1759_));
 sg13g2_nor2_1 _5659_ (.A(net917),
    .B(_1625_),
    .Y(_1812_));
 sg13g2_nand3_1 _5660_ (.B(_1653_),
    .C(_1665_),
    .A(net909),
    .Y(_1813_));
 sg13g2_o21ai_1 _5661_ (.B1(_1620_),
    .Y(_1814_),
    .A1(_1812_),
    .A2(_1813_));
 sg13g2_a21oi_1 _5662_ (.A1(_1741_),
    .A2(_1811_),
    .Y(_1815_),
    .B1(_1814_));
 sg13g2_nand2_1 _5663_ (.Y(_1816_),
    .A(net918),
    .B(_1655_));
 sg13g2_a21oi_1 _5664_ (.A1(net925),
    .A2(_1740_),
    .Y(_1817_),
    .B1(net904));
 sg13g2_a221oi_1 _5665_ (.B2(_1817_),
    .C1(_1616_),
    .B1(_1816_),
    .A1(_1626_),
    .Y(_1818_),
    .A2(_1758_));
 sg13g2_a21oi_1 _5666_ (.A1(_1611_),
    .A2(_1723_),
    .Y(_1819_),
    .B1(_1772_));
 sg13g2_o21ai_1 _5667_ (.B1(net929),
    .Y(_1820_),
    .A1(net909),
    .A2(_1796_));
 sg13g2_a21oi_1 _5668_ (.A1(net909),
    .A2(_1819_),
    .Y(_1821_),
    .B1(_1820_));
 sg13g2_a21oi_1 _5669_ (.A1(_1800_),
    .A2(_1801_),
    .Y(_1822_),
    .B1(net929));
 sg13g2_nor3_1 _5670_ (.A(net932),
    .B(_1821_),
    .C(_1822_),
    .Y(_1823_));
 sg13g2_o21ai_1 _5671_ (.B1(net901),
    .Y(_1824_),
    .A1(_1793_),
    .A2(_1823_));
 sg13g2_nor3_1 _5672_ (.A(net901),
    .B(_1815_),
    .C(_1818_),
    .Y(_1825_));
 sg13g2_nand3_1 _5673_ (.B(_1810_),
    .C(_1825_),
    .A(_1806_),
    .Y(_1826_));
 sg13g2_nand3_1 _5674_ (.B(_1824_),
    .C(_1826_),
    .A(net982),
    .Y(_1827_));
 sg13g2_nand4_1 _5675_ (.B(net982),
    .C(_1824_),
    .A(\i_music.i_sample.sample_acc[1] ),
    .Y(_1828_),
    .D(_1826_));
 sg13g2_nor4_1 _5676_ (.A(net910),
    .B(_1656_),
    .C(_1684_),
    .D(_1771_),
    .Y(_1829_));
 sg13g2_o21ai_1 _5677_ (.B1(_1593_),
    .Y(_1830_),
    .A1(_1654_),
    .A2(_1715_));
 sg13g2_o21ai_1 _5678_ (.B1(_1830_),
    .Y(_1831_),
    .A1(_1670_),
    .A2(_1816_));
 sg13g2_nor2_1 _5679_ (.A(net905),
    .B(_1831_),
    .Y(_1832_));
 sg13g2_o21ai_1 _5680_ (.B1(_1580_),
    .Y(_1833_),
    .A1(_1829_),
    .A2(_1832_));
 sg13g2_nor2_1 _5681_ (.A(_1659_),
    .B(_1797_),
    .Y(_1834_));
 sg13g2_nor3_1 _5682_ (.A(net911),
    .B(_1743_),
    .C(_1834_),
    .Y(_1835_));
 sg13g2_nor2_1 _5683_ (.A(_1685_),
    .B(_1713_),
    .Y(_1836_));
 sg13g2_a21oi_1 _5684_ (.A1(net924),
    .A2(_1696_),
    .Y(_1837_),
    .B1(_1791_));
 sg13g2_nor3_1 _5685_ (.A(net907),
    .B(_1836_),
    .C(_1837_),
    .Y(_1838_));
 sg13g2_nor3_1 _5686_ (.A(_1618_),
    .B(_1835_),
    .C(_1838_),
    .Y(_1839_));
 sg13g2_nor2_1 _5687_ (.A(_1715_),
    .B(_1816_),
    .Y(_1840_));
 sg13g2_a21oi_1 _5688_ (.A1(net900),
    .A2(_1684_),
    .Y(_1841_),
    .B1(net905));
 sg13g2_a21oi_1 _5689_ (.A1(_1778_),
    .A2(_1841_),
    .Y(_1842_),
    .B1(_1616_));
 sg13g2_o21ai_1 _5690_ (.B1(_1842_),
    .Y(_1843_),
    .A1(_1807_),
    .A2(_1840_));
 sg13g2_nor3_1 _5691_ (.A(_1611_),
    .B(_1759_),
    .C(_1795_),
    .Y(_1844_));
 sg13g2_nor2_1 _5692_ (.A(net902),
    .B(_1670_),
    .Y(_1845_));
 sg13g2_nor3_1 _5693_ (.A(net907),
    .B(_1749_),
    .C(_1845_),
    .Y(_1846_));
 sg13g2_o21ai_1 _5694_ (.B1(_1620_),
    .Y(_1847_),
    .A1(_1844_),
    .A2(_1846_));
 sg13g2_nand3_1 _5695_ (.B(_1843_),
    .C(_1847_),
    .A(_1833_),
    .Y(_1848_));
 sg13g2_o21ai_1 _5696_ (.B1(net901),
    .Y(_1849_),
    .A1(_1839_),
    .A2(_1848_));
 sg13g2_a221oi_1 _5697_ (.B2(net919),
    .C1(net907),
    .B1(_1718_),
    .A1(net922),
    .Y(_1850_),
    .A2(_1609_));
 sg13g2_o21ai_1 _5698_ (.B1(net908),
    .Y(_1851_),
    .A1(_1683_),
    .A2(_1695_));
 sg13g2_nor2_1 _5699_ (.A(_1698_),
    .B(_1771_),
    .Y(_1852_));
 sg13g2_nand2_1 _5700_ (.Y(_1853_),
    .A(net911),
    .B(_1739_));
 sg13g2_a21oi_1 _5701_ (.A1(net913),
    .A2(_1717_),
    .Y(_1854_),
    .B1(_1853_));
 sg13g2_mux2_1 _5702_ (.A0(_1703_),
    .A1(_1732_),
    .S(_1665_),
    .X(_1855_));
 sg13g2_o21ai_1 _5703_ (.B1(_1580_),
    .Y(_1856_),
    .A1(_1854_),
    .A2(_1855_));
 sg13g2_o21ai_1 _5704_ (.B1(_1669_),
    .Y(_1857_),
    .A1(net902),
    .A2(_1613_));
 sg13g2_a21oi_1 _5705_ (.A1(net919),
    .A2(_1652_),
    .Y(_1858_),
    .B1(net912));
 sg13g2_a21oi_1 _5706_ (.A1(_1857_),
    .A2(_1858_),
    .Y(_1859_),
    .B1(_1618_));
 sg13g2_o21ai_1 _5707_ (.B1(_1859_),
    .Y(_1860_),
    .A1(_1790_),
    .A2(_1845_));
 sg13g2_o21ai_1 _5708_ (.B1(net927),
    .Y(_1861_),
    .A1(_1812_),
    .A2(_1851_));
 sg13g2_o21ai_1 _5709_ (.B1(net911),
    .Y(_1862_),
    .A1(_1716_),
    .A2(_1852_));
 sg13g2_nor3_1 _5710_ (.A(net911),
    .B(_1738_),
    .C(_1836_),
    .Y(_1863_));
 sg13g2_nor2_1 _5711_ (.A(net927),
    .B(_1863_),
    .Y(_1864_));
 sg13g2_a21oi_1 _5712_ (.A1(_1862_),
    .A2(_1864_),
    .Y(_1865_),
    .B1(net931));
 sg13g2_o21ai_1 _5713_ (.B1(_1865_),
    .Y(_1866_),
    .A1(_1850_),
    .A2(_1861_));
 sg13g2_nand4_1 _5714_ (.B(_1856_),
    .C(_1860_),
    .A(_1600_),
    .Y(_1867_),
    .D(_1866_));
 sg13g2_nand3_1 _5715_ (.B(_1849_),
    .C(_1867_),
    .A(net982),
    .Y(_1868_));
 sg13g2_nand4_1 _5716_ (.B(net982),
    .C(_1849_),
    .A(net334),
    .Y(_1869_),
    .D(_1867_));
 sg13g2_xor2_1 _5717_ (.B(_1827_),
    .A(\i_music.i_sample.sample_acc[1] ),
    .X(_1870_));
 sg13g2_o21ai_1 _5718_ (.B1(_1828_),
    .Y(_1871_),
    .A1(_1869_),
    .A2(_1870_));
 sg13g2_xnor2_1 _5719_ (.Y(_1872_),
    .A(\i_music.i_sample.sample_acc[2] ),
    .B(_1783_));
 sg13g2_nor2b_1 _5720_ (.A(_1872_),
    .B_N(_1871_),
    .Y(_1873_));
 sg13g2_a21o_1 _5721_ (.A2(_1783_),
    .A1(\i_music.i_sample.sample_acc[2] ),
    .B1(_1873_),
    .X(_1874_));
 sg13g2_xnor2_1 _5722_ (.Y(_1875_),
    .A(net371),
    .B(_1737_));
 sg13g2_a22oi_1 _5723_ (.Y(_1876_),
    .B1(_1874_),
    .B2(_1875_),
    .A2(_1737_),
    .A1(\i_music.i_sample.sample_acc[3] ));
 sg13g2_xnor2_1 _5724_ (.Y(_1877_),
    .A(\i_music.i_sample.sample_acc[4] ),
    .B(_1693_));
 sg13g2_o21ai_1 _5725_ (.B1(_1694_),
    .Y(_1878_),
    .A1(_1876_),
    .A2(_1877_));
 sg13g2_a21oi_1 _5726_ (.A1(_1651_),
    .A2(_1878_),
    .Y(_1879_),
    .B1(_1650_));
 sg13g2_xor2_1 _5727_ (.B(_1624_),
    .A(\i_music.i_sample.sample_acc[6] ),
    .X(_1880_));
 sg13g2_nor2b_1 _5728_ (.A(_1879_),
    .B_N(_1880_),
    .Y(_1881_));
 sg13g2_a21o_1 _5729_ (.A2(_1624_),
    .A1(\i_music.i_sample.sample_acc[6] ),
    .B1(_1881_),
    .X(_1882_));
 sg13g2_nor2b_1 _5730_ (.A(net255),
    .B_N(_1882_),
    .Y(_1883_));
 sg13g2_xnor2_1 _5731_ (.Y(_1884_),
    .A(\i_music.i_sample.sample_acc[8] ),
    .B(_1883_));
 sg13g2_nor2_1 _5732_ (.A(_1573_),
    .B(net256),
    .Y(_0106_));
 sg13g2_xor2_1 _5733_ (.B(_1882_),
    .A(net319),
    .X(_1885_));
 sg13g2_and2_1 _5734_ (.A(_0136_),
    .B(_1885_),
    .X(_0107_));
 sg13g2_and2_1 _5735_ (.A(\i_music.i_sample.t1.genblk1[18].state.Q ),
    .B(net1088),
    .X(_0108_));
 sg13g2_a21o_2 _5736_ (.A2(_1533_),
    .A1(net1089),
    .B1(net1156),
    .X(_1886_));
 sg13g2_inv_2 _5737_ (.Y(_1887_),
    .A(_1886_));
 sg13g2_o21ai_1 _5738_ (.B1(_1548_),
    .Y(_1888_),
    .A1(net325),
    .A2(_1545_));
 sg13g2_mux2_1 _5739_ (.A0(net325),
    .A1(_1888_),
    .S(_1886_),
    .X(_0109_));
 sg13g2_nand2_2 _5740_ (.Y(_1889_),
    .A(net1157),
    .B(_2985_));
 sg13g2_nand3_1 _5741_ (.B(\i_music.violin_note_idx[3][0] ),
    .C(\i_music.violin_note_idx[3][2] ),
    .A(\i_music.violin_note_idx[3][1] ),
    .Y(_1890_));
 sg13g2_nor2_1 _5742_ (.A(_2949_),
    .B(_1890_),
    .Y(_1891_));
 sg13g2_nor3_2 _5743_ (.A(_2949_),
    .B(_2951_),
    .C(_1890_),
    .Y(_1892_));
 sg13g2_o21ai_1 _5744_ (.B1(_1544_),
    .Y(_1893_),
    .A1(\i_music.violin_note_idx[3][4] ),
    .A2(_1891_));
 sg13g2_o21ai_1 _5745_ (.B1(_1548_),
    .Y(_1894_),
    .A1(_1892_),
    .A2(_1893_));
 sg13g2_mux2_1 _5746_ (.A0(net336),
    .A1(_1894_),
    .S(_1886_),
    .X(_1895_));
 sg13g2_nand2_1 _5747_ (.Y(_1896_),
    .A(_1889_),
    .B(_1895_));
 sg13g2_inv_1 _5748_ (.Y(_0110_),
    .A(_1896_));
 sg13g2_xnor2_1 _5749_ (.Y(_1897_),
    .A(\i_music.violin_note_idx[3][5] ),
    .B(_1892_));
 sg13g2_nand2_1 _5750_ (.Y(_1898_),
    .A(_1544_),
    .B(_1897_));
 sg13g2_nand3_1 _5751_ (.B(_1886_),
    .C(_1898_),
    .A(_1548_),
    .Y(_1899_));
 sg13g2_a21oi_1 _5752_ (.A1(net343),
    .A2(_1887_),
    .Y(_1900_),
    .B1(_1554_));
 sg13g2_nand2_1 _5753_ (.Y(_0111_),
    .A(_1899_),
    .B(_1900_));
 sg13g2_nand3_1 _5754_ (.B(\i_music.violin_note_idx[3][6] ),
    .C(_1892_),
    .A(\i_music.violin_note_idx[3][5] ),
    .Y(_1901_));
 sg13g2_a21oi_1 _5755_ (.A1(\i_music.violin_note_idx[3][5] ),
    .A2(_1892_),
    .Y(_1902_),
    .B1(net314));
 sg13g2_nand2_1 _5756_ (.Y(_1903_),
    .A(_1546_),
    .B(_1901_));
 sg13g2_o21ai_1 _5757_ (.B1(_1561_),
    .Y(_1904_),
    .A1(_1902_),
    .A2(_1903_));
 sg13g2_mux2_1 _5758_ (.A0(net314),
    .A1(_1904_),
    .S(_1886_),
    .X(_0112_));
 sg13g2_xnor2_1 _5759_ (.Y(_1905_),
    .A(_0043_),
    .B(_1901_));
 sg13g2_o21ai_1 _5760_ (.B1(_1561_),
    .Y(_1906_),
    .A1(_1547_),
    .A2(_1905_));
 sg13g2_mux2_1 _5761_ (.A0(net220),
    .A1(_1906_),
    .S(_1886_),
    .X(_0113_));
 sg13g2_nand4_1 _5762_ (.B(\i_music.violin_note_idx[3][6] ),
    .C(\i_music.violin_note_idx[3][7] ),
    .A(\i_music.violin_note_idx[3][5] ),
    .Y(_1907_),
    .D(_1892_));
 sg13g2_xor2_1 _5763_ (.B(_1907_),
    .A(\i_music.violin_note_idx[3][8] ),
    .X(_1908_));
 sg13g2_a21oi_1 _5764_ (.A1(_1557_),
    .A2(_1908_),
    .Y(_1909_),
    .B1(net1156));
 sg13g2_nor2_1 _5765_ (.A(net265),
    .B(_1886_),
    .Y(_1910_));
 sg13g2_nor2_1 _5766_ (.A(_1554_),
    .B(_1909_),
    .Y(_1911_));
 sg13g2_a21oi_1 _5767_ (.A1(_1886_),
    .A2(_1911_),
    .Y(_0114_),
    .B1(_1910_));
 sg13g2_xnor2_1 _5768_ (.Y(_1912_),
    .A(\i_music.violin_note_idx[3][1] ),
    .B(\i_music.violin_note_idx[3][0] ));
 sg13g2_a221oi_1 _5769_ (.B2(_1912_),
    .C1(_1887_),
    .B1(_1546_),
    .A1(net1170),
    .Y(_1913_),
    .A2(_1541_));
 sg13g2_a21o_1 _5770_ (.A2(_1887_),
    .A1(net308),
    .B1(_1913_),
    .X(_0115_));
 sg13g2_o21ai_1 _5771_ (.B1(_2957_),
    .Y(_1914_),
    .A1(_2954_),
    .A2(_2956_));
 sg13g2_and2_1 _5772_ (.A(_1890_),
    .B(_1914_),
    .X(_1915_));
 sg13g2_nand2_2 _5773_ (.Y(_1916_),
    .A(net1170),
    .B(net1089));
 sg13g2_a21oi_1 _5774_ (.A1(_1557_),
    .A2(_1915_),
    .Y(_1917_),
    .B1(_1916_));
 sg13g2_a22oi_1 _5775_ (.Y(_0116_),
    .B1(_1917_),
    .B2(_1533_),
    .A2(_1887_),
    .A1(_2957_));
 sg13g2_xnor2_1 _5776_ (.Y(_1918_),
    .A(net333),
    .B(_1890_));
 sg13g2_a221oi_1 _5777_ (.B2(_1918_),
    .C1(_1887_),
    .B1(_1546_),
    .A1(net1170),
    .Y(_1919_),
    .A2(_1541_));
 sg13g2_a21oi_1 _5778_ (.A1(_2949_),
    .A2(_1887_),
    .Y(_0117_),
    .B1(_1919_));
 sg13g2_nor3_2 _5779_ (.A(_0847_),
    .B(_0878_),
    .C(_0881_),
    .Y(_0118_));
 sg13g2_nand4_1 _5780_ (.B(\i_music.i_pwm.count[4] ),
    .C(\i_music.i_pwm.count[6] ),
    .A(\i_music.i_pwm.count[5] ),
    .Y(_1920_),
    .D(\i_music.i_pwm.count[7] ));
 sg13g2_nand4_1 _5781_ (.B(\i_music.i_pwm.count[1] ),
    .C(\i_music.i_pwm.count[3] ),
    .A(_2926_),
    .Y(_1921_),
    .D(\i_music.i_pwm.count[2] ));
 sg13g2_o21ai_1 _5782_ (.B1(net1174),
    .Y(_1922_),
    .A1(_1920_),
    .A2(_1921_));
 sg13g2_nor2_1 _5783_ (.A(_2991_),
    .B(_1922_),
    .Y(_0119_));
 sg13g2_a21o_1 _5784_ (.A2(\i_music.i_pwm.count[1] ),
    .A1(net301),
    .B1(_1922_),
    .X(_1923_));
 sg13g2_a21oi_1 _5785_ (.A1(_2926_),
    .A2(_2960_),
    .Y(_0120_),
    .B1(_1923_));
 sg13g2_and3_1 _5786_ (.X(_1924_),
    .A(\i_music.i_pwm.count[0] ),
    .B(\i_music.i_pwm.count[1] ),
    .C(net227));
 sg13g2_a21oi_1 _5787_ (.A1(\i_music.i_pwm.count[0] ),
    .A2(\i_music.i_pwm.count[1] ),
    .Y(_1925_),
    .B1(net227));
 sg13g2_nor3_1 _5788_ (.A(_1922_),
    .B(_1924_),
    .C(net228),
    .Y(_0121_));
 sg13g2_and2_1 _5789_ (.A(net266),
    .B(_1924_),
    .X(_1926_));
 sg13g2_nor2_1 _5790_ (.A(net266),
    .B(_1924_),
    .Y(_1927_));
 sg13g2_nor3_1 _5791_ (.A(_1922_),
    .B(_1926_),
    .C(net267),
    .Y(_0122_));
 sg13g2_nor2_1 _5792_ (.A(net292),
    .B(_1926_),
    .Y(_1928_));
 sg13g2_and2_1 _5793_ (.A(net292),
    .B(_1926_),
    .X(_1929_));
 sg13g2_nor3_1 _5794_ (.A(_1922_),
    .B(_1928_),
    .C(_1929_),
    .Y(_0123_));
 sg13g2_nor2_1 _5795_ (.A(net285),
    .B(_1929_),
    .Y(_1930_));
 sg13g2_and2_1 _5796_ (.A(net285),
    .B(_1929_),
    .X(_1931_));
 sg13g2_nor3_1 _5797_ (.A(_1922_),
    .B(net286),
    .C(_1931_),
    .Y(_0124_));
 sg13g2_nor2_1 _5798_ (.A(net283),
    .B(_1931_),
    .Y(_1932_));
 sg13g2_and2_1 _5799_ (.A(net283),
    .B(_1931_),
    .X(_1933_));
 sg13g2_nor3_1 _5800_ (.A(_1922_),
    .B(net284),
    .C(_1933_),
    .Y(_0125_));
 sg13g2_a21oi_1 _5801_ (.A1(net322),
    .A2(_1933_),
    .Y(_1934_),
    .B1(_1922_));
 sg13g2_o21ai_1 _5802_ (.B1(_1934_),
    .Y(_1935_),
    .A1(net322),
    .A2(_1933_));
 sg13g2_inv_1 _5803_ (.Y(_0126_),
    .A(_1935_));
 sg13g2_xor2_1 _5804_ (.B(_1870_),
    .A(_1869_),
    .X(_1936_));
 sg13g2_mux2_1 _5805_ (.A0(_1936_),
    .A1(net290),
    .S(net1031),
    .X(_0127_));
 sg13g2_xor2_1 _5806_ (.B(_1872_),
    .A(_1871_),
    .X(_1937_));
 sg13g2_nand2_1 _5807_ (.Y(_1938_),
    .A(net257),
    .B(net1031));
 sg13g2_o21ai_1 _5808_ (.B1(_1938_),
    .Y(_0128_),
    .A1(net1031),
    .A2(_1937_));
 sg13g2_xnor2_1 _5809_ (.Y(_1939_),
    .A(_1874_),
    .B(_1875_));
 sg13g2_nand2_1 _5810_ (.Y(_1940_),
    .A(net247),
    .B(net1031));
 sg13g2_o21ai_1 _5811_ (.B1(_1940_),
    .Y(_0129_),
    .A1(net1031),
    .A2(_1939_));
 sg13g2_xor2_1 _5812_ (.B(_1877_),
    .A(_1876_),
    .X(_1941_));
 sg13g2_nor2_1 _5813_ (.A(net1031),
    .B(_1941_),
    .Y(_1942_));
 sg13g2_a21oi_1 _5814_ (.A1(_2989_),
    .A2(net1030),
    .Y(_0130_),
    .B1(_1942_));
 sg13g2_xnor2_1 _5815_ (.Y(_1943_),
    .A(_1651_),
    .B(_1878_));
 sg13g2_nand2_1 _5816_ (.Y(_1944_),
    .A(net232),
    .B(net1030));
 sg13g2_o21ai_1 _5817_ (.B1(_1944_),
    .Y(_0131_),
    .A1(net1030),
    .A2(_1943_));
 sg13g2_xnor2_1 _5818_ (.Y(_1945_),
    .A(_1879_),
    .B(_1880_));
 sg13g2_nor2_1 _5819_ (.A(net1030),
    .B(_1945_),
    .Y(_1946_));
 sg13g2_a21oi_1 _5820_ (.A1(_2987_),
    .A2(net1031),
    .Y(_0132_),
    .B1(_1946_));
 sg13g2_nor2_1 _5821_ (.A(_1885_),
    .B(net1030),
    .Y(_1947_));
 sg13g2_a21oi_1 _5822_ (.A1(_2986_),
    .A2(net1030),
    .Y(_0133_),
    .B1(_1947_));
 sg13g2_nand2_1 _5823_ (.Y(_1948_),
    .A(net243),
    .B(net1030));
 sg13g2_o21ai_1 _5824_ (.B1(_1948_),
    .Y(_0134_),
    .A1(_1884_),
    .A2(net1030));
 sg13g2_nand2b_1 _5825_ (.Y(_0135_),
    .B(net1171),
    .A_N(net209));
 sg13g2_a21oi_1 _5826_ (.A1(net1164),
    .A2(_2996_),
    .Y(_1949_),
    .B1(net217));
 sg13g2_a21oi_1 _5827_ (.A1(net217),
    .A2(_1916_),
    .Y(_0137_),
    .B1(_1949_));
 sg13g2_a21oi_1 _5828_ (.A1(\i_display.i_vga.low_count[2] ),
    .A2(net1088),
    .Y(_1950_),
    .B1(net331));
 sg13g2_nor3_1 _5829_ (.A(net1158),
    .B(_2997_),
    .C(net332),
    .Y(_0138_));
 sg13g2_o21ai_1 _5830_ (.B1(net1165),
    .Y(_1951_),
    .A1(net218),
    .A2(_2998_));
 sg13g2_a21oi_1 _5831_ (.A1(net218),
    .A2(_2998_),
    .Y(_0139_),
    .B1(_1951_));
 sg13g2_a21oi_1 _5832_ (.A1(\i_display.i_vga.low_count[4] ),
    .A2(_2997_),
    .Y(_1952_),
    .B1(net323));
 sg13g2_nor3_1 _5833_ (.A(net1155),
    .B(_3057_),
    .C(net324),
    .Y(_0140_));
 sg13g2_o21ai_1 _5834_ (.B1(net1165),
    .Y(_1953_),
    .A1(net310),
    .A2(_3057_));
 sg13g2_a21oi_1 _5835_ (.A1(net310),
    .A2(_3057_),
    .Y(_0141_),
    .B1(_1953_));
 sg13g2_nor2b_1 _5836_ (.A(net245),
    .B_N(_3057_),
    .Y(_1954_));
 sg13g2_o21ai_1 _5837_ (.B1(net1165),
    .Y(_1955_),
    .A1(net1141),
    .A2(_1954_));
 sg13g2_a21oi_1 _5838_ (.A1(net1141),
    .A2(_1954_),
    .Y(_0142_),
    .B1(_1955_));
 sg13g2_o21ai_1 _5839_ (.B1(net1165),
    .Y(_1956_),
    .A1(net210),
    .A2(_3058_));
 sg13g2_a21oi_1 _5840_ (.A1(net210),
    .A2(_3058_),
    .Y(_0143_),
    .B1(_1956_));
 sg13g2_o21ai_1 _5841_ (.B1(_2929_),
    .Y(_1957_),
    .A1(_2928_),
    .A2(_3058_));
 sg13g2_and3_1 _5842_ (.X(_0144_),
    .A(net1164),
    .B(_3059_),
    .C(_1957_));
 sg13g2_a21oi_1 _5843_ (.A1(_2945_),
    .A2(_3059_),
    .Y(_1958_),
    .B1(net1155));
 sg13g2_nor2b_1 _5844_ (.A(_3060_),
    .B_N(_1958_),
    .Y(_0145_));
 sg13g2_o21ai_1 _5845_ (.B1(net1167),
    .Y(_1959_),
    .A1(net287),
    .A2(_3060_));
 sg13g2_nor2_1 _5846_ (.A(_3061_),
    .B(_1959_),
    .Y(_0146_));
 sg13g2_o21ai_1 _5847_ (.B1(net1167),
    .Y(_1960_),
    .A1(net260),
    .A2(_3061_));
 sg13g2_nor2_1 _5848_ (.A(_3062_),
    .B(net261),
    .Y(_0147_));
 sg13g2_o21ai_1 _5849_ (.B1(net1168),
    .Y(_1961_),
    .A1(net273),
    .A2(_3062_));
 sg13g2_nor2_1 _5850_ (.A(_3063_),
    .B(_1961_),
    .Y(_0148_));
 sg13g2_o21ai_1 _5851_ (.B1(net1167),
    .Y(_1962_),
    .A1(net293),
    .A2(_3063_));
 sg13g2_nor2_1 _5852_ (.A(_3064_),
    .B(_1962_),
    .Y(_0149_));
 sg13g2_o21ai_1 _5853_ (.B1(net1173),
    .Y(_1963_),
    .A1(net296),
    .A2(_3064_));
 sg13g2_nor2_1 _5854_ (.A(_3065_),
    .B(_1963_),
    .Y(_0150_));
 sg13g2_o21ai_1 _5855_ (.B1(net1173),
    .Y(_1964_),
    .A1(net288),
    .A2(_3065_));
 sg13g2_nor2_1 _5856_ (.A(_3066_),
    .B(net289),
    .Y(_0151_));
 sg13g2_o21ai_1 _5857_ (.B1(net1173),
    .Y(_1965_),
    .A1(net300),
    .A2(_3066_));
 sg13g2_nor2_1 _5858_ (.A(_3067_),
    .B(_1965_),
    .Y(_0152_));
 sg13g2_o21ai_1 _5859_ (.B1(net1167),
    .Y(_1966_),
    .A1(net274),
    .A2(_3067_));
 sg13g2_nor2_1 _5860_ (.A(_3068_),
    .B(net275),
    .Y(_0153_));
 sg13g2_o21ai_1 _5861_ (.B1(net1167),
    .Y(_1967_),
    .A1(net353),
    .A2(_3068_));
 sg13g2_nor2_1 _5862_ (.A(_3069_),
    .B(_1967_),
    .Y(_0154_));
 sg13g2_o21ai_1 _5863_ (.B1(net1167),
    .Y(_1968_),
    .A1(net360),
    .A2(_3069_));
 sg13g2_nor2_1 _5864_ (.A(_3070_),
    .B(_1968_),
    .Y(_0155_));
 sg13g2_o21ai_1 _5865_ (.B1(net1167),
    .Y(_1969_),
    .A1(net367),
    .A2(_3070_));
 sg13g2_nor2_1 _5866_ (.A(_3071_),
    .B(_1969_),
    .Y(_0156_));
 sg13g2_o21ai_1 _5867_ (.B1(net1168),
    .Y(_1970_),
    .A1(net347),
    .A2(_3071_));
 sg13g2_nor2_1 _5868_ (.A(_3072_),
    .B(_1970_),
    .Y(_0157_));
 sg13g2_nor2b_1 _5869_ (.A(_0035_),
    .B_N(_3071_),
    .Y(_1971_));
 sg13g2_o21ai_1 _5870_ (.B1(net1168),
    .Y(_1972_),
    .A1(net237),
    .A2(_1971_));
 sg13g2_a21oi_1 _5871_ (.A1(net237),
    .A2(_1971_),
    .Y(_0158_),
    .B1(_1972_));
 sg13g2_a21oi_1 _5872_ (.A1(\i_music.count[23] ),
    .A2(_3072_),
    .Y(_1973_),
    .B1(net225));
 sg13g2_nor3_1 _5873_ (.A(net1157),
    .B(_3073_),
    .C(net226),
    .Y(_0159_));
 sg13g2_and2_1 _5874_ (.A(net346),
    .B(_3076_),
    .X(_1974_));
 sg13g2_o21ai_1 _5875_ (.B1(net1175),
    .Y(_1975_),
    .A1(net346),
    .A2(_3076_));
 sg13g2_nor2_1 _5876_ (.A(_1974_),
    .B(_1975_),
    .Y(_0163_));
 sg13g2_nor2_1 _5877_ (.A(net342),
    .B(_1974_),
    .Y(_1976_));
 sg13g2_a21oi_1 _5878_ (.A1(net342),
    .A2(_1974_),
    .Y(_1977_),
    .B1(net1160));
 sg13g2_nor2b_1 _5879_ (.A(_1976_),
    .B_N(_1977_),
    .Y(_0164_));
 sg13g2_a21oi_1 _5880_ (.A1(\crotchet[4] ),
    .A2(_1974_),
    .Y(_1978_),
    .B1(net312));
 sg13g2_and3_1 _5881_ (.X(_1979_),
    .A(net348),
    .B(net312),
    .C(_1974_));
 sg13g2_nor3_1 _5882_ (.A(net1160),
    .B(net313),
    .C(_1979_),
    .Y(_0165_));
 sg13g2_o21ai_1 _5883_ (.B1(net1175),
    .Y(_1980_),
    .A1(net268),
    .A2(_1979_));
 sg13g2_a21oi_1 _5884_ (.A1(net268),
    .A2(_1979_),
    .Y(_0166_),
    .B1(_1980_));
 sg13g2_nand2_1 _5885_ (.Y(_1981_),
    .A(net1159),
    .B(net215));
 sg13g2_nor2_1 _5886_ (.A(\i_music.i_pwm.count[6] ),
    .B(_2986_),
    .Y(_1982_));
 sg13g2_nand2b_1 _5887_ (.Y(_1983_),
    .B(\i_music.i_pwm.count[2] ),
    .A_N(\i_music.i_pwm.sample[2] ));
 sg13g2_a22oi_1 _5888_ (.Y(_1984_),
    .B1(\i_music.i_pwm.sample[0] ),
    .B2(_2926_),
    .A2(\i_music.i_pwm.sample[1] ),
    .A1(_2960_));
 sg13g2_a21oi_1 _5889_ (.A1(\i_music.i_pwm.count[1] ),
    .A2(_2990_),
    .Y(_1985_),
    .B1(_1984_));
 sg13g2_nand2b_1 _5890_ (.Y(_1986_),
    .B(\i_music.i_pwm.sample[2] ),
    .A_N(\i_music.i_pwm.count[2] ));
 sg13g2_o21ai_1 _5891_ (.B1(_1986_),
    .Y(_1987_),
    .A1(\i_music.i_pwm.count[3] ),
    .A2(_2989_));
 sg13g2_a21oi_1 _5892_ (.A1(_1983_),
    .A2(_1985_),
    .Y(_1988_),
    .B1(_1987_));
 sg13g2_a221oi_1 _5893_ (.B2(\i_music.i_pwm.count[3] ),
    .C1(_1988_),
    .B1(_2989_),
    .A1(\i_music.i_pwm.count[4] ),
    .Y(_1989_),
    .A2(_2988_));
 sg13g2_a21oi_1 _5894_ (.A1(_2961_),
    .A2(\i_music.i_pwm.sample[4] ),
    .Y(_1990_),
    .B1(_1989_));
 sg13g2_o21ai_1 _5895_ (.B1(_1990_),
    .Y(_1991_),
    .A1(\i_music.i_pwm.count[5] ),
    .A2(_2987_));
 sg13g2_a22oi_1 _5896_ (.Y(_1992_),
    .B1(_2987_),
    .B2(\i_music.i_pwm.count[5] ),
    .A2(_2986_),
    .A1(\i_music.i_pwm.count[6] ));
 sg13g2_a221oi_1 _5897_ (.B2(_1992_),
    .C1(_1982_),
    .B1(_1991_),
    .A1(_2962_),
    .Y(_1993_),
    .A2(\i_music.i_pwm.sample[7] ));
 sg13g2_o21ai_1 _5898_ (.B1(net1174),
    .Y(_1994_),
    .A1(_2962_),
    .A2(\i_music.i_pwm.sample[7] ));
 sg13g2_o21ai_1 _5899_ (.B1(_1981_),
    .Y(_0167_),
    .A1(_1993_),
    .A2(_1994_));
 sg13g2_nand2_1 _5900_ (.Y(_1995_),
    .A(net1083),
    .B(_1533_));
 sg13g2_inv_1 _5901_ (.Y(_1996_),
    .A(net981));
 sg13g2_nand2_1 _5902_ (.Y(_1997_),
    .A(\i_music.violin_note_idx[1][1] ),
    .B(\i_music.violin_note_idx[1][0] ));
 sg13g2_nand2_1 _5903_ (.Y(_1998_),
    .A(_1542_),
    .B(_1997_));
 sg13g2_a21oi_1 _5904_ (.A1(net328),
    .A2(net981),
    .Y(_1999_),
    .B1(net1156));
 sg13g2_o21ai_1 _5905_ (.B1(_1999_),
    .Y(_0168_),
    .A1(net981),
    .A2(_1998_));
 sg13g2_o21ai_1 _5906_ (.B1(_1544_),
    .Y(_2000_),
    .A1(_0041_),
    .A2(_1997_));
 sg13g2_a21o_1 _5907_ (.A2(_1997_),
    .A1(_0041_),
    .B1(_2000_),
    .X(_2001_));
 sg13g2_nand2_1 _5908_ (.Y(_2002_),
    .A(net1169),
    .B(net981));
 sg13g2_a21oi_1 _5909_ (.A1(net294),
    .A2(_1995_),
    .Y(_2003_),
    .B1(net1157));
 sg13g2_o21ai_1 _5910_ (.B1(_2003_),
    .Y(_0169_),
    .A1(net981),
    .A2(_2001_));
 sg13g2_a21oi_1 _5911_ (.A1(_1996_),
    .A2(_2000_),
    .Y(_2004_),
    .B1(net262));
 sg13g2_nor4_1 _5912_ (.A(_2944_),
    .B(_0041_),
    .C(net981),
    .D(_1997_),
    .Y(_2005_));
 sg13g2_nor3_1 _5913_ (.A(net1156),
    .B(net263),
    .C(_2005_),
    .Y(_0170_));
 sg13g2_nor2_1 _5914_ (.A(net250),
    .B(net978),
    .Y(_2006_));
 sg13g2_nor2_1 _5915_ (.A(net1156),
    .B(_1534_),
    .Y(_2007_));
 sg13g2_nand2_1 _5916_ (.Y(_2008_),
    .A(_2925_),
    .B(_2955_));
 sg13g2_nand3_1 _5917_ (.B(_1557_),
    .C(_2008_),
    .A(_1549_),
    .Y(_2009_));
 sg13g2_a21oi_1 _5918_ (.A1(_2007_),
    .A2(_2009_),
    .Y(_0171_),
    .B1(_2006_));
 sg13g2_xnor2_1 _5919_ (.Y(_2010_),
    .A(net252),
    .B(_1549_));
 sg13g2_nand2_1 _5920_ (.Y(_2011_),
    .A(_1557_),
    .B(_2010_));
 sg13g2_nor2_1 _5921_ (.A(net252),
    .B(net978),
    .Y(_2012_));
 sg13g2_a21oi_1 _5922_ (.A1(_2007_),
    .A2(_2011_),
    .Y(_0172_),
    .B1(_2012_));
 sg13g2_o21ai_1 _5923_ (.B1(_2950_),
    .Y(_2013_),
    .A1(_2958_),
    .A2(_1549_));
 sg13g2_nand3b_1 _5924_ (.B(_1557_),
    .C(_2013_),
    .Y(_2014_),
    .A_N(_1550_));
 sg13g2_nor2_1 _5925_ (.A(net222),
    .B(net978),
    .Y(_2015_));
 sg13g2_a21oi_1 _5926_ (.A1(_2007_),
    .A2(_2014_),
    .Y(_0173_),
    .B1(_2015_));
 sg13g2_mux2_1 _5927_ (.A0(\crotchet[0] ),
    .A1(net258),
    .S(net1001),
    .X(_0174_));
 sg13g2_mux2_1 _5928_ (.A0(_0793_),
    .A1(net278),
    .S(net1001),
    .X(_0175_));
 sg13g2_mux2_1 _5929_ (.A0(_0782_),
    .A1(net239),
    .S(_3091_),
    .X(_0176_));
 sg13g2_mux2_1 _5930_ (.A0(net1057),
    .A1(net1137),
    .S(_3091_),
    .X(_0177_));
 sg13g2_nand2_1 _5931_ (.Y(_2016_),
    .A(net219),
    .B(net1001));
 sg13g2_o21ai_1 _5932_ (.B1(_2016_),
    .Y(_0178_),
    .A1(net1001),
    .A2(_3096_));
 sg13g2_mux2_1 _5933_ (.A0(net1059),
    .A1(net1134),
    .S(net1001),
    .X(_0179_));
 sg13g2_mux2_1 _5934_ (.A0(_0775_),
    .A1(net351),
    .S(_3091_),
    .X(_0180_));
 sg13g2_nor3_1 _5935_ (.A(net234),
    .B(_1541_),
    .C(_1547_),
    .Y(_2017_));
 sg13g2_nor2_1 _5936_ (.A(\i_music.violin_note_idx[2][0] ),
    .B(net978),
    .Y(_2018_));
 sg13g2_a21oi_1 _5937_ (.A1(net978),
    .A2(_2017_),
    .Y(_0182_),
    .B1(_2018_));
 sg13g2_nand2_1 _5938_ (.Y(_0183_),
    .A(_3077_),
    .B(_0023_));
 sg13g2_nand3_1 _5939_ (.B(_3079_),
    .C(_3082_),
    .A(_3077_),
    .Y(_0186_));
 sg13g2_nand3_1 _5940_ (.B(net304),
    .C(net981),
    .A(net1169),
    .Y(_2019_));
 sg13g2_nand4_1 _5941_ (.B(\i_music.violin_note_idx[1][0] ),
    .C(\i_music.violin_note_idx[1][2] ),
    .A(\i_music.violin_note_idx[1][1] ),
    .Y(_2020_),
    .D(\i_music.violin_note_idx[1][3] ));
 sg13g2_inv_1 _5942_ (.Y(_2021_),
    .A(_2020_));
 sg13g2_nor2_1 _5943_ (.A(_0038_),
    .B(_2020_),
    .Y(_2022_));
 sg13g2_xor2_1 _5944_ (.B(_2020_),
    .A(_0038_),
    .X(_2023_));
 sg13g2_nand3_1 _5945_ (.B(net977),
    .C(_2023_),
    .A(_1546_),
    .Y(_2024_));
 sg13g2_nand3_1 _5946_ (.B(_2019_),
    .C(_2024_),
    .A(_1889_),
    .Y(_0187_));
 sg13g2_nor2_1 _5947_ (.A(net279),
    .B(net977),
    .Y(_2025_));
 sg13g2_xor2_1 _5948_ (.B(_2022_),
    .A(\i_music.violin_note_idx[1][5] ),
    .X(_2026_));
 sg13g2_nor2_2 _5949_ (.A(net2),
    .B(_1889_),
    .Y(_2027_));
 sg13g2_a221oi_1 _5950_ (.B2(net1169),
    .C1(_2027_),
    .B1(_2026_),
    .A1(net2),
    .Y(_2028_),
    .A2(_1536_));
 sg13g2_a21oi_1 _5951_ (.A1(_2002_),
    .A2(_2028_),
    .Y(_0188_),
    .B1(_2025_));
 sg13g2_nand3_1 _5952_ (.B(\i_music.violin_note_idx[1][5] ),
    .C(_2021_),
    .A(\i_music.violin_note_idx[1][4] ),
    .Y(_2029_));
 sg13g2_xor2_1 _5953_ (.B(_2029_),
    .A(\i_music.violin_note_idx[1][6] ),
    .X(_2030_));
 sg13g2_a21oi_1 _5954_ (.A1(_1544_),
    .A2(_2030_),
    .Y(_2031_),
    .B1(net1156));
 sg13g2_nor2_1 _5955_ (.A(_2027_),
    .B(_2031_),
    .Y(_2032_));
 sg13g2_nor2_1 _5956_ (.A(net299),
    .B(net977),
    .Y(_2033_));
 sg13g2_a21oi_1 _5957_ (.A1(net977),
    .A2(_2032_),
    .Y(_0189_),
    .B1(_2033_));
 sg13g2_nor2_1 _5958_ (.A(_0039_),
    .B(_2029_),
    .Y(_2034_));
 sg13g2_xnor2_1 _5959_ (.Y(_2035_),
    .A(\i_music.violin_note_idx[1][7] ),
    .B(_2034_));
 sg13g2_a21oi_1 _5960_ (.A1(_1544_),
    .A2(_2035_),
    .Y(_2036_),
    .B1(net1156));
 sg13g2_nor2_1 _5961_ (.A(_2027_),
    .B(_2036_),
    .Y(_2037_));
 sg13g2_nor2_1 _5962_ (.A(net335),
    .B(_2002_),
    .Y(_2038_));
 sg13g2_a21oi_1 _5963_ (.A1(net977),
    .A2(_2037_),
    .Y(_0190_),
    .B1(_2038_));
 sg13g2_nor2_1 _5964_ (.A(net320),
    .B(net977),
    .Y(_2039_));
 sg13g2_nor2_1 _5965_ (.A(_1539_),
    .B(_2029_),
    .Y(_2040_));
 sg13g2_o21ai_1 _5966_ (.B1(net1169),
    .Y(_2041_),
    .A1(\i_music.violin_note_idx[1][8] ),
    .A2(_2040_));
 sg13g2_a21oi_1 _5967_ (.A1(\i_music.violin_note_idx[1][8] ),
    .A2(_2040_),
    .Y(_2042_),
    .B1(_2041_));
 sg13g2_nor2_1 _5968_ (.A(_2027_),
    .B(_2042_),
    .Y(_2043_));
 sg13g2_a21oi_1 _5969_ (.A1(net977),
    .A2(_2043_),
    .Y(_0191_),
    .B1(_2039_));
 sg13g2_nor2_1 _5970_ (.A(net952),
    .B(net947),
    .Y(_2044_));
 sg13g2_or2_1 _5971_ (.X(_2045_),
    .B(net945),
    .A(net950));
 sg13g2_nor2_1 _5972_ (.A(net958),
    .B(\i_music.i_sample.t1.genblk1[0].state.Q ),
    .Y(_2046_));
 sg13g2_or2_1 _5973_ (.X(_2047_),
    .B(net943),
    .A(net958));
 sg13g2_and2_1 _5974_ (.A(net958),
    .B(net943),
    .X(_2048_));
 sg13g2_nand2_2 _5975_ (.Y(_2049_),
    .A(net953),
    .B(net941));
 sg13g2_nand2_1 _5976_ (.Y(_2050_),
    .A(net955),
    .B(net950));
 sg13g2_a21oi_1 _5977_ (.A1(\i_music.i_sample.t1.genblk1[2].state.Q ),
    .A2(_2048_),
    .Y(_2051_),
    .B1(_2046_));
 sg13g2_mux2_1 _5978_ (.A0(net936),
    .A1(net947),
    .S(_2051_),
    .X(_2052_));
 sg13g2_nor2b_2 _5979_ (.A(net958),
    .B_N(net952),
    .Y(_2053_));
 sg13g2_a21oi_1 _5980_ (.A1(net947),
    .A2(_2053_),
    .Y(_2054_),
    .B1(_2046_));
 sg13g2_nand2_1 _5981_ (.Y(_2055_),
    .A(net965),
    .B(_2054_));
 sg13g2_nand2_2 _5982_ (.Y(_2056_),
    .A(net943),
    .B(net947));
 sg13g2_nand2_2 _5983_ (.Y(_2057_),
    .A(net957),
    .B(net944));
 sg13g2_nand2_2 _5984_ (.Y(_2058_),
    .A(net954),
    .B(_2045_));
 sg13g2_inv_1 _5985_ (.Y(_2059_),
    .A(_2058_));
 sg13g2_nor2b_1 _5986_ (.A(_2058_),
    .B_N(_2056_),
    .Y(_2060_));
 sg13g2_o21ai_1 _5987_ (.B1(net967),
    .Y(_2061_),
    .A1(_2055_),
    .A2(_2060_));
 sg13g2_a21oi_1 _5988_ (.A1(net938),
    .A2(_2052_),
    .Y(_2062_),
    .B1(_2061_));
 sg13g2_nor2_2 _5989_ (.A(net968),
    .B(net939),
    .Y(_2063_));
 sg13g2_nand2_1 _5990_ (.Y(_2064_),
    .A(net940),
    .B(net963));
 sg13g2_nor2_2 _5991_ (.A(net937),
    .B(net949),
    .Y(_2065_));
 sg13g2_nand2b_2 _5992_ (.Y(_2066_),
    .B(net958),
    .A_N(net952));
 sg13g2_nand2b_2 _5993_ (.Y(_2067_),
    .B(net947),
    .A_N(net952));
 sg13g2_nor2_2 _5994_ (.A(net942),
    .B(net945),
    .Y(_2068_));
 sg13g2_or2_1 _5995_ (.X(_2069_),
    .B(net947),
    .A(net943));
 sg13g2_nand2_2 _5996_ (.Y(_2070_),
    .A(net954),
    .B(_2068_));
 sg13g2_nand2b_2 _5997_ (.Y(_2071_),
    .B(net941),
    .A_N(net949));
 sg13g2_o21ai_1 _5998_ (.B1(_2070_),
    .Y(_2072_),
    .A1(net950),
    .A2(_2068_));
 sg13g2_o21ai_1 _5999_ (.B1(_2072_),
    .Y(_2073_),
    .A1(net949),
    .A2(_2057_));
 sg13g2_nor2_2 _6000_ (.A(net969),
    .B(net964),
    .Y(_2074_));
 sg13g2_nand2_2 _6001_ (.Y(_2075_),
    .A(net940),
    .B(net939));
 sg13g2_nor2_2 _6002_ (.A(net953),
    .B(net944),
    .Y(_2076_));
 sg13g2_or2_2 _6003_ (.X(_2077_),
    .B(net944),
    .A(net954));
 sg13g2_nor2_2 _6004_ (.A(net953),
    .B(net949),
    .Y(_2078_));
 sg13g2_or2_1 _6005_ (.X(_2079_),
    .B(net949),
    .A(net957));
 sg13g2_and2_2 _6006_ (.A(net952),
    .B(net947),
    .X(_2080_));
 sg13g2_nand2_2 _6007_ (.Y(_2081_),
    .A(net950),
    .B(net944));
 sg13g2_nor2_1 _6008_ (.A(net955),
    .B(_2080_),
    .Y(_2082_));
 sg13g2_nand2_1 _6009_ (.Y(_2083_),
    .A(_2057_),
    .B(_2066_));
 sg13g2_and2_2 _6010_ (.A(_2056_),
    .B(net935),
    .X(_2084_));
 sg13g2_nand2_2 _6011_ (.Y(_2085_),
    .A(_2056_),
    .B(net935));
 sg13g2_nand2_2 _6012_ (.Y(_2086_),
    .A(_2083_),
    .B(_2084_));
 sg13g2_o21ai_1 _6013_ (.B1(_2086_),
    .Y(_2087_),
    .A1(_2047_),
    .A2(_2080_));
 sg13g2_a221oi_1 _6014_ (.B2(_2087_),
    .C1(net972),
    .B1(_2074_),
    .A1(_2063_),
    .Y(_2088_),
    .A2(_2073_));
 sg13g2_nand2b_1 _6015_ (.Y(_2089_),
    .B(_2088_),
    .A_N(_2062_));
 sg13g2_nor2_2 _6016_ (.A(net942),
    .B(net950),
    .Y(_2090_));
 sg13g2_or2_2 _6017_ (.X(_2091_),
    .B(net949),
    .A(net941));
 sg13g2_nand2_1 _6018_ (.Y(_2092_),
    .A(net959),
    .B(_2091_));
 sg13g2_nand2b_1 _6019_ (.Y(_2093_),
    .B(net947),
    .A_N(net943));
 sg13g2_nand2_2 _6020_ (.Y(_2094_),
    .A(net944),
    .B(_2071_));
 sg13g2_mux2_1 _6021_ (.A0(net944),
    .A1(_2094_),
    .S(_2092_),
    .X(_2095_));
 sg13g2_a221oi_1 _6022_ (.B2(net957),
    .C1(net967),
    .B1(_2095_),
    .A1(_2053_),
    .Y(_2096_),
    .A2(_2093_));
 sg13g2_and2_2 _6023_ (.A(net941),
    .B(net949),
    .X(_2097_));
 sg13g2_nand2_2 _6024_ (.Y(_2098_),
    .A(net941),
    .B(net949));
 sg13g2_a221oi_1 _6025_ (.B2(_2083_),
    .C1(net959),
    .B1(_2098_),
    .A1(_2076_),
    .Y(_2099_),
    .A2(_2091_));
 sg13g2_nor2_1 _6026_ (.A(net941),
    .B(net934),
    .Y(_2100_));
 sg13g2_nand2_1 _6027_ (.Y(_2101_),
    .A(net959),
    .B(_2049_));
 sg13g2_o21ai_1 _6028_ (.B1(net966),
    .Y(_2102_),
    .A1(_2100_),
    .A2(_2101_));
 sg13g2_o21ai_1 _6029_ (.B1(net972),
    .Y(_2103_),
    .A1(_2099_),
    .A2(_2102_));
 sg13g2_o21ai_1 _6030_ (.B1(_2089_),
    .Y(_2104_),
    .A1(_2096_),
    .A2(_2103_));
 sg13g2_nor2_2 _6031_ (.A(net1155),
    .B(net1067),
    .Y(_2105_));
 sg13g2_nor2b_2 _6032_ (.A(net944),
    .B_N(net941),
    .Y(_2106_));
 sg13g2_nor2_1 _6033_ (.A(net936),
    .B(_2106_),
    .Y(_2107_));
 sg13g2_or2_1 _6034_ (.X(_2108_),
    .B(_2106_),
    .A(net936));
 sg13g2_nand2_1 _6035_ (.Y(_2109_),
    .A(net938),
    .B(_2107_));
 sg13g2_o21ai_1 _6036_ (.B1(net961),
    .Y(_2110_),
    .A1(net951),
    .A2(_2077_));
 sg13g2_inv_1 _6037_ (.Y(_2111_),
    .A(_2110_));
 sg13g2_nand2_2 _6038_ (.Y(_2112_),
    .A(net955),
    .B(_2081_));
 sg13g2_nor2_1 _6039_ (.A(_2097_),
    .B(_2112_),
    .Y(_2113_));
 sg13g2_o21ai_1 _6040_ (.B1(_2109_),
    .Y(_2114_),
    .A1(_2110_),
    .A2(_2113_));
 sg13g2_nand2_1 _6041_ (.Y(_2115_),
    .A(_2071_),
    .B(_2081_));
 sg13g2_nand2_2 _6042_ (.Y(_2116_),
    .A(net937),
    .B(_2091_));
 sg13g2_nand2_1 _6043_ (.Y(_2117_),
    .A(net937),
    .B(_2115_));
 sg13g2_nand3_1 _6044_ (.B(_2114_),
    .C(_2117_),
    .A(net966),
    .Y(_2118_));
 sg13g2_and2_2 _6045_ (.A(net945),
    .B(_2097_),
    .X(_2119_));
 sg13g2_nand2_2 _6046_ (.Y(_2120_),
    .A(net945),
    .B(_2097_));
 sg13g2_nor2_2 _6047_ (.A(_2090_),
    .B(_2119_),
    .Y(_2121_));
 sg13g2_o21ai_1 _6048_ (.B1(net964),
    .Y(_2122_),
    .A1(net956),
    .A2(_2056_));
 sg13g2_nand2b_1 _6049_ (.Y(_2123_),
    .B(net940),
    .A_N(_2122_));
 sg13g2_nor2_2 _6050_ (.A(net936),
    .B(_2090_),
    .Y(_2124_));
 sg13g2_a21oi_1 _6051_ (.A1(_2056_),
    .A2(_2065_),
    .Y(_2125_),
    .B1(_2123_));
 sg13g2_nand2_1 _6052_ (.Y(_2126_),
    .A(_2121_),
    .B(_2125_));
 sg13g2_nand3_1 _6053_ (.B(net935),
    .C(_2098_),
    .A(_2057_),
    .Y(_2127_));
 sg13g2_and2_1 _6054_ (.A(net954),
    .B(_2071_),
    .X(_2128_));
 sg13g2_nand2_2 _6055_ (.Y(_2129_),
    .A(net953),
    .B(_2071_));
 sg13g2_nand3_1 _6056_ (.B(_2127_),
    .C(_2129_),
    .A(_2074_),
    .Y(_2130_));
 sg13g2_nand3_1 _6057_ (.B(_2126_),
    .C(_2130_),
    .A(_2118_),
    .Y(_2131_));
 sg13g2_nor2_2 _6058_ (.A(_2966_),
    .B(net971),
    .Y(_2132_));
 sg13g2_o21ai_1 _6059_ (.B1(net938),
    .Y(_2133_),
    .A1(_2046_),
    .A2(_2119_));
 sg13g2_nor2_1 _6060_ (.A(_2044_),
    .B(_2080_),
    .Y(_2134_));
 sg13g2_nand2_1 _6061_ (.Y(_2135_),
    .A(_2045_),
    .B(_2081_));
 sg13g2_o21ai_1 _6062_ (.B1(_2116_),
    .Y(_2136_),
    .A1(_2085_),
    .A2(_2135_));
 sg13g2_nand2_1 _6063_ (.Y(_2137_),
    .A(_2076_),
    .B(_2097_));
 sg13g2_nand3_1 _6064_ (.B(_2136_),
    .C(_2137_),
    .A(net960),
    .Y(_2138_));
 sg13g2_nand2_1 _6065_ (.Y(_2139_),
    .A(_2133_),
    .B(_2138_));
 sg13g2_o21ai_1 _6066_ (.B1(net960),
    .Y(_2140_),
    .A1(net945),
    .A2(_2049_));
 sg13g2_nor2_2 _6067_ (.A(net969),
    .B(net973),
    .Y(_2141_));
 sg13g2_o21ai_1 _6068_ (.B1(_2141_),
    .Y(_2142_),
    .A1(_2047_),
    .A2(_2080_));
 sg13g2_nor2_1 _6069_ (.A(net971),
    .B(_2075_),
    .Y(_2143_));
 sg13g2_nor2_1 _6070_ (.A(net942),
    .B(_2081_),
    .Y(_2144_));
 sg13g2_and2_1 _6071_ (.A(net937),
    .B(_2071_),
    .X(_2145_));
 sg13g2_nand2_1 _6072_ (.Y(_2146_),
    .A(_2081_),
    .B(_2145_));
 sg13g2_o21ai_1 _6073_ (.B1(_2146_),
    .Y(_2147_),
    .A1(_2058_),
    .A2(_2144_));
 sg13g2_a22oi_1 _6074_ (.Y(_2148_),
    .B1(_2143_),
    .B2(_2147_),
    .A2(_2139_),
    .A1(_2132_));
 sg13g2_o21ai_1 _6075_ (.B1(net975),
    .Y(_2149_),
    .A1(_2140_),
    .A2(_2142_));
 sg13g2_a21oi_1 _6076_ (.A1(net972),
    .A2(_2131_),
    .Y(_2150_),
    .B1(_2149_));
 sg13g2_a22oi_1 _6077_ (.Y(_2151_),
    .B1(_2148_),
    .B2(_2150_),
    .A2(_2104_),
    .A1(_2969_));
 sg13g2_nand2_1 _6078_ (.Y(_2152_),
    .A(_2105_),
    .B(_2151_));
 sg13g2_nand2b_1 _6079_ (.Y(_2153_),
    .B(_1868_),
    .A_N(net334));
 sg13g2_nand3_1 _6080_ (.B(_1869_),
    .C(_2153_),
    .A(_0136_),
    .Y(_2154_));
 sg13g2_o21ai_1 _6081_ (.B1(_2154_),
    .Y(_0192_),
    .A1(_1369_),
    .A2(_2152_));
 sg13g2_nand2_1 _6082_ (.Y(_2155_),
    .A(_0136_),
    .B(_1936_));
 sg13g2_nand3_1 _6083_ (.B(_2045_),
    .C(net934),
    .A(net942),
    .Y(_2156_));
 sg13g2_a21oi_1 _6084_ (.A1(net936),
    .A2(_2049_),
    .Y(_2157_),
    .B1(net938));
 sg13g2_and2_1 _6085_ (.A(net938),
    .B(_2071_),
    .X(_2158_));
 sg13g2_a22oi_1 _6086_ (.Y(_2159_),
    .B1(_2158_),
    .B2(_2070_),
    .A2(_2157_),
    .A1(_2156_));
 sg13g2_nor2_1 _6087_ (.A(_2078_),
    .B(_2085_),
    .Y(_2160_));
 sg13g2_a22oi_1 _6088_ (.Y(_2161_),
    .B1(_2091_),
    .B2(_2160_),
    .A2(_2078_),
    .A1(net944));
 sg13g2_o21ai_1 _6089_ (.B1(_2137_),
    .Y(_2162_),
    .A1(net937),
    .A2(_2091_));
 sg13g2_o21ai_1 _6090_ (.B1(net971),
    .Y(_2163_),
    .A1(_2075_),
    .A2(_2162_));
 sg13g2_a221oi_1 _6091_ (.B2(_2063_),
    .C1(_2163_),
    .B1(_2161_),
    .A1(net966),
    .Y(_2164_),
    .A2(_2159_));
 sg13g2_nand2_1 _6092_ (.Y(_2165_),
    .A(net951),
    .B(_2085_));
 sg13g2_nand3_1 _6093_ (.B(_2098_),
    .C(_2115_),
    .A(net953),
    .Y(_2166_));
 sg13g2_a21oi_1 _6094_ (.A1(_2145_),
    .A2(_2165_),
    .Y(_2167_),
    .B1(net938));
 sg13g2_a21oi_2 _6095_ (.B1(net960),
    .Y(_2168_),
    .A2(_2048_),
    .A1(\i_music.i_sample.t1.genblk1[2].state.Q ));
 sg13g2_a22oi_1 _6096_ (.Y(_2169_),
    .B1(_2168_),
    .B2(_2127_),
    .A2(_2167_),
    .A1(_2166_));
 sg13g2_nand2b_2 _6097_ (.Y(_2170_),
    .B(_2090_),
    .A_N(net946));
 sg13g2_nand3_1 _6098_ (.B(_2120_),
    .C(_2170_),
    .A(net956),
    .Y(_2171_));
 sg13g2_a21oi_1 _6099_ (.A1(net942),
    .A2(_2134_),
    .Y(_2172_),
    .B1(net938));
 sg13g2_a221oi_1 _6100_ (.B2(net953),
    .C1(net959),
    .B1(_2115_),
    .A1(_2076_),
    .Y(_2173_),
    .A2(_2098_));
 sg13g2_a21oi_1 _6101_ (.A1(_2171_),
    .A2(_2172_),
    .Y(_2174_),
    .B1(_2173_));
 sg13g2_a221oi_1 _6102_ (.B2(_2141_),
    .C1(_2164_),
    .B1(_2174_),
    .A1(_2132_),
    .Y(_2175_),
    .A2(_2169_));
 sg13g2_nand2_2 _6103_ (.Y(_2176_),
    .A(net962),
    .B(_2077_));
 sg13g2_a21oi_1 _6104_ (.A1(net946),
    .A2(_2128_),
    .Y(_2177_),
    .B1(_2176_));
 sg13g2_nand2_2 _6105_ (.Y(_2178_),
    .A(net956),
    .B(_2124_));
 sg13g2_a221oi_1 _6106_ (.B2(_2079_),
    .C1(net962),
    .B1(_2178_),
    .A1(_2066_),
    .Y(_2179_),
    .A2(_2085_));
 sg13g2_o21ai_1 _6107_ (.B1(net966),
    .Y(_2180_),
    .A1(_2177_),
    .A2(_2179_));
 sg13g2_nor2_1 _6108_ (.A(net946),
    .B(_2050_),
    .Y(_2181_));
 sg13g2_nor2_1 _6109_ (.A(net955),
    .B(_2121_),
    .Y(_2182_));
 sg13g2_o21ai_1 _6110_ (.B1(_2074_),
    .Y(_2183_),
    .A1(_2181_),
    .A2(_2182_));
 sg13g2_nand2_1 _6111_ (.Y(_2184_),
    .A(_2063_),
    .B(_2086_));
 sg13g2_nand4_1 _6112_ (.B(_2180_),
    .C(_2183_),
    .A(net972),
    .Y(_2185_),
    .D(_2184_));
 sg13g2_nand2_1 _6113_ (.Y(_2186_),
    .A(net935),
    .B(_2134_));
 sg13g2_a21oi_1 _6114_ (.A1(_2070_),
    .A2(_2186_),
    .Y(_2187_),
    .B1(net960));
 sg13g2_a22oi_1 _6115_ (.Y(_2188_),
    .B1(_2119_),
    .B2(net954),
    .A2(_2084_),
    .A1(_2065_));
 sg13g2_nand2b_1 _6116_ (.Y(_2189_),
    .B(_2188_),
    .A_N(_2055_));
 sg13g2_nor2b_1 _6117_ (.A(_2187_),
    .B_N(_2189_),
    .Y(_2190_));
 sg13g2_o21ai_1 _6118_ (.B1(net960),
    .Y(_2191_),
    .A1(_2084_),
    .A2(_2116_));
 sg13g2_nor2_1 _6119_ (.A(net959),
    .B(_2100_),
    .Y(_2192_));
 sg13g2_nand3_1 _6120_ (.B(_2129_),
    .C(_2192_),
    .A(_2057_),
    .Y(_2193_));
 sg13g2_a22oi_1 _6121_ (.Y(_2194_),
    .B1(_2191_),
    .B2(_2193_),
    .A2(_2134_),
    .A1(_2128_));
 sg13g2_a221oi_1 _6122_ (.B2(_2132_),
    .C1(_2969_),
    .B1(_2194_),
    .A1(_2141_),
    .Y(_2195_),
    .A2(_2190_));
 sg13g2_o21ai_1 _6123_ (.B1(_2105_),
    .Y(_2196_),
    .A1(net975),
    .A2(_2175_));
 sg13g2_a21o_1 _6124_ (.A2(_2195_),
    .A1(_2185_),
    .B1(_2196_),
    .X(_2197_));
 sg13g2_o21ai_1 _6125_ (.B1(_2155_),
    .Y(_0193_),
    .A1(_1369_),
    .A2(_2197_));
 sg13g2_o21ai_1 _6126_ (.B1(_2050_),
    .Y(_2198_),
    .A1(_2078_),
    .A2(_2085_));
 sg13g2_nor2_1 _6127_ (.A(net963),
    .B(_2121_),
    .Y(_2199_));
 sg13g2_o21ai_1 _6128_ (.B1(net968),
    .Y(_2200_),
    .A1(net939),
    .A2(_2198_));
 sg13g2_a21oi_1 _6129_ (.A1(_2198_),
    .A2(_2199_),
    .Y(_2201_),
    .B1(_2200_));
 sg13g2_a21oi_1 _6130_ (.A1(net951),
    .A2(_2085_),
    .Y(_2202_),
    .B1(net937));
 sg13g2_nand2_1 _6131_ (.Y(_2203_),
    .A(net955),
    .B(_2165_));
 sg13g2_a22oi_1 _6132_ (.Y(_2204_),
    .B1(_2192_),
    .B2(_2203_),
    .A2(_2171_),
    .A1(_2111_));
 sg13g2_nor2_1 _6133_ (.A(net966),
    .B(_2204_),
    .Y(_2205_));
 sg13g2_o21ai_1 _6134_ (.B1(net972),
    .Y(_2206_),
    .A1(_2201_),
    .A2(_2205_));
 sg13g2_nor2_1 _6135_ (.A(_2077_),
    .B(_2091_),
    .Y(_2207_));
 sg13g2_nand3_1 _6136_ (.B(_2094_),
    .C(_2107_),
    .A(net954),
    .Y(_2208_));
 sg13g2_nand2b_1 _6137_ (.Y(_2209_),
    .B(_2208_),
    .A_N(_2207_));
 sg13g2_o21ai_1 _6138_ (.B1(_2049_),
    .Y(_2210_),
    .A1(net936),
    .A2(_2097_));
 sg13g2_o21ai_1 _6139_ (.B1(net966),
    .Y(_2211_),
    .A1(net959),
    .A2(_2210_));
 sg13g2_a21oi_1 _6140_ (.A1(net961),
    .A2(_2209_),
    .Y(_2212_),
    .B1(_2211_));
 sg13g2_a221oi_1 _6141_ (.B2(_2085_),
    .C1(_2075_),
    .B1(_2078_),
    .A1(_2056_),
    .Y(_2213_),
    .A2(_2059_));
 sg13g2_nor2_1 _6142_ (.A(net951),
    .B(_2056_),
    .Y(_2214_));
 sg13g2_nor2_1 _6143_ (.A(_2076_),
    .B(_2214_),
    .Y(_2215_));
 sg13g2_a21oi_1 _6144_ (.A1(_2129_),
    .A2(_2215_),
    .Y(_2216_),
    .B1(_2064_));
 sg13g2_or4_1 _6145_ (.A(net971),
    .B(_2212_),
    .C(_2213_),
    .D(_2216_),
    .X(_2217_));
 sg13g2_nand3_1 _6146_ (.B(_2206_),
    .C(_2217_),
    .A(net975),
    .Y(_2218_));
 sg13g2_nand3_1 _6147_ (.B(_2077_),
    .C(_2090_),
    .A(net962),
    .Y(_2219_));
 sg13g2_a21o_1 _6148_ (.A2(_2145_),
    .A1(net935),
    .B1(net961),
    .X(_2220_));
 sg13g2_a22oi_1 _6149_ (.Y(_2221_),
    .B1(_2220_),
    .B2(_2176_),
    .A2(_2219_),
    .A1(_2202_));
 sg13g2_nand3_1 _6150_ (.B(net950),
    .C(net946),
    .A(net955),
    .Y(_2222_));
 sg13g2_nor2b_1 _6151_ (.A(_2082_),
    .B_N(_2222_),
    .Y(_2223_));
 sg13g2_o21ai_1 _6152_ (.B1(_2049_),
    .Y(_2224_),
    .A1(_2106_),
    .A2(_2223_));
 sg13g2_o21ai_1 _6153_ (.B1(net966),
    .Y(_2225_),
    .A1(net962),
    .A2(_2059_));
 sg13g2_nand3_1 _6154_ (.B(_2082_),
    .C(_2084_),
    .A(net966),
    .Y(_2226_));
 sg13g2_a22oi_1 _6155_ (.Y(_2227_),
    .B1(_2225_),
    .B2(_2226_),
    .A2(_2224_),
    .A1(net962));
 sg13g2_nor2_1 _6156_ (.A(net971),
    .B(_2227_),
    .Y(_2228_));
 sg13g2_o21ai_1 _6157_ (.B1(_2228_),
    .Y(_2229_),
    .A1(net968),
    .A2(_2221_));
 sg13g2_nor3_1 _6158_ (.A(_2068_),
    .B(_2182_),
    .C(_2214_),
    .Y(_2230_));
 sg13g2_o21ai_1 _6159_ (.B1(_2063_),
    .Y(_2231_),
    .A1(_2207_),
    .A2(_2230_));
 sg13g2_nor2_1 _6160_ (.A(_2080_),
    .B(_2178_),
    .Y(_2232_));
 sg13g2_nor2_1 _6161_ (.A(_2078_),
    .B(_2092_),
    .Y(_2233_));
 sg13g2_a21oi_1 _6162_ (.A1(_2085_),
    .A2(_2233_),
    .Y(_2234_),
    .B1(net940));
 sg13g2_o21ai_1 _6163_ (.B1(_2234_),
    .Y(_2235_),
    .A1(_2220_),
    .A2(_2232_));
 sg13g2_nor2_1 _6164_ (.A(_2075_),
    .B(_2182_),
    .Y(_2236_));
 sg13g2_o21ai_1 _6165_ (.B1(_2236_),
    .Y(_2237_),
    .A1(net941),
    .A2(_2222_));
 sg13g2_nand4_1 _6166_ (.B(_2231_),
    .C(_2235_),
    .A(net971),
    .Y(_2238_),
    .D(_2237_));
 sg13g2_nand3_1 _6167_ (.B(_2229_),
    .C(_2238_),
    .A(_2969_),
    .Y(_2239_));
 sg13g2_nand4_1 _6168_ (.B(_2105_),
    .C(_2218_),
    .A(net982),
    .Y(_2240_),
    .D(_2239_));
 sg13g2_o21ai_1 _6169_ (.B1(_2240_),
    .Y(_0194_),
    .A1(_1573_),
    .A2(_1937_));
 sg13g2_nand3_1 _6170_ (.B(net934),
    .C(_2188_),
    .A(net960),
    .Y(_2241_));
 sg13g2_nand3_1 _6171_ (.B(_2116_),
    .C(_2168_),
    .A(_2077_),
    .Y(_2242_));
 sg13g2_nand3_1 _6172_ (.B(_2241_),
    .C(_2242_),
    .A(net967),
    .Y(_2243_));
 sg13g2_a21o_1 _6173_ (.A2(_2108_),
    .A1(net953),
    .B1(_2220_),
    .X(_2244_));
 sg13g2_a21oi_1 _6174_ (.A1(net937),
    .A2(_2097_),
    .Y(_2245_),
    .B1(_2080_));
 sg13g2_nand3_1 _6175_ (.B(_2070_),
    .C(_2245_),
    .A(net959),
    .Y(_2246_));
 sg13g2_nand3_1 _6176_ (.B(_2244_),
    .C(_2246_),
    .A(net940),
    .Y(_2247_));
 sg13g2_nand3_1 _6177_ (.B(_2243_),
    .C(_2247_),
    .A(net971),
    .Y(_2248_));
 sg13g2_nand2b_1 _6178_ (.Y(_2249_),
    .B(_2066_),
    .A_N(_2053_));
 sg13g2_nor4_1 _6179_ (.A(net961),
    .B(_2068_),
    .C(_2119_),
    .D(_2249_),
    .Y(_2250_));
 sg13g2_o21ai_1 _6180_ (.B1(_2067_),
    .Y(_2251_),
    .A1(_2065_),
    .A2(net935));
 sg13g2_nor2_1 _6181_ (.A(_2140_),
    .B(_2251_),
    .Y(_2252_));
 sg13g2_nor2_1 _6182_ (.A(_2250_),
    .B(_2252_),
    .Y(_2253_));
 sg13g2_nand3_1 _6183_ (.B(_2056_),
    .C(_2067_),
    .A(net954),
    .Y(_2254_));
 sg13g2_nor2_2 _6184_ (.A(net956),
    .B(net936),
    .Y(_2255_));
 sg13g2_o21ai_1 _6185_ (.B1(_2254_),
    .Y(_2256_),
    .A1(_2044_),
    .A2(_2116_));
 sg13g2_o21ai_1 _6186_ (.B1(_2077_),
    .Y(_2257_),
    .A1(_2058_),
    .A2(_2144_));
 sg13g2_a221oi_1 _6187_ (.B2(_2063_),
    .C1(net972),
    .B1(_2257_),
    .A1(net967),
    .Y(_2258_),
    .A2(_2253_));
 sg13g2_o21ai_1 _6188_ (.B1(_2258_),
    .Y(_2259_),
    .A1(_2075_),
    .A2(_2256_));
 sg13g2_nand3_1 _6189_ (.B(_2248_),
    .C(_2259_),
    .A(_2969_),
    .Y(_2260_));
 sg13g2_nor2b_1 _6190_ (.A(_2121_),
    .B_N(_2249_),
    .Y(_2261_));
 sg13g2_nor2_1 _6191_ (.A(net936),
    .B(_2261_),
    .Y(_2262_));
 sg13g2_nand2_1 _6192_ (.Y(_2263_),
    .A(net963),
    .B(_2262_));
 sg13g2_nor2_1 _6193_ (.A(_2181_),
    .B(_2263_),
    .Y(_2264_));
 sg13g2_a221oi_1 _6194_ (.B2(_2165_),
    .C1(net962),
    .B1(_2145_),
    .A1(net955),
    .Y(_2265_),
    .A2(_2120_));
 sg13g2_o21ai_1 _6195_ (.B1(_2132_),
    .Y(_2266_),
    .A1(_2264_),
    .A2(_2265_));
 sg13g2_a21oi_1 _6196_ (.A1(net948),
    .A2(_2065_),
    .Y(_2267_),
    .B1(net961));
 sg13g2_o21ai_1 _6197_ (.B1(_2267_),
    .Y(_2268_),
    .A1(_2069_),
    .A2(_2249_));
 sg13g2_nand3b_1 _6198_ (.B(_2178_),
    .C(net964),
    .Y(_2269_),
    .A_N(_2144_));
 sg13g2_a21oi_1 _6199_ (.A1(_2268_),
    .A2(_2269_),
    .Y(_2270_),
    .B1(_2966_));
 sg13g2_nor3_1 _6200_ (.A(_2075_),
    .B(_2113_),
    .C(_2255_),
    .Y(_2271_));
 sg13g2_o21ai_1 _6201_ (.B1(net971),
    .Y(_2272_),
    .A1(_2270_),
    .A2(_2271_));
 sg13g2_nand3_1 _6202_ (.B(_2094_),
    .C(_2107_),
    .A(net937),
    .Y(_2273_));
 sg13g2_nand2_1 _6203_ (.Y(_2274_),
    .A(_2067_),
    .B(_2128_));
 sg13g2_a21oi_1 _6204_ (.A1(_2273_),
    .A2(_2274_),
    .Y(_2275_),
    .B1(net939));
 sg13g2_a21oi_1 _6205_ (.A1(_2091_),
    .A2(_2255_),
    .Y(_2276_),
    .B1(net960));
 sg13g2_o21ai_1 _6206_ (.B1(_2276_),
    .Y(_2277_),
    .A1(_2068_),
    .A2(_2129_));
 sg13g2_nand3b_1 _6207_ (.B(_2277_),
    .C(_2141_),
    .Y(_2278_),
    .A_N(_2275_));
 sg13g2_nand4_1 _6208_ (.B(_2266_),
    .C(_2272_),
    .A(net975),
    .Y(_2279_),
    .D(_2278_));
 sg13g2_nand4_1 _6209_ (.B(_2105_),
    .C(_2260_),
    .A(net982),
    .Y(_2280_),
    .D(_2279_));
 sg13g2_o21ai_1 _6210_ (.B1(_2280_),
    .Y(_0195_),
    .A1(_1573_),
    .A2(_1939_));
 sg13g2_nand2_1 _6211_ (.Y(_2281_),
    .A(_2120_),
    .B(_2255_));
 sg13g2_o21ai_1 _6212_ (.B1(_2281_),
    .Y(_2282_),
    .A1(_2080_),
    .A2(_2178_));
 sg13g2_a21oi_1 _6213_ (.A1(_2048_),
    .A2(_2080_),
    .Y(_2283_),
    .B1(net960));
 sg13g2_a22oi_1 _6214_ (.Y(_2284_),
    .B1(_2283_),
    .B2(_2281_),
    .A2(_2282_),
    .A1(net964));
 sg13g2_a21oi_1 _6215_ (.A1(net956),
    .A2(_2170_),
    .Y(_2285_),
    .B1(_2123_));
 sg13g2_a221oi_1 _6216_ (.B2(net969),
    .C1(_2285_),
    .B1(_2284_),
    .A1(_2074_),
    .Y(_2286_),
    .A2(_2124_));
 sg13g2_nor2_1 _6217_ (.A(net973),
    .B(_2286_),
    .Y(_2287_));
 sg13g2_nor2_1 _6218_ (.A(_2078_),
    .B(_2176_),
    .Y(_2288_));
 sg13g2_inv_1 _6219_ (.Y(_2289_),
    .A(_2288_));
 sg13g2_a21oi_1 _6220_ (.A1(_2178_),
    .A2(_2288_),
    .Y(_2290_),
    .B1(_2225_));
 sg13g2_o21ai_1 _6221_ (.B1(_2074_),
    .Y(_2291_),
    .A1(net946),
    .A2(net934));
 sg13g2_nor2b_1 _6222_ (.A(_2290_),
    .B_N(net974),
    .Y(_2292_));
 sg13g2_a21oi_1 _6223_ (.A1(_2291_),
    .A2(_2292_),
    .Y(_2293_),
    .B1(_2287_));
 sg13g2_nor2_1 _6224_ (.A(net963),
    .B(_2112_),
    .Y(_2294_));
 sg13g2_nor2b_1 _6225_ (.A(_2122_),
    .B_N(_2124_),
    .Y(_2295_));
 sg13g2_o21ai_1 _6226_ (.B1(net969),
    .Y(_2296_),
    .A1(_2294_),
    .A2(_2295_));
 sg13g2_nand3_1 _6227_ (.B(_2112_),
    .C(_2273_),
    .A(_2074_),
    .Y(_2297_));
 sg13g2_a21oi_1 _6228_ (.A1(net950),
    .A2(net935),
    .Y(_2298_),
    .B1(net955));
 sg13g2_o21ai_1 _6229_ (.B1(_2063_),
    .Y(_2299_),
    .A1(_2181_),
    .A2(_2298_));
 sg13g2_nand4_1 _6230_ (.B(_2296_),
    .C(_2297_),
    .A(net974),
    .Y(_2300_),
    .D(_2299_));
 sg13g2_o21ai_1 _6231_ (.B1(net967),
    .Y(_2301_),
    .A1(_2065_),
    .A2(_2255_));
 sg13g2_nand2_1 _6232_ (.Y(_2302_),
    .A(net940),
    .B(_2066_));
 sg13g2_or2_1 _6233_ (.X(_2303_),
    .B(_2302_),
    .A(_2135_));
 sg13g2_nand3_1 _6234_ (.B(_2301_),
    .C(_2303_),
    .A(net964),
    .Y(_2304_));
 sg13g2_nand3_1 _6235_ (.B(_2120_),
    .C(_2302_),
    .A(net956),
    .Y(_2305_));
 sg13g2_a21oi_1 _6236_ (.A1(_2276_),
    .A2(_2305_),
    .Y(_2306_),
    .B1(net973));
 sg13g2_a21oi_1 _6237_ (.A1(_2304_),
    .A2(_2306_),
    .Y(_2307_),
    .B1(net975));
 sg13g2_a22oi_1 _6238_ (.Y(_2308_),
    .B1(_2300_),
    .B2(_2307_),
    .A2(_2293_),
    .A1(net976));
 sg13g2_nor2b_1 _6239_ (.A(_2308_),
    .B_N(_2105_),
    .Y(_2309_));
 sg13g2_a22oi_1 _6240_ (.Y(_2310_),
    .B1(_2309_),
    .B2(net983),
    .A2(_1941_),
    .A1(_0136_));
 sg13g2_inv_1 _6241_ (.Y(_0196_),
    .A(_2310_));
 sg13g2_or2_1 _6242_ (.X(_2311_),
    .B(_1943_),
    .A(_1573_));
 sg13g2_a21o_1 _6243_ (.A2(_2178_),
    .A1(net934),
    .B1(net938),
    .X(_2312_));
 sg13g2_o21ai_1 _6244_ (.B1(_2312_),
    .Y(_2313_),
    .A1(net963),
    .A2(_2968_));
 sg13g2_nand3_1 _6245_ (.B(_2063_),
    .C(net935),
    .A(_2053_),
    .Y(_2314_));
 sg13g2_nor2_1 _6246_ (.A(net968),
    .B(_2112_),
    .Y(_2315_));
 sg13g2_a21oi_1 _6247_ (.A1(net968),
    .A2(_2313_),
    .Y(_2316_),
    .B1(_2315_));
 sg13g2_nand3_1 _6248_ (.B(_2314_),
    .C(_2316_),
    .A(net972),
    .Y(_2317_));
 sg13g2_o21ai_1 _6249_ (.B1(net940),
    .Y(_2318_),
    .A1(net962),
    .A2(_2050_));
 sg13g2_nand2_1 _6250_ (.Y(_2319_),
    .A(_2110_),
    .B(_2318_));
 sg13g2_o21ai_1 _6251_ (.B1(_2319_),
    .Y(_2320_),
    .A1(_2064_),
    .A2(_2223_));
 sg13g2_o21ai_1 _6252_ (.B1(_2317_),
    .Y(_2321_),
    .A1(net973),
    .A2(_2320_));
 sg13g2_o21ai_1 _6253_ (.B1(_2262_),
    .Y(_2322_),
    .A1(net963),
    .A2(_2968_));
 sg13g2_a21oi_1 _6254_ (.A1(net968),
    .A2(_2288_),
    .Y(_2323_),
    .B1(_2074_));
 sg13g2_nand4_1 _6255_ (.B(net934),
    .C(_2141_),
    .A(net964),
    .Y(_2324_),
    .D(_2170_));
 sg13g2_nand3_1 _6256_ (.B(_2141_),
    .C(_2178_),
    .A(net939),
    .Y(_2325_));
 sg13g2_nand3_1 _6257_ (.B(_2324_),
    .C(_2325_),
    .A(net976),
    .Y(_2326_));
 sg13g2_a221oi_1 _6258_ (.B2(net973),
    .C1(_2326_),
    .B1(_2323_),
    .A1(_2132_),
    .Y(_2327_),
    .A2(_2322_));
 sg13g2_a21oi_1 _6259_ (.A1(_2969_),
    .A2(_2321_),
    .Y(_2328_),
    .B1(_2327_));
 sg13g2_nand2b_1 _6260_ (.Y(_2329_),
    .B(_2105_),
    .A_N(_2328_));
 sg13g2_o21ai_1 _6261_ (.B1(_2311_),
    .Y(_0197_),
    .A1(_1369_),
    .A2(_2329_));
 sg13g2_a22oi_1 _6262_ (.Y(_2330_),
    .B1(_2063_),
    .B2(net934),
    .A2(net973),
    .A1(net962));
 sg13g2_nand2_1 _6263_ (.Y(_2331_),
    .A(net975),
    .B(_2330_));
 sg13g2_a21oi_1 _6264_ (.A1(net968),
    .A2(_2263_),
    .Y(_2332_),
    .B1(_2331_));
 sg13g2_a21oi_1 _6265_ (.A1(net963),
    .A2(net934),
    .Y(_2333_),
    .B1(net940));
 sg13g2_nor2_1 _6266_ (.A(_2315_),
    .B(_2333_),
    .Y(_2334_));
 sg13g2_o21ai_1 _6267_ (.B1(_2334_),
    .Y(_2335_),
    .A1(_2064_),
    .A2(_2298_));
 sg13g2_a221oi_1 _6268_ (.B2(net973),
    .C1(net975),
    .B1(_2335_),
    .A1(_2141_),
    .Y(_2336_),
    .A2(_2289_));
 sg13g2_o21ai_1 _6269_ (.B1(net982),
    .Y(_2337_),
    .A1(_2332_),
    .A2(_2336_));
 sg13g2_a22oi_1 _6270_ (.Y(_2338_),
    .B1(_2105_),
    .B2(_2337_),
    .A2(_1945_),
    .A1(_0136_));
 sg13g2_inv_1 _6271_ (.Y(_0198_),
    .A(_2338_));
 sg13g2_nor2_1 _6272_ (.A(\i_music.violin_note_idx[1][0] ),
    .B(net977),
    .Y(_2339_));
 sg13g2_nor3_1 _6273_ (.A(net230),
    .B(_1547_),
    .C(net981),
    .Y(_2340_));
 sg13g2_nor2_1 _6274_ (.A(_2339_),
    .B(_2340_),
    .Y(_0199_));
 sg13g2_nor2_1 _6275_ (.A(net366),
    .B(_3000_),
    .Y(_2341_));
 sg13g2_nand3_1 _6276_ (.B(net1130),
    .C(_3088_),
    .A(\i_display.i_vga.timing_ver.counter[2] ),
    .Y(_2342_));
 sg13g2_nor4_1 _6277_ (.A(\i_display.i_vga.timing_ver.counter[10] ),
    .B(_2920_),
    .C(\i_display.i_vga.timing_ver.counter[8] ),
    .D(\i_display.i_vga.timing_ver.counter[7] ),
    .Y(_2343_));
 sg13g2_nand4_1 _6278_ (.B(\i_display.i_vga.timing_ver.counter[4] ),
    .C(_1426_),
    .A(\i_display.i_vga.timing_ver.counter[6] ),
    .Y(_2344_),
    .D(_2343_));
 sg13g2_nor2_1 _6279_ (.A(_2342_),
    .B(_2344_),
    .Y(_2345_));
 sg13g2_nor2b_1 _6280_ (.A(_2345_),
    .B_N(_3088_),
    .Y(_2346_));
 sg13g2_o21ai_1 _6281_ (.B1(net1174),
    .Y(_0200_),
    .A1(_2341_),
    .A2(_2346_));
 sg13g2_a21oi_1 _6282_ (.A1(_2922_),
    .A2(_3088_),
    .Y(_2347_),
    .B1(net1159));
 sg13g2_o21ai_1 _6283_ (.B1(_2347_),
    .Y(_0201_),
    .A1(_2922_),
    .A2(_2346_));
 sg13g2_a21o_1 _6284_ (.A2(_3088_),
    .A1(net1130),
    .B1(net270),
    .X(_2348_));
 sg13g2_nand2b_1 _6285_ (.Y(_2349_),
    .B(_2344_),
    .A_N(_2342_));
 sg13g2_a21o_1 _6286_ (.A2(_2349_),
    .A1(_2348_),
    .B1(net1159),
    .X(_0202_));
 sg13g2_and4_1 _6287_ (.A(net212),
    .B(\i_display.i_vga.timing_ver.counter[2] ),
    .C(net1130),
    .D(_3092_),
    .X(_2350_));
 sg13g2_nor2_2 _6288_ (.A(net1159),
    .B(_2345_),
    .Y(_2351_));
 sg13g2_inv_1 _6289_ (.Y(_2352_),
    .A(_2351_));
 sg13g2_nor2b_1 _6290_ (.A(net212),
    .B_N(_2342_),
    .Y(_2353_));
 sg13g2_nor3_1 _6291_ (.A(_2350_),
    .B(_2352_),
    .C(_2353_),
    .Y(_0203_));
 sg13g2_nand2_1 _6292_ (.Y(_2354_),
    .A(\i_display.i_vga.timing_ver.counter[4] ),
    .B(\i_display.i_vga.timing_ver.counter[3] ));
 sg13g2_nor2_1 _6293_ (.A(_2342_),
    .B(_2354_),
    .Y(_2355_));
 sg13g2_xnor2_1 _6294_ (.Y(_2356_),
    .A(net340),
    .B(_2350_));
 sg13g2_nor2_1 _6295_ (.A(_2352_),
    .B(_2356_),
    .Y(_0204_));
 sg13g2_or2_1 _6296_ (.X(_2357_),
    .B(_2355_),
    .A(net378));
 sg13g2_nand2_1 _6297_ (.Y(_2358_),
    .A(net378),
    .B(_2355_));
 sg13g2_a21o_1 _6298_ (.A2(_2358_),
    .A1(_2357_),
    .B1(_2352_),
    .X(_0205_));
 sg13g2_and4_1 _6299_ (.A(\i_display.i_vga.timing_ver.counter[6] ),
    .B(\i_display.i_vga.timing_ver.counter[5] ),
    .C(\i_display.i_vga.timing_ver.counter[4] ),
    .D(_2350_),
    .X(_2359_));
 sg13g2_xor2_1 _6300_ (.B(_2358_),
    .A(net362),
    .X(_2360_));
 sg13g2_nand2_1 _6301_ (.Y(_0206_),
    .A(net1174),
    .B(net363));
 sg13g2_nand2_1 _6302_ (.Y(_2361_),
    .A(net379),
    .B(_2359_));
 sg13g2_or2_1 _6303_ (.X(_2362_),
    .B(_2359_),
    .A(net379));
 sg13g2_a21o_1 _6304_ (.A2(_2362_),
    .A1(_2361_),
    .B1(_2352_),
    .X(_0207_));
 sg13g2_xnor2_1 _6305_ (.Y(_2363_),
    .A(_2921_),
    .B(_2361_));
 sg13g2_nand2_1 _6306_ (.Y(_0208_),
    .A(_2351_),
    .B(_2363_));
 sg13g2_o21ai_1 _6307_ (.B1(_2920_),
    .Y(_2364_),
    .A1(_2921_),
    .A2(_2361_));
 sg13g2_nand4_1 _6308_ (.B(\i_display.i_vga.timing_ver.counter[8] ),
    .C(\i_display.i_vga.timing_ver.counter[7] ),
    .A(net368),
    .Y(_2365_),
    .D(_2359_));
 sg13g2_a21o_1 _6309_ (.A2(net369),
    .A1(_2364_),
    .B1(net1159),
    .X(_0209_));
 sg13g2_xor2_1 _6310_ (.B(_2365_),
    .A(net315),
    .X(_2366_));
 sg13g2_nand2_1 _6311_ (.Y(_0210_),
    .A(_2351_),
    .B(net316));
 sg13g2_nor2_1 _6312_ (.A(net1163),
    .B(net1005),
    .Y(_2367_));
 sg13g2_nand2_1 _6313_ (.Y(_2368_),
    .A(net241),
    .B(net994));
 sg13g2_xnor2_1 _6314_ (.Y(_2369_),
    .A(_0052_),
    .B(_0793_));
 sg13g2_xnor2_1 _6315_ (.Y(_2370_),
    .A(_0049_),
    .B(net1059));
 sg13g2_xnor2_1 _6316_ (.Y(_2371_),
    .A(_0050_),
    .B(_3096_));
 sg13g2_xnor2_1 _6317_ (.Y(_2372_),
    .A(\crotchet[0] ),
    .B(\i_display.frame_crotchet[0] ));
 sg13g2_o21ai_1 _6318_ (.B1(_2372_),
    .Y(_2373_),
    .A1(_0048_),
    .A2(_0775_));
 sg13g2_nand2b_1 _6319_ (.Y(_2374_),
    .B(_0778_),
    .A_N(_0053_));
 sg13g2_xnor2_1 _6320_ (.Y(_2375_),
    .A(_0051_),
    .B(_0781_));
 sg13g2_a22oi_1 _6321_ (.Y(_2376_),
    .B1(net1057),
    .B2(_0053_),
    .A2(_0775_),
    .A1(_0048_));
 sg13g2_nand4_1 _6322_ (.B(_2374_),
    .C(_2375_),
    .A(_2371_),
    .Y(_2377_),
    .D(_2376_));
 sg13g2_nor4_2 _6323_ (.A(_2369_),
    .B(_2370_),
    .C(_2373_),
    .Y(_2378_),
    .D(_2377_));
 sg13g2_nor2_1 _6324_ (.A(net1129),
    .B(_2378_),
    .Y(_2379_));
 sg13g2_a21oi_1 _6325_ (.A1(_0079_),
    .A2(_2378_),
    .Y(_2380_),
    .B1(_2379_));
 sg13g2_o21ai_1 _6326_ (.B1(_0786_),
    .Y(_2381_),
    .A1(_3097_),
    .A2(net1058));
 sg13g2_nand2_1 _6327_ (.Y(_2382_),
    .A(net1058),
    .B(_0812_));
 sg13g2_a21oi_1 _6328_ (.A1(_2381_),
    .A2(_2382_),
    .Y(_2383_),
    .B1(_0841_));
 sg13g2_nor2_1 _6329_ (.A(_0774_),
    .B(_2383_),
    .Y(_2384_));
 sg13g2_a21oi_1 _6330_ (.A1(_0788_),
    .A2(_2381_),
    .Y(_2385_),
    .B1(_0792_));
 sg13g2_o21ai_1 _6331_ (.B1(_0794_),
    .Y(_2386_),
    .A1(_2384_),
    .A2(_2385_));
 sg13g2_o21ai_1 _6332_ (.B1(\crotchet[0] ),
    .Y(_2387_),
    .A1(_3097_),
    .A2(net1058));
 sg13g2_nor4_1 _6333_ (.A(_0775_),
    .B(net1057),
    .C(_0782_),
    .D(_0793_),
    .Y(_2388_));
 sg13g2_nand2_1 _6334_ (.Y(_2389_),
    .A(_2387_),
    .B(_2388_));
 sg13g2_a21oi_2 _6335_ (.B1(_2378_),
    .Y(_2390_),
    .A2(_2389_),
    .A1(_2386_));
 sg13g2_or2_2 _6336_ (.X(_2391_),
    .B(_2390_),
    .A(net1001));
 sg13g2_o21ai_1 _6337_ (.B1(_2368_),
    .Y(_0211_),
    .A1(_2380_),
    .A2(_2391_));
 sg13g2_a21o_1 _6338_ (.A2(_2390_),
    .A1(net1005),
    .B1(net1163),
    .X(_2392_));
 sg13g2_a21oi_1 _6339_ (.A1(net1129),
    .A2(net1005),
    .Y(_2393_),
    .B1(net1128));
 sg13g2_nand2_2 _6340_ (.Y(_2394_),
    .A(net1128),
    .B(net241));
 sg13g2_nor2_1 _6341_ (.A(_3090_),
    .B(_2394_),
    .Y(_2395_));
 sg13g2_nor3_1 _6342_ (.A(_2392_),
    .B(_2393_),
    .C(_2395_),
    .Y(_0212_));
 sg13g2_nand2_1 _6343_ (.Y(_2396_),
    .A(net1125),
    .B(net994));
 sg13g2_nor2_1 _6344_ (.A(_0081_),
    .B(_2394_),
    .Y(_2397_));
 sg13g2_xnor2_1 _6345_ (.Y(_2398_),
    .A(net357),
    .B(_2394_));
 sg13g2_o21ai_1 _6346_ (.B1(_2396_),
    .Y(_0213_),
    .A1(_2391_),
    .A2(_2398_));
 sg13g2_nand2_1 _6347_ (.Y(_2399_),
    .A(net1124),
    .B(net994));
 sg13g2_xnor2_1 _6348_ (.Y(_2400_),
    .A(_2933_),
    .B(_2397_));
 sg13g2_o21ai_1 _6349_ (.B1(_2399_),
    .Y(_0214_),
    .A1(_2391_),
    .A2(_2400_));
 sg13g2_nand3_1 _6350_ (.B(net1126),
    .C(_2395_),
    .A(net1124),
    .Y(_2401_));
 sg13g2_nor2_1 _6351_ (.A(_2916_),
    .B(_2917_),
    .Y(_2402_));
 sg13g2_nor4_2 _6352_ (.A(_2916_),
    .B(_2917_),
    .C(_2918_),
    .Y(_2403_),
    .D(_2394_));
 sg13g2_a221oi_1 _6353_ (.B2(net1005),
    .C1(_2392_),
    .B1(_2403_),
    .A1(_2916_),
    .Y(_0215_),
    .A2(_2401_));
 sg13g2_nand2_1 _6354_ (.Y(_2404_),
    .A(net1119),
    .B(net994));
 sg13g2_xnor2_1 _6355_ (.Y(_2405_),
    .A(_2932_),
    .B(_2403_));
 sg13g2_o21ai_1 _6356_ (.B1(_2404_),
    .Y(_0216_),
    .A1(_2391_),
    .A2(_2405_));
 sg13g2_nand2_1 _6357_ (.Y(_2406_),
    .A(net1117),
    .B(net994));
 sg13g2_nand2_1 _6358_ (.Y(_2407_),
    .A(net1119),
    .B(_2403_));
 sg13g2_nor2_1 _6359_ (.A(net349),
    .B(_2407_),
    .Y(_2408_));
 sg13g2_xnor2_1 _6360_ (.Y(_2409_),
    .A(net349),
    .B(_2407_));
 sg13g2_o21ai_1 _6361_ (.B1(_2406_),
    .Y(_0217_),
    .A1(_2391_),
    .A2(_2409_));
 sg13g2_nand2_1 _6362_ (.Y(_2410_),
    .A(net1116),
    .B(net994));
 sg13g2_xnor2_1 _6363_ (.Y(_2411_),
    .A(_2939_),
    .B(_2408_));
 sg13g2_o21ai_1 _6364_ (.B1(_2410_),
    .Y(_0218_),
    .A1(_2391_),
    .A2(_2411_));
 sg13g2_nand2_1 _6365_ (.Y(_2412_),
    .A(net337),
    .B(net994));
 sg13g2_nand4_1 _6366_ (.B(net1117),
    .C(net1120),
    .A(\i_display.frame[7] ),
    .Y(_2413_),
    .D(_2403_));
 sg13g2_nor2_1 _6367_ (.A(_0095_),
    .B(_2413_),
    .Y(_2414_));
 sg13g2_xnor2_1 _6368_ (.Y(_2415_),
    .A(_0095_),
    .B(_2413_));
 sg13g2_o21ai_1 _6369_ (.B1(_2412_),
    .Y(_0219_),
    .A1(_2391_),
    .A2(_2415_));
 sg13g2_nand2_1 _6370_ (.Y(_2416_),
    .A(net317),
    .B(net994));
 sg13g2_xnor2_1 _6371_ (.Y(_2417_),
    .A(_2942_),
    .B(_2414_));
 sg13g2_o21ai_1 _6372_ (.B1(_2416_),
    .Y(_0220_),
    .A1(_2391_),
    .A2(_2417_));
 sg13g2_nor2b_2 _6373_ (.A(net1135),
    .B_N(net1133),
    .Y(_2418_));
 sg13g2_nor2b_2 _6374_ (.A(net1136),
    .B_N(_2418_),
    .Y(_2419_));
 sg13g2_nand2b_2 _6375_ (.Y(_2420_),
    .B(_2418_),
    .A_N(net1136));
 sg13g2_nor2_2 _6376_ (.A(net1134),
    .B(_0050_),
    .Y(_2421_));
 sg13g2_nor2_1 _6377_ (.A(_2419_),
    .B(_2421_),
    .Y(_2422_));
 sg13g2_or2_2 _6378_ (.X(_2423_),
    .B(_2421_),
    .A(_2419_));
 sg13g2_nand3_1 _6379_ (.B(_0740_),
    .C(_2423_),
    .A(net1123),
    .Y(_2424_));
 sg13g2_a21o_1 _6380_ (.A2(_2423_),
    .A1(net1123),
    .B1(_0740_),
    .X(_2425_));
 sg13g2_and2_1 _6381_ (.A(_2424_),
    .B(_2425_),
    .X(_2426_));
 sg13g2_nor2b_1 _6382_ (.A(net1134),
    .B_N(net219),
    .Y(_2427_));
 sg13g2_nand3_1 _6383_ (.B(net1137),
    .C(_2427_),
    .A(net1138),
    .Y(_2428_));
 sg13g2_and2_1 _6384_ (.A(_0049_),
    .B(net1028),
    .X(_2429_));
 sg13g2_nand2_2 _6385_ (.Y(_2430_),
    .A(_0049_),
    .B(net1028));
 sg13g2_o21ai_1 _6386_ (.B1(net1117),
    .Y(_2431_),
    .A1(net1119),
    .A2(_2402_));
 sg13g2_nor2_1 _6387_ (.A(net1138),
    .B(_2420_),
    .Y(_2432_));
 sg13g2_xnor2_1 _6388_ (.Y(_2433_),
    .A(net1116),
    .B(_2431_));
 sg13g2_nand2_1 _6389_ (.Y(_2434_),
    .A(_2432_),
    .B(_2433_));
 sg13g2_o21ai_1 _6390_ (.B1(net1117),
    .Y(_2435_),
    .A1(net1119),
    .A2(net1122));
 sg13g2_xor2_1 _6391_ (.B(_2435_),
    .A(net1116),
    .X(_2436_));
 sg13g2_nand3_1 _6392_ (.B(_2419_),
    .C(_2436_),
    .A(net1138),
    .Y(_2437_));
 sg13g2_nand3_1 _6393_ (.B(_2434_),
    .C(_2437_),
    .A(net1028),
    .Y(_2438_));
 sg13g2_o21ai_1 _6394_ (.B1(_2438_),
    .Y(_2439_),
    .A1(_0092_),
    .A2(_2428_));
 sg13g2_and2_1 _6395_ (.A(net1123),
    .B(net1029),
    .X(_2440_));
 sg13g2_nand2_1 _6396_ (.Y(_2441_),
    .A(net1126),
    .B(net1029));
 sg13g2_nor2_1 _6397_ (.A(_0716_),
    .B(_2441_),
    .Y(_2442_));
 sg13g2_nand2_1 _6398_ (.Y(_2443_),
    .A(net1127),
    .B(net1029));
 sg13g2_nand4_1 _6399_ (.B(net1148),
    .C(net1065),
    .A(net1127),
    .Y(_2444_),
    .D(net1029));
 sg13g2_nand3_1 _6400_ (.B(_0730_),
    .C(net1029),
    .A(net1129),
    .Y(_2445_));
 sg13g2_a22oi_1 _6401_ (.Y(_2446_),
    .B1(net1029),
    .B2(net1127),
    .A2(net1065),
    .A1(net1148));
 sg13g2_xnor2_1 _6402_ (.Y(_2447_),
    .A(_0720_),
    .B(_2443_));
 sg13g2_o21ai_1 _6403_ (.B1(_2444_),
    .Y(_2448_),
    .A1(_2445_),
    .A2(_2446_));
 sg13g2_xor2_1 _6404_ (.B(_2441_),
    .A(_0716_),
    .X(_2449_));
 sg13g2_a21oi_1 _6405_ (.A1(_2448_),
    .A2(_2449_),
    .Y(_2450_),
    .B1(_2442_));
 sg13g2_xnor2_1 _6406_ (.Y(_2451_),
    .A(_0711_),
    .B(_2440_));
 sg13g2_nor2_1 _6407_ (.A(_2450_),
    .B(_2451_),
    .Y(_2452_));
 sg13g2_a21oi_1 _6408_ (.A1(_0711_),
    .A2(_2440_),
    .Y(_2453_),
    .B1(_2452_));
 sg13g2_nand2_1 _6409_ (.Y(_2454_),
    .A(net1122),
    .B(net1029));
 sg13g2_xor2_1 _6410_ (.B(_2454_),
    .A(_0704_),
    .X(_2455_));
 sg13g2_xor2_1 _6411_ (.B(_2455_),
    .A(_2453_),
    .X(_2456_));
 sg13g2_xor2_1 _6412_ (.B(_2451_),
    .A(_2450_),
    .X(_2457_));
 sg13g2_a21o_1 _6413_ (.A2(net1029),
    .A1(net1129),
    .B1(_0730_),
    .X(_2458_));
 sg13g2_and2_1 _6414_ (.A(_2445_),
    .B(_2458_),
    .X(_2459_));
 sg13g2_xor2_1 _6415_ (.B(_2459_),
    .A(_2457_),
    .X(_2460_));
 sg13g2_xnor2_1 _6416_ (.Y(_2461_),
    .A(_2457_),
    .B(_2459_));
 sg13g2_xnor2_1 _6417_ (.Y(_2462_),
    .A(_2445_),
    .B(_2447_));
 sg13g2_xnor2_1 _6418_ (.Y(_2463_),
    .A(_2457_),
    .B(_2462_));
 sg13g2_xor2_1 _6419_ (.B(_2462_),
    .A(_2457_),
    .X(_2464_));
 sg13g2_xor2_1 _6420_ (.B(_2449_),
    .A(_2448_),
    .X(_2465_));
 sg13g2_xor2_1 _6421_ (.B(_2465_),
    .A(_2457_),
    .X(_2466_));
 sg13g2_xnor2_1 _6422_ (.Y(_2467_),
    .A(_2457_),
    .B(_2465_));
 sg13g2_o21ai_1 _6423_ (.B1(_2467_),
    .Y(_2468_),
    .A1(_2461_),
    .A2(_2464_));
 sg13g2_xnor2_1 _6424_ (.Y(_2469_),
    .A(net988),
    .B(_2468_));
 sg13g2_nand2_1 _6425_ (.Y(_2470_),
    .A(_2439_),
    .B(_2469_));
 sg13g2_inv_1 _6426_ (.Y(_2471_),
    .A(_2470_));
 sg13g2_nand2_2 _6427_ (.Y(_2472_),
    .A(_2461_),
    .B(_2463_));
 sg13g2_o21ai_1 _6428_ (.B1(_2460_),
    .Y(_2473_),
    .A1(_2464_),
    .A2(_2466_));
 sg13g2_nor2_1 _6429_ (.A(_2917_),
    .B(net1138),
    .Y(_2474_));
 sg13g2_xnor2_1 _6430_ (.Y(_2475_),
    .A(net1122),
    .B(_2474_));
 sg13g2_nand2_1 _6431_ (.Y(_2476_),
    .A(_2420_),
    .B(net1028));
 sg13g2_o21ai_1 _6432_ (.B1(_2476_),
    .Y(_2477_),
    .A1(_0074_),
    .A2(net1028));
 sg13g2_a21o_2 _6433_ (.A2(_2475_),
    .A1(net1028),
    .B1(_2477_),
    .X(_2478_));
 sg13g2_o21ai_1 _6434_ (.B1(_2466_),
    .Y(_2479_),
    .A1(_2461_),
    .A2(_2463_));
 sg13g2_nand3_1 _6435_ (.B(_2472_),
    .C(_2479_),
    .A(net988),
    .Y(_2480_));
 sg13g2_a21o_1 _6436_ (.A2(_2479_),
    .A1(_2472_),
    .B1(net988),
    .X(_2481_));
 sg13g2_and2_1 _6437_ (.A(_2480_),
    .B(_2481_),
    .X(_2482_));
 sg13g2_nand2_1 _6438_ (.Y(_2483_),
    .A(_2478_),
    .B(_2482_));
 sg13g2_nand2_1 _6439_ (.Y(_2484_),
    .A(net989),
    .B(_2478_));
 sg13g2_nand3_1 _6440_ (.B(_2480_),
    .C(_2481_),
    .A(_2439_),
    .Y(_2485_));
 sg13g2_or2_1 _6441_ (.X(_2486_),
    .B(_2485_),
    .A(_2484_));
 sg13g2_a21o_1 _6442_ (.A2(_2473_),
    .A1(_2472_),
    .B1(_2486_),
    .X(_2487_));
 sg13g2_nand2_1 _6443_ (.Y(_2488_),
    .A(net1119),
    .B(net1122));
 sg13g2_a21oi_1 _6444_ (.A1(_2915_),
    .A2(_2916_),
    .Y(_2489_),
    .B1(_2432_));
 sg13g2_xnor2_1 _6445_ (.Y(_2490_),
    .A(_0069_),
    .B(_2402_));
 sg13g2_o21ai_1 _6446_ (.B1(_2419_),
    .Y(_2491_),
    .A1(net1138),
    .A2(_2490_));
 sg13g2_a21o_1 _6447_ (.A2(_2489_),
    .A1(_2488_),
    .B1(_2491_),
    .X(_2492_));
 sg13g2_o21ai_1 _6448_ (.B1(_2492_),
    .Y(_2493_),
    .A1(_0069_),
    .A2(net1028));
 sg13g2_nand2_1 _6449_ (.Y(_2494_),
    .A(net989),
    .B(_2493_));
 sg13g2_nand3_1 _6450_ (.B(_2472_),
    .C(_2473_),
    .A(net988),
    .Y(_2495_));
 sg13g2_a21o_1 _6451_ (.A2(_2473_),
    .A1(_2472_),
    .B1(net989),
    .X(_2496_));
 sg13g2_and2_2 _6452_ (.A(_2495_),
    .B(_2496_),
    .X(_2497_));
 sg13g2_inv_1 _6453_ (.Y(_2498_),
    .A(_2497_));
 sg13g2_nand2_1 _6454_ (.Y(_2499_),
    .A(_2439_),
    .B(_2497_));
 sg13g2_nand2_1 _6455_ (.Y(_2500_),
    .A(_2486_),
    .B(_2499_));
 sg13g2_nand2_1 _6456_ (.Y(_2501_),
    .A(_2487_),
    .B(_2500_));
 sg13g2_o21ai_1 _6457_ (.B1(_2487_),
    .Y(_2502_),
    .A1(_2494_),
    .A2(_2501_));
 sg13g2_nor4_1 _6458_ (.A(_2932_),
    .B(net1138),
    .C(_2402_),
    .D(_2420_),
    .Y(_2503_));
 sg13g2_o21ai_1 _6459_ (.B1(_2428_),
    .Y(_2504_),
    .A1(_2489_),
    .A2(_2503_));
 sg13g2_o21ai_1 _6460_ (.B1(_2476_),
    .Y(_2505_),
    .A1(_2938_),
    .A2(_2504_));
 sg13g2_a21o_2 _6461_ (.A2(_2504_),
    .A1(_2938_),
    .B1(_2505_),
    .X(_2506_));
 sg13g2_nand2_1 _6462_ (.Y(_2507_),
    .A(net988),
    .B(_2506_));
 sg13g2_xnor2_1 _6463_ (.Y(_2508_),
    .A(_2471_),
    .B(_2502_));
 sg13g2_nor2_1 _6464_ (.A(_2507_),
    .B(_2508_),
    .Y(_2509_));
 sg13g2_a21oi_1 _6465_ (.A1(_2471_),
    .A2(_2502_),
    .Y(_2510_),
    .B1(_2509_));
 sg13g2_nand3_1 _6466_ (.B(net988),
    .C(_2510_),
    .A(_2439_),
    .Y(_2511_));
 sg13g2_xor2_1 _6467_ (.B(_2508_),
    .A(_2507_),
    .X(_2512_));
 sg13g2_xor2_1 _6468_ (.B(_2485_),
    .A(_2484_),
    .X(_2513_));
 sg13g2_nand3_1 _6469_ (.B(_2463_),
    .C(_2466_),
    .A(_2461_),
    .Y(_2514_));
 sg13g2_nand3_1 _6470_ (.B(_2464_),
    .C(_2467_),
    .A(_2460_),
    .Y(_2515_));
 sg13g2_a21oi_1 _6471_ (.A1(_2514_),
    .A2(_2515_),
    .Y(_2516_),
    .B1(net988));
 sg13g2_and3_1 _6472_ (.X(_2517_),
    .A(net988),
    .B(_2514_),
    .C(_2515_));
 sg13g2_nor2_1 _6473_ (.A(_2516_),
    .B(_2517_),
    .Y(_2518_));
 sg13g2_o21ai_1 _6474_ (.B1(_2439_),
    .Y(_2519_),
    .A1(_2516_),
    .A2(_2517_));
 sg13g2_a21oi_2 _6475_ (.B1(_0075_),
    .Y(_2520_),
    .A2(net1028),
    .A1(_2420_));
 sg13g2_nand2_1 _6476_ (.Y(_2521_),
    .A(net989),
    .B(_2520_));
 sg13g2_nand2_1 _6477_ (.Y(_2522_),
    .A(_2519_),
    .B(_2521_));
 sg13g2_nand2_1 _6478_ (.Y(_2523_),
    .A(_2469_),
    .B(_2478_));
 sg13g2_o21ai_1 _6479_ (.B1(_2523_),
    .Y(_2524_),
    .A1(_2519_),
    .A2(_2521_));
 sg13g2_nand3_1 _6480_ (.B(_2522_),
    .C(_2524_),
    .A(_2513_),
    .Y(_2525_));
 sg13g2_nand2_1 _6481_ (.Y(_2526_),
    .A(_2469_),
    .B(_2493_));
 sg13g2_inv_1 _6482_ (.Y(_2527_),
    .A(_2526_));
 sg13g2_a21o_1 _6483_ (.A2(_2524_),
    .A1(_2522_),
    .B1(_2513_),
    .X(_2528_));
 sg13g2_nand3_1 _6484_ (.B(_2527_),
    .C(_2528_),
    .A(_2525_),
    .Y(_2529_));
 sg13g2_nand2_1 _6485_ (.Y(_2530_),
    .A(_2525_),
    .B(_2529_));
 sg13g2_xor2_1 _6486_ (.B(_2501_),
    .A(_2494_),
    .X(_2531_));
 sg13g2_nand2_1 _6487_ (.Y(_2532_),
    .A(_2469_),
    .B(_2506_));
 sg13g2_xnor2_1 _6488_ (.Y(_2533_),
    .A(_2530_),
    .B(_2531_));
 sg13g2_nor2_1 _6489_ (.A(_2532_),
    .B(_2533_),
    .Y(_2534_));
 sg13g2_a21oi_1 _6490_ (.A1(_2530_),
    .A2(_2531_),
    .Y(_2535_),
    .B1(_2534_));
 sg13g2_nor2b_1 _6491_ (.A(_2535_),
    .B_N(_2512_),
    .Y(_2536_));
 sg13g2_xor2_1 _6492_ (.B(_2533_),
    .A(_2532_),
    .X(_2537_));
 sg13g2_nand2_1 _6493_ (.Y(_2538_),
    .A(_2493_),
    .B(_2497_));
 sg13g2_xor2_1 _6494_ (.B(_2521_),
    .A(_2519_),
    .X(_2539_));
 sg13g2_nand2_1 _6495_ (.Y(_2540_),
    .A(_2497_),
    .B(_2520_));
 sg13g2_a21oi_1 _6496_ (.A1(_2497_),
    .A2(_2520_),
    .Y(_2541_),
    .B1(_2523_));
 sg13g2_xnor2_1 _6497_ (.Y(_2542_),
    .A(_2539_),
    .B(_2541_));
 sg13g2_nand3_1 _6498_ (.B(_2495_),
    .C(_2496_),
    .A(_2478_),
    .Y(_2543_));
 sg13g2_nand2_1 _6499_ (.Y(_2544_),
    .A(_2469_),
    .B(_2520_));
 sg13g2_or3_1 _6500_ (.A(_2523_),
    .B(_2539_),
    .C(_2540_),
    .X(_2545_));
 sg13g2_o21ai_1 _6501_ (.B1(_2545_),
    .Y(_2546_),
    .A1(_2538_),
    .A2(_2542_));
 sg13g2_a21o_1 _6502_ (.A2(_2528_),
    .A1(_2525_),
    .B1(_2527_),
    .X(_2547_));
 sg13g2_and3_1 _6503_ (.X(_2548_),
    .A(_2529_),
    .B(_2546_),
    .C(_2547_));
 sg13g2_nand3_1 _6504_ (.B(_2546_),
    .C(_2547_),
    .A(_2529_),
    .Y(_2549_));
 sg13g2_a21o_1 _6505_ (.A2(_2547_),
    .A1(_2529_),
    .B1(_2546_),
    .X(_2550_));
 sg13g2_and4_1 _6506_ (.A(_2497_),
    .B(_2506_),
    .C(_2549_),
    .D(_2550_),
    .X(_2551_));
 sg13g2_or2_1 _6507_ (.X(_2552_),
    .B(_2551_),
    .A(_2548_));
 sg13g2_nand2_1 _6508_ (.Y(_2553_),
    .A(_2537_),
    .B(_2552_));
 sg13g2_xnor2_1 _6509_ (.Y(_2554_),
    .A(_2537_),
    .B(_2552_));
 sg13g2_a22oi_1 _6510_ (.Y(_2555_),
    .B1(_2549_),
    .B2(_2550_),
    .A2(_2506_),
    .A1(_2497_));
 sg13g2_xor2_1 _6511_ (.B(_2542_),
    .A(_2538_),
    .X(_2556_));
 sg13g2_xnor2_1 _6512_ (.Y(_2557_),
    .A(_2543_),
    .B(_2544_));
 sg13g2_nand4_1 _6513_ (.B(_2482_),
    .C(_2497_),
    .A(_2478_),
    .Y(_2558_),
    .D(_2520_));
 sg13g2_or2_1 _6514_ (.X(_2559_),
    .B(_2558_),
    .A(_2557_));
 sg13g2_nand2_1 _6515_ (.Y(_2560_),
    .A(_2482_),
    .B(_2493_));
 sg13g2_xnor2_1 _6516_ (.Y(_2561_),
    .A(_2557_),
    .B(_2558_));
 sg13g2_o21ai_1 _6517_ (.B1(_2559_),
    .Y(_2562_),
    .A1(_2560_),
    .A2(_2561_));
 sg13g2_and2_1 _6518_ (.A(_2556_),
    .B(_2562_),
    .X(_2563_));
 sg13g2_and2_1 _6519_ (.A(_2482_),
    .B(_2506_),
    .X(_2564_));
 sg13g2_xor2_1 _6520_ (.B(_2562_),
    .A(_2556_),
    .X(_2565_));
 sg13g2_a21oi_1 _6521_ (.A1(_2564_),
    .A2(_2565_),
    .Y(_2566_),
    .B1(_2563_));
 sg13g2_nor3_1 _6522_ (.A(_2551_),
    .B(_2555_),
    .C(_2566_),
    .Y(_2567_));
 sg13g2_or3_1 _6523_ (.A(_2551_),
    .B(_2555_),
    .C(_2566_),
    .X(_2568_));
 sg13g2_or2_1 _6524_ (.X(_2569_),
    .B(_2565_),
    .A(_2564_));
 sg13g2_a21oi_1 _6525_ (.A1(_2498_),
    .A2(_2520_),
    .Y(_2570_),
    .B1(_2493_));
 sg13g2_a21oi_1 _6526_ (.A1(_2483_),
    .A2(_2540_),
    .Y(_2571_),
    .B1(_2570_));
 sg13g2_nand2_1 _6527_ (.Y(_2572_),
    .A(_2506_),
    .B(_2571_));
 sg13g2_xnor2_1 _6528_ (.Y(_2573_),
    .A(_2560_),
    .B(_2561_));
 sg13g2_or2_1 _6529_ (.X(_2574_),
    .B(_2571_),
    .A(_2506_));
 sg13g2_a221oi_1 _6530_ (.B2(_2573_),
    .C1(_2518_),
    .B1(_2572_),
    .A1(_2564_),
    .Y(_2575_),
    .A2(_2565_));
 sg13g2_and3_1 _6531_ (.X(_2576_),
    .A(_2569_),
    .B(_2574_),
    .C(_2575_));
 sg13g2_o21ai_1 _6532_ (.B1(_2566_),
    .Y(_2577_),
    .A1(_2551_),
    .A2(_2555_));
 sg13g2_nand3_1 _6533_ (.B(_2576_),
    .C(_2577_),
    .A(_2568_),
    .Y(_2578_));
 sg13g2_a21oi_1 _6534_ (.A1(_2576_),
    .A2(_2577_),
    .Y(_2579_),
    .B1(_2567_));
 sg13g2_o21ai_1 _6535_ (.B1(_2553_),
    .Y(_2580_),
    .A1(_2554_),
    .A2(_2579_));
 sg13g2_xnor2_1 _6536_ (.Y(_2581_),
    .A(_2512_),
    .B(_2535_));
 sg13g2_nand2_1 _6537_ (.Y(_2582_),
    .A(_2580_),
    .B(_2581_));
 sg13g2_a21oi_1 _6538_ (.A1(_2580_),
    .A2(_2581_),
    .Y(_2583_),
    .B1(_2536_));
 sg13g2_o21ai_1 _6539_ (.B1(_2510_),
    .Y(_2584_),
    .A1(_2511_),
    .A2(_2583_));
 sg13g2_nand2_1 _6540_ (.Y(_2585_),
    .A(_2430_),
    .B(_2584_));
 sg13g2_nand4_1 _6541_ (.B(_2423_),
    .C(_2430_),
    .A(_2935_),
    .Y(_2586_),
    .D(_2584_));
 sg13g2_o21ai_1 _6542_ (.B1(_2585_),
    .Y(_2587_),
    .A1(_0081_),
    .A2(_2422_));
 sg13g2_nand2_1 _6543_ (.Y(_2588_),
    .A(_2586_),
    .B(_2587_));
 sg13g2_o21ai_1 _6544_ (.B1(_2586_),
    .Y(_2589_),
    .A1(_0703_),
    .A2(_2588_));
 sg13g2_nand2_1 _6545_ (.Y(_2590_),
    .A(_2426_),
    .B(_2589_));
 sg13g2_nand2_1 _6546_ (.Y(_2591_),
    .A(_2934_),
    .B(_2423_));
 sg13g2_xnor2_1 _6547_ (.Y(_2592_),
    .A(_2511_),
    .B(_2583_));
 sg13g2_or3_1 _6548_ (.A(_2429_),
    .B(_2591_),
    .C(_2592_),
    .X(_2593_));
 sg13g2_o21ai_1 _6549_ (.B1(_2591_),
    .Y(_2594_),
    .A1(_2429_),
    .A2(_2592_));
 sg13g2_nand3_1 _6550_ (.B(_2593_),
    .C(_2594_),
    .A(_0709_),
    .Y(_2595_));
 sg13g2_and2_1 _6551_ (.A(_2593_),
    .B(_2595_),
    .X(_2596_));
 sg13g2_xnor2_1 _6552_ (.Y(_2597_),
    .A(_0703_),
    .B(_2588_));
 sg13g2_nor2_1 _6553_ (.A(_2596_),
    .B(_2597_),
    .Y(_2598_));
 sg13g2_nor2_1 _6554_ (.A(_0079_),
    .B(_2422_),
    .Y(_2599_));
 sg13g2_or2_1 _6555_ (.X(_2600_),
    .B(_2581_),
    .A(_2580_));
 sg13g2_nand3_1 _6556_ (.B(_2582_),
    .C(_2600_),
    .A(_2430_),
    .Y(_2601_));
 sg13g2_nand4_1 _6557_ (.B(_2582_),
    .C(_2599_),
    .A(_2430_),
    .Y(_2602_),
    .D(_2600_));
 sg13g2_xor2_1 _6558_ (.B(_2601_),
    .A(_2599_),
    .X(_2603_));
 sg13g2_o21ai_1 _6559_ (.B1(_2602_),
    .Y(_2604_),
    .A1(_0717_),
    .A2(_2603_));
 sg13g2_a21o_1 _6560_ (.A2(_2594_),
    .A1(_2593_),
    .B1(_0709_),
    .X(_2605_));
 sg13g2_and2_1 _6561_ (.A(_2595_),
    .B(_2605_),
    .X(_2606_));
 sg13g2_nand2_1 _6562_ (.Y(_2607_),
    .A(_2604_),
    .B(_2606_));
 sg13g2_a21oi_1 _6563_ (.A1(_2568_),
    .A2(_2577_),
    .Y(_2608_),
    .B1(_2576_));
 sg13g2_nand3_1 _6564_ (.B(_2430_),
    .C(_2578_),
    .A(_0727_),
    .Y(_2609_));
 sg13g2_nor2_1 _6565_ (.A(_2608_),
    .B(_2609_),
    .Y(_2610_));
 sg13g2_or2_1 _6566_ (.X(_2611_),
    .B(_2610_),
    .A(_0721_));
 sg13g2_nand2_1 _6567_ (.Y(_2612_),
    .A(_0721_),
    .B(_2610_));
 sg13g2_xor2_1 _6568_ (.B(_2579_),
    .A(_2554_),
    .X(_2613_));
 sg13g2_nand3_1 _6569_ (.B(_2611_),
    .C(_2613_),
    .A(_2430_),
    .Y(_2614_));
 sg13g2_a22oi_1 _6570_ (.Y(_2615_),
    .B1(_2612_),
    .B2(_2614_),
    .A2(_2603_),
    .A1(_0717_));
 sg13g2_o21ai_1 _6571_ (.B1(_2615_),
    .Y(_2616_),
    .A1(_0717_),
    .A2(_2603_));
 sg13g2_xnor2_1 _6572_ (.Y(_2617_),
    .A(_2604_),
    .B(_2606_));
 sg13g2_o21ai_1 _6573_ (.B1(_2607_),
    .Y(_2618_),
    .A1(_2616_),
    .A2(_2617_));
 sg13g2_xor2_1 _6574_ (.B(_2597_),
    .A(_2596_),
    .X(_2619_));
 sg13g2_a21oi_1 _6575_ (.A1(_2618_),
    .A2(_2619_),
    .Y(_2620_),
    .B1(_2598_));
 sg13g2_xnor2_1 _6576_ (.Y(_2621_),
    .A(_2426_),
    .B(_2589_));
 sg13g2_o21ai_1 _6577_ (.B1(_2590_),
    .Y(_2622_),
    .A1(_2620_),
    .A2(_2621_));
 sg13g2_nand2_1 _6578_ (.Y(_2623_),
    .A(net1122),
    .B(_2423_));
 sg13g2_xnor2_1 _6579_ (.Y(_2624_),
    .A(_0697_),
    .B(_2623_));
 sg13g2_xnor2_1 _6580_ (.Y(_2625_),
    .A(_2424_),
    .B(_2624_));
 sg13g2_xnor2_1 _6581_ (.Y(_2626_),
    .A(_2622_),
    .B(_2625_));
 sg13g2_xor2_1 _6582_ (.B(_2621_),
    .A(_2620_),
    .X(_2627_));
 sg13g2_xnor2_1 _6583_ (.Y(_2628_),
    .A(_2616_),
    .B(_2617_));
 sg13g2_inv_1 _6584_ (.Y(_2629_),
    .A(_2628_));
 sg13g2_xor2_1 _6585_ (.B(_2619_),
    .A(_2618_),
    .X(_2630_));
 sg13g2_nand2_1 _6586_ (.Y(_2631_),
    .A(_2629_),
    .B(_2630_));
 sg13g2_nand3_1 _6587_ (.B(_2629_),
    .C(_2630_),
    .A(_2627_),
    .Y(_2632_));
 sg13g2_xor2_1 _6588_ (.B(_2632_),
    .A(_2626_),
    .X(_2633_));
 sg13g2_nor4_2 _6589_ (.A(net1133),
    .B(net1135),
    .C(net1140),
    .Y(_2634_),
    .D(net1136));
 sg13g2_inv_1 _6590_ (.Y(_2635_),
    .A(_2634_));
 sg13g2_nor2_1 _6591_ (.A(_2909_),
    .B(_2635_),
    .Y(_2636_));
 sg13g2_nand2_1 _6592_ (.Y(_2637_),
    .A(net1091),
    .B(_2634_));
 sg13g2_and2_1 _6593_ (.A(net1133),
    .B(net1135),
    .X(_2638_));
 sg13g2_nand2_1 _6594_ (.Y(_2639_),
    .A(net1133),
    .B(net1137));
 sg13g2_xnor2_1 _6595_ (.Y(_2640_),
    .A(_2908_),
    .B(_2639_));
 sg13g2_o21ai_1 _6596_ (.B1(_2635_),
    .Y(_2641_),
    .A1(_2638_),
    .A2(_2640_));
 sg13g2_nand2_1 _6597_ (.Y(_2642_),
    .A(_2637_),
    .B(_2641_));
 sg13g2_nand2b_1 _6598_ (.Y(_2643_),
    .B(_2633_),
    .A_N(_2642_));
 sg13g2_nand2_1 _6599_ (.Y(_2644_),
    .A(\i_display.i_vga.timing_ver.counter[0] ),
    .B(_0730_));
 sg13g2_nand2_1 _6600_ (.Y(_2645_),
    .A(\i_display.i_vga.timing_ver.counter[2] ),
    .B(_0709_));
 sg13g2_nand2_1 _6601_ (.Y(_2646_),
    .A(_0703_),
    .B(_2645_));
 sg13g2_nand2_2 _6602_ (.Y(_2647_),
    .A(\i_display.i_vga.timing_ver.counter[5] ),
    .B(_2646_));
 sg13g2_and3_1 _6603_ (.X(_2648_),
    .A(_0691_),
    .B(_0697_),
    .C(_2647_));
 sg13g2_nor2_1 _6604_ (.A(_0684_),
    .B(_2648_),
    .Y(_2649_));
 sg13g2_mux2_1 _6605_ (.A0(_0678_),
    .A1(_2920_),
    .S(_2649_),
    .X(_2650_));
 sg13g2_nor2_1 _6606_ (.A(_0728_),
    .B(_2650_),
    .Y(_2651_));
 sg13g2_nand2_1 _6607_ (.Y(_2652_),
    .A(net1130),
    .B(_2651_));
 sg13g2_o21ai_1 _6608_ (.B1(_2652_),
    .Y(_2653_),
    .A1(_0721_),
    .A2(_2651_));
 sg13g2_nand2_1 _6609_ (.Y(_2654_),
    .A(net1141),
    .B(_1527_));
 sg13g2_nor3_1 _6610_ (.A(net1132),
    .B(\i_display.i_vga.hblank ),
    .C(_2654_),
    .Y(_2655_));
 sg13g2_nand2_1 _6611_ (.Y(_2656_),
    .A(\i_display.i_vga.low_count[8] ),
    .B(_2655_));
 sg13g2_nand2_1 _6612_ (.Y(_2657_),
    .A(_0679_),
    .B(_2656_));
 sg13g2_o21ai_1 _6613_ (.B1(_2657_),
    .Y(_2658_),
    .A1(_2929_),
    .A2(_2656_));
 sg13g2_nand2_1 _6614_ (.Y(_2659_),
    .A(_0730_),
    .B(_2658_));
 sg13g2_mux2_1 _6615_ (.A0(net1148),
    .A1(_0720_),
    .S(_2659_),
    .X(_2660_));
 sg13g2_or2_1 _6616_ (.X(_2661_),
    .B(_2660_),
    .A(_2653_));
 sg13g2_xnor2_1 _6617_ (.Y(_2662_),
    .A(_2653_),
    .B(_2660_));
 sg13g2_xor2_1 _6618_ (.B(_2662_),
    .A(_2644_),
    .X(_2663_));
 sg13g2_nand3_1 _6619_ (.B(_2628_),
    .C(_2630_),
    .A(_2627_),
    .Y(_2664_));
 sg13g2_nand2_1 _6620_ (.Y(_2665_),
    .A(net1091),
    .B(net1135));
 sg13g2_and2_1 _6621_ (.A(net1091),
    .B(_2638_),
    .X(_2666_));
 sg13g2_nor2_1 _6622_ (.A(_2634_),
    .B(_2638_),
    .Y(_2667_));
 sg13g2_a21o_2 _6623_ (.A2(_2667_),
    .A1(_2640_),
    .B1(_2666_),
    .X(_2668_));
 sg13g2_xor2_1 _6624_ (.B(_2664_),
    .A(_2626_),
    .X(_2669_));
 sg13g2_a221oi_1 _6625_ (.B2(_2669_),
    .C1(_2964_),
    .B1(_2668_),
    .A1(_2636_),
    .Y(_2670_),
    .A2(_2663_));
 sg13g2_nor3_1 _6626_ (.A(\i_display.i_vga.timing_ver.counter[1] ),
    .B(\i_display.i_vga.timing_ver.counter[0] ),
    .C(_2645_),
    .Y(_2671_));
 sg13g2_nor2b_1 _6627_ (.A(\i_display.i_vga.timing_ver.counter[4] ),
    .B_N(_2671_),
    .Y(_2672_));
 sg13g2_nor2_1 _6628_ (.A(net990),
    .B(_2672_),
    .Y(_2673_));
 sg13g2_o21ai_1 _6629_ (.B1(_2647_),
    .Y(_2674_),
    .A1(_0740_),
    .A2(_2646_));
 sg13g2_xor2_1 _6630_ (.B(_2674_),
    .A(_2673_),
    .X(_2675_));
 sg13g2_o21ai_1 _6631_ (.B1(net1063),
    .Y(_2676_),
    .A1(\i_display.i_vga.low_count[2] ),
    .A2(net1067));
 sg13g2_nand2_1 _6632_ (.Y(_2677_),
    .A(_0710_),
    .B(_2676_));
 sg13g2_a21oi_1 _6633_ (.A1(_2658_),
    .A2(_2677_),
    .Y(_2678_),
    .B1(_0704_));
 sg13g2_a21o_1 _6634_ (.A2(net991),
    .A1(_0704_),
    .B1(_2678_),
    .X(_2679_));
 sg13g2_xnor2_1 _6635_ (.Y(_2680_),
    .A(_0739_),
    .B(_2679_));
 sg13g2_nor2_1 _6636_ (.A(_2675_),
    .B(_2680_),
    .Y(_2681_));
 sg13g2_nand3_1 _6637_ (.B(net991),
    .C(_2677_),
    .A(_0704_),
    .Y(_2682_));
 sg13g2_nand2b_1 _6638_ (.Y(_2683_),
    .B(_2682_),
    .A_N(_2678_));
 sg13g2_o21ai_1 _6639_ (.B1(_2646_),
    .Y(_2684_),
    .A1(_0717_),
    .A2(_2354_));
 sg13g2_nor2_1 _6640_ (.A(net990),
    .B(_2671_),
    .Y(_2685_));
 sg13g2_xnor2_1 _6641_ (.Y(_2686_),
    .A(_2684_),
    .B(_2685_));
 sg13g2_nor2b_1 _6642_ (.A(_2676_),
    .B_N(net991),
    .Y(_2687_));
 sg13g2_xnor2_1 _6643_ (.Y(_2688_),
    .A(_0711_),
    .B(_2687_));
 sg13g2_a21oi_1 _6644_ (.A1(_0722_),
    .A2(_0728_),
    .Y(_2689_),
    .B1(net990));
 sg13g2_nand2b_1 _6645_ (.Y(_2690_),
    .B(_0717_),
    .A_N(net990));
 sg13g2_o21ai_1 _6646_ (.B1(_2690_),
    .Y(_2691_),
    .A1(_0717_),
    .A2(_2689_));
 sg13g2_xnor2_1 _6647_ (.Y(_2692_),
    .A(_0709_),
    .B(_2691_));
 sg13g2_nor2_1 _6648_ (.A(_2688_),
    .B(_2692_),
    .Y(_2693_));
 sg13g2_xor2_1 _6649_ (.B(_2692_),
    .A(_2688_),
    .X(_2694_));
 sg13g2_xnor2_1 _6650_ (.Y(_2695_),
    .A(_0717_),
    .B(_2689_));
 sg13g2_nand3_1 _6651_ (.B(net1063),
    .C(net991),
    .A(net1067),
    .Y(_2696_));
 sg13g2_mux2_1 _6652_ (.A0(\i_display.i_vga.low_count[2] ),
    .A1(_0716_),
    .S(_2696_),
    .X(_2697_));
 sg13g2_o21ai_1 _6653_ (.B1(_2661_),
    .Y(_2698_),
    .A1(_2644_),
    .A2(_2662_));
 sg13g2_xor2_1 _6654_ (.B(_2697_),
    .A(_2695_),
    .X(_2699_));
 sg13g2_nand2_1 _6655_ (.Y(_2700_),
    .A(_2698_),
    .B(_2699_));
 sg13g2_o21ai_1 _6656_ (.B1(_2700_),
    .Y(_2701_),
    .A1(_2695_),
    .A2(_2697_));
 sg13g2_a21oi_1 _6657_ (.A1(_2694_),
    .A2(_2701_),
    .Y(_2702_),
    .B1(_2693_));
 sg13g2_xor2_1 _6658_ (.B(_2686_),
    .A(_2683_),
    .X(_2703_));
 sg13g2_nand2b_1 _6659_ (.Y(_2704_),
    .B(_2703_),
    .A_N(_2702_));
 sg13g2_o21ai_1 _6660_ (.B1(_2704_),
    .Y(_2705_),
    .A1(_2683_),
    .A2(_2686_));
 sg13g2_xor2_1 _6661_ (.B(_2680_),
    .A(_2675_),
    .X(_2706_));
 sg13g2_a21oi_1 _6662_ (.A1(_2705_),
    .A2(_2706_),
    .Y(_2707_),
    .B1(_2681_));
 sg13g2_and2_1 _6663_ (.A(_0740_),
    .B(_2672_),
    .X(_2708_));
 sg13g2_nor2_1 _6664_ (.A(net990),
    .B(_2708_),
    .Y(_2709_));
 sg13g2_xor2_1 _6665_ (.B(_2647_),
    .A(_0697_),
    .X(_2710_));
 sg13g2_xnor2_1 _6666_ (.Y(_2711_),
    .A(_2709_),
    .B(_2710_));
 sg13g2_o21ai_1 _6667_ (.B1(\i_display.i_vga.low_count[6] ),
    .Y(_2712_),
    .A1(\i_display.i_vga.low_count[5] ),
    .A2(\i_display.i_vga.low_count[4] ));
 sg13g2_nand3_1 _6668_ (.B(_1527_),
    .C(_2712_),
    .A(net1064),
    .Y(_2713_));
 sg13g2_nor3_1 _6669_ (.A(\i_display.i_vga.low_count[5] ),
    .B(_0704_),
    .C(_2677_),
    .Y(_2714_));
 sg13g2_nand2b_1 _6670_ (.Y(_2715_),
    .B(net991),
    .A_N(_2714_));
 sg13g2_xnor2_1 _6671_ (.Y(_2716_),
    .A(_2713_),
    .B(_2715_));
 sg13g2_nand2_1 _6672_ (.Y(_2717_),
    .A(_2711_),
    .B(_2716_));
 sg13g2_xnor2_1 _6673_ (.Y(_2718_),
    .A(_2711_),
    .B(_2716_));
 sg13g2_xor2_1 _6674_ (.B(_2718_),
    .A(_2707_),
    .X(_2719_));
 sg13g2_inv_1 _6675_ (.Y(_2720_),
    .A(_2719_));
 sg13g2_nand2_1 _6676_ (.Y(_2721_),
    .A(net1116),
    .B(_2720_));
 sg13g2_xor2_1 _6677_ (.B(_2701_),
    .A(_2694_),
    .X(_2722_));
 sg13g2_nor2_1 _6678_ (.A(_2916_),
    .B(net980),
    .Y(_2723_));
 sg13g2_xnor2_1 _6679_ (.Y(_2724_),
    .A(_2698_),
    .B(_2699_));
 sg13g2_xnor2_1 _6680_ (.Y(_2725_),
    .A(_2933_),
    .B(net984));
 sg13g2_xnor2_1 _6681_ (.Y(_2726_),
    .A(_2916_),
    .B(net980));
 sg13g2_nor2_1 _6682_ (.A(_2725_),
    .B(_2726_),
    .Y(_2727_));
 sg13g2_o21ai_1 _6683_ (.B1(_2644_),
    .Y(_2728_),
    .A1(_0727_),
    .A2(_0730_));
 sg13g2_xnor2_1 _6684_ (.Y(_2729_),
    .A(_2935_),
    .B(_2663_));
 sg13g2_o21ai_1 _6685_ (.B1(_2729_),
    .Y(_2730_),
    .A1(net1127),
    .A2(_2728_));
 sg13g2_o21ai_1 _6686_ (.B1(_2730_),
    .Y(_2731_),
    .A1(_2918_),
    .A2(_2663_));
 sg13g2_a21oi_1 _6687_ (.A1(net1123),
    .A2(net984),
    .Y(_2732_),
    .B1(_2723_));
 sg13g2_a21oi_1 _6688_ (.A1(_2916_),
    .A2(net980),
    .Y(_2733_),
    .B1(_2732_));
 sg13g2_a21o_1 _6689_ (.A2(_2731_),
    .A1(_2727_),
    .B1(_2733_),
    .X(_2734_));
 sg13g2_xnor2_1 _6690_ (.Y(_2735_),
    .A(_2705_),
    .B(_2706_));
 sg13g2_xnor2_1 _6691_ (.Y(_2736_),
    .A(_2938_),
    .B(net933));
 sg13g2_xnor2_1 _6692_ (.Y(_2737_),
    .A(_2702_),
    .B(_2703_));
 sg13g2_xnor2_1 _6693_ (.Y(_2738_),
    .A(_0069_),
    .B(_2737_));
 sg13g2_nor2_1 _6694_ (.A(_2736_),
    .B(_2738_),
    .Y(_2739_));
 sg13g2_nor3_1 _6695_ (.A(_0069_),
    .B(_2736_),
    .C(_2737_),
    .Y(_2740_));
 sg13g2_a221oi_1 _6696_ (.B2(_2734_),
    .C1(_2740_),
    .B1(_2739_),
    .A1(net1117),
    .Y(_2741_),
    .A2(net933));
 sg13g2_xnor2_1 _6697_ (.Y(_2742_),
    .A(_2939_),
    .B(_2719_));
 sg13g2_nand2b_1 _6698_ (.Y(_2743_),
    .B(_2742_),
    .A_N(_2741_));
 sg13g2_o21ai_1 _6699_ (.B1(_2717_),
    .Y(_2744_),
    .A1(_2707_),
    .A2(_2718_));
 sg13g2_a21oi_1 _6700_ (.A1(_0697_),
    .A2(_2647_),
    .Y(_2745_),
    .B1(_0691_));
 sg13g2_nor2_1 _6701_ (.A(_2648_),
    .B(_2745_),
    .Y(_2746_));
 sg13g2_a21oi_1 _6702_ (.A1(_2708_),
    .A2(_2710_),
    .Y(_2747_),
    .B1(net990));
 sg13g2_xnor2_1 _6703_ (.Y(_2748_),
    .A(_2746_),
    .B(_2747_));
 sg13g2_nor2b_1 _6704_ (.A(_2713_),
    .B_N(_2714_),
    .Y(_2749_));
 sg13g2_nor2b_1 _6705_ (.A(_2749_),
    .B_N(net991),
    .Y(_2750_));
 sg13g2_o21ai_1 _6706_ (.B1(net1064),
    .Y(_2751_),
    .A1(net1141),
    .A2(_1527_));
 sg13g2_nand2b_1 _6707_ (.Y(_2752_),
    .B(_2654_),
    .A_N(_2751_));
 sg13g2_xnor2_1 _6708_ (.Y(_2753_),
    .A(_2750_),
    .B(_2752_));
 sg13g2_and2_1 _6709_ (.A(_2748_),
    .B(_2753_),
    .X(_2754_));
 sg13g2_xor2_1 _6710_ (.B(_2753_),
    .A(_2748_),
    .X(_2755_));
 sg13g2_xnor2_1 _6711_ (.Y(_2756_),
    .A(_2744_),
    .B(_2755_));
 sg13g2_xnor2_1 _6712_ (.Y(_2757_),
    .A(_2934_),
    .B(_2728_));
 sg13g2_nor3_1 _6713_ (.A(_2725_),
    .B(_2726_),
    .C(_2757_),
    .Y(_2758_));
 sg13g2_nand4_1 _6714_ (.B(_2739_),
    .C(_2742_),
    .A(_2729_),
    .Y(_2759_),
    .D(_2758_));
 sg13g2_o21ai_1 _6715_ (.B1(_2759_),
    .Y(_2760_),
    .A1(\i_display.frame[8] ),
    .A2(_2756_));
 sg13g2_a21oi_1 _6716_ (.A1(_2721_),
    .A2(_2743_),
    .Y(_2761_),
    .B1(_2760_));
 sg13g2_a21oi_1 _6717_ (.A1(_2744_),
    .A2(_2755_),
    .Y(_2762_),
    .B1(_2754_));
 sg13g2_xor2_1 _6718_ (.B(_2648_),
    .A(_0684_),
    .X(_2763_));
 sg13g2_nand2_1 _6719_ (.Y(_2764_),
    .A(_1424_),
    .B(_2708_));
 sg13g2_nor2b_1 _6720_ (.A(net990),
    .B_N(_2764_),
    .Y(_2765_));
 sg13g2_xor2_1 _6721_ (.B(_2765_),
    .A(_2763_),
    .X(_2766_));
 sg13g2_o21ai_1 _6722_ (.B1(_2656_),
    .Y(_2767_),
    .A1(_0685_),
    .A2(_2655_));
 sg13g2_nand2_1 _6723_ (.Y(_2768_),
    .A(net1141),
    .B(_2749_));
 sg13g2_nand2_1 _6724_ (.Y(_2769_),
    .A(net991),
    .B(_2768_));
 sg13g2_xor2_1 _6725_ (.B(_2769_),
    .A(_2767_),
    .X(_2770_));
 sg13g2_xnor2_1 _6726_ (.Y(_2771_),
    .A(_2766_),
    .B(_2770_));
 sg13g2_xnor2_1 _6727_ (.Y(_2772_),
    .A(_2762_),
    .B(_2771_));
 sg13g2_a221oi_1 _6728_ (.B2(_2942_),
    .C1(_2761_),
    .B1(_2772_),
    .A1(\i_display.frame[8] ),
    .Y(_2773_),
    .A2(_2756_));
 sg13g2_nand4_1 _6729_ (.B(net1141),
    .C(net991),
    .A(\i_display.i_vga.low_count[8] ),
    .Y(_2774_),
    .D(_2749_));
 sg13g2_nor3_1 _6730_ (.A(net990),
    .B(_2763_),
    .C(_2764_),
    .Y(_2775_));
 sg13g2_xnor2_1 _6731_ (.Y(_2776_),
    .A(_2774_),
    .B(_2775_));
 sg13g2_a21oi_1 _6732_ (.A1(_2766_),
    .A2(_2770_),
    .Y(_2777_),
    .B1(_2776_));
 sg13g2_o21ai_1 _6733_ (.B1(_2777_),
    .Y(_2778_),
    .A1(_2762_),
    .A2(_2771_));
 sg13g2_nor2_1 _6734_ (.A(_2942_),
    .B(_2772_),
    .Y(_2779_));
 sg13g2_nor3_1 _6735_ (.A(_2773_),
    .B(_2778_),
    .C(_2779_),
    .Y(_2780_));
 sg13g2_and2_1 _6736_ (.A(net1135),
    .B(_2780_),
    .X(_2781_));
 sg13g2_a21oi_1 _6737_ (.A1(_2909_),
    .A2(_0024_),
    .Y(_2782_),
    .B1(net1133));
 sg13g2_nor2b_1 _6738_ (.A(_2724_),
    .B_N(_2781_),
    .Y(_2783_));
 sg13g2_nand2_1 _6739_ (.Y(_2784_),
    .A(\i_display.frame_crotchet[1] ),
    .B(_2783_));
 sg13g2_o21ai_1 _6740_ (.B1(_2784_),
    .Y(_2785_),
    .A1(_2781_),
    .A2(_2782_));
 sg13g2_a21oi_1 _6741_ (.A1(_2720_),
    .A2(_2735_),
    .Y(_2786_),
    .B1(_2756_));
 sg13g2_nor2b_1 _6742_ (.A(_2772_),
    .B_N(_2786_),
    .Y(_2787_));
 sg13g2_nor2_2 _6743_ (.A(_2778_),
    .B(_2787_),
    .Y(_2788_));
 sg13g2_o21ai_1 _6744_ (.B1(net1133),
    .Y(_2789_),
    .A1(net1135),
    .A2(_2788_));
 sg13g2_nand2_1 _6745_ (.Y(_2790_),
    .A(net1128),
    .B(net1138));
 sg13g2_xnor2_1 _6746_ (.Y(_2791_),
    .A(_2663_),
    .B(_2790_));
 sg13g2_nor2_1 _6747_ (.A(_0077_),
    .B(_2663_),
    .Y(_2792_));
 sg13g2_xnor2_1 _6748_ (.Y(_2793_),
    .A(_2935_),
    .B(net984));
 sg13g2_nor2_1 _6749_ (.A(_2792_),
    .B(_2793_),
    .Y(_2794_));
 sg13g2_xnor2_1 _6750_ (.Y(_2795_),
    .A(_2792_),
    .B(_2793_));
 sg13g2_inv_1 _6751_ (.Y(_2796_),
    .A(_2795_));
 sg13g2_nand3_1 _6752_ (.B(_2418_),
    .C(_2788_),
    .A(\i_display.frame_crotchet[1] ),
    .Y(_2797_));
 sg13g2_inv_1 _6753_ (.Y(_2798_),
    .A(_2797_));
 sg13g2_nor2_1 _6754_ (.A(_2795_),
    .B(_2797_),
    .Y(_2799_));
 sg13g2_a221oi_1 _6755_ (.B2(_2666_),
    .C1(_2799_),
    .B1(_2791_),
    .A1(_2785_),
    .Y(_2800_),
    .A2(_2789_));
 sg13g2_a221oi_1 _6756_ (.B2(_2964_),
    .C1(net1159),
    .B1(_2800_),
    .A1(_2643_),
    .Y(_0221_),
    .A2(_2670_));
 sg13g2_nor2_1 _6757_ (.A(_0026_),
    .B(_2635_),
    .Y(_2801_));
 sg13g2_a22oi_1 _6758_ (.Y(_2802_),
    .B1(net984),
    .B2(_2801_),
    .A2(_2668_),
    .A1(_2633_));
 sg13g2_nand4_1 _6759_ (.B(_2427_),
    .C(_2722_),
    .A(_2965_),
    .Y(_2803_),
    .D(_2780_));
 sg13g2_nor2_1 _6760_ (.A(net1126),
    .B(net984),
    .Y(_2804_));
 sg13g2_nor2_1 _6761_ (.A(_2794_),
    .B(_2804_),
    .Y(_2805_));
 sg13g2_xnor2_1 _6762_ (.Y(_2806_),
    .A(_0075_),
    .B(net980));
 sg13g2_xor2_1 _6763_ (.B(_2806_),
    .A(_2805_),
    .X(_2807_));
 sg13g2_nand2_1 _6764_ (.Y(_2808_),
    .A(net1139),
    .B(_2796_));
 sg13g2_o21ai_1 _6765_ (.B1(_2808_),
    .Y(_2809_),
    .A1(net1139),
    .A2(net984));
 sg13g2_a221oi_1 _6766_ (.B2(_2666_),
    .C1(\i_display.frame_crotchet[6] ),
    .B1(_2809_),
    .A1(_2798_),
    .Y(_2810_),
    .A2(_2807_));
 sg13g2_a221oi_1 _6767_ (.B2(_2810_),
    .C1(net1159),
    .B1(net281),
    .A1(\i_display.frame_crotchet[6] ),
    .Y(_0222_),
    .A2(_2802_));
 sg13g2_nand2b_1 _6768_ (.Y(_2811_),
    .B(_2628_),
    .A_N(_2627_));
 sg13g2_nor2_1 _6769_ (.A(_2627_),
    .B(_2630_),
    .Y(_2812_));
 sg13g2_or2_1 _6770_ (.X(_2813_),
    .B(_2812_),
    .A(_2626_));
 sg13g2_nand3_1 _6771_ (.B(_2811_),
    .C(_2813_),
    .A(_2668_),
    .Y(_2814_));
 sg13g2_o21ai_1 _6772_ (.B1(_2812_),
    .Y(_2815_),
    .A1(_2626_),
    .A2(_2629_));
 sg13g2_nor2b_1 _6773_ (.A(_2722_),
    .B_N(net984),
    .Y(_2816_));
 sg13g2_xnor2_1 _6774_ (.Y(_2817_),
    .A(net980),
    .B(net984));
 sg13g2_nand3_1 _6775_ (.B(_2634_),
    .C(_2817_),
    .A(net1091),
    .Y(_2818_));
 sg13g2_a21oi_1 _6776_ (.A1(net1091),
    .A2(_2817_),
    .Y(_2819_),
    .B1(_2635_));
 sg13g2_nand4_1 _6777_ (.B(_2813_),
    .C(_2815_),
    .A(_2641_),
    .Y(_2820_),
    .D(_2818_));
 sg13g2_a21oi_1 _6778_ (.A1(net1091),
    .A2(_2819_),
    .Y(_2821_),
    .B1(_2964_));
 sg13g2_nand3_1 _6779_ (.B(_2820_),
    .C(_2821_),
    .A(_2814_),
    .Y(_2822_));
 sg13g2_nand2_1 _6780_ (.Y(_2823_),
    .A(net1139),
    .B(_2807_));
 sg13g2_nand2b_1 _6781_ (.Y(_2824_),
    .B(net980),
    .A_N(net1139));
 sg13g2_a21oi_1 _6782_ (.A1(_2823_),
    .A2(_2824_),
    .Y(_2825_),
    .B1(_2665_));
 sg13g2_or2_1 _6783_ (.X(_2826_),
    .B(_2825_),
    .A(_2788_));
 sg13g2_nor2_1 _6784_ (.A(_2909_),
    .B(_0024_),
    .Y(_2827_));
 sg13g2_nor2_1 _6785_ (.A(\i_display.in_line ),
    .B(_0025_),
    .Y(_2828_));
 sg13g2_nor4_2 _6786_ (.A(net1133),
    .B(_2781_),
    .C(_2827_),
    .Y(_2829_),
    .D(_2828_));
 sg13g2_a221oi_1 _6787_ (.B2(net1134),
    .C1(_2829_),
    .B1(_2826_),
    .A1(net1139),
    .Y(_2830_),
    .A2(_2783_));
 sg13g2_nor2_1 _6788_ (.A(net1135),
    .B(_2808_),
    .Y(_2831_));
 sg13g2_nor3_1 _6789_ (.A(_2789_),
    .B(_2825_),
    .C(_2831_),
    .Y(_2832_));
 sg13g2_o21ai_1 _6790_ (.B1(_2964_),
    .Y(_2833_),
    .A1(_2830_),
    .A2(_2832_));
 sg13g2_and3_1 _6791_ (.X(_0223_),
    .A(net1174),
    .B(_2822_),
    .C(_2833_));
 sg13g2_nand3_1 _6792_ (.B(_2813_),
    .C(_2815_),
    .A(_2668_),
    .Y(_2834_));
 sg13g2_nand2b_1 _6793_ (.Y(_2835_),
    .B(_2816_),
    .A_N(_2737_));
 sg13g2_xnor2_1 _6794_ (.Y(_2836_),
    .A(_2737_),
    .B(_2816_));
 sg13g2_o21ai_1 _6795_ (.B1(net381),
    .Y(_2837_),
    .A1(_2637_),
    .A2(_2836_));
 sg13g2_nand2b_1 _6796_ (.Y(_2838_),
    .B(_2834_),
    .A_N(_2837_));
 sg13g2_and2_1 _6797_ (.A(net980),
    .B(_2781_),
    .X(_2839_));
 sg13g2_nand2_1 _6798_ (.Y(_2840_),
    .A(_2917_),
    .B(net980));
 sg13g2_o21ai_1 _6799_ (.B1(_2840_),
    .Y(_2841_),
    .A1(_2805_),
    .A2(_2806_));
 sg13g2_xor2_1 _6800_ (.B(_2737_),
    .A(_0074_),
    .X(_2842_));
 sg13g2_xnor2_1 _6801_ (.Y(_2843_),
    .A(_2841_),
    .B(_2842_));
 sg13g2_xor2_1 _6802_ (.B(_2737_),
    .A(net1136),
    .X(_2844_));
 sg13g2_a21oi_1 _6803_ (.A1(net1140),
    .A2(_2843_),
    .Y(_2845_),
    .B1(_2665_));
 sg13g2_o21ai_1 _6804_ (.B1(_2845_),
    .Y(_2846_),
    .A1(net1139),
    .A2(_2844_));
 sg13g2_o21ai_1 _6805_ (.B1(_2846_),
    .Y(_2847_),
    .A1(_2778_),
    .A2(_2787_));
 sg13g2_a221oi_1 _6806_ (.B2(net1133),
    .C1(_2829_),
    .B1(_2847_),
    .A1(net1140),
    .Y(_2848_),
    .A2(_2839_));
 sg13g2_o21ai_1 _6807_ (.B1(_2846_),
    .Y(_2849_),
    .A1(net1135),
    .A2(_2823_));
 sg13g2_nor2_1 _6808_ (.A(_2789_),
    .B(_2849_),
    .Y(_2850_));
 sg13g2_o21ai_1 _6809_ (.B1(_2964_),
    .Y(_2851_),
    .A1(_2848_),
    .A2(_2850_));
 sg13g2_and3_1 _6810_ (.X(_0224_),
    .A(net1174),
    .B(_2838_),
    .C(_2851_));
 sg13g2_o21ai_1 _6811_ (.B1(_2627_),
    .Y(_2852_),
    .A1(_2629_),
    .A2(_2630_));
 sg13g2_and3_1 _6812_ (.X(_2853_),
    .A(_2626_),
    .B(_2631_),
    .C(_2852_));
 sg13g2_o21ai_1 _6813_ (.B1(_2627_),
    .Y(_2854_),
    .A1(_2628_),
    .A2(_2630_));
 sg13g2_nor2_1 _6814_ (.A(_2626_),
    .B(_2854_),
    .Y(_2855_));
 sg13g2_o21ai_1 _6815_ (.B1(_2668_),
    .Y(_2856_),
    .A1(_2853_),
    .A2(_2855_));
 sg13g2_nand2b_1 _6816_ (.Y(_2857_),
    .B(net933),
    .A_N(_2835_));
 sg13g2_nand2b_1 _6817_ (.Y(_2858_),
    .B(_2835_),
    .A_N(net933));
 sg13g2_nand4_1 _6818_ (.B(_2634_),
    .C(_2857_),
    .A(net1091),
    .Y(_2859_),
    .D(_2858_));
 sg13g2_mux2_1 _6819_ (.A0(_2852_),
    .A1(_2627_),
    .S(_2626_),
    .X(_2860_));
 sg13g2_inv_1 _6820_ (.Y(_2861_),
    .A(_2860_));
 sg13g2_or2_1 _6821_ (.X(_2862_),
    .B(_2860_),
    .A(_2642_));
 sg13g2_and4_1 _6822_ (.A(net351),
    .B(_2856_),
    .C(_2859_),
    .D(_2862_),
    .X(_2863_));
 sg13g2_and2_1 _6823_ (.A(net1136),
    .B(_2783_),
    .X(_2864_));
 sg13g2_o21ai_1 _6824_ (.B1(_2789_),
    .Y(_2865_),
    .A1(_2829_),
    .A2(_2864_));
 sg13g2_mux2_1 _6825_ (.A0(_2796_),
    .A1(_2807_),
    .S(_0053_),
    .X(_2866_));
 sg13g2_nand3_1 _6826_ (.B(_2788_),
    .C(_2866_),
    .A(_2418_),
    .Y(_2867_));
 sg13g2_nor2_1 _6827_ (.A(_0053_),
    .B(_2737_),
    .Y(_2868_));
 sg13g2_nand2_1 _6828_ (.Y(_2869_),
    .A(net933),
    .B(_2868_));
 sg13g2_xor2_1 _6829_ (.B(_2868_),
    .A(net933),
    .X(_2870_));
 sg13g2_a22oi_1 _6830_ (.Y(_2871_),
    .B1(_2841_),
    .B2(_2842_),
    .A2(_2737_),
    .A1(_2916_));
 sg13g2_xnor2_1 _6831_ (.Y(_2872_),
    .A(_2915_),
    .B(net933));
 sg13g2_nand2b_1 _6832_ (.Y(_2873_),
    .B(_2871_),
    .A_N(_2872_));
 sg13g2_nand2b_1 _6833_ (.Y(_2874_),
    .B(_2872_),
    .A_N(_2871_));
 sg13g2_nand3_1 _6834_ (.B(_2873_),
    .C(_2874_),
    .A(net1138),
    .Y(_2875_));
 sg13g2_o21ai_1 _6835_ (.B1(_2875_),
    .Y(_2876_),
    .A1(net1140),
    .A2(_2870_));
 sg13g2_nand2_1 _6836_ (.Y(_2877_),
    .A(_2666_),
    .B(_2876_));
 sg13g2_nand3_1 _6837_ (.B(_2867_),
    .C(_2877_),
    .A(_2865_),
    .Y(_2878_));
 sg13g2_o21ai_1 _6838_ (.B1(net1174),
    .Y(_2879_),
    .A1(net351),
    .A2(_2878_));
 sg13g2_nor2_1 _6839_ (.A(_2863_),
    .B(_2879_),
    .Y(_0225_));
 sg13g2_a21oi_1 _6840_ (.A1(net326),
    .A2(_2638_),
    .Y(_2880_),
    .B1(_2641_));
 sg13g2_xnor2_1 _6841_ (.Y(_2881_),
    .A(_2719_),
    .B(_2858_));
 sg13g2_o21ai_1 _6842_ (.B1(net351),
    .Y(_2882_),
    .A1(_2637_),
    .A2(_2881_));
 sg13g2_a21oi_1 _6843_ (.A1(_2861_),
    .A2(_2880_),
    .Y(_2883_),
    .B1(_2882_));
 sg13g2_a21o_1 _6844_ (.A2(_2839_),
    .A1(net1136),
    .B1(_2829_),
    .X(_2884_));
 sg13g2_nand4_1 _6845_ (.B(_2418_),
    .C(_2788_),
    .A(net1136),
    .Y(_2885_),
    .D(_2807_));
 sg13g2_o21ai_1 _6846_ (.B1(_2874_),
    .Y(_2886_),
    .A1(net1119),
    .A2(net933));
 sg13g2_xnor2_1 _6847_ (.Y(_2887_),
    .A(net1117),
    .B(_2719_));
 sg13g2_xnor2_1 _6848_ (.Y(_2888_),
    .A(_2886_),
    .B(_2887_));
 sg13g2_xnor2_1 _6849_ (.Y(_2889_),
    .A(net1136),
    .B(_2869_));
 sg13g2_xnor2_1 _6850_ (.Y(_2890_),
    .A(_2720_),
    .B(_2889_));
 sg13g2_o21ai_1 _6851_ (.B1(_2666_),
    .Y(_2891_),
    .A1(net1139),
    .A2(_2890_));
 sg13g2_a21o_1 _6852_ (.A2(_2888_),
    .A1(net1139),
    .B1(_2891_),
    .X(_2892_));
 sg13g2_nand3_1 _6853_ (.B(_2885_),
    .C(_2892_),
    .A(_2964_),
    .Y(_2893_));
 sg13g2_a21oi_1 _6854_ (.A1(_2789_),
    .A2(_2884_),
    .Y(_2894_),
    .B1(_2893_));
 sg13g2_nor3_1 _6855_ (.A(net1159),
    .B(_2883_),
    .C(_2894_),
    .Y(_0226_));
 sg13g2_nand2_1 _6856_ (.Y(_2895_),
    .A(net1115),
    .B(_0769_));
 sg13g2_a21oi_1 _6857_ (.A1(_0871_),
    .A2(_2895_),
    .Y(_0227_),
    .B1(net1161));
 sg13g2_mux2_1 _6858_ (.A0(_0857_),
    .A1(_2913_),
    .S(_0769_),
    .X(_2896_));
 sg13g2_nor2_1 _6859_ (.A(net1160),
    .B(_2896_),
    .Y(_0228_));
 sg13g2_nand2_1 _6860_ (.Y(_2897_),
    .A(net1110),
    .B(_0769_));
 sg13g2_a21oi_1 _6861_ (.A1(_0802_),
    .A2(_2897_),
    .Y(_0229_),
    .B1(net1160));
 sg13g2_nand2_1 _6862_ (.Y(_2898_),
    .A(net1106),
    .B(_0769_));
 sg13g2_a21oi_1 _6863_ (.A1(_0845_),
    .A2(_2898_),
    .Y(_0230_),
    .B1(net1160));
 sg13g2_nand2_1 _6864_ (.Y(_2899_),
    .A(net1099),
    .B(_0769_));
 sg13g2_a21oi_1 _6865_ (.A1(_0826_),
    .A2(_2899_),
    .Y(_0231_),
    .B1(net1160));
 sg13g2_nand2_1 _6866_ (.Y(_2900_),
    .A(net1098),
    .B(_0769_));
 sg13g2_a21oi_1 _6867_ (.A1(_0816_),
    .A2(_2900_),
    .Y(_0232_),
    .B1(net1161));
 sg13g2_nor3_1 _6868_ (.A(_3118_),
    .B(_3164_),
    .C(_0769_),
    .Y(_2901_));
 sg13g2_o21ai_1 _6869_ (.B1(_2367_),
    .Y(_2902_),
    .A1(net224),
    .A2(_2901_));
 sg13g2_a21oi_1 _6870_ (.A1(net224),
    .A2(_2901_),
    .Y(_0233_),
    .B1(_2902_));
 sg13g2_nor2_2 _6871_ (.A(net1161),
    .B(net1022),
    .Y(_2903_));
 sg13g2_o21ai_1 _6872_ (.B1(_2903_),
    .Y(_2904_),
    .A1(net297),
    .A2(_0766_));
 sg13g2_a21oi_1 _6873_ (.A1(_2910_),
    .A2(_0766_),
    .Y(_0234_),
    .B1(_2904_));
 sg13g2_nor2_1 _6874_ (.A(net1093),
    .B(_0766_),
    .Y(_2905_));
 sg13g2_and3_1 _6875_ (.X(_2906_),
    .A(_3109_),
    .B(_3188_),
    .C(_0766_));
 sg13g2_nor4_1 _6876_ (.A(net1161),
    .B(net1025),
    .C(_2905_),
    .D(_2906_),
    .Y(_0235_));
 sg13g2_o21ai_1 _6877_ (.B1(_2903_),
    .Y(_2907_),
    .A1(net1091),
    .A2(_0766_));
 sg13g2_a21oi_1 _6878_ (.A1(_2908_),
    .A2(_0766_),
    .Y(_0236_),
    .B1(_2907_));
 sg13g2_dfrbp_1 _6879_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net25),
    .D(_0000_),
    .Q_N(_0082_),
    .Q(\i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[0] ));
 sg13g2_dfrbp_1 _6880_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net26),
    .D(_0001_),
    .Q_N(_0091_),
    .Q(\i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[1] ));
 sg13g2_dfrbp_1 _6881_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net27),
    .D(_0002_),
    .Q_N(_0094_),
    .Q(\i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[2] ));
 sg13g2_dfrbp_1 _6882_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net28),
    .D(_0003_),
    .Q_N(_0027_),
    .Q(\i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[3] ));
 sg13g2_dfrbp_1 _6883_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net29),
    .D(_0004_),
    .Q_N(_0029_),
    .Q(\i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[4] ));
 sg13g2_dfrbp_1 _6884_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net30),
    .D(_0005_),
    .Q_N(_0030_),
    .Q(\i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[5] ));
 sg13g2_dfrbp_1 _6885_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net31),
    .D(_0006_),
    .Q_N(_0031_),
    .Q(\i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[6] ));
 sg13g2_dfrbp_1 _6886_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net50),
    .D(_0007_),
    .Q_N(_0032_),
    .Q(\i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[7] ));
 sg13g2_dfrbp_1 _6887_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net24),
    .D(_0008_),
    .Q_N(_0033_),
    .Q(\i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[8] ));
 sg13g2_dfrbp_1 _6888_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net109),
    .D(_0101_),
    .Q_N(_3401_),
    .Q(\i_music.violin_note_idx[2][4] ));
 sg13g2_dfrbp_1 _6889_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net108),
    .D(_0102_),
    .Q_N(_3400_),
    .Q(\i_music.violin_note_idx[2][5] ));
 sg13g2_dfrbp_1 _6890_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net107),
    .D(_0103_),
    .Q_N(_3399_),
    .Q(\i_music.violin_note_idx[2][6] ));
 sg13g2_dfrbp_1 _6891_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net106),
    .D(net277),
    .Q_N(_3398_),
    .Q(\i_music.violin_note_idx[2][7] ));
 sg13g2_dfrbp_1 _6892_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net105),
    .D(_0105_),
    .Q_N(_3397_),
    .Q(\i_music.violin_note_idx[2][8] ));
 sg13g2_dfrbp_1 _6893_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net104),
    .D(_0106_),
    .Q_N(_3396_),
    .Q(\i_music.i_sample.sample_acc[8] ));
 sg13g2_dfrbp_1 _6894_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net103),
    .D(_0107_),
    .Q_N(_0060_),
    .Q(\i_music.i_sample.sample_acc[7] ));
 sg13g2_dfrbp_1 _6895_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net102),
    .D(_0108_),
    .Q_N(_3395_),
    .Q(\i_music.i_sample.thresh[10] ));
 sg13g2_dfrbp_1 _6896_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net101),
    .D(_0109_),
    .Q_N(_3394_),
    .Q(\i_music.violin_note_idx[3][0] ));
 sg13g2_dfrbp_1 _6897_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net99),
    .D(_0110_),
    .Q_N(_3393_),
    .Q(\i_music.violin_note_idx[3][4] ));
 sg13g2_dfrbp_1 _6898_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net98),
    .D(_0111_),
    .Q_N(_3392_),
    .Q(\i_music.violin_note_idx[3][5] ));
 sg13g2_dfrbp_1 _6899_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net97),
    .D(_0112_),
    .Q_N(_3391_),
    .Q(\i_music.violin_note_idx[3][6] ));
 sg13g2_dfrbp_1 _6900_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net96),
    .D(net221),
    .Q_N(_0043_),
    .Q(\i_music.violin_note_idx[3][7] ));
 sg13g2_dfrbp_1 _6901_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net95),
    .D(_0114_),
    .Q_N(_3390_),
    .Q(\i_music.violin_note_idx[3][8] ));
 sg13g2_dfrbp_1 _6902_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net94),
    .D(net309),
    .Q_N(_3389_),
    .Q(\i_music.violin_note_idx[3][1] ));
 sg13g2_dfrbp_1 _6903_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net74),
    .D(net307),
    .Q_N(_3388_),
    .Q(\i_music.violin_note_idx[3][2] ));
 sg13g2_dfrbp_1 _6904_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net72),
    .D(_0117_),
    .Q_N(_3387_),
    .Q(\i_music.violin_note_idx[3][3] ));
 sg13g2_dfrbp_1 _6905_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net51),
    .D(_0118_),
    .Q_N(_3402_),
    .Q(\i_display.y_value$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:567$12.$result[9] ));
 sg13g2_dfrbp_1 _6906_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net52),
    .D(_0018_),
    .Q_N(_3403_),
    .Q(_0025_));
 sg13g2_dfrbp_1 _6907_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net53),
    .D(_0017_),
    .Q_N(_3404_),
    .Q(_0024_));
 sg13g2_dfrbp_1 _6908_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net54),
    .D(_0009_),
    .Q_N(_0070_),
    .Q(\i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[-5] ));
 sg13g2_dfrbp_1 _6909_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net55),
    .D(_0010_),
    .Q_N(_0072_),
    .Q(\i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[-4] ));
 sg13g2_dfrbp_1 _6910_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net56),
    .D(_0011_),
    .Q_N(_0076_),
    .Q(\i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[-3] ));
 sg13g2_dfrbp_1 _6911_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net57),
    .D(_0012_),
    .Q_N(_0073_),
    .Q(\i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[-2] ));
 sg13g2_dfrbp_1 _6912_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net58),
    .D(_0013_),
    .Q_N(_0078_),
    .Q(\i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[-1] ));
 sg13g2_dfrbp_1 _6913_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net59),
    .D(_0014_),
    .Q_N(_0080_),
    .Q(\i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[0] ));
 sg13g2_dfrbp_1 _6914_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net76),
    .D(_0015_),
    .Q_N(_0090_),
    .Q(\i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[1] ));
 sg13g2_dfrbp_1 _6915_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net70),
    .D(_0016_),
    .Q_N(_0093_),
    .Q(\i_display.y_offset$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/display.sv:565$10.$result[2] ));
 sg13g2_dfrbp_1 _6916_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net69),
    .D(_0119_),
    .Q_N(_0098_),
    .Q(\i_music.i_pwm.count[0] ));
 sg13g2_dfrbp_1 _6917_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net68),
    .D(net302),
    .Q_N(_3386_),
    .Q(\i_music.i_pwm.count[1] ));
 sg13g2_dfrbp_1 _6918_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net67),
    .D(net229),
    .Q_N(_3385_),
    .Q(\i_music.i_pwm.count[2] ));
 sg13g2_dfrbp_1 _6919_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net66),
    .D(_0122_),
    .Q_N(_3384_),
    .Q(\i_music.i_pwm.count[3] ));
 sg13g2_dfrbp_1 _6920_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net65),
    .D(_0123_),
    .Q_N(_3383_),
    .Q(\i_music.i_pwm.count[4] ));
 sg13g2_dfrbp_1 _6921_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net64),
    .D(_0124_),
    .Q_N(_3382_),
    .Q(\i_music.i_pwm.count[5] ));
 sg13g2_dfrbp_1 _6922_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net63),
    .D(_0125_),
    .Q_N(_3381_),
    .Q(\i_music.i_pwm.count[6] ));
 sg13g2_dfrbp_1 _6923_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net62),
    .D(_0126_),
    .Q_N(_3380_),
    .Q(\i_music.i_pwm.count[7] ));
 sg13g2_dfrbp_1 _6924_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net61),
    .D(net291),
    .Q_N(_3379_),
    .Q(\i_music.i_pwm.sample[0] ));
 sg13g2_dfrbp_1 _6925_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net60),
    .D(_0128_),
    .Q_N(_3378_),
    .Q(\i_music.i_pwm.sample[1] ));
 sg13g2_dfrbp_1 _6926_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net49),
    .D(net248),
    .Q_N(_3377_),
    .Q(\i_music.i_pwm.sample[2] ));
 sg13g2_dfrbp_1 _6927_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net48),
    .D(_0130_),
    .Q_N(_3376_),
    .Q(\i_music.i_pwm.sample[3] ));
 sg13g2_dfrbp_1 _6928_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net47),
    .D(net233),
    .Q_N(_3375_),
    .Q(\i_music.i_pwm.sample[4] ));
 sg13g2_dfrbp_1 _6929_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net46),
    .D(_0132_),
    .Q_N(_3374_),
    .Q(\i_music.i_pwm.sample[5] ));
 sg13g2_dfrbp_1 _6930_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net45),
    .D(net272),
    .Q_N(_3373_),
    .Q(\i_music.i_pwm.sample[6] ));
 sg13g2_dfrbp_1 _6931_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net77),
    .D(net244),
    .Q_N(_3405_),
    .Q(\i_music.i_pwm.sample[7] ));
 sg13g2_dfrbp_1 _6932_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net78),
    .D(_0237_),
    .Q_N(_3406_),
    .Q(\i_music.i_sample.sample_idx[0] ));
 sg13g2_dfrbp_1 _6933_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net79),
    .D(_0238_),
    .Q_N(_3407_),
    .Q(\i_music.i_sample.sample_idx[1] ));
 sg13g2_dfrbp_1 _6934_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net80),
    .D(_0239_),
    .Q_N(_3408_),
    .Q(\i_music.i_sample.sample_idx[2] ));
 sg13g2_dfrbp_1 _6935_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net81),
    .D(_0240_),
    .Q_N(_3409_),
    .Q(\i_music.i_sample.sample_idx[3] ));
 sg13g2_dfrbp_1 _6936_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net82),
    .D(_0241_),
    .Q_N(_3410_),
    .Q(\i_music.i_sample.sample_idx[4] ));
 sg13g2_dfrbp_1 _6937_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net83),
    .D(_0242_),
    .Q_N(_3411_),
    .Q(\i_music.i_sample.sample_idx[5] ));
 sg13g2_dfrbp_1 _6938_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net84),
    .D(_0243_),
    .Q_N(_3412_),
    .Q(\i_music.i_sample.sample_idx[6] ));
 sg13g2_dfrbp_1 _6939_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net85),
    .D(_0244_),
    .Q_N(_3413_),
    .Q(\i_music.i_sample.sample_idx[7] ));
 sg13g2_dfrbp_1 _6940_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net86),
    .D(_0245_),
    .Q_N(_0068_),
    .Q(\i_music.i_sample.thresh[0] ));
 sg13g2_dfrbp_1 _6941_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net87),
    .D(_0246_),
    .Q_N(_0056_),
    .Q(\i_music.i_sample.thresh[1] ));
 sg13g2_dfrbp_1 _6942_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net88),
    .D(_0247_),
    .Q_N(_0057_),
    .Q(\i_music.i_sample.thresh[2] ));
 sg13g2_dfrbp_1 _6943_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net89),
    .D(_0248_),
    .Q_N(_0058_),
    .Q(\i_music.i_sample.thresh[3] ));
 sg13g2_dfrbp_1 _6944_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net90),
    .D(_0249_),
    .Q_N(_0065_),
    .Q(\i_music.i_sample.thresh[4] ));
 sg13g2_dfrbp_1 _6945_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net91),
    .D(_0250_),
    .Q_N(_0059_),
    .Q(\i_music.i_sample.thresh[5] ));
 sg13g2_dfrbp_1 _6946_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net92),
    .D(_0251_),
    .Q_N(_3414_),
    .Q(\i_music.i_sample.thresh[6] ));
 sg13g2_dfrbp_1 _6947_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net93),
    .D(_0252_),
    .Q_N(_3415_),
    .Q(\i_music.i_sample.thresh[7] ));
 sg13g2_dfrbp_1 _6948_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net142),
    .D(_0253_),
    .Q_N(_3416_),
    .Q(\i_music.i_sample.thresh[8] ));
 sg13g2_dfrbp_1 _6949_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net44),
    .D(_0254_),
    .Q_N(_3372_),
    .Q(\i_music.i_sample.thresh[9] ));
 sg13g2_dlhq_1 _6950_ (.D(\i_music.i_sample.t1.genblk1[18].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[18].state.Q ));
 sg13g2_dlhq_1 _6951_ (.D(\i_music.i_sample.t1.genblk1[17].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[17].state.Q ));
 sg13g2_dlhq_1 _6952_ (.D(\i_music.i_sample.t1.genblk1[16].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[16].state.Q ));
 sg13g2_dlhq_1 _6953_ (.D(\i_music.i_sample.t1.genblk1[15].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[15].state.Q ));
 sg13g2_dlhq_1 _6954_ (.D(\i_music.i_sample.t1.genblk1[14].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[14].state.Q ));
 sg13g2_dlhq_1 _6955_ (.D(\i_music.i_sample.t1.genblk1[13].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[13].state.Q ));
 sg13g2_dlhq_1 _6956_ (.D(\i_music.i_sample.t1.genblk1[12].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[12].state.Q ));
 sg13g2_dlhq_1 _6957_ (.D(\i_music.i_sample.t1.genblk1[11].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[11].state.Q ));
 sg13g2_dlhq_1 _6958_ (.D(\i_music.i_sample.t1.genblk1[10].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[10].state.Q ));
 sg13g2_dlhq_1 _6959_ (.D(\i_music.i_sample.t1.genblk1[9].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[9].state.Q ));
 sg13g2_dlhq_1 _6960_ (.D(\i_music.i_sample.t1.genblk1[8].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[8].state.Q ));
 sg13g2_dlhq_1 _6961_ (.D(\i_music.i_sample.t1.genblk1[7].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[7].state.Q ));
 sg13g2_dlhq_1 _6962_ (.D(\i_music.i_sample.t1.genblk1[6].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[6].state.Q ));
 sg13g2_dlhq_1 _6963_ (.D(\i_music.i_sample.t1.genblk1[5].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[5].state.Q ));
 sg13g2_dlhq_1 _6964_ (.D(\i_music.i_sample.t1.genblk1[4].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[4].state.Q ));
 sg13g2_dlhq_1 _6965_ (.D(\i_music.i_sample.t1.genblk1[3].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[3].state.Q ));
 sg13g2_dlhq_1 _6966_ (.D(\i_music.i_sample.t1.genblk1[2].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[2].state.Q ));
 sg13g2_dlhq_1 _6967_ (.D(\i_music.i_sample.t1.genblk1[1].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[1].state.Q ));
 sg13g2_dlhq_1 _6968_ (.D(\i_music.i_sample.t1.genblk1[0].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[0].state.Q ));
 sg13g2_dlhq_1 _6969_ (.D(\i_music.i_sample.t1.genblk1[17].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[17].state.Q ));
 sg13g2_dlhq_1 _6970_ (.D(\i_music.i_sample.t1.genblk1[16].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[16].state.Q ));
 sg13g2_dlhq_1 _6971_ (.D(\i_music.i_sample.t1.genblk1[15].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[15].state.Q ));
 sg13g2_dlhq_1 _6972_ (.D(\i_music.i_sample.t1.genblk1[14].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[14].state.Q ));
 sg13g2_dlhq_1 _6973_ (.D(\i_music.i_sample.t1.genblk1[13].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[13].state.Q ));
 sg13g2_dlhq_1 _6974_ (.D(\i_music.i_sample.t1.genblk1[12].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[12].state.Q ));
 sg13g2_dlhq_1 _6975_ (.D(\i_music.i_sample.t1.genblk1[11].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[11].state.Q ));
 sg13g2_dlhq_1 _6976_ (.D(\i_music.i_sample.t1.genblk1[10].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[10].state.Q ));
 sg13g2_dlhq_1 _6977_ (.D(\i_music.i_sample.t1.genblk1[9].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[9].state.Q ));
 sg13g2_dlhq_1 _6978_ (.D(\i_music.i_sample.t1.genblk1[8].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[8].state.Q ));
 sg13g2_dlhq_1 _6979_ (.D(\i_music.i_sample.t1.genblk1[7].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[7].state.Q ));
 sg13g2_dlhq_1 _6980_ (.D(\i_music.i_sample.t1.genblk1[6].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[6].state.Q ));
 sg13g2_dlhq_1 _6981_ (.D(\i_music.i_sample.t1.genblk1[5].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[5].state.Q ));
 sg13g2_dlhq_1 _6982_ (.D(\i_music.i_sample.t1.genblk1[4].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[4].state.Q ));
 sg13g2_dlhq_1 _6983_ (.D(\i_music.i_sample.t1.genblk1[3].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[3].state.Q ));
 sg13g2_dlhq_1 _6984_ (.D(\i_music.i_sample.t1.genblk1[2].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[2].state.Q ));
 sg13g2_dlhq_1 _6985_ (.D(\i_music.i_sample.t1.genblk1[1].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[1].state.Q ));
 sg13g2_dlhq_1 _6986_ (.D(\i_music.i_sample.t1.genblk1[0].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[0].state.Q ));
 sg13g2_dlhq_1 _6987_ (.D(\i_music.i_sample.t1.genblk1[17].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[17].state.Q ));
 sg13g2_dlhq_1 _6988_ (.D(\i_music.i_sample.t1.genblk1[16].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[16].state.Q ));
 sg13g2_dlhq_1 _6989_ (.D(\i_music.i_sample.t1.genblk1[15].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[15].state.Q ));
 sg13g2_dlhq_1 _6990_ (.D(\i_music.i_sample.t1.genblk1[14].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[14].state.Q ));
 sg13g2_dlhq_1 _6991_ (.D(\i_music.i_sample.t1.genblk1[13].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[13].state.Q ));
 sg13g2_dlhq_1 _6992_ (.D(\i_music.i_sample.t1.genblk1[12].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[12].state.Q ));
 sg13g2_dlhq_1 _6993_ (.D(\i_music.i_sample.t1.genblk1[11].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[11].state.Q ));
 sg13g2_dlhq_1 _6994_ (.D(\i_music.i_sample.t1.genblk1[10].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[10].state.Q ));
 sg13g2_dlhq_1 _6995_ (.D(\i_music.i_sample.t1.genblk1[9].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[9].state.Q ));
 sg13g2_dlhq_1 _6996_ (.D(\i_music.i_sample.t1.genblk1[8].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[8].state.Q ));
 sg13g2_dlhq_1 _6997_ (.D(\i_music.i_sample.t1.genblk1[7].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[7].state.Q ));
 sg13g2_dlhq_1 _6998_ (.D(\i_music.i_sample.t1.genblk1[6].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[6].state.Q ));
 sg13g2_dlhq_1 _6999_ (.D(\i_music.i_sample.t1.genblk1[5].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[5].state.Q ));
 sg13g2_dlhq_1 _7000_ (.D(\i_music.i_sample.t1.genblk1[4].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[4].state.Q ));
 sg13g2_dlhq_1 _7001_ (.D(\i_music.i_sample.t1.genblk1[3].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[3].state.Q ));
 sg13g2_dlhq_1 _7002_ (.D(\i_music.i_sample.t1.genblk1[2].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[2].state.Q ));
 sg13g2_dlhq_1 _7003_ (.D(\i_music.i_sample.t1.genblk1[1].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[1].state.Q ));
 sg13g2_dlhq_1 _7004_ (.D(\i_music.i_sample.t1.genblk1[0].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[0].state.Q ));
 sg13g2_dlhq_1 _7005_ (.D(\i_music.i_sample.t1.genblk1[17].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[17].state.Q ));
 sg13g2_dlhq_1 _7006_ (.D(\i_music.i_sample.t1.genblk1[16].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[16].state.Q ));
 sg13g2_dlhq_1 _7007_ (.D(\i_music.i_sample.t1.genblk1[15].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[15].state.Q ));
 sg13g2_dlhq_1 _7008_ (.D(\i_music.i_sample.t1.genblk1[14].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[14].state.Q ));
 sg13g2_dlhq_1 _7009_ (.D(\i_music.i_sample.t1.genblk1[13].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[13].state.Q ));
 sg13g2_dlhq_1 _7010_ (.D(\i_music.i_sample.t1.genblk1[12].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[12].state.Q ));
 sg13g2_dlhq_1 _7011_ (.D(\i_music.i_sample.t1.genblk1[11].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[11].state.Q ));
 sg13g2_dlhq_1 _7012_ (.D(\i_music.i_sample.t1.genblk1[10].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[10].state.Q ));
 sg13g2_dlhq_1 _7013_ (.D(\i_music.i_sample.t1.genblk1[9].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[9].state.Q ));
 sg13g2_dlhq_1 _7014_ (.D(\i_music.i_sample.t1.genblk1[8].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[8].state.Q ));
 sg13g2_dlhq_1 _7015_ (.D(\i_music.i_sample.t1.genblk1[7].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[7].state.Q ));
 sg13g2_dlhq_1 _7016_ (.D(\i_music.i_sample.t1.genblk1[6].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[6].state.Q ));
 sg13g2_dlhq_1 _7017_ (.D(\i_music.i_sample.t1.genblk1[5].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[5].state.Q ));
 sg13g2_dlhq_1 _7018_ (.D(\i_music.i_sample.t1.genblk1[4].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[4].state.Q ));
 sg13g2_dlhq_1 _7019_ (.D(\i_music.i_sample.t1.genblk1[3].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[3].state.Q ));
 sg13g2_dlhq_1 _7020_ (.D(\i_music.i_sample.t1.genblk1[2].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[2].state.Q ));
 sg13g2_dlhq_1 _7021_ (.D(\i_music.i_sample.t1.genblk1[1].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[1].state.Q ));
 sg13g2_dlhq_1 _7022_ (.D(\i_music.i_sample.t1.genblk1[0].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[0].state.Q ));
 sg13g2_dfrbp_1 _7023_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net43),
    .D(_0135_),
    .Q_N(_0097_),
    .Q(\i_display.i_vga.low_count[0] ));
 sg13g2_dfrbp_1 _7024_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net42),
    .D(_0136_),
    .Q_N(_0067_),
    .Q(\i_display.i_vga.low_count[1] ));
 sg13g2_dfrbp_1 _7025_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net41),
    .D(_0137_),
    .Q_N(_0061_),
    .Q(\i_display.i_vga.low_count[2] ));
 sg13g2_dfrbp_1 _7026_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net40),
    .D(_0138_),
    .Q_N(_0066_),
    .Q(\i_display.i_vga.low_count[3] ));
 sg13g2_dfrbp_1 _7027_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net39),
    .D(_0139_),
    .Q_N(_0062_),
    .Q(\i_display.i_vga.low_count[4] ));
 sg13g2_dfrbp_1 _7028_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net38),
    .D(_0140_),
    .Q_N(_0064_),
    .Q(\i_display.i_vga.low_count[5] ));
 sg13g2_dfrbp_1 _7029_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net37),
    .D(_0141_),
    .Q_N(_0046_),
    .Q(\i_display.i_vga.low_count[6] ));
 sg13g2_dfrbp_1 _7030_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net36),
    .D(_0142_),
    .Q_N(_0063_),
    .Q(\i_display.i_vga.low_count[7] ));
 sg13g2_dfrbp_1 _7031_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net35),
    .D(net211),
    .Q_N(_0045_),
    .Q(\i_display.i_vga.low_count[8] ));
 sg13g2_dfrbp_1 _7032_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net34),
    .D(_0144_),
    .Q_N(_3371_),
    .Q(\i_display.i_vga.low_count[9] ));
 sg13g2_dfrbp_1 _7033_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net33),
    .D(_0145_),
    .Q_N(_3370_),
    .Q(\i_music.count[10] ));
 sg13g2_dfrbp_1 _7034_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net32),
    .D(_0146_),
    .Q_N(_3369_),
    .Q(\i_music.count[11] ));
 sg13g2_dfrbp_1 _7035_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net23),
    .D(_0147_),
    .Q_N(_3368_),
    .Q(\i_music.count[12] ));
 sg13g2_dfrbp_1 _7036_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net204),
    .D(_0148_),
    .Q_N(_3367_),
    .Q(\i_music.count[13] ));
 sg13g2_dfrbp_1 _7037_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net203),
    .D(_0149_),
    .Q_N(_3366_),
    .Q(\i_music.count[14] ));
 sg13g2_dfrbp_1 _7038_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net202),
    .D(_0150_),
    .Q_N(_3365_),
    .Q(\i_music.count[15] ));
 sg13g2_dfrbp_1 _7039_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net201),
    .D(_0151_),
    .Q_N(_3364_),
    .Q(\i_music.count[16] ));
 sg13g2_dfrbp_1 _7040_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net200),
    .D(_0152_),
    .Q_N(_3363_),
    .Q(\i_music.count[17] ));
 sg13g2_dfrbp_1 _7041_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net199),
    .D(_0153_),
    .Q_N(_3362_),
    .Q(\i_music.count[18] ));
 sg13g2_dfrbp_1 _7042_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net198),
    .D(_0154_),
    .Q_N(_3361_),
    .Q(\i_music.count[19] ));
 sg13g2_dfrbp_1 _7043_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net197),
    .D(_0155_),
    .Q_N(_3360_),
    .Q(\i_music.count[20] ));
 sg13g2_dfrbp_1 _7044_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net196),
    .D(_0156_),
    .Q_N(_3359_),
    .Q(\i_music.count[21] ));
 sg13g2_dfrbp_1 _7045_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net195),
    .D(_0157_),
    .Q_N(_0035_),
    .Q(\i_music.count[22] ));
 sg13g2_dfrbp_1 _7046_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net194),
    .D(net238),
    .Q_N(_3358_),
    .Q(\i_music.count[23] ));
 sg13g2_dfrbp_1 _7047_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net193),
    .D(_0159_),
    .Q_N(_3357_),
    .Q(\i_music.count[24] ));
 sg13g2_dfrbp_1 _7048_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net192),
    .D(_0160_),
    .Q_N(_0047_),
    .Q(\crotchet[0] ));
 sg13g2_dfrbp_1 _7049_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net191),
    .D(_0161_),
    .Q_N(_3356_),
    .Q(\crotchet[1] ));
 sg13g2_dfrbp_1 _7050_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net190),
    .D(_0162_),
    .Q_N(_3355_),
    .Q(\crotchet[2] ));
 sg13g2_dfrbp_1 _7051_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net189),
    .D(_0163_),
    .Q_N(_3354_),
    .Q(\crotchet[3] ));
 sg13g2_dfrbp_1 _7052_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net188),
    .D(_0164_),
    .Q_N(_3353_),
    .Q(\crotchet[4] ));
 sg13g2_dfrbp_1 _7053_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net187),
    .D(_0165_),
    .Q_N(_3352_),
    .Q(\crotchet[5] ));
 sg13g2_dfrbp_1 _7054_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net186),
    .D(net269),
    .Q_N(_3351_),
    .Q(\crotchet[6] ));
 sg13g2_dfrbp_1 _7055_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net185),
    .D(net216),
    .Q_N(_3350_),
    .Q(\i_music.i_pwm.pwm ));
 sg13g2_dfrbp_1 _7056_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net184),
    .D(net329),
    .Q_N(_0040_),
    .Q(\i_music.violin_note_idx[1][1] ));
 sg13g2_dfrbp_1 _7057_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net182),
    .D(net295),
    .Q_N(_0041_),
    .Q(\i_music.violin_note_idx[1][2] ));
 sg13g2_dfrbp_1 _7058_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net180),
    .D(net264),
    .Q_N(_0037_),
    .Q(\i_music.violin_note_idx[1][3] ));
 sg13g2_dfrbp_1 _7059_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net178),
    .D(net251),
    .Q_N(_3349_),
    .Q(\i_music.violin_note_idx[2][1] ));
 sg13g2_dfrbp_1 _7060_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net176),
    .D(net253),
    .Q_N(_3348_),
    .Q(\i_music.violin_note_idx[2][2] ));
 sg13g2_dfrbp_1 _7061_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net174),
    .D(net223),
    .Q_N(_3347_),
    .Q(\i_music.violin_note_idx[2][3] ));
 sg13g2_dfrbp_1 _7062_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net172),
    .D(net259),
    .Q_N(_3346_),
    .Q(\i_display.frame_crotchet[0] ));
 sg13g2_dfrbp_1 _7063_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net171),
    .D(_0175_),
    .Q_N(_0052_),
    .Q(\i_display.frame_crotchet[1] ));
 sg13g2_dfrbp_1 _7064_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net170),
    .D(_0176_),
    .Q_N(_0051_),
    .Q(\i_display.frame_crotchet[2] ));
 sg13g2_dfrbp_1 _7065_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net169),
    .D(_0177_),
    .Q_N(_0053_),
    .Q(\i_display.frame_crotchet[3] ));
 sg13g2_dfrbp_1 _7066_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net168),
    .D(_0178_),
    .Q_N(_0050_),
    .Q(\i_display.frame_crotchet[4] ));
 sg13g2_dfrbp_1 _7067_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net163),
    .D(_0179_),
    .Q_N(_0049_),
    .Q(\i_display.frame_crotchet[5] ));
 sg13g2_dfrbp_1 _7068_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net162),
    .D(_0180_),
    .Q_N(_0048_),
    .Q(\i_display.frame_crotchet[6] ));
 sg13g2_dfrbp_1 _7069_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net161),
    .D(_0181_),
    .Q_N(_3345_),
    .Q(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[5] ));
 sg13g2_dfrbp_1 _7070_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net143),
    .D(net235),
    .Q_N(_0099_),
    .Q(\i_music.violin_note_idx[2][0] ));
 sg13g2_dfrbp_1 _7071_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net144),
    .D(_0019_),
    .Q_N(_3417_),
    .Q(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[0] ));
 sg13g2_dfrbp_1 _7072_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net145),
    .D(_0020_),
    .Q_N(_3418_),
    .Q(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[2] ));
 sg13g2_dfrbp_1 _7073_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net146),
    .D(_0021_),
    .Q_N(_3419_),
    .Q(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[6] ));
 sg13g2_dfrbp_1 _7074_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net164),
    .D(_0022_),
    .Q_N(_3420_),
    .Q(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[7] ));
 sg13g2_dfrbp_1 _7075_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net160),
    .D(_0023_),
    .Q_N(_3344_),
    .Q(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[8] ));
 sg13g2_dfrbp_1 _7076_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net158),
    .D(_0183_),
    .Q_N(_3343_),
    .Q(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[1] ));
 sg13g2_dfrbp_1 _7077_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net157),
    .D(_0184_),
    .Q_N(_3342_),
    .Q(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[3] ));
 sg13g2_dfrbp_1 _7078_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net156),
    .D(_0185_),
    .Q_N(_3341_),
    .Q(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[4] ));
 sg13g2_dfrbp_1 _7079_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net155),
    .D(_0186_),
    .Q_N(_3340_),
    .Q(\i_music.cello_rom$func$/home/runner/work/tinytapeout-ihp-25a-sources/tinytapeout-ihp-25a-sources/tt08-hdl/tt_um_MichaelBell_canon/src/music.v:430$166.$result[10] ));
 sg13g2_dfrbp_1 _7080_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net154),
    .D(net305),
    .Q_N(_0038_),
    .Q(\i_music.violin_note_idx[1][4] ));
 sg13g2_dfrbp_1 _7081_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net153),
    .D(_0188_),
    .Q_N(_0036_),
    .Q(\i_music.violin_note_idx[1][5] ));
 sg13g2_dfrbp_1 _7082_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net152),
    .D(_0189_),
    .Q_N(_0039_),
    .Q(\i_music.violin_note_idx[1][6] ));
 sg13g2_dfrbp_1 _7083_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net151),
    .D(_0190_),
    .Q_N(_0042_),
    .Q(\i_music.violin_note_idx[1][7] ));
 sg13g2_dfrbp_1 _7084_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net150),
    .D(net321),
    .Q_N(_0044_),
    .Q(\i_music.violin_note_idx[1][8] ));
 sg13g2_dfrbp_1 _7085_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net149),
    .D(_0192_),
    .Q_N(_3339_),
    .Q(\i_music.i_sample.sample_acc[0] ));
 sg13g2_dfrbp_1 _7086_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net148),
    .D(_0193_),
    .Q_N(_3338_),
    .Q(\i_music.i_sample.sample_acc[1] ));
 sg13g2_dfrbp_1 _7087_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net147),
    .D(_0194_),
    .Q_N(_3337_),
    .Q(\i_music.i_sample.sample_acc[2] ));
 sg13g2_dfrbp_1 _7088_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net141),
    .D(_0195_),
    .Q_N(_0054_),
    .Q(\i_music.i_sample.sample_acc[3] ));
 sg13g2_dfrbp_1 _7089_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net140),
    .D(_0196_),
    .Q_N(_3336_),
    .Q(\i_music.i_sample.sample_acc[4] ));
 sg13g2_dfrbp_1 _7090_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net139),
    .D(_0197_),
    .Q_N(_0055_),
    .Q(\i_music.i_sample.sample_acc[5] ));
 sg13g2_dfrbp_1 _7091_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net138),
    .D(_0198_),
    .Q_N(_3335_),
    .Q(\i_music.i_sample.sample_acc[6] ));
 sg13g2_dfrbp_1 _7092_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net165),
    .D(net231),
    .Q_N(_0100_),
    .Q(\i_music.violin_note_idx[1][0] ));
 sg13g2_dfrbp_1 _7093_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net166),
    .D(net246),
    .Q_N(_3421_),
    .Q(\i_display.hsync ));
 sg13g2_dfrbp_1 _7094_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net167),
    .D(net208),
    .Q_N(_3422_),
    .Q(\i_display.i_vga.vblank ));
 sg13g2_dfrbp_1 _7095_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net181),
    .D(\i_display.i_vga.hblank_tmp ),
    .Q_N(_3423_),
    .Q(\i_display.i_vga.hblank ));
 sg13g2_dfrbp_1 _7096_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net137),
    .D(net214),
    .Q_N(_3334_),
    .Q(\i_display.i_vga.timing_ver.sync ));
 sg13g2_dfrbp_1 _7097_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net135),
    .D(_0200_),
    .Q_N(_3333_),
    .Q(\i_display.i_vga.timing_ver.counter[0] ));
 sg13g2_dfrbp_1 _7098_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net133),
    .D(_0201_),
    .Q_N(_3332_),
    .Q(\i_display.i_vga.timing_ver.counter[1] ));
 sg13g2_dfrbp_1 _7099_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net131),
    .D(_0202_),
    .Q_N(_3331_),
    .Q(\i_display.i_vga.timing_ver.counter[2] ));
 sg13g2_dfrbp_1 _7100_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net129),
    .D(_0203_),
    .Q_N(_3330_),
    .Q(\i_display.i_vga.timing_ver.counter[3] ));
 sg13g2_dfrbp_1 _7101_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net127),
    .D(_0204_),
    .Q_N(_3329_),
    .Q(\i_display.i_vga.timing_ver.counter[4] ));
 sg13g2_dfrbp_1 _7102_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net125),
    .D(_0205_),
    .Q_N(_3328_),
    .Q(\i_display.i_vga.timing_ver.counter[5] ));
 sg13g2_dfrbp_1 _7103_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net123),
    .D(_0206_),
    .Q_N(_3327_),
    .Q(\i_display.i_vga.timing_ver.counter[6] ));
 sg13g2_dfrbp_1 _7104_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net121),
    .D(_0207_),
    .Q_N(_3326_),
    .Q(\i_display.i_vga.timing_ver.counter[7] ));
 sg13g2_dfrbp_1 _7105_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net119),
    .D(_0208_),
    .Q_N(_3325_),
    .Q(\i_display.i_vga.timing_ver.counter[8] ));
 sg13g2_dfrbp_1 _7106_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net117),
    .D(_0209_),
    .Q_N(_3324_),
    .Q(\i_display.i_vga.timing_ver.counter[9] ));
 sg13g2_dfrbp_1 _7107_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net115),
    .D(_0210_),
    .Q_N(_0034_),
    .Q(\i_display.i_vga.timing_ver.counter[10] ));
 sg13g2_dfrbp_1 _7108_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net113),
    .D(net242),
    .Q_N(_0079_),
    .Q(\i_display.frame[0] ));
 sg13g2_dfrbp_1 _7109_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net111),
    .D(_0212_),
    .Q_N(_0077_),
    .Q(\i_display.frame[1] ));
 sg13g2_dfrbp_1 _7110_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net100),
    .D(_0213_),
    .Q_N(_0081_),
    .Q(\i_display.frame[2] ));
 sg13g2_dfrbp_1 _7111_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net73),
    .D(_0214_),
    .Q_N(_0075_),
    .Q(\i_display.frame[3] ));
 sg13g2_dfrbp_1 _7112_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net183),
    .D(_0215_),
    .Q_N(_0074_),
    .Q(\i_display.frame[4] ));
 sg13g2_dfrbp_1 _7113_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net179),
    .D(_0216_),
    .Q_N(_0069_),
    .Q(\i_display.frame[5] ));
 sg13g2_dfrbp_1 _7114_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net175),
    .D(net350),
    .Q_N(_0089_),
    .Q(\i_display.frame[6] ));
 sg13g2_dfrbp_1 _7115_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net159),
    .D(_0218_),
    .Q_N(_0092_),
    .Q(\i_display.frame[7] ));
 sg13g2_dfrbp_1 _7116_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net134),
    .D(net338),
    .Q_N(_0095_),
    .Q(\i_display.frame[8] ));
 sg13g2_dfrbp_1 _7117_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net130),
    .D(net318),
    .Q_N(_0028_),
    .Q(\i_display.frame[9] ));
 sg13g2_dfrbp_1 _7118_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net126),
    .D(_0221_),
    .Q_N(_3323_),
    .Q(\i_display.colour[0] ));
 sg13g2_dfrbp_1 _7119_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net124),
    .D(net282),
    .Q_N(_3322_),
    .Q(\i_display.colour[1] ));
 sg13g2_dfrbp_1 _7120_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net122),
    .D(_0223_),
    .Q_N(_3321_),
    .Q(\i_display.colour[2] ));
 sg13g2_dfrbp_1 _7121_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net120),
    .D(_0224_),
    .Q_N(_3320_),
    .Q(\i_display.colour[3] ));
 sg13g2_dfrbp_1 _7122_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net118),
    .D(_0225_),
    .Q_N(_3319_),
    .Q(\i_display.colour[4] ));
 sg13g2_dfrbp_1 _7123_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net116),
    .D(_0226_),
    .Q_N(_3318_),
    .Q(\i_display.colour[5] ));
 sg13g2_dfrbp_1 _7124_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net114),
    .D(_0227_),
    .Q_N(_0088_),
    .Q(\i_display.x_idx[2] ));
 sg13g2_dfrbp_1 _7125_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net110),
    .D(_0228_),
    .Q_N(_0087_),
    .Q(\i_display.x_idx[3] ));
 sg13g2_dfrbp_1 _7126_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net71),
    .D(_0229_),
    .Q_N(_0086_),
    .Q(\i_display.x_idx[4] ));
 sg13g2_dfrbp_1 _7127_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net177),
    .D(_0230_),
    .Q_N(_0085_),
    .Q(\i_display.x_idx[5] ));
 sg13g2_dfrbp_1 _7128_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net136),
    .D(_0231_),
    .Q_N(_0084_),
    .Q(\i_display.x_idx[6] ));
 sg13g2_dfrbp_1 _7129_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net128),
    .D(_0232_),
    .Q_N(_0083_),
    .Q(\i_display.x_idx[7] ));
 sg13g2_dfrbp_1 _7130_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net75),
    .D(_0233_),
    .Q_N(_0071_),
    .Q(\i_display.x_idx[8] ));
 sg13g2_dfrbp_1 _7131_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net173),
    .D(net298),
    .Q_N(_0096_),
    .Q(\i_display.x_idx[0] ));
 sg13g2_dfrbp_1 _7132_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net112),
    .D(_0235_),
    .Q_N(_3317_),
    .Q(\i_display.x_idx[1] ));
 sg13g2_dfrbp_1 _7133_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net132),
    .D(net327),
    .Q_N(_0026_),
    .Q(\i_display.in_line ));
 sg13g2_tiehi _6887__24 (.L_HI(net24));
 sg13g2_tiehi _6879__25 (.L_HI(net25));
 sg13g2_tiehi _6880__26 (.L_HI(net26));
 sg13g2_tiehi _6881__27 (.L_HI(net27));
 sg13g2_tiehi _6882__28 (.L_HI(net28));
 sg13g2_tiehi _6883__29 (.L_HI(net29));
 sg13g2_tiehi _6884__30 (.L_HI(net30));
 sg13g2_tiehi _6885__31 (.L_HI(net31));
 sg13g2_tiehi _7034__32 (.L_HI(net32));
 sg13g2_tiehi _7033__33 (.L_HI(net33));
 sg13g2_tiehi _7032__34 (.L_HI(net34));
 sg13g2_tiehi _7031__35 (.L_HI(net35));
 sg13g2_tiehi _7030__36 (.L_HI(net36));
 sg13g2_tiehi _7029__37 (.L_HI(net37));
 sg13g2_tiehi _7028__38 (.L_HI(net38));
 sg13g2_tiehi _7027__39 (.L_HI(net39));
 sg13g2_tiehi _7026__40 (.L_HI(net40));
 sg13g2_tiehi _7025__41 (.L_HI(net41));
 sg13g2_tiehi _7024__42 (.L_HI(net42));
 sg13g2_tiehi _7023__43 (.L_HI(net43));
 sg13g2_tiehi _6949__44 (.L_HI(net44));
 sg13g2_tiehi _6930__45 (.L_HI(net45));
 sg13g2_tiehi _6929__46 (.L_HI(net46));
 sg13g2_tiehi _6928__47 (.L_HI(net47));
 sg13g2_tiehi _6927__48 (.L_HI(net48));
 sg13g2_tiehi _6926__49 (.L_HI(net49));
 sg13g2_tiehi _6886__50 (.L_HI(net50));
 sg13g2_tiehi _6905__51 (.L_HI(net51));
 sg13g2_tiehi _6906__52 (.L_HI(net52));
 sg13g2_tiehi _6907__53 (.L_HI(net53));
 sg13g2_tiehi _6908__54 (.L_HI(net54));
 sg13g2_tiehi _6909__55 (.L_HI(net55));
 sg13g2_tiehi _6910__56 (.L_HI(net56));
 sg13g2_tiehi _6911__57 (.L_HI(net57));
 sg13g2_tiehi _6912__58 (.L_HI(net58));
 sg13g2_tiehi _6913__59 (.L_HI(net59));
 sg13g2_tiehi _6925__60 (.L_HI(net60));
 sg13g2_tiehi _6924__61 (.L_HI(net61));
 sg13g2_tiehi _6923__62 (.L_HI(net62));
 sg13g2_tiehi _6922__63 (.L_HI(net63));
 sg13g2_tiehi _6921__64 (.L_HI(net64));
 sg13g2_tiehi _6920__65 (.L_HI(net65));
 sg13g2_tiehi _6919__66 (.L_HI(net66));
 sg13g2_tiehi _6918__67 (.L_HI(net67));
 sg13g2_tiehi _6917__68 (.L_HI(net68));
 sg13g2_tiehi _6916__69 (.L_HI(net69));
 sg13g2_tiehi _6915__70 (.L_HI(net70));
 sg13g2_tiehi _7126__71 (.L_HI(net71));
 sg13g2_tiehi _6904__72 (.L_HI(net72));
 sg13g2_tiehi _7111__73 (.L_HI(net73));
 sg13g2_tiehi _6903__74 (.L_HI(net74));
 sg13g2_tiehi _7130__75 (.L_HI(net75));
 sg13g2_tiehi _6914__76 (.L_HI(net76));
 sg13g2_tiehi _6931__77 (.L_HI(net77));
 sg13g2_tiehi _6932__78 (.L_HI(net78));
 sg13g2_tiehi _6933__79 (.L_HI(net79));
 sg13g2_tiehi _6934__80 (.L_HI(net80));
 sg13g2_tiehi _6935__81 (.L_HI(net81));
 sg13g2_tiehi _6936__82 (.L_HI(net82));
 sg13g2_tiehi _6937__83 (.L_HI(net83));
 sg13g2_tiehi _6938__84 (.L_HI(net84));
 sg13g2_tiehi _6939__85 (.L_HI(net85));
 sg13g2_tiehi _6940__86 (.L_HI(net86));
 sg13g2_tiehi _6941__87 (.L_HI(net87));
 sg13g2_tiehi _6942__88 (.L_HI(net88));
 sg13g2_tiehi _6943__89 (.L_HI(net89));
 sg13g2_tiehi _6944__90 (.L_HI(net90));
 sg13g2_tiehi _6945__91 (.L_HI(net91));
 sg13g2_tiehi _6946__92 (.L_HI(net92));
 sg13g2_tiehi _6947__93 (.L_HI(net93));
 sg13g2_tiehi _6902__94 (.L_HI(net94));
 sg13g2_tiehi _6901__95 (.L_HI(net95));
 sg13g2_tiehi _6900__96 (.L_HI(net96));
 sg13g2_tiehi _6899__97 (.L_HI(net97));
 sg13g2_tiehi _6898__98 (.L_HI(net98));
 sg13g2_tiehi _6897__99 (.L_HI(net99));
 sg13g2_tiehi _7110__100 (.L_HI(net100));
 sg13g2_tiehi _6896__101 (.L_HI(net101));
 sg13g2_tiehi _6895__102 (.L_HI(net102));
 sg13g2_tiehi _6894__103 (.L_HI(net103));
 sg13g2_tiehi _6893__104 (.L_HI(net104));
 sg13g2_tiehi _6892__105 (.L_HI(net105));
 sg13g2_tiehi _6891__106 (.L_HI(net106));
 sg13g2_tiehi _6890__107 (.L_HI(net107));
 sg13g2_tiehi _6889__108 (.L_HI(net108));
 sg13g2_tiehi _6888__109 (.L_HI(net109));
 sg13g2_tiehi _7125__110 (.L_HI(net110));
 sg13g2_tiehi _7109__111 (.L_HI(net111));
 sg13g2_tiehi _7132__112 (.L_HI(net112));
 sg13g2_tiehi _7108__113 (.L_HI(net113));
 sg13g2_tiehi _7124__114 (.L_HI(net114));
 sg13g2_tiehi _7107__115 (.L_HI(net115));
 sg13g2_tiehi _7123__116 (.L_HI(net116));
 sg13g2_tiehi _7106__117 (.L_HI(net117));
 sg13g2_tiehi _7122__118 (.L_HI(net118));
 sg13g2_tiehi _7105__119 (.L_HI(net119));
 sg13g2_tiehi _7121__120 (.L_HI(net120));
 sg13g2_tiehi _7104__121 (.L_HI(net121));
 sg13g2_tiehi _7120__122 (.L_HI(net122));
 sg13g2_tiehi _7103__123 (.L_HI(net123));
 sg13g2_tiehi _7119__124 (.L_HI(net124));
 sg13g2_tiehi _7102__125 (.L_HI(net125));
 sg13g2_tiehi _7118__126 (.L_HI(net126));
 sg13g2_tiehi _7101__127 (.L_HI(net127));
 sg13g2_tiehi _7129__128 (.L_HI(net128));
 sg13g2_tiehi _7100__129 (.L_HI(net129));
 sg13g2_tiehi _7117__130 (.L_HI(net130));
 sg13g2_tiehi _7099__131 (.L_HI(net131));
 sg13g2_tiehi _7133__132 (.L_HI(net132));
 sg13g2_tiehi _7098__133 (.L_HI(net133));
 sg13g2_tiehi _7116__134 (.L_HI(net134));
 sg13g2_tiehi _7097__135 (.L_HI(net135));
 sg13g2_tiehi _7128__136 (.L_HI(net136));
 sg13g2_tiehi _7096__137 (.L_HI(net137));
 sg13g2_tiehi _7091__138 (.L_HI(net138));
 sg13g2_tiehi _7090__139 (.L_HI(net139));
 sg13g2_tiehi _7089__140 (.L_HI(net140));
 sg13g2_tiehi _7088__141 (.L_HI(net141));
 sg13g2_tiehi _6948__142 (.L_HI(net142));
 sg13g2_tiehi _7070__143 (.L_HI(net143));
 sg13g2_tiehi _7071__144 (.L_HI(net144));
 sg13g2_tiehi _7072__145 (.L_HI(net145));
 sg13g2_tiehi _7073__146 (.L_HI(net146));
 sg13g2_tiehi _7087__147 (.L_HI(net147));
 sg13g2_tiehi _7086__148 (.L_HI(net148));
 sg13g2_tiehi _7085__149 (.L_HI(net149));
 sg13g2_tiehi _7084__150 (.L_HI(net150));
 sg13g2_tiehi _7083__151 (.L_HI(net151));
 sg13g2_tiehi _7082__152 (.L_HI(net152));
 sg13g2_tiehi _7081__153 (.L_HI(net153));
 sg13g2_tiehi _7080__154 (.L_HI(net154));
 sg13g2_tiehi _7079__155 (.L_HI(net155));
 sg13g2_tiehi _7078__156 (.L_HI(net156));
 sg13g2_tiehi _7077__157 (.L_HI(net157));
 sg13g2_tiehi _7076__158 (.L_HI(net158));
 sg13g2_tiehi _7115__159 (.L_HI(net159));
 sg13g2_tiehi _7075__160 (.L_HI(net160));
 sg13g2_tiehi _7069__161 (.L_HI(net161));
 sg13g2_tiehi _7068__162 (.L_HI(net162));
 sg13g2_tiehi _7067__163 (.L_HI(net163));
 sg13g2_tiehi _7074__164 (.L_HI(net164));
 sg13g2_tiehi _7092__165 (.L_HI(net165));
 sg13g2_tiehi _7093__166 (.L_HI(net166));
 sg13g2_tiehi _7094__167 (.L_HI(net167));
 sg13g2_tiehi _7066__168 (.L_HI(net168));
 sg13g2_tiehi _7065__169 (.L_HI(net169));
 sg13g2_tiehi _7064__170 (.L_HI(net170));
 sg13g2_tiehi _7063__171 (.L_HI(net171));
 sg13g2_tiehi _7062__172 (.L_HI(net172));
 sg13g2_tiehi _7131__173 (.L_HI(net173));
 sg13g2_tiehi _7061__174 (.L_HI(net174));
 sg13g2_tiehi _7114__175 (.L_HI(net175));
 sg13g2_tiehi _7060__176 (.L_HI(net176));
 sg13g2_tiehi _7127__177 (.L_HI(net177));
 sg13g2_tiehi _7059__178 (.L_HI(net178));
 sg13g2_tiehi _7113__179 (.L_HI(net179));
 sg13g2_tiehi _7058__180 (.L_HI(net180));
 sg13g2_tiehi _7095__181 (.L_HI(net181));
 sg13g2_tiehi _7057__182 (.L_HI(net182));
 sg13g2_tiehi _7112__183 (.L_HI(net183));
 sg13g2_tiehi _7056__184 (.L_HI(net184));
 sg13g2_tiehi _7055__185 (.L_HI(net185));
 sg13g2_tiehi _7054__186 (.L_HI(net186));
 sg13g2_tiehi _7053__187 (.L_HI(net187));
 sg13g2_tiehi _7052__188 (.L_HI(net188));
 sg13g2_tiehi _7051__189 (.L_HI(net189));
 sg13g2_tiehi _7050__190 (.L_HI(net190));
 sg13g2_tiehi _7049__191 (.L_HI(net191));
 sg13g2_tiehi _7048__192 (.L_HI(net192));
 sg13g2_tiehi _7047__193 (.L_HI(net193));
 sg13g2_tiehi _7046__194 (.L_HI(net194));
 sg13g2_tiehi _7045__195 (.L_HI(net195));
 sg13g2_tiehi _7044__196 (.L_HI(net196));
 sg13g2_tiehi _7043__197 (.L_HI(net197));
 sg13g2_tiehi _7042__198 (.L_HI(net198));
 sg13g2_tiehi _7041__199 (.L_HI(net199));
 sg13g2_tiehi _7040__200 (.L_HI(net200));
 sg13g2_tiehi _7039__201 (.L_HI(net201));
 sg13g2_tiehi _7038__202 (.L_HI(net202));
 sg13g2_tiehi _7037__203 (.L_HI(net203));
 sg13g2_tiehi _7036__204 (.L_HI(net204));
 sg13g2_tiehi tt_um_MichaelBell_canon_205 (.L_HI(net205));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_tielo tt_um_MichaelBell_canon_10 (.L_LO(net10));
 sg13g2_tielo tt_um_MichaelBell_canon_11 (.L_LO(net11));
 sg13g2_tielo tt_um_MichaelBell_canon_12 (.L_LO(net12));
 sg13g2_tielo tt_um_MichaelBell_canon_13 (.L_LO(net13));
 sg13g2_tielo tt_um_MichaelBell_canon_14 (.L_LO(net14));
 sg13g2_tielo tt_um_MichaelBell_canon_15 (.L_LO(net15));
 sg13g2_tielo tt_um_MichaelBell_canon_16 (.L_LO(net16));
 sg13g2_tielo tt_um_MichaelBell_canon_17 (.L_LO(net17));
 sg13g2_tielo tt_um_MichaelBell_canon_18 (.L_LO(net18));
 sg13g2_tielo tt_um_MichaelBell_canon_19 (.L_LO(net19));
 sg13g2_tielo tt_um_MichaelBell_canon_20 (.L_LO(net20));
 sg13g2_tielo tt_um_MichaelBell_canon_21 (.L_LO(net21));
 sg13g2_tielo tt_um_MichaelBell_canon_22 (.L_LO(net22));
 sg13g2_tiehi _7035__23 (.L_HI(net23));
 sg13g2_buf_2 _7331_ (.A(\i_music.i_pwm.pwm ),
    .X(uio_out[7]));
 sg13g2_buf_1 _7332_ (.A(\i_display.i_vga.timing_ver.sync ),
    .X(uo_out[3]));
 sg13g2_buf_2 _7333_ (.A(\i_display.hsync ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout884 (.A(_0865_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_0849_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_0830_),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(net888),
    .X(net887));
 sg13g2_buf_1 fanout888 (.A(_0873_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(_0864_),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(net891),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_0860_),
    .X(net891));
 sg13g2_buf_4 fanout892 (.X(net892),
    .A(_0859_));
 sg13g2_buf_2 fanout893 (.A(net894),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_0848_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_0846_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(net898),
    .X(net896));
 sg13g2_buf_1 fanout897 (.A(net898),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_0828_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(_0803_),
    .X(net899));
 sg13g2_buf_4 fanout900 (.X(net900),
    .A(_1628_));
 sg13g2_buf_2 fanout901 (.A(_1599_),
    .X(net901));
 sg13g2_buf_4 fanout902 (.X(net902),
    .A(_1608_));
 sg13g2_buf_4 fanout903 (.X(net903),
    .A(_1607_));
 sg13g2_buf_2 fanout904 (.A(net905),
    .X(net904));
 sg13g2_buf_1 fanout905 (.A(net908),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(net907),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(net908),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(_1596_),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(net910),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(_1595_),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(net912),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_1595_),
    .X(net912));
 sg13g2_buf_4 fanout913 (.X(net913),
    .A(net915));
 sg13g2_buf_4 fanout914 (.X(net914),
    .A(_1592_));
 sg13g2_buf_2 fanout915 (.A(_1592_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(net918),
    .X(net916));
 sg13g2_buf_4 fanout917 (.X(net917),
    .A(net918));
 sg13g2_buf_1 fanout918 (.A(_1591_),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(net920),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_1591_),
    .X(net920));
 sg13g2_buf_4 fanout921 (.X(net921),
    .A(_1587_));
 sg13g2_buf_2 fanout922 (.A(_1587_),
    .X(net922));
 sg13g2_buf_4 fanout923 (.X(net923),
    .A(_1586_));
 sg13g2_buf_4 fanout924 (.X(net924),
    .A(_1586_));
 sg13g2_buf_4 fanout925 (.X(net925),
    .A(_1584_));
 sg13g2_buf_4 fanout926 (.X(net926),
    .A(_1583_));
 sg13g2_buf_2 fanout927 (.A(_1579_),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(_1579_),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(_1578_),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(_1578_),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(net932),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(_1575_),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(_2735_),
    .X(net933));
 sg13g2_buf_4 fanout934 (.X(net934),
    .A(_2079_));
 sg13g2_buf_4 fanout935 (.X(net935),
    .A(_2069_));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(_2044_));
 sg13g2_buf_2 fanout937 (.A(_2968_),
    .X(net937));
 sg13g2_buf_4 fanout938 (.X(net938),
    .A(_2967_));
 sg13g2_buf_2 fanout939 (.A(_2967_),
    .X(net939));
 sg13g2_buf_4 fanout940 (.X(net940),
    .A(_2966_));
 sg13g2_buf_4 fanout941 (.X(net941),
    .A(net943));
 sg13g2_buf_2 fanout942 (.A(net943),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(\i_music.i_sample.t1.genblk1[0].state.Q ),
    .X(net943));
 sg13g2_buf_4 fanout944 (.X(net944),
    .A(net946));
 sg13g2_buf_2 fanout945 (.A(net946),
    .X(net945));
 sg13g2_buf_4 fanout946 (.X(net946),
    .A(net948));
 sg13g2_buf_2 fanout947 (.A(net948),
    .X(net947));
 sg13g2_buf_1 fanout948 (.A(\i_music.i_sample.t1.genblk1[1].state.Q ),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(net950),
    .X(net949));
 sg13g2_buf_4 fanout950 (.X(net950),
    .A(net952));
 sg13g2_buf_1 fanout951 (.A(net952),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(\i_music.i_sample.t1.genblk1[2].state.Q ),
    .X(net952));
 sg13g2_buf_4 fanout953 (.X(net953),
    .A(net954));
 sg13g2_buf_4 fanout954 (.X(net954),
    .A(net957));
 sg13g2_buf_2 fanout955 (.A(net957),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(net957),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(net958),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(\i_music.i_sample.t1.genblk1[3].state.Q ),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(net961),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(net961),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(net965),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(net964),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(net964),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(net965),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(\i_music.i_sample.t1.genblk1[4].state.Q ),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(net970),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(net970),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(net970),
    .X(net968));
 sg13g2_buf_1 fanout969 (.A(net970),
    .X(net969));
 sg13g2_buf_1 fanout970 (.A(\i_music.i_sample.t1.genblk1[5].state.Q ),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(net972),
    .X(net971));
 sg13g2_buf_4 fanout972 (.X(net972),
    .A(net973));
 sg13g2_buf_2 fanout973 (.A(net974),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(\i_music.i_sample.t1.genblk1[6].state.Q ),
    .X(net974));
 sg13g2_buf_4 fanout975 (.X(net975),
    .A(net976));
 sg13g2_buf_2 fanout976 (.A(\i_music.i_sample.t1.genblk1[7].state.Q ),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_2002_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_1535_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_1535_),
    .X(net979));
 sg13g2_buf_4 fanout980 (.X(net980),
    .A(_2722_));
 sg13g2_buf_2 fanout981 (.A(_1995_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(net983),
    .X(net982));
 sg13g2_buf_4 fanout983 (.X(net983),
    .A(_1368_));
 sg13g2_buf_4 fanout984 (.X(net984),
    .A(_2724_));
 sg13g2_buf_2 fanout985 (.A(_1170_),
    .X(net985));
 sg13g2_buf_1 fanout986 (.A(_1170_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_1108_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(net989),
    .X(net988));
 sg13g2_buf_1 fanout989 (.A(_2456_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_2650_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(_2658_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_3266_),
    .X(net992));
 sg13g2_buf_4 fanout993 (.X(net993),
    .A(_3231_));
 sg13g2_buf_2 fanout994 (.A(_2367_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(net996),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_3241_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(net998),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_3238_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_3214_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_3178_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_3091_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_3139_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_3090_),
    .X(net1003));
 sg13g2_buf_1 fanout1004 (.A(_3090_),
    .X(net1004));
 sg13g2_buf_4 fanout1005 (.X(net1005),
    .A(_3089_));
 sg13g2_buf_4 fanout1006 (.X(net1006),
    .A(_1083_));
 sg13g2_buf_4 fanout1007 (.X(net1007),
    .A(_1071_));
 sg13g2_buf_2 fanout1008 (.A(net1011),
    .X(net1008));
 sg13g2_buf_1 fanout1009 (.A(net1011),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(net1011),
    .X(net1010));
 sg13g2_buf_1 fanout1011 (.A(_1012_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(net1013),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(net1015),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(net1015),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_1001_),
    .X(net1015));
 sg13g2_buf_4 fanout1016 (.X(net1016),
    .A(net1017));
 sg13g2_buf_2 fanout1017 (.A(_0991_),
    .X(net1017));
 sg13g2_buf_4 fanout1018 (.X(net1018),
    .A(_0987_));
 sg13g2_buf_2 fanout1019 (.A(net1020),
    .X(net1019));
 sg13g2_buf_1 fanout1020 (.A(net1022),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_4 fanout1022 (.X(net1022),
    .A(_3099_));
 sg13g2_buf_2 fanout1023 (.A(net1024),
    .X(net1023));
 sg13g2_buf_4 fanout1024 (.X(net1024),
    .A(_3099_));
 sg13g2_buf_2 fanout1025 (.A(_3099_),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(net1027),
    .X(net1026));
 sg13g2_buf_4 fanout1027 (.X(net1027),
    .A(_3098_));
 sg13g2_buf_2 fanout1028 (.A(_2428_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_2428_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(net1031),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_1916_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(net1033),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(net1034),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(net1036),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(net1036),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_1021_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(net1039),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(net1041),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(net1041),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_1014_),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(net1043),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(net1045),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(_1011_),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(_1011_),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(net1047),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_1011_),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(net1049),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(net1050),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(net1051),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(_1000_),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(net1055),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(net1055),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(net1055),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_0997_),
    .X(net1055));
 sg13g2_buf_4 fanout1056 (.X(net1056),
    .A(_0990_));
 sg13g2_buf_2 fanout1057 (.A(_0779_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(net1059),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_0777_),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_3141_),
    .X(net1060));
 sg13g2_buf_4 fanout1061 (.X(net1061),
    .A(_3128_));
 sg13g2_buf_2 fanout1062 (.A(_3101_),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(net1065),
    .X(net1063));
 sg13g2_buf_1 fanout1064 (.A(net1065),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(net1066),
    .X(net1065));
 sg13g2_buf_4 fanout1066 (.X(net1066),
    .A(_3056_));
 sg13g2_buf_4 fanout1067 (.X(net1067),
    .A(net1069));
 sg13g2_buf_4 fanout1068 (.X(net1068),
    .A(_3036_));
 sg13g2_buf_1 fanout1069 (.A(_3036_),
    .X(net1069));
 sg13g2_buf_4 fanout1070 (.X(net1070),
    .A(net1073));
 sg13g2_buf_1 fanout1071 (.A(net1073),
    .X(net1071));
 sg13g2_buf_4 fanout1072 (.X(net1072),
    .A(net1073));
 sg13g2_buf_2 fanout1073 (.A(net1074),
    .X(net1073));
 sg13g2_buf_4 fanout1074 (.X(net1074),
    .A(_3035_));
 sg13g2_buf_2 fanout1075 (.A(net1076),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(net1077),
    .X(net1076));
 sg13g2_buf_1 fanout1077 (.A(net1078),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(net1079),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(_3033_),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(net1081),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(_3032_),
    .X(net1081));
 sg13g2_buf_4 fanout1082 (.X(net1082),
    .A(net1083));
 sg13g2_buf_4 fanout1083 (.X(net1083),
    .A(_3008_));
 sg13g2_buf_2 fanout1084 (.A(net1085),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(net1086),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(net1089),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(net1088),
    .X(net1087));
 sg13g2_buf_4 fanout1088 (.X(net1088),
    .A(net1089));
 sg13g2_buf_4 fanout1089 (.X(net1089),
    .A(_2995_));
 sg13g2_buf_4 fanout1090 (.X(net1090),
    .A(_2912_));
 sg13g2_buf_2 fanout1091 (.A(\i_display.in_line ),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(net1095),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(net1095),
    .X(net1093));
 sg13g2_buf_1 fanout1094 (.A(net1095),
    .X(net1094));
 sg13g2_buf_1 fanout1095 (.A(\i_display.x_idx[1] ),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(\i_display.x_idx[0] ),
    .X(net1096));
 sg13g2_buf_4 fanout1097 (.X(net1097),
    .A(net1098));
 sg13g2_buf_2 fanout1098 (.A(net345),
    .X(net1098));
 sg13g2_buf_4 fanout1099 (.X(net1099),
    .A(net359));
 sg13g2_buf_2 fanout1100 (.A(\i_display.x_idx[6] ),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(net1103),
    .X(net1101));
 sg13g2_buf_1 fanout1102 (.A(net1103),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(net1106),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(net1105),
    .X(net1104));
 sg13g2_buf_1 fanout1105 (.A(net1106),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(net355),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(net1108),
    .X(net1107));
 sg13g2_buf_1 fanout1108 (.A(net1109),
    .X(net1108));
 sg13g2_buf_4 fanout1109 (.X(net1109),
    .A(\i_display.x_idx[4] ));
 sg13g2_buf_2 fanout1110 (.A(net1111),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(\i_display.x_idx[4] ),
    .X(net1111));
 sg13g2_buf_4 fanout1112 (.X(net1112),
    .A(\i_display.x_idx[3] ));
 sg13g2_buf_4 fanout1113 (.X(net1113),
    .A(\i_display.x_idx[3] ));
 sg13g2_buf_4 fanout1114 (.X(net1114),
    .A(net1115));
 sg13g2_buf_2 fanout1115 (.A(net356),
    .X(net1115));
 sg13g2_buf_4 fanout1116 (.X(net1116),
    .A(net361));
 sg13g2_buf_2 fanout1117 (.A(\i_display.frame[6] ),
    .X(net1117));
 sg13g2_buf_1 fanout1118 (.A(\i_display.frame[6] ),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(net358),
    .X(net1119));
 sg13g2_buf_2 fanout1120 (.A(\i_display.frame[5] ),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(net1122),
    .X(net1121));
 sg13g2_buf_4 fanout1122 (.X(net1122),
    .A(\i_display.frame[4] ));
 sg13g2_buf_2 fanout1123 (.A(\i_display.frame[3] ),
    .X(net1123));
 sg13g2_buf_2 fanout1124 (.A(net339),
    .X(net1124));
 sg13g2_buf_2 fanout1125 (.A(net1126),
    .X(net1125));
 sg13g2_buf_2 fanout1126 (.A(net364),
    .X(net1126));
 sg13g2_buf_2 fanout1127 (.A(net1128),
    .X(net1127));
 sg13g2_buf_2 fanout1128 (.A(net365),
    .X(net1128));
 sg13g2_buf_4 fanout1129 (.X(net1129),
    .A(net241));
 sg13g2_buf_2 fanout1130 (.A(\i_display.i_vga.timing_ver.counter[1] ),
    .X(net1130));
 sg13g2_buf_2 fanout1131 (.A(net1132),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(\i_display.i_vga.vblank ),
    .X(net1132));
 sg13g2_buf_2 fanout1133 (.A(net1134),
    .X(net1133));
 sg13g2_buf_2 fanout1134 (.A(net354),
    .X(net1134));
 sg13g2_buf_2 fanout1135 (.A(\i_display.frame_crotchet[4] ),
    .X(net1135));
 sg13g2_buf_4 fanout1136 (.X(net1136),
    .A(net1137));
 sg13g2_buf_2 fanout1137 (.A(net352),
    .X(net1137));
 sg13g2_buf_2 fanout1138 (.A(net1140),
    .X(net1138));
 sg13g2_buf_2 fanout1139 (.A(net1140),
    .X(net1139));
 sg13g2_buf_2 fanout1140 (.A(\i_display.frame_crotchet[2] ),
    .X(net1140));
 sg13g2_buf_2 fanout1141 (.A(net1142),
    .X(net1141));
 sg13g2_buf_2 fanout1142 (.A(\i_display.i_vga.low_count[7] ),
    .X(net1142));
 sg13g2_buf_4 fanout1143 (.X(net1143),
    .A(net1145));
 sg13g2_buf_2 fanout1144 (.A(net1145),
    .X(net1144));
 sg13g2_buf_4 fanout1145 (.X(net1145),
    .A(net1147));
 sg13g2_buf_4 fanout1146 (.X(net1146),
    .A(net1147));
 sg13g2_buf_2 fanout1147 (.A(net1149),
    .X(net1147));
 sg13g2_buf_4 fanout1148 (.X(net1148),
    .A(net1149));
 sg13g2_buf_2 fanout1149 (.A(\i_display.i_vga.low_count[1] ),
    .X(net1149));
 sg13g2_buf_4 fanout1150 (.X(net1150),
    .A(net1152));
 sg13g2_buf_2 fanout1151 (.A(net1152),
    .X(net1151));
 sg13g2_buf_2 fanout1152 (.A(net1154),
    .X(net1152));
 sg13g2_buf_4 fanout1153 (.X(net1153),
    .A(net1154));
 sg13g2_buf_2 fanout1154 (.A(net380),
    .X(net1154));
 sg13g2_buf_4 fanout1155 (.X(net1155),
    .A(net1158));
 sg13g2_buf_2 fanout1156 (.A(net1157),
    .X(net1156));
 sg13g2_buf_2 fanout1157 (.A(net1158),
    .X(net1157));
 sg13g2_buf_4 fanout1158 (.X(net1158),
    .A(_2923_));
 sg13g2_buf_4 fanout1159 (.X(net1159),
    .A(net1163));
 sg13g2_buf_2 fanout1160 (.A(net1161),
    .X(net1160));
 sg13g2_buf_2 fanout1161 (.A(net1162),
    .X(net1161));
 sg13g2_buf_2 fanout1162 (.A(net1163),
    .X(net1162));
 sg13g2_buf_4 fanout1163 (.X(net1163),
    .A(_2923_));
 sg13g2_buf_2 fanout1164 (.A(net1166),
    .X(net1164));
 sg13g2_buf_1 fanout1165 (.A(net1166),
    .X(net1165));
 sg13g2_buf_4 fanout1166 (.X(net1166),
    .A(net1175));
 sg13g2_buf_2 fanout1167 (.A(net1168),
    .X(net1167));
 sg13g2_buf_2 fanout1168 (.A(net1175),
    .X(net1168));
 sg13g2_buf_2 fanout1169 (.A(net1170),
    .X(net1169));
 sg13g2_buf_2 fanout1170 (.A(net1171),
    .X(net1170));
 sg13g2_buf_4 fanout1171 (.X(net1171),
    .A(net1175));
 sg13g2_buf_4 fanout1172 (.X(net1172),
    .A(net1173));
 sg13g2_buf_2 fanout1173 (.A(net1175),
    .X(net1173));
 sg13g2_buf_4 fanout1174 (.X(net1174),
    .A(net1175));
 sg13g2_buf_4 fanout1175 (.X(net1175),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[1]));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_MichaelBell_canon_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_5_13__leaf_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_5_15__leaf_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_5_19__leaf_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_5_23__leaf_clk_regs));
 sg13g2_inv_1 clkload7 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_inv_1 clkload8 (.A(clknet_5_29__leaf_clk_regs));
 sg13g2_inv_1 clkload9 (.A(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_0__1501_ (.A(_1501_),
    .X(clknet_0__1501_));
 sg13g2_buf_2 clkbuf_1_0__f__1501_ (.A(clknet_0__1501_),
    .X(clknet_1_0__leaf__1501_));
 sg13g2_buf_2 clkbuf_1_1__f__1501_ (.A(clknet_0__1501_),
    .X(clknet_1_1__leaf__1501_));
 sg13g2_buf_2 \clkbuf_0_i_music.i_sample.t4.CG.GCLK  (.A(\i_music.i_sample.t4.CG.GCLK ),
    .X(\clknet_0_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_0__f_i_music.i_sample.t4.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t4.CG.GCLK ),
    .X(\clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_1__f_i_music.i_sample.t4.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t4.CG.GCLK ),
    .X(\clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_2__f_i_music.i_sample.t4.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t4.CG.GCLK ),
    .X(\clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_3__f_i_music.i_sample.t4.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t4.CG.GCLK ),
    .X(\clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_inv_1 clkload10 (.A(\clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_inv_1 clkload11 (.A(\clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_0_i_music.i_sample.t3.CG.GCLK  (.A(\i_music.i_sample.t3.CG.GCLK ),
    .X(\clknet_0_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_0__f_i_music.i_sample.t3.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t3.CG.GCLK ),
    .X(\clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_1__f_i_music.i_sample.t3.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t3.CG.GCLK ),
    .X(\clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_2__f_i_music.i_sample.t3.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t3.CG.GCLK ),
    .X(\clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_3__f_i_music.i_sample.t3.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t3.CG.GCLK ),
    .X(\clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_inv_1 clkload12 (.A(\clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_inv_1 clkload13 (.A(\clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_0_i_music.i_sample.t2.CG.GCLK  (.A(\i_music.i_sample.t2.CG.GCLK ),
    .X(\clknet_0_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_0__f_i_music.i_sample.t2.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t2.CG.GCLK ),
    .X(\clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_1__f_i_music.i_sample.t2.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t2.CG.GCLK ),
    .X(\clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_2__f_i_music.i_sample.t2.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t2.CG.GCLK ),
    .X(\clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_3__f_i_music.i_sample.t2.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t2.CG.GCLK ),
    .X(\clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_inv_1 clkload14 (.A(\clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_inv_1 clkload15 (.A(\clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_0_i_music.i_sample.t1.CG.GCLK  (.A(\i_music.i_sample.t1.CG.GCLK ),
    .X(\clknet_0_i_music.i_sample.t1.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_0__f_i_music.i_sample.t1.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t1.CG.GCLK ),
    .X(\clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_1__f_i_music.i_sample.t1.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t1.CG.GCLK ),
    .X(\clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_2__f_i_music.i_sample.t1.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t1.CG.GCLK ),
    .X(\clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ));
 sg13g2_buf_2 \clkbuf_2_3__f_i_music.i_sample.t1.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t1.CG.GCLK ),
    .X(\clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ));
 sg13g2_inv_1 clkload16 (.A(\clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(delaynet_1_clk));
 sg13g2_buf_2 delaybuf_1_clk (.A(delaynet_1_clk),
    .X(delaynet_2_clk));
 sg13g2_buf_2 delaybuf_2_clk (.A(delaynet_2_clk),
    .X(clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0098_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0034_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold3 (.A(\i_display.i_vga.timing_ver.blank ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0097_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0045_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0143_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold7 (.A(\i_display.i_vga.timing_ver.counter[3] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold8 (.A(_3003_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold9 (.A(\i_display.i_vga.timing_ver.sync_tmp ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold10 (.A(\i_music.i_pwm.pwm ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0167_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0061_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0062_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_display.frame_crotchet[4] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold15 (.A(\i_music.violin_note_idx[3][7] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0113_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold17 (.A(\i_music.violin_note_idx[2][3] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0173_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold19 (.A(\i_display.x_idx[8] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_music.count[24] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold21 (.A(_1973_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold22 (.A(\i_music.i_pwm.count[2] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold23 (.A(_1925_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0121_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0100_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0199_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold27 (.A(\i_music.i_pwm.sample[4] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0131_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0099_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0182_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold31 (.A(\i_music.violin_note_idx[2][8] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_music.count[23] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0158_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold34 (.A(\i_display.frame_crotchet[2] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold35 (.A(\i_music.i_pwm.sample[5] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold36 (.A(\i_display.frame[0] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0211_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold38 (.A(\i_music.i_pwm.sample[7] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0134_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0046_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold41 (.A(\i_display.i_vga.hsync_tmp ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold42 (.A(\i_music.i_pwm.sample[2] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0129_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold44 (.A(\i_music.violin_note_idx[2][6] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold45 (.A(\i_music.violin_note_idx[2][1] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0171_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold47 (.A(\i_music.violin_note_idx[2][2] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0172_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold49 (.A(\i_music.i_pwm.sample[3] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0060_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold51 (.A(_1884_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold52 (.A(\i_music.i_pwm.sample[1] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold53 (.A(\i_display.frame_crotchet[0] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0174_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold55 (.A(\i_music.count[12] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold56 (.A(_1960_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold57 (.A(\i_music.violin_note_idx[1][3] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold58 (.A(_2004_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0170_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold60 (.A(\i_music.violin_note_idx[3][8] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold61 (.A(\i_music.i_pwm.count[3] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold62 (.A(_1927_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold63 (.A(\crotchet[6] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0166_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold65 (.A(\i_display.i_vga.timing_ver.counter[2] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold66 (.A(\i_music.i_pwm.sample[6] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0133_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold68 (.A(\i_music.count[13] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold69 (.A(\i_music.count[18] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold70 (.A(_1966_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold71 (.A(\i_music.violin_note_idx[2][7] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0104_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold73 (.A(\i_display.frame_crotchet[1] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold74 (.A(\i_music.violin_note_idx[1][5] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0052_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold76 (.A(_2803_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0222_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold78 (.A(\i_music.i_pwm.count[6] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold79 (.A(_1932_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold80 (.A(\i_music.i_pwm.count[5] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold81 (.A(_1930_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_music.count[11] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold83 (.A(\i_music.count[16] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold84 (.A(_1964_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold85 (.A(\i_music.i_pwm.sample[0] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0127_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold87 (.A(\i_music.i_pwm.count[4] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold88 (.A(\i_music.count[14] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold89 (.A(\i_music.violin_note_idx[1][2] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0169_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold91 (.A(\i_music.count[15] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold92 (.A(\i_display.x_idx[0] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0234_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold94 (.A(\i_music.violin_note_idx[1][6] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold95 (.A(\i_music.count[17] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold96 (.A(\i_music.i_pwm.count[0] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0120_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold98 (.A(\i_music.violin_note_idx[2][5] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_music.violin_note_idx[1][4] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0187_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold101 (.A(\i_music.violin_note_idx[3][2] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0116_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold103 (.A(\i_music.violin_note_idx[3][1] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0115_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold105 (.A(\i_display.i_vga.low_count[6] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold106 (.A(\i_music.violin_note_idx[2][4] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold107 (.A(\crotchet[5] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold108 (.A(_1978_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold109 (.A(\i_music.violin_note_idx[3][6] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold110 (.A(\i_display.i_vga.timing_ver.counter[10] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold111 (.A(_2366_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold112 (.A(\i_display.frame[9] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0220_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold114 (.A(\i_music.i_sample.sample_acc[7] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold115 (.A(\i_music.violin_note_idx[1][8] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0191_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold117 (.A(\i_music.i_pwm.count[7] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_display.i_vga.low_count[5] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold119 (.A(_1952_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold120 (.A(\i_music.violin_note_idx[3][0] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0026_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0236_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold123 (.A(\i_music.violin_note_idx[1][1] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0168_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold125 (.A(\i_display.i_vga.low_count[9] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold126 (.A(\i_display.i_vga.low_count[3] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold127 (.A(_1950_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold128 (.A(\i_music.violin_note_idx[3][3] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold129 (.A(\i_music.i_sample.sample_acc[0] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold130 (.A(\i_music.violin_note_idx[1][7] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold131 (.A(\i_music.violin_note_idx[3][4] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold132 (.A(\i_display.frame[8] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0219_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold134 (.A(\i_display.frame[3] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold135 (.A(\i_display.i_vga.timing_ver.counter[4] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0050_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold137 (.A(\crotchet[4] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold138 (.A(\i_music.violin_note_idx[3][5] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold139 (.A(\i_music.count[10] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold140 (.A(\i_display.x_idx[7] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold141 (.A(\crotchet[3] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold142 (.A(\i_music.count[22] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold143 (.A(\crotchet[4] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0089_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0217_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold146 (.A(\i_display.frame_crotchet[6] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold147 (.A(\i_display.frame_crotchet[3] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold148 (.A(\i_music.count[19] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold149 (.A(\i_display.frame_crotchet[5] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold150 (.A(\i_display.x_idx[5] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_display.x_idx[2] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0081_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold153 (.A(\i_display.frame[5] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold154 (.A(\i_display.x_idx[6] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold155 (.A(\i_music.count[20] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold156 (.A(\i_display.frame[7] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold157 (.A(\i_display.i_vga.timing_ver.counter[6] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold158 (.A(_2360_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold159 (.A(\i_display.frame[2] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold160 (.A(\i_display.frame[1] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold161 (.A(\i_display.i_vga.timing_ver.counter[0] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold162 (.A(\i_music.count[21] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold163 (.A(\i_display.i_vga.timing_ver.counter[9] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold164 (.A(_2365_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold165 (.A(\i_music.i_sample.sample_idx[6] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0054_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold167 (.A(\i_music.i_sample.sample_idx[7] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold168 (.A(\i_music.i_sample.sample_idx[2] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold169 (.A(\i_music.i_sample.sample_idx[0] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold170 (.A(\i_display.i_vga.timing_ver.counter[8] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold171 (.A(\i_music.i_sample.sample_idx[3] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold172 (.A(\i_music.i_sample.sample_idx[1] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold173 (.A(\i_display.i_vga.timing_ver.counter[5] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold174 (.A(\i_display.i_vga.timing_ver.counter[7] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold175 (.A(\i_display.i_vga.low_count[0] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold176 (.A(\i_display.frame_crotchet[6] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold177 (.A(\i_music.count[23] ),
    .X(net382));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_4 FILLER_0_14 ();
 sg13g2_fill_1 FILLER_0_18 ();
 sg13g2_fill_2 FILLER_0_24 ();
 sg13g2_fill_1 FILLER_0_26 ();
 sg13g2_fill_2 FILLER_0_32 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_fill_1 FILLER_0_81 ();
 sg13g2_decap_8 FILLER_0_87 ();
 sg13g2_decap_4 FILLER_0_94 ();
 sg13g2_fill_1 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_109 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_fill_2 FILLER_0_137 ();
 sg13g2_decap_8 FILLER_0_143 ();
 sg13g2_decap_8 FILLER_0_150 ();
 sg13g2_fill_2 FILLER_0_157 ();
 sg13g2_decap_8 FILLER_0_176 ();
 sg13g2_fill_1 FILLER_0_183 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_decap_8 FILLER_0_208 ();
 sg13g2_decap_4 FILLER_0_215 ();
 sg13g2_decap_8 FILLER_0_225 ();
 sg13g2_decap_8 FILLER_0_232 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_decap_8 FILLER_0_246 ();
 sg13g2_decap_4 FILLER_0_253 ();
 sg13g2_fill_2 FILLER_0_274 ();
 sg13g2_fill_1 FILLER_0_276 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_4 FILLER_0_322 ();
 sg13g2_fill_2 FILLER_0_330 ();
 sg13g2_fill_1 FILLER_0_332 ();
 sg13g2_fill_1 FILLER_0_337 ();
 sg13g2_fill_2 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_348 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_4 FILLER_0_369 ();
 sg13g2_fill_1 FILLER_0_381 ();
 sg13g2_fill_2 FILLER_0_403 ();
 sg13g2_fill_2 FILLER_1_0 ();
 sg13g2_fill_1 FILLER_1_2 ();
 sg13g2_fill_2 FILLER_1_22 ();
 sg13g2_fill_1 FILLER_1_24 ();
 sg13g2_fill_2 FILLER_1_58 ();
 sg13g2_fill_2 FILLER_1_121 ();
 sg13g2_decap_4 FILLER_1_149 ();
 sg13g2_fill_1 FILLER_1_153 ();
 sg13g2_fill_2 FILLER_1_159 ();
 sg13g2_fill_1 FILLER_1_184 ();
 sg13g2_fill_2 FILLER_1_206 ();
 sg13g2_fill_1 FILLER_1_208 ();
 sg13g2_fill_1 FILLER_1_273 ();
 sg13g2_fill_1 FILLER_1_317 ();
 sg13g2_fill_2 FILLER_1_336 ();
 sg13g2_fill_1 FILLER_1_338 ();
 sg13g2_fill_2 FILLER_1_344 ();
 sg13g2_fill_1 FILLER_1_346 ();
 sg13g2_fill_1 FILLER_1_392 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_fill_1 FILLER_2_0 ();
 sg13g2_decap_4 FILLER_2_29 ();
 sg13g2_fill_1 FILLER_2_41 ();
 sg13g2_fill_2 FILLER_2_67 ();
 sg13g2_fill_1 FILLER_2_69 ();
 sg13g2_decap_4 FILLER_2_104 ();
 sg13g2_fill_1 FILLER_2_154 ();
 sg13g2_fill_1 FILLER_2_160 ();
 sg13g2_fill_1 FILLER_2_208 ();
 sg13g2_fill_2 FILLER_2_311 ();
 sg13g2_fill_1 FILLER_2_313 ();
 sg13g2_fill_2 FILLER_2_321 ();
 sg13g2_fill_1 FILLER_2_323 ();
 sg13g2_fill_2 FILLER_2_329 ();
 sg13g2_fill_2 FILLER_2_361 ();
 sg13g2_fill_1 FILLER_2_363 ();
 sg13g2_fill_2 FILLER_2_385 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_fill_1 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_36 ();
 sg13g2_fill_2 FILLER_3_53 ();
 sg13g2_fill_1 FILLER_3_55 ();
 sg13g2_fill_1 FILLER_3_64 ();
 sg13g2_fill_2 FILLER_3_156 ();
 sg13g2_fill_1 FILLER_3_158 ();
 sg13g2_fill_1 FILLER_3_207 ();
 sg13g2_fill_2 FILLER_3_231 ();
 sg13g2_fill_1 FILLER_3_253 ();
 sg13g2_fill_2 FILLER_3_300 ();
 sg13g2_fill_2 FILLER_3_306 ();
 sg13g2_fill_1 FILLER_3_308 ();
 sg13g2_fill_1 FILLER_3_345 ();
 sg13g2_fill_1 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_27 ();
 sg13g2_fill_2 FILLER_4_34 ();
 sg13g2_fill_1 FILLER_4_36 ();
 sg13g2_decap_8 FILLER_4_87 ();
 sg13g2_decap_8 FILLER_4_94 ();
 sg13g2_decap_8 FILLER_4_101 ();
 sg13g2_fill_1 FILLER_4_108 ();
 sg13g2_fill_1 FILLER_4_129 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_fill_1 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_206 ();
 sg13g2_decap_4 FILLER_4_216 ();
 sg13g2_decap_8 FILLER_4_253 ();
 sg13g2_decap_8 FILLER_4_260 ();
 sg13g2_decap_8 FILLER_4_276 ();
 sg13g2_decap_8 FILLER_4_283 ();
 sg13g2_decap_8 FILLER_4_290 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_4 FILLER_4_308 ();
 sg13g2_fill_2 FILLER_4_324 ();
 sg13g2_fill_1 FILLER_4_326 ();
 sg13g2_fill_2 FILLER_4_365 ();
 sg13g2_fill_1 FILLER_4_385 ();
 sg13g2_fill_2 FILLER_4_392 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_2 ();
 sg13g2_fill_2 FILLER_5_38 ();
 sg13g2_fill_1 FILLER_5_40 ();
 sg13g2_fill_2 FILLER_5_66 ();
 sg13g2_fill_1 FILLER_5_68 ();
 sg13g2_decap_4 FILLER_5_83 ();
 sg13g2_fill_1 FILLER_5_87 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_4 FILLER_5_119 ();
 sg13g2_fill_1 FILLER_5_142 ();
 sg13g2_fill_2 FILLER_5_164 ();
 sg13g2_fill_1 FILLER_5_166 ();
 sg13g2_fill_2 FILLER_5_184 ();
 sg13g2_fill_2 FILLER_5_191 ();
 sg13g2_decap_4 FILLER_5_203 ();
 sg13g2_fill_1 FILLER_5_207 ();
 sg13g2_decap_4 FILLER_5_227 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_4 FILLER_5_287 ();
 sg13g2_fill_1 FILLER_5_291 ();
 sg13g2_decap_4 FILLER_5_315 ();
 sg13g2_fill_2 FILLER_5_324 ();
 sg13g2_fill_2 FILLER_5_336 ();
 sg13g2_fill_1 FILLER_5_338 ();
 sg13g2_fill_1 FILLER_5_361 ();
 sg13g2_fill_2 FILLER_5_384 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_29 ();
 sg13g2_fill_1 FILLER_6_35 ();
 sg13g2_fill_2 FILLER_6_52 ();
 sg13g2_fill_2 FILLER_6_71 ();
 sg13g2_fill_1 FILLER_6_73 ();
 sg13g2_fill_1 FILLER_6_82 ();
 sg13g2_fill_1 FILLER_6_183 ();
 sg13g2_fill_1 FILLER_6_201 ();
 sg13g2_fill_2 FILLER_6_238 ();
 sg13g2_fill_1 FILLER_6_240 ();
 sg13g2_fill_2 FILLER_6_280 ();
 sg13g2_decap_4 FILLER_6_321 ();
 sg13g2_fill_2 FILLER_6_325 ();
 sg13g2_fill_1 FILLER_6_332 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_30 ();
 sg13g2_fill_2 FILLER_7_40 ();
 sg13g2_fill_2 FILLER_7_47 ();
 sg13g2_fill_2 FILLER_7_74 ();
 sg13g2_fill_1 FILLER_7_116 ();
 sg13g2_fill_2 FILLER_7_168 ();
 sg13g2_fill_1 FILLER_7_187 ();
 sg13g2_fill_1 FILLER_7_226 ();
 sg13g2_fill_2 FILLER_7_251 ();
 sg13g2_fill_1 FILLER_7_284 ();
 sg13g2_fill_2 FILLER_7_290 ();
 sg13g2_fill_1 FILLER_7_292 ();
 sg13g2_fill_2 FILLER_7_322 ();
 sg13g2_fill_2 FILLER_7_329 ();
 sg13g2_fill_2 FILLER_7_336 ();
 sg13g2_fill_1 FILLER_7_343 ();
 sg13g2_fill_1 FILLER_7_387 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_19 ();
 sg13g2_fill_2 FILLER_8_37 ();
 sg13g2_fill_1 FILLER_8_44 ();
 sg13g2_fill_1 FILLER_8_55 ();
 sg13g2_fill_1 FILLER_8_61 ();
 sg13g2_fill_2 FILLER_8_93 ();
 sg13g2_decap_4 FILLER_8_99 ();
 sg13g2_fill_1 FILLER_8_103 ();
 sg13g2_fill_1 FILLER_8_155 ();
 sg13g2_fill_1 FILLER_8_297 ();
 sg13g2_fill_1 FILLER_8_320 ();
 sg13g2_fill_1 FILLER_8_334 ();
 sg13g2_fill_2 FILLER_8_377 ();
 sg13g2_fill_1 FILLER_8_379 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_112 ();
 sg13g2_fill_1 FILLER_9_123 ();
 sg13g2_decap_8 FILLER_9_136 ();
 sg13g2_decap_4 FILLER_9_143 ();
 sg13g2_fill_1 FILLER_9_147 ();
 sg13g2_fill_2 FILLER_9_157 ();
 sg13g2_fill_1 FILLER_9_165 ();
 sg13g2_decap_4 FILLER_9_171 ();
 sg13g2_fill_1 FILLER_9_175 ();
 sg13g2_fill_1 FILLER_9_181 ();
 sg13g2_decap_4 FILLER_9_195 ();
 sg13g2_fill_2 FILLER_9_199 ();
 sg13g2_fill_2 FILLER_9_205 ();
 sg13g2_fill_1 FILLER_9_207 ();
 sg13g2_fill_2 FILLER_9_275 ();
 sg13g2_fill_1 FILLER_9_277 ();
 sg13g2_fill_2 FILLER_9_288 ();
 sg13g2_fill_1 FILLER_9_320 ();
 sg13g2_fill_2 FILLER_9_360 ();
 sg13g2_fill_1 FILLER_9_362 ();
 sg13g2_fill_2 FILLER_9_375 ();
 sg13g2_fill_2 FILLER_9_388 ();
 sg13g2_fill_1 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_29 ();
 sg13g2_fill_2 FILLER_10_36 ();
 sg13g2_fill_1 FILLER_10_65 ();
 sg13g2_fill_2 FILLER_10_75 ();
 sg13g2_fill_1 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_83 ();
 sg13g2_decap_4 FILLER_10_90 ();
 sg13g2_fill_1 FILLER_10_94 ();
 sg13g2_fill_2 FILLER_10_100 ();
 sg13g2_decap_4 FILLER_10_138 ();
 sg13g2_fill_2 FILLER_10_142 ();
 sg13g2_fill_2 FILLER_10_172 ();
 sg13g2_decap_4 FILLER_10_200 ();
 sg13g2_fill_2 FILLER_10_204 ();
 sg13g2_decap_4 FILLER_10_216 ();
 sg13g2_fill_2 FILLER_10_254 ();
 sg13g2_fill_1 FILLER_10_261 ();
 sg13g2_fill_2 FILLER_10_329 ();
 sg13g2_fill_1 FILLER_10_342 ();
 sg13g2_fill_1 FILLER_10_364 ();
 sg13g2_fill_2 FILLER_10_387 ();
 sg13g2_fill_1 FILLER_10_389 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_24 ();
 sg13g2_fill_1 FILLER_11_31 ();
 sg13g2_fill_2 FILLER_11_68 ();
 sg13g2_fill_1 FILLER_11_75 ();
 sg13g2_decap_4 FILLER_11_86 ();
 sg13g2_decap_4 FILLER_11_106 ();
 sg13g2_fill_1 FILLER_11_174 ();
 sg13g2_fill_2 FILLER_11_215 ();
 sg13g2_fill_1 FILLER_11_217 ();
 sg13g2_fill_2 FILLER_11_229 ();
 sg13g2_decap_8 FILLER_11_235 ();
 sg13g2_decap_4 FILLER_11_242 ();
 sg13g2_fill_1 FILLER_11_246 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_fill_1 FILLER_11_273 ();
 sg13g2_fill_2 FILLER_11_319 ();
 sg13g2_fill_1 FILLER_11_321 ();
 sg13g2_fill_1 FILLER_11_332 ();
 sg13g2_fill_1 FILLER_11_343 ();
 sg13g2_fill_1 FILLER_11_349 ();
 sg13g2_fill_1 FILLER_11_356 ();
 sg13g2_fill_1 FILLER_11_376 ();
 sg13g2_fill_2 FILLER_11_391 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_2 ();
 sg13g2_fill_2 FILLER_12_12 ();
 sg13g2_fill_2 FILLER_12_19 ();
 sg13g2_decap_4 FILLER_12_35 ();
 sg13g2_fill_2 FILLER_12_39 ();
 sg13g2_fill_2 FILLER_12_45 ();
 sg13g2_fill_1 FILLER_12_47 ();
 sg13g2_decap_8 FILLER_12_53 ();
 sg13g2_fill_2 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_72 ();
 sg13g2_decap_8 FILLER_12_83 ();
 sg13g2_decap_8 FILLER_12_90 ();
 sg13g2_fill_1 FILLER_12_97 ();
 sg13g2_fill_1 FILLER_12_106 ();
 sg13g2_fill_1 FILLER_12_120 ();
 sg13g2_fill_2 FILLER_12_142 ();
 sg13g2_decap_4 FILLER_12_218 ();
 sg13g2_fill_1 FILLER_12_222 ();
 sg13g2_decap_4 FILLER_12_243 ();
 sg13g2_fill_1 FILLER_12_247 ();
 sg13g2_decap_4 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_267 ();
 sg13g2_decap_4 FILLER_12_274 ();
 sg13g2_fill_1 FILLER_12_278 ();
 sg13g2_fill_2 FILLER_12_284 ();
 sg13g2_fill_1 FILLER_12_286 ();
 sg13g2_fill_2 FILLER_12_307 ();
 sg13g2_fill_1 FILLER_12_309 ();
 sg13g2_fill_2 FILLER_12_314 ();
 sg13g2_fill_2 FILLER_12_328 ();
 sg13g2_fill_1 FILLER_12_330 ();
 sg13g2_fill_2 FILLER_12_387 ();
 sg13g2_fill_2 FILLER_12_394 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_2 ();
 sg13g2_fill_2 FILLER_13_42 ();
 sg13g2_fill_2 FILLER_13_50 ();
 sg13g2_fill_2 FILLER_13_60 ();
 sg13g2_fill_1 FILLER_13_62 ();
 sg13g2_fill_2 FILLER_13_67 ();
 sg13g2_decap_8 FILLER_13_74 ();
 sg13g2_decap_4 FILLER_13_81 ();
 sg13g2_fill_2 FILLER_13_85 ();
 sg13g2_fill_2 FILLER_13_96 ();
 sg13g2_fill_2 FILLER_13_104 ();
 sg13g2_decap_4 FILLER_13_110 ();
 sg13g2_decap_8 FILLER_13_120 ();
 sg13g2_fill_2 FILLER_13_127 ();
 sg13g2_decap_4 FILLER_13_134 ();
 sg13g2_fill_1 FILLER_13_138 ();
 sg13g2_decap_4 FILLER_13_153 ();
 sg13g2_fill_1 FILLER_13_204 ();
 sg13g2_decap_4 FILLER_13_224 ();
 sg13g2_fill_2 FILLER_13_228 ();
 sg13g2_decap_4 FILLER_13_241 ();
 sg13g2_fill_1 FILLER_13_271 ();
 sg13g2_decap_8 FILLER_13_289 ();
 sg13g2_decap_8 FILLER_13_300 ();
 sg13g2_decap_8 FILLER_13_307 ();
 sg13g2_fill_2 FILLER_13_314 ();
 sg13g2_fill_1 FILLER_13_324 ();
 sg13g2_fill_1 FILLER_13_354 ();
 sg13g2_fill_2 FILLER_13_360 ();
 sg13g2_fill_1 FILLER_13_362 ();
 sg13g2_fill_1 FILLER_13_381 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_fill_2 FILLER_14_17 ();
 sg13g2_fill_1 FILLER_14_77 ();
 sg13g2_fill_2 FILLER_14_92 ();
 sg13g2_fill_2 FILLER_14_106 ();
 sg13g2_fill_1 FILLER_14_108 ();
 sg13g2_fill_1 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_146 ();
 sg13g2_decap_8 FILLER_14_153 ();
 sg13g2_decap_8 FILLER_14_160 ();
 sg13g2_fill_2 FILLER_14_167 ();
 sg13g2_fill_2 FILLER_14_230 ();
 sg13g2_decap_4 FILLER_14_251 ();
 sg13g2_fill_1 FILLER_14_255 ();
 sg13g2_fill_2 FILLER_14_297 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_4 FILLER_14_315 ();
 sg13g2_fill_1 FILLER_14_319 ();
 sg13g2_fill_1 FILLER_14_329 ();
 sg13g2_fill_2 FILLER_14_366 ();
 sg13g2_fill_1 FILLER_14_373 ();
 sg13g2_fill_2 FILLER_14_379 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_4 ();
 sg13g2_fill_1 FILLER_15_15 ();
 sg13g2_fill_2 FILLER_15_80 ();
 sg13g2_fill_1 FILLER_15_82 ();
 sg13g2_fill_2 FILLER_15_111 ();
 sg13g2_fill_2 FILLER_15_141 ();
 sg13g2_fill_1 FILLER_15_143 ();
 sg13g2_fill_1 FILLER_15_149 ();
 sg13g2_fill_2 FILLER_15_167 ();
 sg13g2_fill_1 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_197 ();
 sg13g2_fill_1 FILLER_15_208 ();
 sg13g2_fill_1 FILLER_15_243 ();
 sg13g2_decap_4 FILLER_15_249 ();
 sg13g2_decap_8 FILLER_15_257 ();
 sg13g2_fill_1 FILLER_15_264 ();
 sg13g2_fill_1 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_312 ();
 sg13g2_fill_2 FILLER_15_319 ();
 sg13g2_decap_4 FILLER_15_326 ();
 sg13g2_fill_2 FILLER_15_345 ();
 sg13g2_fill_1 FILLER_15_347 ();
 sg13g2_fill_2 FILLER_15_386 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_4 ();
 sg13g2_fill_2 FILLER_16_25 ();
 sg13g2_decap_4 FILLER_16_36 ();
 sg13g2_fill_1 FILLER_16_40 ();
 sg13g2_fill_1 FILLER_16_50 ();
 sg13g2_fill_1 FILLER_16_105 ();
 sg13g2_fill_2 FILLER_16_123 ();
 sg13g2_fill_2 FILLER_16_131 ();
 sg13g2_fill_2 FILLER_16_170 ();
 sg13g2_fill_2 FILLER_16_219 ();
 sg13g2_decap_4 FILLER_16_238 ();
 sg13g2_decap_4 FILLER_16_268 ();
 sg13g2_fill_2 FILLER_16_277 ();
 sg13g2_fill_1 FILLER_16_279 ();
 sg13g2_decap_4 FILLER_16_297 ();
 sg13g2_fill_2 FILLER_16_319 ();
 sg13g2_fill_1 FILLER_16_321 ();
 sg13g2_fill_2 FILLER_16_342 ();
 sg13g2_fill_1 FILLER_16_344 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_17 ();
 sg13g2_fill_1 FILLER_17_40 ();
 sg13g2_decap_4 FILLER_17_68 ();
 sg13g2_fill_1 FILLER_17_72 ();
 sg13g2_fill_2 FILLER_17_77 ();
 sg13g2_fill_1 FILLER_17_79 ();
 sg13g2_fill_1 FILLER_17_94 ();
 sg13g2_fill_2 FILLER_17_103 ();
 sg13g2_fill_1 FILLER_17_105 ();
 sg13g2_decap_4 FILLER_17_110 ();
 sg13g2_fill_1 FILLER_17_123 ();
 sg13g2_fill_2 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_137 ();
 sg13g2_fill_1 FILLER_17_139 ();
 sg13g2_fill_1 FILLER_17_177 ();
 sg13g2_decap_8 FILLER_17_212 ();
 sg13g2_decap_4 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_223 ();
 sg13g2_decap_4 FILLER_17_229 ();
 sg13g2_decap_4 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_268 ();
 sg13g2_decap_4 FILLER_17_275 ();
 sg13g2_fill_1 FILLER_17_292 ();
 sg13g2_fill_2 FILLER_17_300 ();
 sg13g2_fill_2 FILLER_17_313 ();
 sg13g2_fill_1 FILLER_17_315 ();
 sg13g2_fill_2 FILLER_17_329 ();
 sg13g2_fill_2 FILLER_17_349 ();
 sg13g2_fill_2 FILLER_17_366 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_13 ();
 sg13g2_fill_2 FILLER_18_26 ();
 sg13g2_decap_8 FILLER_18_55 ();
 sg13g2_decap_8 FILLER_18_66 ();
 sg13g2_decap_4 FILLER_18_73 ();
 sg13g2_fill_2 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_89 ();
 sg13g2_fill_1 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_97 ();
 sg13g2_fill_2 FILLER_18_121 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_fill_1 FILLER_18_140 ();
 sg13g2_fill_1 FILLER_18_150 ();
 sg13g2_fill_2 FILLER_18_182 ();
 sg13g2_decap_4 FILLER_18_218 ();
 sg13g2_fill_2 FILLER_18_248 ();
 sg13g2_fill_2 FILLER_18_280 ();
 sg13g2_fill_1 FILLER_18_282 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_fill_2 FILLER_18_344 ();
 sg13g2_fill_1 FILLER_18_357 ();
 sg13g2_fill_2 FILLER_18_402 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_fill_2 FILLER_19_19 ();
 sg13g2_fill_2 FILLER_19_56 ();
 sg13g2_fill_1 FILLER_19_58 ();
 sg13g2_fill_1 FILLER_19_75 ();
 sg13g2_fill_1 FILLER_19_98 ();
 sg13g2_fill_1 FILLER_19_114 ();
 sg13g2_fill_2 FILLER_19_121 ();
 sg13g2_fill_1 FILLER_19_123 ();
 sg13g2_decap_4 FILLER_19_156 ();
 sg13g2_fill_1 FILLER_19_160 ();
 sg13g2_fill_2 FILLER_19_173 ();
 sg13g2_fill_1 FILLER_19_175 ();
 sg13g2_decap_4 FILLER_19_193 ();
 sg13g2_fill_2 FILLER_19_197 ();
 sg13g2_decap_4 FILLER_19_224 ();
 sg13g2_fill_1 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_fill_1 FILLER_19_245 ();
 sg13g2_fill_2 FILLER_19_290 ();
 sg13g2_fill_2 FILLER_19_297 ();
 sg13g2_decap_8 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_321 ();
 sg13g2_fill_1 FILLER_19_326 ();
 sg13g2_fill_1 FILLER_19_343 ();
 sg13g2_fill_2 FILLER_19_381 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_fill_2 FILLER_20_34 ();
 sg13g2_fill_1 FILLER_20_36 ();
 sg13g2_fill_1 FILLER_20_49 ();
 sg13g2_fill_1 FILLER_20_55 ();
 sg13g2_fill_2 FILLER_20_74 ();
 sg13g2_fill_2 FILLER_20_101 ();
 sg13g2_fill_2 FILLER_20_108 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_fill_2 FILLER_20_142 ();
 sg13g2_fill_1 FILLER_20_144 ();
 sg13g2_decap_8 FILLER_20_157 ();
 sg13g2_decap_8 FILLER_20_164 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_182 ();
 sg13g2_fill_1 FILLER_20_184 ();
 sg13g2_decap_4 FILLER_20_193 ();
 sg13g2_fill_1 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_272 ();
 sg13g2_fill_1 FILLER_20_313 ();
 sg13g2_fill_1 FILLER_20_322 ();
 sg13g2_fill_2 FILLER_20_340 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_fill_1 FILLER_21_20 ();
 sg13g2_fill_1 FILLER_21_35 ();
 sg13g2_fill_2 FILLER_21_51 ();
 sg13g2_fill_1 FILLER_21_53 ();
 sg13g2_fill_2 FILLER_21_68 ();
 sg13g2_fill_1 FILLER_21_70 ();
 sg13g2_decap_4 FILLER_21_101 ();
 sg13g2_fill_2 FILLER_21_112 ();
 sg13g2_fill_1 FILLER_21_114 ();
 sg13g2_fill_2 FILLER_21_142 ();
 sg13g2_decap_4 FILLER_21_184 ();
 sg13g2_decap_4 FILLER_21_193 ();
 sg13g2_fill_2 FILLER_21_197 ();
 sg13g2_fill_2 FILLER_21_226 ();
 sg13g2_fill_1 FILLER_21_228 ();
 sg13g2_decap_4 FILLER_21_234 ();
 sg13g2_decap_8 FILLER_21_270 ();
 sg13g2_decap_4 FILLER_21_277 ();
 sg13g2_fill_1 FILLER_21_281 ();
 sg13g2_fill_1 FILLER_21_345 ();
 sg13g2_fill_2 FILLER_21_372 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_12 ();
 sg13g2_fill_2 FILLER_22_59 ();
 sg13g2_fill_2 FILLER_22_73 ();
 sg13g2_fill_1 FILLER_22_75 ();
 sg13g2_fill_1 FILLER_22_100 ();
 sg13g2_fill_2 FILLER_22_110 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_fill_2 FILLER_22_210 ();
 sg13g2_fill_1 FILLER_22_217 ();
 sg13g2_fill_2 FILLER_22_248 ();
 sg13g2_fill_2 FILLER_22_303 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_67 ();
 sg13g2_fill_2 FILLER_23_118 ();
 sg13g2_fill_1 FILLER_23_120 ();
 sg13g2_decap_4 FILLER_23_136 ();
 sg13g2_fill_1 FILLER_23_140 ();
 sg13g2_fill_2 FILLER_23_232 ();
 sg13g2_fill_1 FILLER_23_234 ();
 sg13g2_decap_4 FILLER_23_280 ();
 sg13g2_fill_1 FILLER_23_284 ();
 sg13g2_fill_2 FILLER_23_393 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_2 ();
 sg13g2_fill_1 FILLER_24_50 ();
 sg13g2_decap_4 FILLER_24_56 ();
 sg13g2_fill_2 FILLER_24_110 ();
 sg13g2_fill_1 FILLER_24_112 ();
 sg13g2_fill_2 FILLER_24_154 ();
 sg13g2_fill_1 FILLER_24_191 ();
 sg13g2_fill_2 FILLER_24_197 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_209 ();
 sg13g2_fill_2 FILLER_24_259 ();
 sg13g2_decap_4 FILLER_24_287 ();
 sg13g2_fill_1 FILLER_24_334 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_11 ();
 sg13g2_decap_4 FILLER_25_20 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_4 FILLER_25_64 ();
 sg13g2_fill_1 FILLER_25_68 ();
 sg13g2_fill_1 FILLER_25_113 ();
 sg13g2_decap_4 FILLER_25_118 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_decap_4 FILLER_25_132 ();
 sg13g2_fill_1 FILLER_25_136 ();
 sg13g2_decap_8 FILLER_25_141 ();
 sg13g2_fill_1 FILLER_25_148 ();
 sg13g2_fill_2 FILLER_25_154 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_fill_2 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_163 ();
 sg13g2_fill_2 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_243 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_fill_2 FILLER_25_292 ();
 sg13g2_fill_2 FILLER_25_307 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_63 ();
 sg13g2_decap_4 FILLER_26_70 ();
 sg13g2_fill_1 FILLER_26_74 ();
 sg13g2_fill_2 FILLER_26_105 ();
 sg13g2_fill_2 FILLER_26_117 ();
 sg13g2_fill_2 FILLER_26_124 ();
 sg13g2_fill_1 FILLER_26_126 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_167 ();
 sg13g2_decap_8 FILLER_26_187 ();
 sg13g2_decap_4 FILLER_26_194 ();
 sg13g2_decap_8 FILLER_26_207 ();
 sg13g2_fill_1 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_223 ();
 sg13g2_fill_2 FILLER_26_241 ();
 sg13g2_fill_1 FILLER_26_243 ();
 sg13g2_decap_8 FILLER_26_274 ();
 sg13g2_fill_1 FILLER_26_315 ();
 sg13g2_fill_2 FILLER_26_331 ();
 sg13g2_fill_2 FILLER_26_347 ();
 sg13g2_fill_2 FILLER_26_398 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_15 ();
 sg13g2_fill_1 FILLER_27_19 ();
 sg13g2_decap_8 FILLER_27_30 ();
 sg13g2_fill_2 FILLER_27_37 ();
 sg13g2_decap_4 FILLER_27_45 ();
 sg13g2_fill_1 FILLER_27_49 ();
 sg13g2_decap_4 FILLER_27_54 ();
 sg13g2_fill_1 FILLER_27_74 ();
 sg13g2_fill_1 FILLER_27_86 ();
 sg13g2_fill_2 FILLER_27_92 ();
 sg13g2_fill_1 FILLER_27_94 ();
 sg13g2_fill_1 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_decap_4 FILLER_27_192 ();
 sg13g2_fill_2 FILLER_27_196 ();
 sg13g2_fill_2 FILLER_27_226 ();
 sg13g2_fill_2 FILLER_27_336 ();
 sg13g2_fill_2 FILLER_27_397 ();
 sg13g2_fill_1 FILLER_28_73 ();
 sg13g2_fill_2 FILLER_28_89 ();
 sg13g2_fill_1 FILLER_28_91 ();
 sg13g2_fill_2 FILLER_28_106 ();
 sg13g2_fill_1 FILLER_28_108 ();
 sg13g2_fill_2 FILLER_28_124 ();
 sg13g2_decap_4 FILLER_28_135 ();
 sg13g2_fill_1 FILLER_28_139 ();
 sg13g2_decap_4 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_182 ();
 sg13g2_decap_4 FILLER_28_193 ();
 sg13g2_fill_2 FILLER_28_197 ();
 sg13g2_fill_2 FILLER_28_220 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_fill_2 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_decap_8 FILLER_28_254 ();
 sg13g2_fill_1 FILLER_29_75 ();
 sg13g2_fill_2 FILLER_29_86 ();
 sg13g2_fill_1 FILLER_29_88 ();
 sg13g2_decap_4 FILLER_29_95 ();
 sg13g2_fill_2 FILLER_29_111 ();
 sg13g2_fill_1 FILLER_29_113 ();
 sg13g2_fill_2 FILLER_29_138 ();
 sg13g2_fill_1 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_150 ();
 sg13g2_decap_8 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_fill_2 FILLER_29_178 ();
 sg13g2_fill_1 FILLER_29_192 ();
 sg13g2_decap_4 FILLER_29_256 ();
 sg13g2_fill_2 FILLER_29_260 ();
 sg13g2_fill_1 FILLER_29_327 ();
 sg13g2_fill_1 FILLER_29_333 ();
 sg13g2_fill_2 FILLER_29_344 ();
 sg13g2_fill_2 FILLER_29_352 ();
 sg13g2_fill_1 FILLER_29_373 ();
 sg13g2_fill_1 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_36 ();
 sg13g2_fill_1 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_95 ();
 sg13g2_fill_1 FILLER_30_102 ();
 sg13g2_fill_2 FILLER_30_108 ();
 sg13g2_fill_1 FILLER_30_110 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_decap_8 FILLER_30_142 ();
 sg13g2_decap_8 FILLER_30_149 ();
 sg13g2_decap_4 FILLER_30_156 ();
 sg13g2_fill_2 FILLER_30_165 ();
 sg13g2_decap_4 FILLER_30_219 ();
 sg13g2_fill_1 FILLER_30_268 ();
 sg13g2_fill_1 FILLER_30_369 ();
 sg13g2_fill_1 FILLER_31_53 ();
 sg13g2_fill_2 FILLER_31_75 ();
 sg13g2_decap_4 FILLER_31_96 ();
 sg13g2_fill_2 FILLER_31_129 ();
 sg13g2_fill_2 FILLER_31_176 ();
 sg13g2_decap_8 FILLER_31_230 ();
 sg13g2_decap_4 FILLER_31_237 ();
 sg13g2_fill_2 FILLER_31_241 ();
 sg13g2_fill_2 FILLER_31_270 ();
 sg13g2_fill_2 FILLER_31_298 ();
 sg13g2_fill_1 FILLER_31_340 ();
 sg13g2_fill_2 FILLER_31_393 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_41 ();
 sg13g2_fill_1 FILLER_32_51 ();
 sg13g2_fill_1 FILLER_32_66 ();
 sg13g2_fill_2 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_108 ();
 sg13g2_fill_1 FILLER_32_143 ();
 sg13g2_fill_2 FILLER_32_174 ();
 sg13g2_fill_1 FILLER_32_176 ();
 sg13g2_fill_1 FILLER_32_213 ();
 sg13g2_decap_8 FILLER_32_239 ();
 sg13g2_fill_1 FILLER_32_246 ();
 sg13g2_fill_2 FILLER_32_274 ();
 sg13g2_fill_1 FILLER_32_276 ();
 sg13g2_fill_2 FILLER_32_287 ();
 sg13g2_fill_1 FILLER_32_289 ();
 sg13g2_fill_2 FILLER_32_303 ();
 sg13g2_fill_1 FILLER_32_305 ();
 sg13g2_fill_2 FILLER_32_329 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_fill_1 FILLER_33_26 ();
 sg13g2_fill_2 FILLER_33_75 ();
 sg13g2_fill_2 FILLER_33_101 ();
 sg13g2_fill_2 FILLER_33_107 ();
 sg13g2_fill_1 FILLER_33_109 ();
 sg13g2_fill_1 FILLER_33_122 ();
 sg13g2_fill_2 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_188 ();
 sg13g2_decap_8 FILLER_33_195 ();
 sg13g2_fill_2 FILLER_33_202 ();
 sg13g2_fill_1 FILLER_33_208 ();
 sg13g2_fill_2 FILLER_33_214 ();
 sg13g2_fill_2 FILLER_33_231 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_decap_8 FILLER_33_267 ();
 sg13g2_decap_4 FILLER_33_274 ();
 sg13g2_fill_2 FILLER_33_278 ();
 sg13g2_fill_1 FILLER_33_328 ();
 sg13g2_fill_1 FILLER_33_357 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_64 ();
 sg13g2_fill_1 FILLER_34_66 ();
 sg13g2_fill_1 FILLER_34_97 ();
 sg13g2_decap_4 FILLER_34_120 ();
 sg13g2_fill_1 FILLER_34_124 ();
 sg13g2_fill_2 FILLER_34_130 ();
 sg13g2_fill_2 FILLER_34_138 ();
 sg13g2_fill_1 FILLER_34_140 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_decap_4 FILLER_34_178 ();
 sg13g2_fill_1 FILLER_34_182 ();
 sg13g2_fill_2 FILLER_34_191 ();
 sg13g2_fill_1 FILLER_34_193 ();
 sg13g2_fill_2 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_277 ();
 sg13g2_fill_1 FILLER_34_288 ();
 sg13g2_fill_2 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_31 ();
 sg13g2_fill_2 FILLER_35_54 ();
 sg13g2_fill_2 FILLER_35_85 ();
 sg13g2_fill_2 FILLER_35_103 ();
 sg13g2_fill_2 FILLER_35_110 ();
 sg13g2_fill_1 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_121 ();
 sg13g2_decap_4 FILLER_35_135 ();
 sg13g2_fill_1 FILLER_35_139 ();
 sg13g2_fill_2 FILLER_35_169 ();
 sg13g2_fill_2 FILLER_35_207 ();
 sg13g2_fill_1 FILLER_35_209 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_fill_1 FILLER_35_222 ();
 sg13g2_fill_2 FILLER_35_235 ();
 sg13g2_fill_1 FILLER_35_237 ();
 sg13g2_fill_2 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_310 ();
 sg13g2_fill_2 FILLER_35_316 ();
 sg13g2_fill_1 FILLER_35_318 ();
 sg13g2_fill_1 FILLER_35_354 ();
 sg13g2_fill_2 FILLER_35_382 ();
 sg13g2_decap_4 FILLER_36_140 ();
 sg13g2_fill_2 FILLER_36_144 ();
 sg13g2_fill_2 FILLER_36_203 ();
 sg13g2_fill_1 FILLER_36_214 ();
 sg13g2_decap_4 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_fill_2 FILLER_36_263 ();
 sg13g2_fill_2 FILLER_36_271 ();
 sg13g2_fill_2 FILLER_36_313 ();
 sg13g2_fill_2 FILLER_36_354 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_32 ();
 sg13g2_fill_2 FILLER_37_75 ();
 sg13g2_fill_1 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_107 ();
 sg13g2_fill_1 FILLER_37_109 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_2 FILLER_37_154 ();
 sg13g2_fill_2 FILLER_37_182 ();
 sg13g2_fill_1 FILLER_37_198 ();
 sg13g2_fill_2 FILLER_37_209 ();
 sg13g2_fill_1 FILLER_37_251 ();
 sg13g2_fill_2 FILLER_37_277 ();
 sg13g2_fill_2 FILLER_37_364 ();
 sg13g2_fill_1 FILLER_37_381 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_75 ();
 sg13g2_fill_2 FILLER_38_96 ();
 sg13g2_fill_1 FILLER_38_98 ();
 sg13g2_fill_1 FILLER_38_109 ();
 sg13g2_decap_8 FILLER_38_115 ();
 sg13g2_decap_8 FILLER_38_122 ();
 sg13g2_fill_2 FILLER_38_129 ();
 sg13g2_fill_1 FILLER_38_131 ();
 sg13g2_fill_2 FILLER_38_141 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_fill_2 FILLER_38_190 ();
 sg13g2_fill_1 FILLER_38_192 ();
 sg13g2_fill_2 FILLER_38_233 ();
 sg13g2_fill_1 FILLER_38_235 ();
 sg13g2_fill_2 FILLER_38_277 ();
 sg13g2_fill_2 FILLER_38_289 ();
 sg13g2_fill_2 FILLER_38_300 ();
 sg13g2_fill_1 FILLER_38_302 ();
 sg13g2_fill_2 FILLER_38_380 ();
 sg13g2_fill_1 FILLER_38_382 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_decap_4 FILLER_39_48 ();
 sg13g2_fill_1 FILLER_39_52 ();
 sg13g2_decap_8 FILLER_39_64 ();
 sg13g2_decap_8 FILLER_39_71 ();
 sg13g2_decap_8 FILLER_39_78 ();
 sg13g2_decap_8 FILLER_39_85 ();
 sg13g2_fill_1 FILLER_39_92 ();
 sg13g2_decap_8 FILLER_39_97 ();
 sg13g2_decap_8 FILLER_39_104 ();
 sg13g2_decap_8 FILLER_39_111 ();
 sg13g2_decap_8 FILLER_39_118 ();
 sg13g2_fill_2 FILLER_39_125 ();
 sg13g2_fill_1 FILLER_39_159 ();
 sg13g2_fill_2 FILLER_39_213 ();
 sg13g2_fill_2 FILLER_39_287 ();
 sg13g2_fill_1 FILLER_39_289 ();
 sg13g2_fill_1 FILLER_39_340 ();
 sg13g2_fill_2 FILLER_39_356 ();
 sg13g2_fill_2 FILLER_39_364 ();
 sg13g2_fill_2 FILLER_39_381 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_4 FILLER_40_50 ();
 sg13g2_fill_1 FILLER_40_70 ();
 sg13g2_fill_2 FILLER_40_79 ();
 sg13g2_fill_1 FILLER_40_81 ();
 sg13g2_fill_2 FILLER_40_95 ();
 sg13g2_decap_8 FILLER_40_102 ();
 sg13g2_decap_8 FILLER_40_109 ();
 sg13g2_fill_2 FILLER_40_116 ();
 sg13g2_fill_2 FILLER_40_144 ();
 sg13g2_fill_2 FILLER_40_207 ();
 sg13g2_fill_1 FILLER_40_209 ();
 sg13g2_fill_2 FILLER_40_267 ();
 sg13g2_fill_2 FILLER_40_279 ();
 sg13g2_fill_1 FILLER_40_370 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_fill_1 FILLER_41_26 ();
 sg13g2_fill_2 FILLER_41_59 ();
 sg13g2_fill_1 FILLER_41_61 ();
 sg13g2_fill_2 FILLER_41_97 ();
 sg13g2_fill_1 FILLER_41_99 ();
 sg13g2_fill_2 FILLER_41_105 ();
 sg13g2_fill_1 FILLER_41_107 ();
 sg13g2_fill_2 FILLER_41_134 ();
 sg13g2_fill_1 FILLER_41_136 ();
 sg13g2_fill_1 FILLER_41_147 ();
 sg13g2_fill_2 FILLER_41_158 ();
 sg13g2_fill_1 FILLER_41_160 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_4 FILLER_41_175 ();
 sg13g2_fill_1 FILLER_41_179 ();
 sg13g2_fill_1 FILLER_41_215 ();
 sg13g2_decap_8 FILLER_41_221 ();
 sg13g2_decap_8 FILLER_41_228 ();
 sg13g2_fill_1 FILLER_41_235 ();
 sg13g2_decap_4 FILLER_41_240 ();
 sg13g2_fill_1 FILLER_41_251 ();
 sg13g2_fill_1 FILLER_41_257 ();
 sg13g2_fill_2 FILLER_41_284 ();
 sg13g2_decap_8 FILLER_41_312 ();
 sg13g2_fill_2 FILLER_41_319 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_86 ();
 sg13g2_fill_2 FILLER_42_113 ();
 sg13g2_fill_2 FILLER_42_128 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_4 FILLER_42_154 ();
 sg13g2_fill_1 FILLER_42_158 ();
 sg13g2_decap_8 FILLER_42_164 ();
 sg13g2_decap_4 FILLER_42_171 ();
 sg13g2_fill_1 FILLER_42_175 ();
 sg13g2_fill_1 FILLER_42_208 ();
 sg13g2_fill_2 FILLER_42_225 ();
 sg13g2_fill_2 FILLER_42_240 ();
 sg13g2_decap_4 FILLER_42_246 ();
 sg13g2_fill_1 FILLER_42_250 ();
 sg13g2_decap_8 FILLER_42_255 ();
 sg13g2_fill_2 FILLER_42_294 ();
 sg13g2_fill_2 FILLER_42_348 ();
 sg13g2_fill_1 FILLER_42_350 ();
 sg13g2_fill_2 FILLER_42_381 ();
 sg13g2_fill_2 FILLER_43_90 ();
 sg13g2_decap_8 FILLER_43_134 ();
 sg13g2_fill_1 FILLER_43_141 ();
 sg13g2_fill_1 FILLER_43_172 ();
 sg13g2_fill_1 FILLER_43_194 ();
 sg13g2_fill_1 FILLER_43_200 ();
 sg13g2_fill_1 FILLER_43_213 ();
 sg13g2_decap_8 FILLER_43_256 ();
 sg13g2_fill_1 FILLER_43_263 ();
 sg13g2_decap_8 FILLER_43_320 ();
 sg13g2_fill_1 FILLER_43_327 ();
 sg13g2_fill_2 FILLER_43_332 ();
 sg13g2_fill_1 FILLER_43_334 ();
 sg13g2_fill_2 FILLER_43_339 ();
 sg13g2_fill_1 FILLER_43_341 ();
 sg13g2_decap_8 FILLER_43_346 ();
 sg13g2_decap_8 FILLER_43_353 ();
 sg13g2_fill_2 FILLER_43_360 ();
 sg13g2_fill_1 FILLER_43_370 ();
 sg13g2_fill_2 FILLER_44_35 ();
 sg13g2_fill_1 FILLER_44_73 ();
 sg13g2_fill_2 FILLER_44_83 ();
 sg13g2_fill_1 FILLER_44_102 ();
 sg13g2_decap_8 FILLER_44_128 ();
 sg13g2_fill_1 FILLER_44_135 ();
 sg13g2_fill_2 FILLER_44_146 ();
 sg13g2_fill_2 FILLER_44_174 ();
 sg13g2_fill_1 FILLER_44_176 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_fill_2 FILLER_44_196 ();
 sg13g2_fill_1 FILLER_44_198 ();
 sg13g2_fill_1 FILLER_44_261 ();
 sg13g2_fill_1 FILLER_44_275 ();
 sg13g2_fill_1 FILLER_44_280 ();
 sg13g2_fill_2 FILLER_44_291 ();
 sg13g2_fill_1 FILLER_44_293 ();
 sg13g2_fill_2 FILLER_44_324 ();
 sg13g2_fill_1 FILLER_44_326 ();
 sg13g2_fill_2 FILLER_44_332 ();
 sg13g2_fill_1 FILLER_44_337 ();
 sg13g2_decap_4 FILLER_44_345 ();
 sg13g2_decap_8 FILLER_44_362 ();
 sg13g2_fill_1 FILLER_44_369 ();
 sg13g2_fill_2 FILLER_44_384 ();
 sg13g2_fill_2 FILLER_44_407 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_69 ();
 sg13g2_fill_1 FILLER_45_92 ();
 sg13g2_fill_2 FILLER_45_125 ();
 sg13g2_fill_1 FILLER_45_151 ();
 sg13g2_fill_2 FILLER_45_156 ();
 sg13g2_decap_4 FILLER_45_162 ();
 sg13g2_fill_2 FILLER_45_166 ();
 sg13g2_decap_8 FILLER_45_205 ();
 sg13g2_decap_8 FILLER_45_212 ();
 sg13g2_decap_8 FILLER_45_219 ();
 sg13g2_fill_2 FILLER_45_278 ();
 sg13g2_fill_2 FILLER_45_336 ();
 sg13g2_fill_1 FILLER_45_338 ();
 sg13g2_decap_8 FILLER_45_354 ();
 sg13g2_decap_8 FILLER_45_365 ();
 sg13g2_fill_1 FILLER_45_376 ();
 sg13g2_fill_1 FILLER_45_382 ();
 sg13g2_fill_2 FILLER_45_393 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_fill_1 FILLER_46_17 ();
 sg13g2_fill_1 FILLER_46_25 ();
 sg13g2_fill_1 FILLER_46_39 ();
 sg13g2_fill_2 FILLER_46_55 ();
 sg13g2_fill_2 FILLER_46_116 ();
 sg13g2_fill_2 FILLER_46_123 ();
 sg13g2_fill_2 FILLER_46_140 ();
 sg13g2_fill_1 FILLER_46_166 ();
 sg13g2_fill_2 FILLER_46_180 ();
 sg13g2_decap_8 FILLER_46_187 ();
 sg13g2_fill_1 FILLER_46_194 ();
 sg13g2_fill_2 FILLER_46_205 ();
 sg13g2_decap_8 FILLER_46_215 ();
 sg13g2_decap_8 FILLER_46_226 ();
 sg13g2_fill_1 FILLER_46_241 ();
 sg13g2_fill_2 FILLER_46_291 ();
 sg13g2_fill_1 FILLER_46_333 ();
 sg13g2_fill_1 FILLER_46_364 ();
 sg13g2_fill_2 FILLER_46_393 ();
 sg13g2_fill_1 FILLER_46_395 ();
 sg13g2_fill_2 FILLER_47_86 ();
 sg13g2_fill_2 FILLER_47_108 ();
 sg13g2_fill_1 FILLER_47_110 ();
 sg13g2_fill_1 FILLER_47_123 ();
 sg13g2_fill_2 FILLER_47_154 ();
 sg13g2_fill_2 FILLER_47_185 ();
 sg13g2_fill_1 FILLER_47_187 ();
 sg13g2_fill_2 FILLER_47_204 ();
 sg13g2_fill_2 FILLER_47_244 ();
 sg13g2_fill_1 FILLER_47_246 ();
 sg13g2_fill_2 FILLER_47_275 ();
 sg13g2_fill_1 FILLER_47_355 ();
 sg13g2_fill_1 FILLER_47_383 ();
 sg13g2_fill_1 FILLER_48_61 ();
 sg13g2_fill_1 FILLER_48_89 ();
 sg13g2_fill_1 FILLER_48_109 ();
 sg13g2_fill_2 FILLER_48_126 ();
 sg13g2_fill_1 FILLER_48_128 ();
 sg13g2_fill_1 FILLER_48_142 ();
 sg13g2_decap_4 FILLER_48_148 ();
 sg13g2_fill_2 FILLER_48_152 ();
 sg13g2_decap_4 FILLER_48_159 ();
 sg13g2_fill_1 FILLER_48_163 ();
 sg13g2_fill_1 FILLER_48_218 ();
 sg13g2_fill_1 FILLER_48_227 ();
 sg13g2_decap_8 FILLER_48_255 ();
 sg13g2_fill_1 FILLER_48_262 ();
 sg13g2_decap_8 FILLER_48_275 ();
 sg13g2_fill_1 FILLER_48_286 ();
 sg13g2_decap_4 FILLER_48_291 ();
 sg13g2_fill_2 FILLER_48_295 ();
 sg13g2_fill_2 FILLER_48_306 ();
 sg13g2_fill_1 FILLER_48_308 ();
 sg13g2_fill_2 FILLER_48_313 ();
 sg13g2_fill_1 FILLER_48_315 ();
 sg13g2_decap_4 FILLER_48_346 ();
 sg13g2_fill_2 FILLER_48_350 ();
 sg13g2_fill_2 FILLER_48_366 ();
 sg13g2_fill_1 FILLER_48_379 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_83 ();
 sg13g2_fill_2 FILLER_49_130 ();
 sg13g2_fill_1 FILLER_49_132 ();
 sg13g2_fill_2 FILLER_49_141 ();
 sg13g2_fill_1 FILLER_49_143 ();
 sg13g2_decap_8 FILLER_49_149 ();
 sg13g2_decap_8 FILLER_49_156 ();
 sg13g2_fill_1 FILLER_49_163 ();
 sg13g2_decap_8 FILLER_49_173 ();
 sg13g2_decap_4 FILLER_49_180 ();
 sg13g2_fill_2 FILLER_49_184 ();
 sg13g2_decap_4 FILLER_49_194 ();
 sg13g2_fill_2 FILLER_49_215 ();
 sg13g2_fill_1 FILLER_49_217 ();
 sg13g2_fill_2 FILLER_49_241 ();
 sg13g2_fill_1 FILLER_49_243 ();
 sg13g2_fill_2 FILLER_49_264 ();
 sg13g2_fill_1 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_271 ();
 sg13g2_decap_8 FILLER_49_278 ();
 sg13g2_decap_4 FILLER_49_337 ();
 sg13g2_decap_8 FILLER_49_345 ();
 sg13g2_decap_4 FILLER_49_352 ();
 sg13g2_fill_2 FILLER_49_368 ();
 sg13g2_fill_2 FILLER_49_380 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_2 ();
 sg13g2_fill_1 FILLER_50_31 ();
 sg13g2_fill_1 FILLER_50_132 ();
 sg13g2_fill_2 FILLER_50_149 ();
 sg13g2_fill_1 FILLER_50_151 ();
 sg13g2_fill_1 FILLER_50_168 ();
 sg13g2_decap_4 FILLER_50_177 ();
 sg13g2_fill_2 FILLER_50_181 ();
 sg13g2_decap_8 FILLER_50_201 ();
 sg13g2_decap_8 FILLER_50_208 ();
 sg13g2_decap_8 FILLER_50_215 ();
 sg13g2_decap_8 FILLER_50_222 ();
 sg13g2_decap_8 FILLER_50_229 ();
 sg13g2_decap_8 FILLER_50_236 ();
 sg13g2_decap_4 FILLER_50_243 ();
 sg13g2_fill_2 FILLER_50_247 ();
 sg13g2_decap_4 FILLER_50_257 ();
 sg13g2_decap_8 FILLER_50_281 ();
 sg13g2_decap_8 FILLER_50_304 ();
 sg13g2_decap_8 FILLER_50_311 ();
 sg13g2_fill_2 FILLER_50_318 ();
 sg13g2_fill_1 FILLER_50_320 ();
 sg13g2_fill_2 FILLER_50_325 ();
 sg13g2_fill_1 FILLER_50_357 ();
 sg13g2_fill_2 FILLER_50_382 ();
 sg13g2_fill_2 FILLER_50_389 ();
 sg13g2_fill_1 FILLER_50_391 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_fill_2 FILLER_51_40 ();
 sg13g2_fill_2 FILLER_51_90 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_fill_2 FILLER_51_133 ();
 sg13g2_fill_1 FILLER_51_135 ();
 sg13g2_fill_1 FILLER_51_173 ();
 sg13g2_fill_2 FILLER_51_186 ();
 sg13g2_fill_1 FILLER_51_188 ();
 sg13g2_fill_2 FILLER_51_193 ();
 sg13g2_fill_1 FILLER_51_195 ();
 sg13g2_fill_1 FILLER_51_208 ();
 sg13g2_fill_1 FILLER_51_226 ();
 sg13g2_fill_2 FILLER_51_243 ();
 sg13g2_fill_1 FILLER_51_245 ();
 sg13g2_decap_8 FILLER_51_305 ();
 sg13g2_decap_8 FILLER_51_312 ();
 sg13g2_decap_8 FILLER_51_319 ();
 sg13g2_decap_8 FILLER_51_326 ();
 sg13g2_decap_8 FILLER_51_333 ();
 sg13g2_decap_8 FILLER_51_340 ();
 sg13g2_decap_8 FILLER_51_347 ();
 sg13g2_decap_4 FILLER_51_354 ();
 sg13g2_fill_1 FILLER_51_358 ();
 sg13g2_fill_2 FILLER_51_406 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_12 ();
 sg13g2_fill_2 FILLER_52_82 ();
 sg13g2_fill_1 FILLER_52_84 ();
 sg13g2_fill_1 FILLER_52_102 ();
 sg13g2_fill_1 FILLER_52_156 ();
 sg13g2_decap_4 FILLER_52_162 ();
 sg13g2_decap_8 FILLER_52_247 ();
 sg13g2_fill_2 FILLER_52_254 ();
 sg13g2_decap_4 FILLER_52_259 ();
 sg13g2_fill_2 FILLER_52_263 ();
 sg13g2_decap_8 FILLER_52_281 ();
 sg13g2_fill_1 FILLER_52_288 ();
 sg13g2_fill_2 FILLER_52_295 ();
 sg13g2_fill_1 FILLER_52_297 ();
 sg13g2_decap_8 FILLER_52_302 ();
 sg13g2_fill_1 FILLER_52_309 ();
 sg13g2_fill_2 FILLER_52_318 ();
 sg13g2_fill_1 FILLER_52_320 ();
 sg13g2_decap_8 FILLER_52_330 ();
 sg13g2_fill_1 FILLER_52_337 ();
 sg13g2_decap_8 FILLER_52_351 ();
 sg13g2_decap_8 FILLER_52_358 ();
 sg13g2_fill_1 FILLER_52_380 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_fill_2 FILLER_53_54 ();
 sg13g2_fill_1 FILLER_53_71 ();
 sg13g2_fill_1 FILLER_53_113 ();
 sg13g2_fill_1 FILLER_53_145 ();
 sg13g2_fill_1 FILLER_53_167 ();
 sg13g2_fill_1 FILLER_53_189 ();
 sg13g2_fill_1 FILLER_53_213 ();
 sg13g2_fill_2 FILLER_53_219 ();
 sg13g2_fill_1 FILLER_53_221 ();
 sg13g2_fill_1 FILLER_53_232 ();
 sg13g2_fill_1 FILLER_53_262 ();
 sg13g2_fill_1 FILLER_53_273 ();
 sg13g2_fill_2 FILLER_53_290 ();
 sg13g2_fill_1 FILLER_53_326 ();
 sg13g2_fill_2 FILLER_53_348 ();
 sg13g2_decap_4 FILLER_53_362 ();
 sg13g2_fill_2 FILLER_53_366 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_fill_1 FILLER_54_104 ();
 sg13g2_fill_2 FILLER_54_114 ();
 sg13g2_fill_1 FILLER_54_116 ();
 sg13g2_fill_1 FILLER_54_125 ();
 sg13g2_decap_8 FILLER_54_152 ();
 sg13g2_fill_1 FILLER_54_159 ();
 sg13g2_fill_1 FILLER_54_170 ();
 sg13g2_decap_8 FILLER_54_204 ();
 sg13g2_decap_8 FILLER_54_211 ();
 sg13g2_decap_4 FILLER_54_218 ();
 sg13g2_fill_2 FILLER_54_222 ();
 sg13g2_decap_4 FILLER_54_245 ();
 sg13g2_fill_2 FILLER_54_303 ();
 sg13g2_decap_4 FILLER_54_317 ();
 sg13g2_fill_2 FILLER_54_359 ();
 sg13g2_fill_1 FILLER_54_361 ();
 sg13g2_fill_1 FILLER_54_395 ();
 sg13g2_fill_2 FILLER_55_44 ();
 sg13g2_fill_1 FILLER_55_123 ();
 sg13g2_decap_8 FILLER_55_129 ();
 sg13g2_decap_8 FILLER_55_136 ();
 sg13g2_decap_8 FILLER_55_143 ();
 sg13g2_decap_8 FILLER_55_150 ();
 sg13g2_fill_1 FILLER_55_157 ();
 sg13g2_fill_1 FILLER_55_164 ();
 sg13g2_fill_2 FILLER_55_175 ();
 sg13g2_fill_2 FILLER_55_181 ();
 sg13g2_decap_8 FILLER_55_200 ();
 sg13g2_fill_1 FILLER_55_240 ();
 sg13g2_decap_4 FILLER_55_246 ();
 sg13g2_fill_2 FILLER_55_257 ();
 sg13g2_fill_2 FILLER_55_264 ();
 sg13g2_fill_1 FILLER_55_303 ();
 sg13g2_fill_1 FILLER_55_316 ();
 sg13g2_fill_2 FILLER_55_322 ();
 sg13g2_fill_1 FILLER_55_324 ();
 sg13g2_fill_1 FILLER_55_368 ();
 sg13g2_fill_1 FILLER_55_387 ();
 sg13g2_fill_1 FILLER_55_393 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_fill_2 FILLER_56_97 ();
 sg13g2_fill_1 FILLER_56_99 ();
 sg13g2_decap_4 FILLER_56_104 ();
 sg13g2_fill_2 FILLER_56_108 ();
 sg13g2_decap_4 FILLER_56_132 ();
 sg13g2_fill_2 FILLER_56_136 ();
 sg13g2_decap_4 FILLER_56_181 ();
 sg13g2_decap_8 FILLER_56_190 ();
 sg13g2_fill_1 FILLER_56_197 ();
 sg13g2_fill_2 FILLER_56_233 ();
 sg13g2_fill_1 FILLER_56_235 ();
 sg13g2_decap_8 FILLER_56_241 ();
 sg13g2_decap_4 FILLER_56_248 ();
 sg13g2_fill_1 FILLER_56_252 ();
 sg13g2_fill_2 FILLER_56_258 ();
 sg13g2_fill_1 FILLER_56_260 ();
 sg13g2_fill_2 FILLER_56_307 ();
 sg13g2_fill_2 FILLER_56_336 ();
 sg13g2_fill_1 FILLER_56_338 ();
 sg13g2_fill_2 FILLER_56_360 ();
 sg13g2_fill_1 FILLER_56_380 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_fill_2 FILLER_57_59 ();
 sg13g2_fill_1 FILLER_57_65 ();
 sg13g2_decap_4 FILLER_57_75 ();
 sg13g2_fill_1 FILLER_57_79 ();
 sg13g2_decap_8 FILLER_57_90 ();
 sg13g2_decap_8 FILLER_57_97 ();
 sg13g2_decap_4 FILLER_57_202 ();
 sg13g2_fill_1 FILLER_57_206 ();
 sg13g2_fill_2 FILLER_57_275 ();
 sg13g2_fill_2 FILLER_57_288 ();
 sg13g2_fill_1 FILLER_57_290 ();
 sg13g2_decap_8 FILLER_57_353 ();
 sg13g2_fill_2 FILLER_57_360 ();
 sg13g2_fill_2 FILLER_57_387 ();
 sg13g2_fill_1 FILLER_57_389 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_fill_2 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_69 ();
 sg13g2_decap_8 FILLER_58_76 ();
 sg13g2_fill_2 FILLER_58_83 ();
 sg13g2_fill_2 FILLER_58_97 ();
 sg13g2_fill_2 FILLER_58_107 ();
 sg13g2_fill_1 FILLER_58_109 ();
 sg13g2_fill_1 FILLER_58_114 ();
 sg13g2_fill_2 FILLER_58_128 ();
 sg13g2_fill_1 FILLER_58_130 ();
 sg13g2_fill_1 FILLER_58_135 ();
 sg13g2_fill_1 FILLER_58_141 ();
 sg13g2_decap_4 FILLER_58_155 ();
 sg13g2_fill_1 FILLER_58_159 ();
 sg13g2_fill_2 FILLER_58_179 ();
 sg13g2_fill_1 FILLER_58_194 ();
 sg13g2_fill_2 FILLER_58_208 ();
 sg13g2_fill_2 FILLER_58_219 ();
 sg13g2_fill_1 FILLER_58_221 ();
 sg13g2_fill_1 FILLER_58_282 ();
 sg13g2_fill_2 FILLER_58_295 ();
 sg13g2_fill_2 FILLER_58_305 ();
 sg13g2_fill_1 FILLER_58_307 ();
 sg13g2_fill_2 FILLER_58_314 ();
 sg13g2_fill_2 FILLER_58_321 ();
 sg13g2_fill_1 FILLER_58_323 ();
 sg13g2_fill_2 FILLER_58_334 ();
 sg13g2_fill_1 FILLER_58_348 ();
 sg13g2_fill_2 FILLER_58_362 ();
 sg13g2_fill_2 FILLER_58_376 ();
 sg13g2_fill_2 FILLER_58_388 ();
 sg13g2_fill_2 FILLER_59_44 ();
 sg13g2_fill_2 FILLER_59_62 ();
 sg13g2_fill_1 FILLER_59_69 ();
 sg13g2_fill_1 FILLER_59_74 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_fill_1 FILLER_59_133 ();
 sg13g2_decap_8 FILLER_59_143 ();
 sg13g2_decap_4 FILLER_59_150 ();
 sg13g2_fill_1 FILLER_59_154 ();
 sg13g2_fill_2 FILLER_59_164 ();
 sg13g2_fill_1 FILLER_59_166 ();
 sg13g2_fill_1 FILLER_59_171 ();
 sg13g2_fill_2 FILLER_59_180 ();
 sg13g2_fill_1 FILLER_59_182 ();
 sg13g2_fill_2 FILLER_59_191 ();
 sg13g2_fill_1 FILLER_59_193 ();
 sg13g2_fill_2 FILLER_59_208 ();
 sg13g2_fill_1 FILLER_59_210 ();
 sg13g2_fill_1 FILLER_59_221 ();
 sg13g2_fill_2 FILLER_59_253 ();
 sg13g2_fill_2 FILLER_59_268 ();
 sg13g2_fill_2 FILLER_59_296 ();
 sg13g2_fill_1 FILLER_59_298 ();
 sg13g2_fill_2 FILLER_59_318 ();
 sg13g2_fill_1 FILLER_59_320 ();
 sg13g2_fill_1 FILLER_59_345 ();
 sg13g2_fill_2 FILLER_59_361 ();
 sg13g2_fill_1 FILLER_59_391 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_fill_2 FILLER_60_4 ();
 sg13g2_fill_1 FILLER_60_6 ();
 sg13g2_fill_2 FILLER_60_12 ();
 sg13g2_fill_1 FILLER_60_14 ();
 sg13g2_fill_2 FILLER_60_28 ();
 sg13g2_fill_2 FILLER_60_36 ();
 sg13g2_fill_1 FILLER_60_46 ();
 sg13g2_fill_1 FILLER_60_86 ();
 sg13g2_fill_2 FILLER_60_96 ();
 sg13g2_fill_2 FILLER_60_106 ();
 sg13g2_fill_2 FILLER_60_116 ();
 sg13g2_fill_1 FILLER_60_122 ();
 sg13g2_fill_1 FILLER_60_128 ();
 sg13g2_decap_4 FILLER_60_145 ();
 sg13g2_fill_2 FILLER_60_157 ();
 sg13g2_fill_2 FILLER_60_168 ();
 sg13g2_fill_1 FILLER_60_170 ();
 sg13g2_fill_2 FILLER_60_183 ();
 sg13g2_fill_1 FILLER_60_185 ();
 sg13g2_fill_2 FILLER_60_196 ();
 sg13g2_fill_1 FILLER_60_198 ();
 sg13g2_decap_4 FILLER_60_210 ();
 sg13g2_fill_1 FILLER_60_222 ();
 sg13g2_fill_2 FILLER_60_236 ();
 sg13g2_decap_8 FILLER_60_243 ();
 sg13g2_decap_8 FILLER_60_250 ();
 sg13g2_decap_8 FILLER_60_257 ();
 sg13g2_fill_1 FILLER_60_264 ();
 sg13g2_fill_2 FILLER_60_277 ();
 sg13g2_fill_1 FILLER_60_321 ();
 sg13g2_fill_2 FILLER_60_350 ();
 sg13g2_fill_2 FILLER_60_367 ();
 sg13g2_fill_2 FILLER_60_389 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_fill_2 FILLER_61_24 ();
 sg13g2_fill_1 FILLER_61_26 ();
 sg13g2_decap_4 FILLER_61_47 ();
 sg13g2_fill_1 FILLER_61_81 ();
 sg13g2_fill_1 FILLER_61_88 ();
 sg13g2_fill_2 FILLER_61_115 ();
 sg13g2_decap_4 FILLER_61_205 ();
 sg13g2_fill_1 FILLER_61_214 ();
 sg13g2_decap_4 FILLER_61_223 ();
 sg13g2_fill_1 FILLER_61_227 ();
 sg13g2_decap_8 FILLER_61_241 ();
 sg13g2_fill_1 FILLER_61_256 ();
 sg13g2_fill_1 FILLER_61_270 ();
 sg13g2_fill_2 FILLER_61_284 ();
 sg13g2_fill_1 FILLER_61_286 ();
 sg13g2_fill_1 FILLER_61_301 ();
 sg13g2_decap_4 FILLER_61_315 ();
 sg13g2_fill_2 FILLER_61_319 ();
 sg13g2_fill_1 FILLER_61_340 ();
 sg13g2_fill_1 FILLER_61_345 ();
 sg13g2_fill_2 FILLER_61_371 ();
 sg13g2_fill_1 FILLER_61_373 ();
 sg13g2_fill_1 FILLER_61_388 ();
 sg13g2_fill_1 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_18 ();
 sg13g2_fill_2 FILLER_62_27 ();
 sg13g2_fill_2 FILLER_62_38 ();
 sg13g2_fill_1 FILLER_62_71 ();
 sg13g2_fill_2 FILLER_62_89 ();
 sg13g2_fill_1 FILLER_62_108 ();
 sg13g2_fill_2 FILLER_62_118 ();
 sg13g2_fill_1 FILLER_62_120 ();
 sg13g2_fill_2 FILLER_62_126 ();
 sg13g2_fill_1 FILLER_62_128 ();
 sg13g2_fill_1 FILLER_62_146 ();
 sg13g2_fill_1 FILLER_62_155 ();
 sg13g2_fill_2 FILLER_62_214 ();
 sg13g2_fill_2 FILLER_62_221 ();
 sg13g2_fill_1 FILLER_62_223 ();
 sg13g2_fill_1 FILLER_62_273 ();
 sg13g2_decap_8 FILLER_62_278 ();
 sg13g2_decap_8 FILLER_62_285 ();
 sg13g2_fill_1 FILLER_62_304 ();
 sg13g2_fill_2 FILLER_62_309 ();
 sg13g2_decap_8 FILLER_62_315 ();
 sg13g2_fill_2 FILLER_62_322 ();
 sg13g2_decap_8 FILLER_62_364 ();
 sg13g2_decap_4 FILLER_62_378 ();
 sg13g2_decap_4 FILLER_62_389 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_21 ();
 sg13g2_fill_1 FILLER_63_33 ();
 sg13g2_fill_2 FILLER_63_59 ();
 sg13g2_fill_2 FILLER_63_76 ();
 sg13g2_fill_1 FILLER_63_78 ();
 sg13g2_fill_2 FILLER_63_103 ();
 sg13g2_fill_1 FILLER_63_105 ();
 sg13g2_fill_1 FILLER_63_125 ();
 sg13g2_decap_4 FILLER_63_131 ();
 sg13g2_fill_1 FILLER_63_135 ();
 sg13g2_fill_1 FILLER_63_169 ();
 sg13g2_fill_1 FILLER_63_199 ();
 sg13g2_decap_4 FILLER_63_218 ();
 sg13g2_fill_1 FILLER_63_244 ();
 sg13g2_decap_8 FILLER_63_283 ();
 sg13g2_decap_4 FILLER_63_290 ();
 sg13g2_fill_1 FILLER_63_294 ();
 sg13g2_fill_2 FILLER_63_314 ();
 sg13g2_fill_1 FILLER_63_339 ();
 sg13g2_fill_1 FILLER_63_364 ();
 sg13g2_fill_2 FILLER_63_388 ();
 sg13g2_fill_1 FILLER_63_390 ();
 sg13g2_fill_1 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_60 ();
 sg13g2_fill_1 FILLER_64_62 ();
 sg13g2_fill_1 FILLER_64_108 ();
 sg13g2_decap_4 FILLER_64_118 ();
 sg13g2_fill_2 FILLER_64_163 ();
 sg13g2_fill_2 FILLER_64_188 ();
 sg13g2_fill_1 FILLER_64_228 ();
 sg13g2_fill_1 FILLER_64_277 ();
 sg13g2_decap_8 FILLER_64_287 ();
 sg13g2_decap_8 FILLER_64_294 ();
 sg13g2_decap_8 FILLER_64_301 ();
 sg13g2_decap_4 FILLER_64_312 ();
 sg13g2_fill_1 FILLER_64_316 ();
 sg13g2_fill_2 FILLER_64_322 ();
 sg13g2_fill_1 FILLER_64_329 ();
 sg13g2_fill_1 FILLER_64_360 ();
 sg13g2_decap_4 FILLER_64_379 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_22 ();
 sg13g2_decap_4 FILLER_65_30 ();
 sg13g2_fill_1 FILLER_65_83 ();
 sg13g2_fill_2 FILLER_65_92 ();
 sg13g2_fill_1 FILLER_65_94 ();
 sg13g2_fill_2 FILLER_65_122 ();
 sg13g2_decap_4 FILLER_65_137 ();
 sg13g2_fill_2 FILLER_65_175 ();
 sg13g2_fill_1 FILLER_65_177 ();
 sg13g2_fill_1 FILLER_65_183 ();
 sg13g2_decap_4 FILLER_65_196 ();
 sg13g2_fill_1 FILLER_65_200 ();
 sg13g2_fill_1 FILLER_65_217 ();
 sg13g2_fill_2 FILLER_65_229 ();
 sg13g2_fill_1 FILLER_65_231 ();
 sg13g2_decap_8 FILLER_65_244 ();
 sg13g2_decap_8 FILLER_65_251 ();
 sg13g2_decap_8 FILLER_65_258 ();
 sg13g2_decap_4 FILLER_65_265 ();
 sg13g2_fill_2 FILLER_65_301 ();
 sg13g2_fill_1 FILLER_65_320 ();
 sg13g2_fill_1 FILLER_65_326 ();
 sg13g2_fill_1 FILLER_65_332 ();
 sg13g2_fill_1 FILLER_65_346 ();
 sg13g2_fill_1 FILLER_65_370 ();
 sg13g2_fill_1 FILLER_65_383 ();
 sg13g2_decap_8 FILLER_65_398 ();
 sg13g2_decap_4 FILLER_65_405 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_25 ();
 sg13g2_fill_1 FILLER_66_47 ();
 sg13g2_fill_2 FILLER_66_72 ();
 sg13g2_fill_2 FILLER_66_82 ();
 sg13g2_decap_4 FILLER_66_88 ();
 sg13g2_fill_2 FILLER_66_126 ();
 sg13g2_fill_1 FILLER_66_128 ();
 sg13g2_decap_8 FILLER_66_145 ();
 sg13g2_fill_1 FILLER_66_152 ();
 sg13g2_decap_8 FILLER_66_202 ();
 sg13g2_decap_8 FILLER_66_209 ();
 sg13g2_fill_2 FILLER_66_220 ();
 sg13g2_fill_1 FILLER_66_242 ();
 sg13g2_fill_2 FILLER_66_256 ();
 sg13g2_fill_1 FILLER_66_278 ();
 sg13g2_fill_2 FILLER_66_325 ();
 sg13g2_fill_2 FILLER_66_332 ();
 sg13g2_fill_1 FILLER_66_334 ();
 sg13g2_fill_1 FILLER_66_361 ();
 sg13g2_decap_4 FILLER_66_367 ();
 sg13g2_fill_2 FILLER_66_381 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_2 ();
 sg13g2_decap_4 FILLER_67_27 ();
 sg13g2_fill_2 FILLER_67_31 ();
 sg13g2_fill_2 FILLER_67_41 ();
 sg13g2_fill_1 FILLER_67_43 ();
 sg13g2_fill_2 FILLER_67_49 ();
 sg13g2_fill_1 FILLER_67_51 ();
 sg13g2_fill_2 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_67 ();
 sg13g2_decap_8 FILLER_67_74 ();
 sg13g2_fill_1 FILLER_67_81 ();
 sg13g2_decap_8 FILLER_67_87 ();
 sg13g2_decap_4 FILLER_67_94 ();
 sg13g2_decap_4 FILLER_67_106 ();
 sg13g2_decap_4 FILLER_67_121 ();
 sg13g2_fill_2 FILLER_67_144 ();
 sg13g2_fill_2 FILLER_67_163 ();
 sg13g2_fill_1 FILLER_67_165 ();
 sg13g2_fill_2 FILLER_67_178 ();
 sg13g2_fill_1 FILLER_67_180 ();
 sg13g2_fill_2 FILLER_67_187 ();
 sg13g2_decap_4 FILLER_67_193 ();
 sg13g2_fill_1 FILLER_67_210 ();
 sg13g2_decap_4 FILLER_67_214 ();
 sg13g2_fill_1 FILLER_67_218 ();
 sg13g2_fill_1 FILLER_67_244 ();
 sg13g2_decap_4 FILLER_67_282 ();
 sg13g2_fill_2 FILLER_67_286 ();
 sg13g2_fill_1 FILLER_67_335 ();
 sg13g2_fill_2 FILLER_67_341 ();
 sg13g2_fill_1 FILLER_67_343 ();
 sg13g2_fill_2 FILLER_67_361 ();
 sg13g2_fill_1 FILLER_67_363 ();
 sg13g2_fill_1 FILLER_67_389 ();
 sg13g2_fill_2 FILLER_67_406 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_7 ();
 sg13g2_fill_2 FILLER_68_12 ();
 sg13g2_fill_2 FILLER_68_26 ();
 sg13g2_fill_1 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_55 ();
 sg13g2_decap_8 FILLER_68_62 ();
 sg13g2_decap_8 FILLER_68_69 ();
 sg13g2_fill_1 FILLER_68_76 ();
 sg13g2_decap_4 FILLER_68_95 ();
 sg13g2_fill_1 FILLER_68_116 ();
 sg13g2_decap_4 FILLER_68_144 ();
 sg13g2_fill_2 FILLER_68_153 ();
 sg13g2_fill_2 FILLER_68_164 ();
 sg13g2_fill_1 FILLER_68_166 ();
 sg13g2_fill_1 FILLER_68_175 ();
 sg13g2_fill_1 FILLER_68_210 ();
 sg13g2_fill_1 FILLER_68_215 ();
 sg13g2_fill_2 FILLER_68_223 ();
 sg13g2_decap_8 FILLER_68_282 ();
 sg13g2_fill_2 FILLER_68_306 ();
 sg13g2_fill_1 FILLER_68_339 ();
 sg13g2_fill_2 FILLER_68_361 ();
 sg13g2_fill_2 FILLER_68_375 ();
 sg13g2_decap_4 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_40 ();
 sg13g2_fill_2 FILLER_69_51 ();
 sg13g2_fill_1 FILLER_69_53 ();
 sg13g2_decap_4 FILLER_69_67 ();
 sg13g2_decap_4 FILLER_69_85 ();
 sg13g2_fill_2 FILLER_69_97 ();
 sg13g2_fill_1 FILLER_69_132 ();
 sg13g2_fill_2 FILLER_69_146 ();
 sg13g2_fill_2 FILLER_69_228 ();
 sg13g2_fill_2 FILLER_69_248 ();
 sg13g2_fill_1 FILLER_69_258 ();
 sg13g2_fill_2 FILLER_69_277 ();
 sg13g2_fill_2 FILLER_69_285 ();
 sg13g2_fill_1 FILLER_69_287 ();
 sg13g2_fill_1 FILLER_69_336 ();
 sg13g2_fill_1 FILLER_69_361 ();
 sg13g2_fill_1 FILLER_69_376 ();
 sg13g2_fill_1 FILLER_69_382 ();
 sg13g2_fill_2 FILLER_70_20 ();
 sg13g2_fill_1 FILLER_70_37 ();
 sg13g2_fill_2 FILLER_70_78 ();
 sg13g2_fill_1 FILLER_70_80 ();
 sg13g2_fill_1 FILLER_70_96 ();
 sg13g2_fill_2 FILLER_70_115 ();
 sg13g2_fill_1 FILLER_70_117 ();
 sg13g2_fill_2 FILLER_70_135 ();
 sg13g2_fill_2 FILLER_70_165 ();
 sg13g2_fill_1 FILLER_70_167 ();
 sg13g2_fill_2 FILLER_70_191 ();
 sg13g2_fill_1 FILLER_70_205 ();
 sg13g2_decap_4 FILLER_70_214 ();
 sg13g2_fill_2 FILLER_70_232 ();
 sg13g2_fill_1 FILLER_70_234 ();
 sg13g2_decap_4 FILLER_70_239 ();
 sg13g2_fill_2 FILLER_70_247 ();
 sg13g2_fill_1 FILLER_70_254 ();
 sg13g2_fill_1 FILLER_70_314 ();
 sg13g2_fill_2 FILLER_70_343 ();
 sg13g2_fill_1 FILLER_70_351 ();
 sg13g2_fill_1 FILLER_70_361 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_decap_4 FILLER_71_40 ();
 sg13g2_fill_2 FILLER_71_44 ();
 sg13g2_fill_1 FILLER_71_55 ();
 sg13g2_fill_1 FILLER_71_90 ();
 sg13g2_fill_2 FILLER_71_94 ();
 sg13g2_fill_2 FILLER_71_118 ();
 sg13g2_fill_1 FILLER_71_120 ();
 sg13g2_fill_2 FILLER_71_126 ();
 sg13g2_fill_1 FILLER_71_175 ();
 sg13g2_fill_1 FILLER_71_209 ();
 sg13g2_fill_2 FILLER_71_215 ();
 sg13g2_fill_1 FILLER_71_222 ();
 sg13g2_fill_1 FILLER_71_240 ();
 sg13g2_decap_8 FILLER_71_249 ();
 sg13g2_decap_4 FILLER_71_260 ();
 sg13g2_fill_2 FILLER_71_264 ();
 sg13g2_fill_1 FILLER_71_284 ();
 sg13g2_fill_2 FILLER_71_317 ();
 sg13g2_fill_2 FILLER_71_324 ();
 sg13g2_decap_4 FILLER_71_336 ();
 sg13g2_fill_2 FILLER_71_340 ();
 sg13g2_fill_2 FILLER_71_366 ();
 sg13g2_fill_2 FILLER_71_391 ();
 sg13g2_fill_1 FILLER_71_393 ();
 sg13g2_fill_2 FILLER_71_406 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_fill_2 FILLER_72_43 ();
 sg13g2_fill_1 FILLER_72_45 ();
 sg13g2_fill_1 FILLER_72_59 ();
 sg13g2_fill_2 FILLER_72_99 ();
 sg13g2_fill_1 FILLER_72_101 ();
 sg13g2_decap_8 FILLER_72_116 ();
 sg13g2_fill_2 FILLER_72_141 ();
 sg13g2_fill_1 FILLER_72_143 ();
 sg13g2_fill_1 FILLER_72_228 ();
 sg13g2_fill_1 FILLER_72_257 ();
 sg13g2_decap_8 FILLER_72_266 ();
 sg13g2_decap_4 FILLER_72_273 ();
 sg13g2_fill_1 FILLER_72_277 ();
 sg13g2_fill_2 FILLER_72_340 ();
 sg13g2_fill_1 FILLER_72_342 ();
 sg13g2_decap_4 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_4 ();
 sg13g2_fill_1 FILLER_73_16 ();
 sg13g2_fill_1 FILLER_73_27 ();
 sg13g2_decap_4 FILLER_73_33 ();
 sg13g2_fill_1 FILLER_73_37 ();
 sg13g2_fill_2 FILLER_73_68 ();
 sg13g2_fill_2 FILLER_73_75 ();
 sg13g2_fill_1 FILLER_73_116 ();
 sg13g2_decap_4 FILLER_73_137 ();
 sg13g2_fill_1 FILLER_73_145 ();
 sg13g2_fill_2 FILLER_73_169 ();
 sg13g2_fill_2 FILLER_73_179 ();
 sg13g2_fill_1 FILLER_73_181 ();
 sg13g2_fill_1 FILLER_73_238 ();
 sg13g2_decap_8 FILLER_73_270 ();
 sg13g2_decap_4 FILLER_73_277 ();
 sg13g2_fill_1 FILLER_73_281 ();
 sg13g2_fill_2 FILLER_73_286 ();
 sg13g2_fill_1 FILLER_73_288 ();
 sg13g2_fill_2 FILLER_73_293 ();
 sg13g2_fill_1 FILLER_73_295 ();
 sg13g2_fill_1 FILLER_73_312 ();
 sg13g2_fill_2 FILLER_73_319 ();
 sg13g2_fill_2 FILLER_73_355 ();
 sg13g2_fill_1 FILLER_73_369 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_4 FILLER_74_28 ();
 sg13g2_fill_2 FILLER_74_32 ();
 sg13g2_fill_1 FILLER_74_53 ();
 sg13g2_fill_1 FILLER_74_60 ();
 sg13g2_fill_2 FILLER_74_97 ();
 sg13g2_fill_1 FILLER_74_123 ();
 sg13g2_fill_1 FILLER_74_151 ();
 sg13g2_fill_2 FILLER_74_174 ();
 sg13g2_fill_1 FILLER_74_176 ();
 sg13g2_fill_1 FILLER_74_208 ();
 sg13g2_decap_8 FILLER_74_254 ();
 sg13g2_fill_1 FILLER_74_261 ();
 sg13g2_fill_1 FILLER_74_271 ();
 sg13g2_fill_2 FILLER_74_286 ();
 sg13g2_fill_1 FILLER_74_288 ();
 sg13g2_fill_2 FILLER_74_298 ();
 sg13g2_fill_1 FILLER_74_300 ();
 sg13g2_fill_1 FILLER_74_315 ();
 sg13g2_fill_2 FILLER_74_327 ();
 sg13g2_fill_2 FILLER_74_341 ();
 sg13g2_fill_1 FILLER_74_343 ();
 sg13g2_fill_2 FILLER_74_360 ();
 sg13g2_fill_2 FILLER_74_393 ();
 sg13g2_fill_1 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_27 ();
 sg13g2_decap_8 FILLER_75_34 ();
 sg13g2_fill_1 FILLER_75_75 ();
 sg13g2_fill_2 FILLER_75_85 ();
 sg13g2_fill_1 FILLER_75_87 ();
 sg13g2_fill_1 FILLER_75_182 ();
 sg13g2_fill_2 FILLER_75_189 ();
 sg13g2_fill_1 FILLER_75_200 ();
 sg13g2_fill_1 FILLER_75_209 ();
 sg13g2_decap_4 FILLER_75_244 ();
 sg13g2_fill_2 FILLER_75_248 ();
 sg13g2_fill_2 FILLER_75_262 ();
 sg13g2_fill_1 FILLER_75_283 ();
 sg13g2_fill_1 FILLER_75_316 ();
 sg13g2_fill_2 FILLER_75_338 ();
 sg13g2_fill_1 FILLER_75_340 ();
 sg13g2_fill_2 FILLER_75_346 ();
 sg13g2_fill_2 FILLER_75_366 ();
 sg13g2_fill_2 FILLER_75_388 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_7 ();
 sg13g2_fill_1 FILLER_76_9 ();
 sg13g2_fill_2 FILLER_76_45 ();
 sg13g2_fill_1 FILLER_76_70 ();
 sg13g2_fill_2 FILLER_76_79 ();
 sg13g2_fill_1 FILLER_76_96 ();
 sg13g2_fill_1 FILLER_76_120 ();
 sg13g2_decap_8 FILLER_76_212 ();
 sg13g2_fill_2 FILLER_76_219 ();
 sg13g2_decap_4 FILLER_76_229 ();
 sg13g2_decap_4 FILLER_76_237 ();
 sg13g2_fill_1 FILLER_76_241 ();
 sg13g2_fill_2 FILLER_76_299 ();
 sg13g2_fill_2 FILLER_76_329 ();
 sg13g2_fill_1 FILLER_76_331 ();
 sg13g2_fill_2 FILLER_76_342 ();
 sg13g2_fill_1 FILLER_76_375 ();
 sg13g2_fill_2 FILLER_76_383 ();
 sg13g2_fill_2 FILLER_76_394 ();
 sg13g2_fill_1 FILLER_76_396 ();
 sg13g2_fill_2 FILLER_77_0 ();
 sg13g2_decap_4 FILLER_77_32 ();
 sg13g2_decap_4 FILLER_77_39 ();
 sg13g2_fill_2 FILLER_77_58 ();
 sg13g2_fill_1 FILLER_77_60 ();
 sg13g2_fill_1 FILLER_77_71 ();
 sg13g2_fill_2 FILLER_77_172 ();
 sg13g2_fill_1 FILLER_77_174 ();
 sg13g2_fill_1 FILLER_77_216 ();
 sg13g2_fill_2 FILLER_77_234 ();
 sg13g2_fill_1 FILLER_77_236 ();
 sg13g2_fill_1 FILLER_77_245 ();
 sg13g2_fill_1 FILLER_77_281 ();
 sg13g2_fill_2 FILLER_77_348 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_27 ();
 sg13g2_fill_1 FILLER_78_33 ();
 sg13g2_fill_2 FILLER_78_60 ();
 sg13g2_fill_2 FILLER_78_75 ();
 sg13g2_fill_1 FILLER_78_77 ();
 sg13g2_fill_1 FILLER_78_93 ();
 sg13g2_fill_2 FILLER_78_113 ();
 sg13g2_fill_1 FILLER_78_146 ();
 sg13g2_fill_2 FILLER_78_157 ();
 sg13g2_fill_1 FILLER_78_159 ();
 sg13g2_fill_1 FILLER_78_196 ();
 sg13g2_fill_2 FILLER_78_254 ();
 sg13g2_fill_2 FILLER_78_277 ();
 sg13g2_fill_1 FILLER_78_279 ();
 sg13g2_fill_2 FILLER_78_304 ();
 sg13g2_fill_1 FILLER_78_382 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_4 FILLER_79_7 ();
 sg13g2_fill_2 FILLER_79_11 ();
 sg13g2_fill_2 FILLER_79_21 ();
 sg13g2_fill_1 FILLER_79_23 ();
 sg13g2_decap_4 FILLER_79_29 ();
 sg13g2_decap_4 FILLER_79_84 ();
 sg13g2_fill_2 FILLER_79_98 ();
 sg13g2_fill_1 FILLER_79_100 ();
 sg13g2_fill_2 FILLER_79_127 ();
 sg13g2_fill_1 FILLER_79_129 ();
 sg13g2_fill_2 FILLER_79_161 ();
 sg13g2_fill_2 FILLER_79_187 ();
 sg13g2_fill_1 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_235 ();
 sg13g2_fill_2 FILLER_79_247 ();
 sg13g2_fill_1 FILLER_79_249 ();
 sg13g2_fill_1 FILLER_79_268 ();
 sg13g2_fill_2 FILLER_79_279 ();
 sg13g2_fill_1 FILLER_79_281 ();
 sg13g2_fill_1 FILLER_79_290 ();
 sg13g2_fill_1 FILLER_79_312 ();
 sg13g2_fill_2 FILLER_79_347 ();
 sg13g2_fill_1 FILLER_79_349 ();
 sg13g2_fill_2 FILLER_79_381 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_4 FILLER_80_28 ();
 sg13g2_fill_2 FILLER_80_32 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_fill_1 FILLER_80_120 ();
 sg13g2_fill_1 FILLER_80_134 ();
 sg13g2_fill_2 FILLER_80_184 ();
 sg13g2_decap_8 FILLER_80_190 ();
 sg13g2_decap_8 FILLER_80_197 ();
 sg13g2_fill_1 FILLER_80_204 ();
 sg13g2_fill_1 FILLER_80_218 ();
 sg13g2_decap_8 FILLER_80_232 ();
 sg13g2_decap_8 FILLER_80_239 ();
 sg13g2_decap_8 FILLER_80_246 ();
 sg13g2_decap_4 FILLER_80_253 ();
 sg13g2_fill_2 FILLER_80_261 ();
 sg13g2_fill_1 FILLER_80_263 ();
 sg13g2_fill_2 FILLER_80_290 ();
 sg13g2_fill_1 FILLER_80_331 ();
 sg13g2_fill_2 FILLER_80_344 ();
 sg13g2_fill_1 FILLER_80_373 ();
 sg13g2_fill_1 FILLER_80_383 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net205;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[2] = net18;
 assign uio_out[3] = net19;
 assign uio_out[4] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
endmodule

module tt_um_rkarl_Spiral (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire clknet_0_clk;
 wire \angleOffset[0] ;
 wire \angleOffset[1] ;
 wire \angleOffset[2] ;
 wire \angleOffset[3] ;
 wire \angleOffset[4] ;
 wire \angle[0] ;
 wire \angle[1] ;
 wire \angle[2] ;
 wire \angle[3] ;
 wire \cordicAlg.ph[1][1] ;
 wire \cordicAlg.ph[1][2] ;
 wire \cordicAlg.ph[1][3] ;
 wire \cordicAlg.ph[2][1] ;
 wire \cordicAlg.ph[2][2] ;
 wire \cordicAlg.ph[2][3] ;
 wire \cordicAlg.ph[3][0] ;
 wire \cordicAlg.ph[3][1] ;
 wire \cordicAlg.ph[3][2] ;
 wire \cordicAlg.ph[3][3] ;
 wire \cordicAlg.xv[0][1] ;
 wire \cordicAlg.xv[0][2] ;
 wire \cordicAlg.xv[0][3] ;
 wire \cordicAlg.xv[0][4] ;
 wire \cordicAlg.xv[0][5] ;
 wire \cordicAlg.xv[0][6] ;
 wire \cordicAlg.yv[0][0] ;
 wire \cordicAlg.yv[0][1] ;
 wire \cordicAlg.yv[0][2] ;
 wire \cordicAlg.yv[0][3] ;
 wire \cordicAlg.yv[0][4] ;
 wire \cordicAlg.yv[0][5] ;
 wire \cordicAlg.yv[0][6] ;
 wire \cordicAlg.yv[1][6] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \hypotenuse.multSignal[0] ;
 wire \hypotenuse.multX[10] ;
 wire \hypotenuse.multX[11] ;
 wire \hypotenuse.multX[12] ;
 wire \hypotenuse.multX[2] ;
 wire \hypotenuse.multX[3] ;
 wire \hypotenuse.multX[4] ;
 wire \hypotenuse.multX[5] ;
 wire \hypotenuse.multX[6] ;
 wire \hypotenuse.multX[7] ;
 wire \hypotenuse.multX[8] ;
 wire \hypotenuse.multX[9] ;
 wire \hypotenuse.multY[10] ;
 wire \hypotenuse.multY[11] ;
 wire \hypotenuse.multY[12] ;
 wire \hypotenuse.multY[2] ;
 wire \hypotenuse.multY[3] ;
 wire \hypotenuse.multY[4] ;
 wire \hypotenuse.multY[5] ;
 wire \hypotenuse.multY[6] ;
 wire \hypotenuse.multY[7] ;
 wire \hypotenuse.multY[8] ;
 wire \hypotenuse.multY[9] ;
 wire \hypotenuse.mutlReg[1] ;
 wire \hypotenuse.mutlReg[2] ;
 wire \hypotenuse.mutlReg[3] ;
 wire \hypotenuse.mutlReg[4] ;
 wire \hypotenuse.mutlReg[5] ;
 wire \hypotenuse.mutlReg[6] ;
 wire \hypotenuse.stateCheck ;
 wire \hypotenuse.x_pos[0] ;
 wire \hypotenuse.y_pos[0] ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;

 sg13g2_inv_1 _0917_ (.Y(_0105_),
    .A(net152));
 sg13g2_inv_1 _0918_ (.Y(_0106_),
    .A(net215));
 sg13g2_inv_1 _0919_ (.Y(_0107_),
    .A(net229));
 sg13g2_inv_1 _0920_ (.Y(_0108_),
    .A(net206));
 sg13g2_inv_1 _0921_ (.Y(_0109_),
    .A(net148));
 sg13g2_inv_1 _0922_ (.Y(_0110_),
    .A(\hypotenuse.multX[5] ));
 sg13g2_inv_1 _0923_ (.Y(_0111_),
    .A(\hypotenuse.multY[5] ));
 sg13g2_inv_1 _0924_ (.Y(_0112_),
    .A(net203));
 sg13g2_inv_1 _0925_ (.Y(_0113_),
    .A(_0012_));
 sg13g2_inv_1 _0926_ (.Y(_0114_),
    .A(_0014_));
 sg13g2_inv_1 _0927_ (.Y(_0115_),
    .A(net145));
 sg13g2_and2_1 _0928_ (.A(\hvsync_gen.vpos[0] ),
    .B(\hvsync_gen.vpos[1] ),
    .X(_0116_));
 sg13g2_nand2_1 _0929_ (.Y(_0117_),
    .A(\hvsync_gen.vpos[0] ),
    .B(\hvsync_gen.vpos[1] ));
 sg13g2_nor3_1 _0930_ (.A(\hvsync_gen.vpos[3] ),
    .B(\hvsync_gen.vpos[2] ),
    .C(_0116_),
    .Y(_0118_));
 sg13g2_nor2b_1 _0931_ (.A(_0118_),
    .B_N(\hvsync_gen.vpos[4] ),
    .Y(_0119_));
 sg13g2_and2_1 _0932_ (.A(\hvsync_gen.vpos[5] ),
    .B(_0119_),
    .X(_0120_));
 sg13g2_nand3_1 _0933_ (.B(\hvsync_gen.vpos[6] ),
    .C(\hvsync_gen.vpos[5] ),
    .A(\hvsync_gen.vpos[7] ),
    .Y(_0121_));
 sg13g2_and3_1 _0934_ (.X(_0122_),
    .A(\hvsync_gen.vpos[7] ),
    .B(\hvsync_gen.vpos[6] ),
    .C(_0120_));
 sg13g2_nand2b_1 _0935_ (.Y(_0123_),
    .B(_0005_),
    .A_N(_0122_));
 sg13g2_xnor2_1 _0936_ (.Y(_0124_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_0123_));
 sg13g2_xor2_1 _0937_ (.B(_0123_),
    .A(\hvsync_gen.vpos[9] ),
    .X(_0125_));
 sg13g2_and2_1 _0938_ (.A(\hvsync_gen.hpos[0] ),
    .B(net190),
    .X(_0126_));
 sg13g2_a21oi_2 _0939_ (.B1(\hvsync_gen.hpos[2] ),
    .Y(_0127_),
    .A2(\hvsync_gen.hpos[1] ),
    .A1(\hvsync_gen.hpos[0] ));
 sg13g2_nand2b_2 _0940_ (.Y(_0128_),
    .B(_0127_),
    .A_N(\hvsync_gen.hpos[3] ));
 sg13g2_nor3_2 _0941_ (.A(\hvsync_gen.hpos[4] ),
    .B(\hvsync_gen.hpos[5] ),
    .C(_0128_),
    .Y(_0129_));
 sg13g2_nand2b_1 _0942_ (.Y(_0130_),
    .B(\hvsync_gen.hpos[6] ),
    .A_N(_0129_));
 sg13g2_o21ai_1 _0943_ (.B1(_0006_),
    .Y(_0131_),
    .A1(\hvsync_gen.hpos[7] ),
    .A2(_0130_));
 sg13g2_nand2_1 _0944_ (.Y(_0132_),
    .A(\hvsync_gen.hpos[8] ),
    .B(_0131_));
 sg13g2_xnor2_1 _0945_ (.Y(_0133_),
    .A(\hvsync_gen.hpos[9] ),
    .B(_0132_));
 sg13g2_xor2_1 _0946_ (.B(_0132_),
    .A(\hvsync_gen.hpos[9] ),
    .X(_0134_));
 sg13g2_nor2_2 _0947_ (.A(_0125_),
    .B(net126),
    .Y(_0135_));
 sg13g2_nand2_2 _0948_ (.Y(_0136_),
    .A(net128),
    .B(net125));
 sg13g2_nor2_1 _0949_ (.A(net128),
    .B(net124),
    .Y(_0137_));
 sg13g2_nand2_1 _0950_ (.Y(_0138_),
    .A(_0125_),
    .B(_0133_));
 sg13g2_nand2_1 _0951_ (.Y(_0139_),
    .A(_0136_),
    .B(net118));
 sg13g2_nor2_1 _0952_ (.A(net149),
    .B(_0139_),
    .Y(_0000_));
 sg13g2_or2_1 _0953_ (.X(_0140_),
    .B(_0121_),
    .A(_0106_));
 sg13g2_nand2b_1 _0954_ (.Y(_0141_),
    .B(net228),
    .A_N(\hvsync_gen.vpos[4] ));
 sg13g2_nor4_1 _0955_ (.A(net199),
    .B(_0108_),
    .C(net233),
    .D(_0141_),
    .Y(_0142_));
 sg13g2_nor2b_2 _0956_ (.A(_0140_),
    .B_N(_0142_),
    .Y(_0004_));
 sg13g2_nand4_1 _0957_ (.B(net147),
    .C(\hvsync_gen.hpos[4] ),
    .A(\hvsync_gen.hpos[7] ),
    .Y(_0143_),
    .D(\hvsync_gen.hpos[5] ));
 sg13g2_nor2b_1 _0958_ (.A(\hvsync_gen.hpos[8] ),
    .B_N(\hvsync_gen.hpos[9] ),
    .Y(_0144_));
 sg13g2_a21oi_1 _0959_ (.A1(_0143_),
    .A2(_0144_),
    .Y(_0145_),
    .B1(net116));
 sg13g2_nand2_1 _0960_ (.Y(_0146_),
    .A(\hvsync_gen.hpos[8] ),
    .B(\hvsync_gen.hpos[9] ));
 sg13g2_or3_1 _0961_ (.A(net147),
    .B(\hvsync_gen.hpos[4] ),
    .C(\hvsync_gen.hpos[5] ),
    .X(_0147_));
 sg13g2_nand3_1 _0962_ (.B(\hvsync_gen.hpos[9] ),
    .C(_0147_),
    .A(\hvsync_gen.hpos[7] ),
    .Y(_0148_));
 sg13g2_a21oi_1 _0963_ (.A1(_0146_),
    .A2(_0148_),
    .Y(_0003_),
    .B1(net117));
 sg13g2_and2_1 _0964_ (.A(\hypotenuse.multX[11] ),
    .B(\hypotenuse.multY[11] ),
    .X(_0149_));
 sg13g2_nand2_1 _0965_ (.Y(_0150_),
    .A(\hypotenuse.multX[11] ),
    .B(\hypotenuse.multY[11] ));
 sg13g2_xnor2_1 _0966_ (.Y(_0151_),
    .A(\hypotenuse.multX[11] ),
    .B(\hypotenuse.multY[11] ));
 sg13g2_nand2_2 _0967_ (.Y(_0152_),
    .A(\hypotenuse.multX[10] ),
    .B(\hypotenuse.multY[10] ));
 sg13g2_and2_1 _0968_ (.A(\hypotenuse.multX[9] ),
    .B(\hypotenuse.multY[9] ),
    .X(_0153_));
 sg13g2_nand2_1 _0969_ (.Y(_0154_),
    .A(\hypotenuse.multX[9] ),
    .B(\hypotenuse.multY[9] ));
 sg13g2_and2_1 _0970_ (.A(\hypotenuse.multX[8] ),
    .B(\hypotenuse.multY[8] ),
    .X(_0155_));
 sg13g2_nand2_1 _0971_ (.Y(_0156_),
    .A(\hypotenuse.multX[8] ),
    .B(\hypotenuse.multY[8] ));
 sg13g2_nand2_1 _0972_ (.Y(_0157_),
    .A(\hypotenuse.multX[7] ),
    .B(\hypotenuse.multY[7] ));
 sg13g2_and2_1 _0973_ (.A(\hypotenuse.multX[6] ),
    .B(\hypotenuse.multY[6] ),
    .X(_0158_));
 sg13g2_a22oi_1 _0974_ (.Y(_0159_),
    .B1(\hypotenuse.multX[2] ),
    .B2(\hypotenuse.multY[2] ),
    .A2(\hypotenuse.multY[3] ),
    .A1(\hypotenuse.multX[3] ));
 sg13g2_nor2_1 _0975_ (.A(\hypotenuse.multX[4] ),
    .B(\hypotenuse.multY[4] ),
    .Y(_0160_));
 sg13g2_nor2_1 _0976_ (.A(\hypotenuse.multX[3] ),
    .B(\hypotenuse.multY[3] ),
    .Y(_0161_));
 sg13g2_or3_1 _0977_ (.A(_0159_),
    .B(_0160_),
    .C(_0161_),
    .X(_0162_));
 sg13g2_a22oi_1 _0978_ (.Y(_0163_),
    .B1(\hypotenuse.multX[4] ),
    .B2(\hypotenuse.multY[4] ),
    .A2(\hypotenuse.multY[5] ),
    .A1(\hypotenuse.multX[5] ));
 sg13g2_a22oi_1 _0979_ (.Y(_0164_),
    .B1(_0162_),
    .B2(_0163_),
    .A2(_0111_),
    .A1(_0110_));
 sg13g2_xnor2_1 _0980_ (.Y(_0165_),
    .A(\hypotenuse.multX[6] ),
    .B(\hypotenuse.multY[6] ));
 sg13g2_a221oi_1 _0981_ (.B2(_0163_),
    .C1(_0165_),
    .B1(_0162_),
    .A1(_0110_),
    .Y(_0166_),
    .A2(_0111_));
 sg13g2_xor2_1 _0982_ (.B(\hypotenuse.multY[7] ),
    .A(\hypotenuse.multX[7] ),
    .X(_0167_));
 sg13g2_o21ai_1 _0983_ (.B1(_0167_),
    .Y(_0168_),
    .A1(_0158_),
    .A2(_0166_));
 sg13g2_xnor2_1 _0984_ (.Y(_0169_),
    .A(\hypotenuse.multX[8] ),
    .B(\hypotenuse.multY[8] ));
 sg13g2_a21oi_2 _0985_ (.B1(_0169_),
    .Y(_0170_),
    .A2(_0168_),
    .A1(_0157_));
 sg13g2_a21o_1 _0986_ (.A2(_0168_),
    .A1(_0157_),
    .B1(_0169_),
    .X(_0171_));
 sg13g2_xor2_1 _0987_ (.B(\hypotenuse.multY[9] ),
    .A(\hypotenuse.multX[9] ),
    .X(_0172_));
 sg13g2_xnor2_1 _0988_ (.Y(_0173_),
    .A(\hypotenuse.multX[9] ),
    .B(\hypotenuse.multY[9] ));
 sg13g2_a21oi_2 _0989_ (.B1(_0173_),
    .Y(_0174_),
    .A2(_0171_),
    .A1(_0156_));
 sg13g2_o21ai_1 _0990_ (.B1(_0172_),
    .Y(_0175_),
    .A1(_0155_),
    .A2(_0170_));
 sg13g2_xor2_1 _0991_ (.B(\hypotenuse.multY[10] ),
    .A(\hypotenuse.multX[10] ),
    .X(_0176_));
 sg13g2_xnor2_1 _0992_ (.Y(_0177_),
    .A(\hypotenuse.multX[10] ),
    .B(\hypotenuse.multY[10] ));
 sg13g2_o21ai_1 _0993_ (.B1(_0176_),
    .Y(_0178_),
    .A1(_0153_),
    .A2(_0174_));
 sg13g2_a21oi_2 _0994_ (.B1(_0151_),
    .Y(_0179_),
    .A2(net123),
    .A1(_0152_));
 sg13g2_a21o_2 _0995_ (.A2(net123),
    .A1(_0152_),
    .B1(_0151_),
    .X(_0180_));
 sg13g2_and3_1 _0996_ (.X(_0181_),
    .A(_0151_),
    .B(_0152_),
    .C(net123));
 sg13g2_nand3_1 _0997_ (.B(_0152_),
    .C(net123),
    .A(_0151_),
    .Y(_0182_));
 sg13g2_nor2_1 _0998_ (.A(_0179_),
    .B(_0181_),
    .Y(_0183_));
 sg13g2_nand2_2 _0999_ (.Y(_0184_),
    .A(_0180_),
    .B(_0182_));
 sg13g2_nand3_1 _1000_ (.B(net129),
    .C(_0177_),
    .A(_0154_),
    .Y(_0185_));
 sg13g2_nand3_1 _1001_ (.B(net129),
    .C(_0176_),
    .A(_0154_),
    .Y(_0186_));
 sg13g2_o21ai_1 _1002_ (.B1(_0177_),
    .Y(_0187_),
    .A1(_0153_),
    .A2(_0174_));
 sg13g2_nand2_2 _1003_ (.Y(_0188_),
    .A(_0186_),
    .B(_0187_));
 sg13g2_nand2_2 _1004_ (.Y(_0189_),
    .A(net122),
    .B(_0185_));
 sg13g2_nor3_2 _1005_ (.A(_0155_),
    .B(_0170_),
    .C(_0172_),
    .Y(_0190_));
 sg13g2_nand3_1 _1006_ (.B(_0171_),
    .C(_0173_),
    .A(_0156_),
    .Y(_0191_));
 sg13g2_nor2_2 _1007_ (.A(_0174_),
    .B(_0190_),
    .Y(_0192_));
 sg13g2_and3_2 _1008_ (.X(_0193_),
    .A(_0157_),
    .B(_0168_),
    .C(_0169_));
 sg13g2_nor2_2 _1009_ (.A(_0170_),
    .B(_0193_),
    .Y(_0194_));
 sg13g2_or2_2 _1010_ (.X(_0195_),
    .B(_0193_),
    .A(_0170_));
 sg13g2_xnor2_1 _1011_ (.Y(_0196_),
    .A(_0164_),
    .B(_0165_));
 sg13g2_inv_1 _1012_ (.Y(_0197_),
    .A(_0196_));
 sg13g2_or3_1 _1013_ (.A(_0158_),
    .B(_0166_),
    .C(_0167_),
    .X(_0198_));
 sg13g2_nand2_2 _1014_ (.Y(_0199_),
    .A(_0168_),
    .B(_0198_));
 sg13g2_nor2_1 _1015_ (.A(_0197_),
    .B(_0199_),
    .Y(_0200_));
 sg13g2_nand3_1 _1016_ (.B(_0196_),
    .C(_0198_),
    .A(_0168_),
    .Y(_0201_));
 sg13g2_o21ai_1 _1017_ (.B1(_0201_),
    .Y(_0202_),
    .A1(_0170_),
    .A2(_0193_));
 sg13g2_and4_1 _1018_ (.A(net123),
    .B(_0185_),
    .C(_0192_),
    .D(_0202_),
    .X(_0203_));
 sg13g2_nor3_2 _1019_ (.A(_0179_),
    .B(_0181_),
    .C(_0203_),
    .Y(_0204_));
 sg13g2_a21oi_2 _1020_ (.B1(_0194_),
    .Y(_0205_),
    .A2(_0191_),
    .A1(net129));
 sg13g2_a21oi_1 _1021_ (.A1(net129),
    .A2(_0191_),
    .Y(_0206_),
    .B1(_0202_));
 sg13g2_nor3_2 _1022_ (.A(_0174_),
    .B(_0190_),
    .C(_0195_),
    .Y(_0207_));
 sg13g2_a22oi_1 _1023_ (.Y(_0208_),
    .B1(_0200_),
    .B2(_0207_),
    .A2(net121),
    .A1(net122));
 sg13g2_nand2b_1 _1024_ (.Y(_0209_),
    .B(_0208_),
    .A_N(_0206_));
 sg13g2_xor2_1 _1025_ (.B(\hypotenuse.multY[12] ),
    .A(\hypotenuse.multX[12] ),
    .X(_0210_));
 sg13g2_xnor2_1 _1026_ (.Y(_0211_),
    .A(\hypotenuse.multX[12] ),
    .B(\hypotenuse.multY[12] ));
 sg13g2_a21oi_1 _1027_ (.A1(_0150_),
    .A2(_0180_),
    .Y(_0212_),
    .B1(_0210_));
 sg13g2_o21ai_1 _1028_ (.B1(_0211_),
    .Y(_0213_),
    .A1(_0149_),
    .A2(_0179_));
 sg13g2_nor3_1 _1029_ (.A(_0149_),
    .B(_0179_),
    .C(_0211_),
    .Y(_0214_));
 sg13g2_nand3_1 _1030_ (.B(_0180_),
    .C(_0210_),
    .A(_0150_),
    .Y(_0215_));
 sg13g2_nand2_2 _1031_ (.Y(_0216_),
    .A(_0213_),
    .B(_0215_));
 sg13g2_nand2_1 _1032_ (.Y(_0217_),
    .A(_0195_),
    .B(_0199_));
 sg13g2_a21o_2 _1033_ (.A2(_0198_),
    .A1(_0168_),
    .B1(_0196_),
    .X(_0218_));
 sg13g2_nand2b_1 _1034_ (.Y(_0219_),
    .B(_0195_),
    .A_N(_0218_));
 sg13g2_and4_1 _1035_ (.A(net123),
    .B(net121),
    .C(_0192_),
    .D(_0219_),
    .X(_0220_));
 sg13g2_a22oi_1 _1036_ (.Y(_0221_),
    .B1(_0194_),
    .B2(_0218_),
    .A2(_0191_),
    .A1(net129));
 sg13g2_inv_1 _1037_ (.Y(_0222_),
    .A(_0221_));
 sg13g2_a21o_1 _1038_ (.A2(_0222_),
    .A1(_0208_),
    .B1(_0220_),
    .X(_0223_));
 sg13g2_a22oi_1 _1039_ (.Y(_0224_),
    .B1(_0223_),
    .B2(_0184_),
    .A2(_0209_),
    .A1(_0204_));
 sg13g2_a21oi_2 _1040_ (.B1(_0195_),
    .Y(_0225_),
    .A2(_0191_),
    .A1(net129));
 sg13g2_a22oi_1 _1041_ (.Y(_0226_),
    .B1(_0218_),
    .B2(_0225_),
    .A2(net121),
    .A1(net122));
 sg13g2_nor3_1 _1042_ (.A(_0170_),
    .B(_0193_),
    .C(_0201_),
    .Y(_0227_));
 sg13g2_nor3_2 _1043_ (.A(_0174_),
    .B(_0190_),
    .C(_0227_),
    .Y(_0228_));
 sg13g2_a22oi_1 _1044_ (.Y(_0229_),
    .B1(_0228_),
    .B2(_0202_),
    .A2(_0205_),
    .A1(_0197_));
 sg13g2_a21o_1 _1045_ (.A2(_0228_),
    .A1(_0219_),
    .B1(_0205_),
    .X(_0230_));
 sg13g2_nand2_1 _1046_ (.Y(_0231_),
    .A(_0188_),
    .B(_0205_));
 sg13g2_a22oi_1 _1047_ (.Y(_0232_),
    .B1(_0230_),
    .B2(_0188_),
    .A2(_0229_),
    .A1(_0226_));
 sg13g2_or2_1 _1048_ (.X(_0233_),
    .B(_0232_),
    .A(_0183_));
 sg13g2_a221oi_1 _1049_ (.B2(net129),
    .C1(_0218_),
    .B1(_0191_),
    .A1(net122),
    .Y(_0234_),
    .A2(net121));
 sg13g2_or2_1 _1050_ (.X(_0235_),
    .B(_0207_),
    .A(_0205_));
 sg13g2_nor4_1 _1051_ (.A(_0179_),
    .B(_0181_),
    .C(_0234_),
    .D(_0235_),
    .Y(_0236_));
 sg13g2_nor3_1 _1052_ (.A(_0212_),
    .B(_0214_),
    .C(_0236_),
    .Y(_0237_));
 sg13g2_a22oi_1 _1053_ (.Y(_0238_),
    .B1(_0233_),
    .B2(_0237_),
    .A2(_0224_),
    .A1(_0216_));
 sg13g2_nand2_1 _1054_ (.Y(_0239_),
    .A(\angleOffset[1] ),
    .B(\angle[0] ));
 sg13g2_nand2_1 _1055_ (.Y(_0240_),
    .A(\angleOffset[2] ),
    .B(\angle[1] ));
 sg13g2_xnor2_1 _1056_ (.Y(_0241_),
    .A(\angleOffset[2] ),
    .B(\angle[1] ));
 sg13g2_xnor2_1 _1057_ (.Y(_0242_),
    .A(_0239_),
    .B(_0241_));
 sg13g2_xnor2_1 _1058_ (.Y(_0243_),
    .A(_0238_),
    .B(_0242_));
 sg13g2_xor2_1 _1059_ (.B(\angle[0] ),
    .A(\angleOffset[1] ),
    .X(_0244_));
 sg13g2_o21ai_1 _1060_ (.B1(_0218_),
    .Y(_0245_),
    .A1(_0170_),
    .A2(_0193_));
 sg13g2_nand3_1 _1061_ (.B(_0191_),
    .C(_0245_),
    .A(_0175_),
    .Y(_0246_));
 sg13g2_a22oi_1 _1062_ (.Y(_0247_),
    .B1(_0245_),
    .B2(_0192_),
    .A2(_0205_),
    .A1(_0199_));
 sg13g2_a22oi_1 _1063_ (.Y(_0248_),
    .B1(_0226_),
    .B2(_0247_),
    .A2(_0195_),
    .A1(_0188_));
 sg13g2_nand2_1 _1064_ (.Y(_0249_),
    .A(_0201_),
    .B(_0218_));
 sg13g2_xnor2_1 _1065_ (.Y(_0250_),
    .A(_0225_),
    .B(_0249_));
 sg13g2_nor3_1 _1066_ (.A(_0174_),
    .B(_0190_),
    .C(_0197_),
    .Y(_0251_));
 sg13g2_a22oi_1 _1067_ (.Y(_0252_),
    .B1(_0195_),
    .B2(_0251_),
    .A2(net121),
    .A1(net122));
 sg13g2_a21o_1 _1068_ (.A2(_0197_),
    .A1(_0194_),
    .B1(_0199_),
    .X(_0253_));
 sg13g2_nand3b_1 _1069_ (.B(_0191_),
    .C(net129),
    .Y(_0254_),
    .A_N(_0253_));
 sg13g2_a22oi_1 _1070_ (.Y(_0255_),
    .B1(_0246_),
    .B2(_0253_),
    .A2(_0187_),
    .A1(_0186_));
 sg13g2_a22oi_1 _1071_ (.Y(_0256_),
    .B1(_0254_),
    .B2(_0255_),
    .A2(_0252_),
    .A1(_0250_));
 sg13g2_mux2_1 _1072_ (.A0(_0248_),
    .A1(_0256_),
    .S(_0184_),
    .X(_0257_));
 sg13g2_a21oi_1 _1073_ (.A1(_0194_),
    .A2(_0199_),
    .Y(_0258_),
    .B1(_0246_));
 sg13g2_or3_1 _1074_ (.A(_0189_),
    .B(_0225_),
    .C(_0258_),
    .X(_0259_));
 sg13g2_a22oi_1 _1075_ (.Y(_0260_),
    .B1(_0228_),
    .B2(_0217_),
    .A2(_0221_),
    .A1(_0219_));
 sg13g2_a22oi_1 _1076_ (.Y(_0261_),
    .B1(_0189_),
    .B2(_0260_),
    .A2(_0182_),
    .A1(_0180_));
 sg13g2_a221oi_1 _1077_ (.B2(_0228_),
    .C1(_0206_),
    .B1(_0219_),
    .A1(net122),
    .Y(_0262_),
    .A2(net121));
 sg13g2_a21oi_1 _1078_ (.A1(_0188_),
    .A2(_0221_),
    .Y(_0263_),
    .B1(_0262_));
 sg13g2_a22oi_1 _1079_ (.Y(_0264_),
    .B1(_0263_),
    .B2(_0204_),
    .A2(_0261_),
    .A1(_0259_));
 sg13g2_mux2_1 _1080_ (.A0(_0257_),
    .A1(_0264_),
    .S(_0216_),
    .X(_0265_));
 sg13g2_xnor2_1 _1081_ (.Y(_0266_),
    .A(_0244_),
    .B(_0265_));
 sg13g2_a21oi_1 _1082_ (.A1(_0180_),
    .A2(_0182_),
    .Y(_0267_),
    .B1(_0208_));
 sg13g2_a21oi_1 _1083_ (.A1(net122),
    .A2(net121),
    .Y(_0268_),
    .B1(_0207_));
 sg13g2_or2_1 _1084_ (.X(_0269_),
    .B(_0207_),
    .A(_0188_));
 sg13g2_o21ai_1 _1085_ (.B1(_0231_),
    .Y(_0270_),
    .A1(_0188_),
    .A2(_0221_));
 sg13g2_mux4_1 _1086_ (.S0(_0184_),
    .A0(_0269_),
    .A1(_0270_),
    .A2(_0203_),
    .A3(_0208_),
    .S1(_0216_),
    .X(_0271_));
 sg13g2_and2_1 _1087_ (.A(\angleOffset[3] ),
    .B(\angle[2] ),
    .X(_0272_));
 sg13g2_o21ai_1 _1088_ (.B1(_0240_),
    .Y(_0273_),
    .A1(_0239_),
    .A2(_0241_));
 sg13g2_xor2_1 _1089_ (.B(\angle[2] ),
    .A(\angleOffset[3] ),
    .X(_0274_));
 sg13g2_a21oi_1 _1090_ (.A1(_0273_),
    .A2(_0274_),
    .Y(_0275_),
    .B1(_0272_));
 sg13g2_xnor2_1 _1091_ (.Y(_0276_),
    .A(\angleOffset[4] ),
    .B(\angle[3] ));
 sg13g2_xnor2_1 _1092_ (.Y(_0277_),
    .A(_0275_),
    .B(_0276_));
 sg13g2_xnor2_1 _1093_ (.Y(_0278_),
    .A(_0271_),
    .B(_0277_));
 sg13g2_a21o_1 _1094_ (.A2(_0206_),
    .A1(_0189_),
    .B1(_0203_),
    .X(_0279_));
 sg13g2_a221oi_1 _1095_ (.B2(_0183_),
    .C1(_0267_),
    .B1(_0279_),
    .A1(_0213_),
    .Y(_0280_),
    .A2(_0215_));
 sg13g2_or3_1 _1096_ (.A(_0189_),
    .B(_0225_),
    .C(_0228_),
    .X(_0281_));
 sg13g2_a22oi_1 _1097_ (.Y(_0282_),
    .B1(_0217_),
    .B2(_0221_),
    .A2(_0202_),
    .A1(_0192_));
 sg13g2_or2_1 _1098_ (.X(_0283_),
    .B(_0282_),
    .A(_0188_));
 sg13g2_nand3_1 _1099_ (.B(_0281_),
    .C(_0283_),
    .A(_0184_),
    .Y(_0284_));
 sg13g2_and4_1 _1100_ (.A(net122),
    .B(net121),
    .C(_0192_),
    .D(_0194_),
    .X(_0285_));
 sg13g2_nor4_1 _1101_ (.A(_0179_),
    .B(_0181_),
    .C(_0268_),
    .D(_0285_),
    .Y(_0286_));
 sg13g2_nor3_1 _1102_ (.A(_0212_),
    .B(_0214_),
    .C(_0286_),
    .Y(_0287_));
 sg13g2_a21oi_1 _1103_ (.A1(_0284_),
    .A2(_0287_),
    .Y(_0288_),
    .B1(_0280_));
 sg13g2_xor2_1 _1104_ (.B(_0274_),
    .A(_0273_),
    .X(_0289_));
 sg13g2_xnor2_1 _1105_ (.Y(_0290_),
    .A(_0288_),
    .B(_0289_));
 sg13g2_nor4_2 _1106_ (.A(_0243_),
    .B(_0266_),
    .C(_0278_),
    .Y(_0291_),
    .D(_0290_));
 sg13g2_nor2_1 _1107_ (.A(\hvsync_gen.hpos[7] ),
    .B(\hvsync_gen.hpos[8] ),
    .Y(_0292_));
 sg13g2_nor2b_1 _1108_ (.A(\hvsync_gen.vpos[9] ),
    .B_N(_0140_),
    .Y(_0293_));
 sg13g2_o21ai_1 _1109_ (.B1(_0293_),
    .Y(_0294_),
    .A1(_0007_),
    .A2(_0292_));
 sg13g2_nor2_1 _1110_ (.A(net3),
    .B(_0291_),
    .Y(_0295_));
 sg13g2_a21oi_1 _1111_ (.A1(net6),
    .A2(_0291_),
    .Y(_0296_),
    .B1(_0294_));
 sg13g2_nor2b_2 _1112_ (.A(_0295_),
    .B_N(_0296_),
    .Y(uo_out[4]));
 sg13g2_nor2_1 _1113_ (.A(net4),
    .B(_0291_),
    .Y(_0297_));
 sg13g2_nor2b_1 _1114_ (.A(net7),
    .B_N(_0291_),
    .Y(_0298_));
 sg13g2_nor3_2 _1115_ (.A(_0294_),
    .B(_0297_),
    .C(_0298_),
    .Y(uo_out[5]));
 sg13g2_nor2_1 _1116_ (.A(net5),
    .B(_0291_),
    .Y(_0299_));
 sg13g2_nor2b_1 _1117_ (.A(net8),
    .B_N(_0291_),
    .Y(_0300_));
 sg13g2_nor3_2 _1118_ (.A(_0294_),
    .B(_0299_),
    .C(_0300_),
    .Y(uo_out[6]));
 sg13g2_nand2b_1 _1119_ (.Y(_0301_),
    .B(\angleOffset[0] ),
    .A_N(net2));
 sg13g2_xnor2_1 _1120_ (.Y(_0020_),
    .A(\angleOffset[0] ),
    .B(net2));
 sg13g2_nand2_1 _1121_ (.Y(_0302_),
    .A(\angleOffset[1] ),
    .B(net1));
 sg13g2_nor2_1 _1122_ (.A(\angleOffset[1] ),
    .B(net1),
    .Y(_0303_));
 sg13g2_xor2_1 _1123_ (.B(net1),
    .A(\angleOffset[1] ),
    .X(_0304_));
 sg13g2_xnor2_1 _1124_ (.Y(_0021_),
    .A(_0301_),
    .B(_0304_));
 sg13g2_o21ai_1 _1125_ (.B1(_0302_),
    .Y(_0305_),
    .A1(_0301_),
    .A2(_0303_));
 sg13g2_xor2_1 _1126_ (.B(_0305_),
    .A(\angleOffset[2] ),
    .X(_0022_));
 sg13g2_nand3_1 _1127_ (.B(\angleOffset[3] ),
    .C(_0305_),
    .A(\angleOffset[2] ),
    .Y(_0306_));
 sg13g2_a21o_1 _1128_ (.A2(_0305_),
    .A1(\angleOffset[2] ),
    .B1(\angleOffset[3] ),
    .X(_0307_));
 sg13g2_and2_1 _1129_ (.A(_0306_),
    .B(_0307_),
    .X(_0023_));
 sg13g2_xnor2_1 _1130_ (.Y(_0024_),
    .A(\angleOffset[4] ),
    .B(_0306_));
 sg13g2_nor2_1 _1131_ (.A(net236),
    .B(net150),
    .Y(_0308_));
 sg13g2_nand2b_1 _1132_ (.Y(_0309_),
    .B(net145),
    .A_N(\hypotenuse.multSignal[0] ));
 sg13g2_nor2_1 _1133_ (.A(net173),
    .B(net136),
    .Y(_0310_));
 sg13g2_a21oi_1 _1134_ (.A1(net137),
    .A2(_0309_),
    .Y(_0027_),
    .B1(_0310_));
 sg13g2_or2_1 _1135_ (.X(_0311_),
    .B(net143),
    .A(net145));
 sg13g2_nand2_1 _1136_ (.Y(_0312_),
    .A(net144),
    .B(\hypotenuse.mutlReg[2] ));
 sg13g2_nand3_1 _1137_ (.B(_0311_),
    .C(_0312_),
    .A(net146),
    .Y(_0313_));
 sg13g2_nor2_1 _1138_ (.A(net180),
    .B(net137),
    .Y(_0314_));
 sg13g2_a21oi_1 _1139_ (.A1(net137),
    .A2(_0313_),
    .Y(_0028_),
    .B1(_0314_));
 sg13g2_and3_1 _1140_ (.X(_0315_),
    .A(net145),
    .B(net146),
    .C(\hypotenuse.mutlReg[2] ));
 sg13g2_nand2_1 _1141_ (.Y(_0316_),
    .A(net146),
    .B(net142));
 sg13g2_and2_1 _1142_ (.A(\hypotenuse.multSignal[0] ),
    .B(\hypotenuse.mutlReg[3] ),
    .X(_0317_));
 sg13g2_nand3b_1 _1143_ (.B(_0317_),
    .C(\hypotenuse.mutlReg[2] ),
    .Y(_0318_),
    .A_N(_0018_));
 sg13g2_nor2b_1 _1144_ (.A(net144),
    .B_N(net143),
    .Y(_0319_));
 sg13g2_nand4_1 _1145_ (.B(net143),
    .C(_0018_),
    .A(_0115_),
    .Y(_0320_),
    .D(_0317_));
 sg13g2_xor2_1 _1146_ (.B(_0319_),
    .A(_0317_),
    .X(_0321_));
 sg13g2_nand2_1 _1147_ (.Y(_0322_),
    .A(_0315_),
    .B(_0321_));
 sg13g2_xnor2_1 _1148_ (.Y(_0323_),
    .A(_0315_),
    .B(_0321_));
 sg13g2_nor2_1 _1149_ (.A(net175),
    .B(net136),
    .Y(_0324_));
 sg13g2_a21oi_1 _1150_ (.A1(net136),
    .A2(_0323_),
    .Y(_0029_),
    .B1(_0324_));
 sg13g2_mux2_1 _1151_ (.A0(_0316_),
    .A1(_0318_),
    .S(_0319_),
    .X(_0325_));
 sg13g2_nand2_2 _1152_ (.Y(_0326_),
    .A(net146),
    .B(net141));
 sg13g2_nor2b_1 _1153_ (.A(_0312_),
    .B_N(_0316_),
    .Y(_0327_));
 sg13g2_nand2_1 _1154_ (.Y(_0328_),
    .A(net145),
    .B(\hypotenuse.mutlReg[3] ));
 sg13g2_and2_2 _1155_ (.A(net143),
    .B(net142),
    .X(_0329_));
 sg13g2_nand2_1 _1156_ (.Y(_0330_),
    .A(net143),
    .B(net142));
 sg13g2_nand2_1 _1157_ (.Y(_0331_),
    .A(net143),
    .B(\hypotenuse.mutlReg[5] ));
 sg13g2_nand2b_1 _1158_ (.Y(_0332_),
    .B(_0329_),
    .A_N(_0326_));
 sg13g2_o21ai_1 _1159_ (.B1(net146),
    .Y(_0333_),
    .A1(net141),
    .A2(_0329_));
 sg13g2_nand2b_1 _1160_ (.Y(_0334_),
    .B(_0332_),
    .A_N(_0333_));
 sg13g2_xor2_1 _1161_ (.B(_0334_),
    .A(_0328_),
    .X(_0335_));
 sg13g2_xnor2_1 _1162_ (.Y(_0336_),
    .A(_0327_),
    .B(_0335_));
 sg13g2_nor2_1 _1163_ (.A(_0326_),
    .B(_0336_),
    .Y(_0337_));
 sg13g2_xnor2_1 _1164_ (.Y(_0338_),
    .A(_0326_),
    .B(_0336_));
 sg13g2_nand2_1 _1165_ (.Y(_0339_),
    .A(_0325_),
    .B(_0338_));
 sg13g2_xnor2_1 _1166_ (.Y(_0340_),
    .A(_0325_),
    .B(_0338_));
 sg13g2_nand2_1 _1167_ (.Y(_0341_),
    .A(_0320_),
    .B(_0322_));
 sg13g2_xor2_1 _1168_ (.B(_0341_),
    .A(_0340_),
    .X(_0342_));
 sg13g2_nor2_1 _1169_ (.A(net178),
    .B(net136),
    .Y(_0343_));
 sg13g2_a21oi_1 _1170_ (.A1(net136),
    .A2(_0342_),
    .Y(_0030_),
    .B1(_0343_));
 sg13g2_nand2_1 _1171_ (.Y(_0344_),
    .A(\hypotenuse.multSignal[0] ),
    .B(net140));
 sg13g2_o21ai_1 _1172_ (.B1(_0332_),
    .Y(_0345_),
    .A1(_0328_),
    .A2(_0333_));
 sg13g2_nand2_1 _1173_ (.Y(_0346_),
    .A(net143),
    .B(\hypotenuse.mutlReg[3] ));
 sg13g2_inv_1 _1174_ (.Y(_0347_),
    .A(_0346_));
 sg13g2_nand2_1 _1175_ (.Y(_0348_),
    .A(net144),
    .B(net142));
 sg13g2_nor2b_1 _1176_ (.A(_0348_),
    .B_N(_0326_),
    .Y(_0349_));
 sg13g2_nand2b_1 _1177_ (.Y(_0350_),
    .B(_0326_),
    .A_N(_0348_));
 sg13g2_nand2_2 _1178_ (.Y(_0351_),
    .A(net144),
    .B(net141));
 sg13g2_xnor2_1 _1179_ (.Y(_0352_),
    .A(\hypotenuse.mutlReg[3] ),
    .B(_0329_));
 sg13g2_nor2_1 _1180_ (.A(_0351_),
    .B(_0352_),
    .Y(_0353_));
 sg13g2_xor2_1 _1181_ (.B(_0352_),
    .A(_0351_),
    .X(_0354_));
 sg13g2_xnor2_1 _1182_ (.Y(_0355_),
    .A(_0351_),
    .B(_0352_));
 sg13g2_nor2_1 _1183_ (.A(_0316_),
    .B(_0351_),
    .Y(_0356_));
 sg13g2_and4_1 _1184_ (.A(net144),
    .B(net146),
    .C(net141),
    .D(net140),
    .X(_0357_));
 sg13g2_nand4_1 _1185_ (.B(net146),
    .C(net141),
    .A(net144),
    .Y(_0358_),
    .D(net140));
 sg13g2_a22oi_1 _1186_ (.Y(_0359_),
    .B1(net140),
    .B2(net146),
    .A2(net141),
    .A1(net144));
 sg13g2_nand3b_1 _1187_ (.B(_0329_),
    .C(_0358_),
    .Y(_0360_),
    .A_N(_0359_));
 sg13g2_o21ai_1 _1188_ (.B1(_0330_),
    .Y(_0361_),
    .A1(_0357_),
    .A2(_0359_));
 sg13g2_and3_1 _1189_ (.X(_0362_),
    .A(_0356_),
    .B(_0360_),
    .C(_0361_));
 sg13g2_nand3_1 _1190_ (.B(_0360_),
    .C(_0361_),
    .A(_0356_),
    .Y(_0363_));
 sg13g2_a21oi_1 _1191_ (.A1(_0360_),
    .A2(_0361_),
    .Y(_0364_),
    .B1(_0356_));
 sg13g2_a21o_1 _1192_ (.A2(_0361_),
    .A1(_0360_),
    .B1(_0356_),
    .X(_0365_));
 sg13g2_nor3_2 _1193_ (.A(_0355_),
    .B(_0362_),
    .C(_0364_),
    .Y(_0366_));
 sg13g2_nand3_1 _1194_ (.B(_0363_),
    .C(_0365_),
    .A(_0354_),
    .Y(_0367_));
 sg13g2_a21oi_1 _1195_ (.A1(_0363_),
    .A2(_0365_),
    .Y(_0368_),
    .B1(_0354_));
 sg13g2_o21ai_1 _1196_ (.B1(_0355_),
    .Y(_0369_),
    .A1(_0362_),
    .A2(_0364_));
 sg13g2_nor3_1 _1197_ (.A(_0350_),
    .B(_0366_),
    .C(_0368_),
    .Y(_0370_));
 sg13g2_nand3_1 _1198_ (.B(_0367_),
    .C(_0369_),
    .A(_0349_),
    .Y(_0371_));
 sg13g2_a21oi_1 _1199_ (.A1(_0367_),
    .A2(_0369_),
    .Y(_0372_),
    .B1(_0349_));
 sg13g2_o21ai_1 _1200_ (.B1(_0350_),
    .Y(_0373_),
    .A1(_0366_),
    .A2(_0368_));
 sg13g2_nor3_1 _1201_ (.A(_0346_),
    .B(_0370_),
    .C(_0372_),
    .Y(_0374_));
 sg13g2_nand3_1 _1202_ (.B(_0371_),
    .C(_0373_),
    .A(_0347_),
    .Y(_0375_));
 sg13g2_a21oi_1 _1203_ (.A1(_0371_),
    .A2(_0373_),
    .Y(_0376_),
    .B1(_0347_));
 sg13g2_o21ai_1 _1204_ (.B1(_0346_),
    .Y(_0377_),
    .A1(_0370_),
    .A2(_0372_));
 sg13g2_nand3_1 _1205_ (.B(_0375_),
    .C(_0377_),
    .A(_0345_),
    .Y(_0378_));
 sg13g2_a21oi_1 _1206_ (.A1(_0375_),
    .A2(_0377_),
    .Y(_0379_),
    .B1(_0345_));
 sg13g2_nor3_1 _1207_ (.A(_0345_),
    .B(_0374_),
    .C(_0376_),
    .Y(_0380_));
 sg13g2_o21ai_1 _1208_ (.B1(_0345_),
    .Y(_0381_),
    .A1(_0374_),
    .A2(_0376_));
 sg13g2_nor2b_1 _1209_ (.A(_0380_),
    .B_N(_0381_),
    .Y(_0382_));
 sg13g2_xnor2_1 _1210_ (.Y(_0383_),
    .A(_0344_),
    .B(_0382_));
 sg13g2_a21oi_2 _1211_ (.B1(_0337_),
    .Y(_0384_),
    .A2(_0335_),
    .A1(_0327_));
 sg13g2_nor2_1 _1212_ (.A(_0383_),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_xor2_1 _1213_ (.B(_0384_),
    .A(_0383_),
    .X(_0386_));
 sg13g2_o21ai_1 _1214_ (.B1(_0320_),
    .Y(_0387_),
    .A1(_0325_),
    .A2(_0338_));
 sg13g2_nand2_1 _1215_ (.Y(_0388_),
    .A(_0339_),
    .B(_0387_));
 sg13g2_o21ai_1 _1216_ (.B1(_0388_),
    .Y(_0389_),
    .A1(_0322_),
    .A2(_0340_));
 sg13g2_xnor2_1 _1217_ (.Y(_0390_),
    .A(_0386_),
    .B(_0389_));
 sg13g2_nor2_1 _1218_ (.A(net182),
    .B(net136),
    .Y(_0391_));
 sg13g2_a21oi_1 _1219_ (.A1(net136),
    .A2(_0390_),
    .Y(_0031_),
    .B1(_0391_));
 sg13g2_o21ai_1 _1220_ (.B1(_0378_),
    .Y(_0392_),
    .A1(_0344_),
    .A2(_0379_));
 sg13g2_a21oi_1 _1221_ (.A1(\hypotenuse.mutlReg[3] ),
    .A2(_0329_),
    .Y(_0393_),
    .B1(_0353_));
 sg13g2_nand2_1 _1222_ (.Y(_0394_),
    .A(_0358_),
    .B(_0360_));
 sg13g2_o21ai_1 _1223_ (.B1(_0394_),
    .Y(_0395_),
    .A1(_0362_),
    .A2(_0366_));
 sg13g2_nand4_1 _1224_ (.B(_0360_),
    .C(_0363_),
    .A(_0358_),
    .Y(_0396_),
    .D(_0367_));
 sg13g2_and2_1 _1225_ (.A(_0395_),
    .B(_0396_),
    .X(_0397_));
 sg13g2_nand2b_1 _1226_ (.Y(_0398_),
    .B(_0397_),
    .A_N(_0393_));
 sg13g2_xor2_1 _1227_ (.B(_0397_),
    .A(_0393_),
    .X(_0399_));
 sg13g2_nand2_1 _1228_ (.Y(_0400_),
    .A(_0371_),
    .B(_0375_));
 sg13g2_nor2b_1 _1229_ (.A(_0399_),
    .B_N(_0400_),
    .Y(_0401_));
 sg13g2_inv_1 _1230_ (.Y(_0402_),
    .A(_0401_));
 sg13g2_xor2_1 _1231_ (.B(_0400_),
    .A(_0399_),
    .X(_0403_));
 sg13g2_nor2b_1 _1232_ (.A(_0403_),
    .B_N(_0392_),
    .Y(_0404_));
 sg13g2_xor2_1 _1233_ (.B(_0403_),
    .A(_0392_),
    .X(_0405_));
 sg13g2_a21oi_1 _1234_ (.A1(_0386_),
    .A2(_0389_),
    .Y(_0406_),
    .B1(_0385_));
 sg13g2_xnor2_1 _1235_ (.Y(_0407_),
    .A(_0405_),
    .B(_0406_));
 sg13g2_nor2_1 _1236_ (.A(net194),
    .B(net137),
    .Y(_0408_));
 sg13g2_a21oi_1 _1237_ (.A1(net137),
    .A2(_0407_),
    .Y(_0032_),
    .B1(_0408_));
 sg13g2_a22oi_1 _1238_ (.Y(_0409_),
    .B1(net140),
    .B2(net144),
    .A2(net142),
    .A1(\hypotenuse.mutlReg[3] ));
 sg13g2_nand2_2 _1239_ (.Y(_0410_),
    .A(\hypotenuse.mutlReg[3] ),
    .B(net140));
 sg13g2_inv_1 _1240_ (.Y(_0411_),
    .A(_0410_));
 sg13g2_or2_1 _1241_ (.X(_0412_),
    .B(_0410_),
    .A(_0348_));
 sg13g2_o21ai_1 _1242_ (.B1(_0412_),
    .Y(_0413_),
    .A1(_0331_),
    .A2(_0409_));
 sg13g2_nor2b_1 _1243_ (.A(_0409_),
    .B_N(_0412_),
    .Y(_0414_));
 sg13g2_xnor2_1 _1244_ (.Y(_0415_),
    .A(_0331_),
    .B(_0414_));
 sg13g2_xor2_1 _1245_ (.B(_0415_),
    .A(_0019_),
    .X(_0416_));
 sg13g2_a21oi_2 _1246_ (.B1(_0416_),
    .Y(_0417_),
    .A2(_0398_),
    .A1(_0395_));
 sg13g2_nand3_1 _1247_ (.B(_0398_),
    .C(_0416_),
    .A(_0395_),
    .Y(_0418_));
 sg13g2_nand2b_1 _1248_ (.Y(_0419_),
    .B(_0418_),
    .A_N(_0417_));
 sg13g2_nor2_1 _1249_ (.A(_0402_),
    .B(_0419_),
    .Y(_0420_));
 sg13g2_xnor2_1 _1250_ (.Y(_0421_),
    .A(_0402_),
    .B(_0419_));
 sg13g2_o21ai_1 _1251_ (.B1(_0388_),
    .Y(_0422_),
    .A1(_0383_),
    .A2(_0384_));
 sg13g2_a21oi_1 _1252_ (.A1(_0383_),
    .A2(_0384_),
    .Y(_0423_),
    .B1(_0405_));
 sg13g2_a221oi_1 _1253_ (.B2(_0423_),
    .C1(_0404_),
    .B1(_0422_),
    .A1(_0315_),
    .Y(_0424_),
    .A2(_0411_));
 sg13g2_nor2_1 _1254_ (.A(_0421_),
    .B(_0424_),
    .Y(_0425_));
 sg13g2_xnor2_1 _1255_ (.Y(_0426_),
    .A(_0421_),
    .B(_0424_));
 sg13g2_nor2_1 _1256_ (.A(net201),
    .B(net136),
    .Y(_0427_));
 sg13g2_a21oi_1 _1257_ (.A1(net137),
    .A2(_0426_),
    .Y(_0033_),
    .B1(_0427_));
 sg13g2_nand2_1 _1258_ (.Y(_0428_),
    .A(\hypotenuse.mutlReg[3] ),
    .B(\hypotenuse.mutlReg[5] ));
 sg13g2_nand2_1 _1259_ (.Y(_0429_),
    .A(net143),
    .B(net140));
 sg13g2_xor2_1 _1260_ (.B(_0429_),
    .A(_0428_),
    .X(_0430_));
 sg13g2_a21oi_1 _1261_ (.A1(\hypotenuse.mutlReg[4] ),
    .A2(_0413_),
    .Y(_0431_),
    .B1(_0430_));
 sg13g2_nand3_1 _1262_ (.B(_0413_),
    .C(_0430_),
    .A(net142),
    .Y(_0432_));
 sg13g2_nand2b_1 _1263_ (.Y(_0433_),
    .B(_0432_),
    .A_N(_0431_));
 sg13g2_mux2_1 _1264_ (.A0(_0415_),
    .A1(_0413_),
    .S(_0019_),
    .X(_0434_));
 sg13g2_nand2b_2 _1265_ (.Y(_0435_),
    .B(_0434_),
    .A_N(_0433_));
 sg13g2_xor2_1 _1266_ (.B(_0434_),
    .A(_0433_),
    .X(_0436_));
 sg13g2_inv_1 _1267_ (.Y(_0437_),
    .A(_0436_));
 sg13g2_xnor2_1 _1268_ (.Y(_0438_),
    .A(_0417_),
    .B(_0437_));
 sg13g2_nor2_1 _1269_ (.A(_0420_),
    .B(_0425_),
    .Y(_0439_));
 sg13g2_xnor2_1 _1270_ (.Y(_0440_),
    .A(_0438_),
    .B(_0439_));
 sg13g2_nor2_1 _1271_ (.A(net208),
    .B(net138),
    .Y(_0441_));
 sg13g2_a21oi_1 _1272_ (.A1(net138),
    .A2(_0440_),
    .Y(_0034_),
    .B1(_0441_));
 sg13g2_nor2_1 _1273_ (.A(net214),
    .B(net138),
    .Y(_0442_));
 sg13g2_nand2b_1 _1274_ (.Y(_0443_),
    .B(net141),
    .A_N(net142));
 sg13g2_nor2_1 _1275_ (.A(_0410_),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_xor2_1 _1276_ (.B(_0443_),
    .A(_0410_),
    .X(_0445_));
 sg13g2_o21ai_1 _1277_ (.B1(_0432_),
    .Y(_0446_),
    .A1(_0428_),
    .A2(_0429_));
 sg13g2_and2_1 _1278_ (.A(_0445_),
    .B(_0446_),
    .X(_0447_));
 sg13g2_inv_1 _1279_ (.Y(_0448_),
    .A(_0447_));
 sg13g2_xor2_1 _1280_ (.B(_0446_),
    .A(_0445_),
    .X(_0449_));
 sg13g2_nor2b_1 _1281_ (.A(_0435_),
    .B_N(_0449_),
    .Y(_0450_));
 sg13g2_nand2b_1 _1282_ (.Y(_0451_),
    .B(_0449_),
    .A_N(_0435_));
 sg13g2_xnor2_1 _1283_ (.Y(_0452_),
    .A(_0435_),
    .B(_0449_));
 sg13g2_xor2_1 _1284_ (.B(_0449_),
    .A(_0435_),
    .X(_0453_));
 sg13g2_or2_1 _1285_ (.X(_0454_),
    .B(_0438_),
    .A(_0421_));
 sg13g2_o21ai_1 _1286_ (.B1(_0437_),
    .Y(_0455_),
    .A1(_0417_),
    .A2(_0420_));
 sg13g2_o21ai_1 _1287_ (.B1(_0455_),
    .Y(_0456_),
    .A1(_0424_),
    .A2(_0454_));
 sg13g2_xnor2_1 _1288_ (.Y(_0457_),
    .A(_0452_),
    .B(_0456_));
 sg13g2_a21oi_1 _1289_ (.A1(net138),
    .A2(_0457_),
    .Y(_0035_),
    .B1(_0442_));
 sg13g2_xor2_1 _1290_ (.B(net140),
    .A(net141),
    .X(_0458_));
 sg13g2_a21oi_1 _1291_ (.A1(net142),
    .A2(_0458_),
    .Y(_0459_),
    .B1(_0444_));
 sg13g2_xor2_1 _1292_ (.B(_0459_),
    .A(_0447_),
    .X(_0460_));
 sg13g2_a21oi_1 _1293_ (.A1(_0452_),
    .A2(_0456_),
    .Y(_0461_),
    .B1(_0450_));
 sg13g2_xnor2_1 _1294_ (.Y(_0462_),
    .A(_0460_),
    .B(_0461_));
 sg13g2_nor2_1 _1295_ (.A(net202),
    .B(net138),
    .Y(_0463_));
 sg13g2_a21oi_1 _1296_ (.A1(net138),
    .A2(_0462_),
    .Y(_0036_),
    .B1(_0463_));
 sg13g2_nor2_1 _1297_ (.A(_0453_),
    .B(_0460_),
    .Y(_0464_));
 sg13g2_a21oi_1 _1298_ (.A1(_0448_),
    .A2(_0451_),
    .Y(_0465_),
    .B1(_0459_));
 sg13g2_a21oi_1 _1299_ (.A1(_0456_),
    .A2(_0464_),
    .Y(_0466_),
    .B1(_0465_));
 sg13g2_nand2_1 _1300_ (.Y(_0467_),
    .A(\hypotenuse.mutlReg[6] ),
    .B(_0443_));
 sg13g2_xor2_1 _1301_ (.B(_0467_),
    .A(_0466_),
    .X(_0468_));
 sg13g2_mux2_1 _1302_ (.A0(net195),
    .A1(_0468_),
    .S(net138),
    .X(_0037_));
 sg13g2_xnor2_1 _1303_ (.Y(_0469_),
    .A(\hvsync_gen.hpos[3] ),
    .B(_0127_));
 sg13g2_nand2_1 _1304_ (.Y(_0470_),
    .A(_0008_),
    .B(_0117_));
 sg13g2_xor2_1 _1305_ (.B(_0470_),
    .A(\hvsync_gen.vpos[3] ),
    .X(_0471_));
 sg13g2_inv_1 _1306_ (.Y(_0472_),
    .A(_0471_));
 sg13g2_nor2_2 _1307_ (.A(_0469_),
    .B(_0471_),
    .Y(_0473_));
 sg13g2_a21oi_1 _1308_ (.A1(_0469_),
    .A2(_0471_),
    .Y(_0474_),
    .B1(net149));
 sg13g2_nor2b_1 _1309_ (.A(_0473_),
    .B_N(_0474_),
    .Y(_0038_));
 sg13g2_xnor2_1 _1310_ (.Y(_0475_),
    .A(\hvsync_gen.vpos[4] ),
    .B(_0118_));
 sg13g2_inv_1 _1311_ (.Y(_0476_),
    .A(_0475_));
 sg13g2_xor2_1 _1312_ (.B(_0128_),
    .A(_0009_),
    .X(_0477_));
 sg13g2_nand2_1 _1313_ (.Y(_0478_),
    .A(_0476_),
    .B(_0477_));
 sg13g2_xnor2_1 _1314_ (.Y(_0479_),
    .A(_0475_),
    .B(_0477_));
 sg13g2_nand2_1 _1315_ (.Y(_0480_),
    .A(_0469_),
    .B(_0472_));
 sg13g2_nor2_1 _1316_ (.A(_0479_),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_nand2_1 _1317_ (.Y(_0482_),
    .A(_0479_),
    .B(_0480_));
 sg13g2_nor2b_1 _1318_ (.A(_0481_),
    .B_N(_0482_),
    .Y(_0483_));
 sg13g2_nor2b_1 _1319_ (.A(_0479_),
    .B_N(_0473_),
    .Y(_0484_));
 sg13g2_xor2_1 _1320_ (.B(_0479_),
    .A(_0473_),
    .X(_0485_));
 sg13g2_a21o_1 _1321_ (.A2(_0485_),
    .A1(net127),
    .B1(net125),
    .X(_0486_));
 sg13g2_nand2_1 _1322_ (.Y(_0487_),
    .A(_0009_),
    .B(_0469_));
 sg13g2_mux2_2 _1323_ (.A0(_0477_),
    .A1(_0009_),
    .S(_0469_),
    .X(_0488_));
 sg13g2_nor2_1 _1324_ (.A(_0475_),
    .B(_0488_),
    .Y(_0489_));
 sg13g2_nor2_1 _1325_ (.A(_0476_),
    .B(_0488_),
    .Y(_0490_));
 sg13g2_nand2_1 _1326_ (.Y(_0491_),
    .A(_0476_),
    .B(_0488_));
 sg13g2_xnor2_1 _1327_ (.Y(_0492_),
    .A(_0476_),
    .B(_0488_));
 sg13g2_and2_1 _1328_ (.A(_0480_),
    .B(_0492_),
    .X(_0493_));
 sg13g2_nor2_1 _1329_ (.A(_0481_),
    .B(_0493_),
    .Y(_0494_));
 sg13g2_a22oi_1 _1330_ (.Y(_0495_),
    .B1(_0494_),
    .B2(_0125_),
    .A2(_0483_),
    .A1(_0135_));
 sg13g2_nor2_1 _1331_ (.A(net128),
    .B(_0133_),
    .Y(_0496_));
 sg13g2_nand2_2 _1332_ (.Y(_0497_),
    .A(_0125_),
    .B(net124));
 sg13g2_xor2_1 _1333_ (.B(_0492_),
    .A(_0473_),
    .X(_0498_));
 sg13g2_a221oi_1 _1334_ (.B2(net119),
    .C1(net149),
    .B1(_0498_),
    .A1(_0486_),
    .Y(_0039_),
    .A2(_0495_));
 sg13g2_xnor2_1 _1335_ (.Y(_0499_),
    .A(\hvsync_gen.vpos[5] ),
    .B(_0119_));
 sg13g2_inv_1 _1336_ (.Y(_0500_),
    .A(_0499_));
 sg13g2_nor2_2 _1337_ (.A(\hvsync_gen.hpos[5] ),
    .B(_0487_),
    .Y(_0501_));
 sg13g2_o21ai_1 _1338_ (.B1(\hvsync_gen.hpos[5] ),
    .Y(_0502_),
    .A1(\hvsync_gen.hpos[4] ),
    .A2(_0128_));
 sg13g2_nor2b_2 _1339_ (.A(_0129_),
    .B_N(_0502_),
    .Y(_0503_));
 sg13g2_a21oi_1 _1340_ (.A1(_0009_),
    .A2(_0469_),
    .Y(_0504_),
    .B1(_0503_));
 sg13g2_nor2_2 _1341_ (.A(_0501_),
    .B(_0504_),
    .Y(_0505_));
 sg13g2_nand2_1 _1342_ (.Y(_0506_),
    .A(_0500_),
    .B(_0505_));
 sg13g2_nor2_1 _1343_ (.A(_0500_),
    .B(_0505_),
    .Y(_0507_));
 sg13g2_nand2_1 _1344_ (.Y(_0508_),
    .A(_0499_),
    .B(_0505_));
 sg13g2_xnor2_1 _1345_ (.Y(_0509_),
    .A(_0499_),
    .B(_0505_));
 sg13g2_nor2_1 _1346_ (.A(_0489_),
    .B(_0493_),
    .Y(_0510_));
 sg13g2_xor2_1 _1347_ (.B(_0510_),
    .A(_0509_),
    .X(_0511_));
 sg13g2_or2_1 _1348_ (.X(_0512_),
    .B(_0503_),
    .A(_0500_));
 sg13g2_nor2_1 _1349_ (.A(_0499_),
    .B(_0503_),
    .Y(_0513_));
 sg13g2_xnor2_1 _1350_ (.Y(_0514_),
    .A(_0499_),
    .B(_0503_));
 sg13g2_xor2_1 _1351_ (.B(_0503_),
    .A(_0499_),
    .X(_0515_));
 sg13g2_a21o_1 _1352_ (.A2(_0482_),
    .A1(_0478_),
    .B1(_0515_),
    .X(_0516_));
 sg13g2_nand3_1 _1353_ (.B(_0482_),
    .C(_0515_),
    .A(_0478_),
    .Y(_0517_));
 sg13g2_and2_1 _1354_ (.A(_0516_),
    .B(_0517_),
    .X(_0518_));
 sg13g2_a21oi_1 _1355_ (.A1(_0475_),
    .A2(_0477_),
    .Y(_0519_),
    .B1(_0484_));
 sg13g2_or2_1 _1356_ (.X(_0520_),
    .B(_0519_),
    .A(_0514_));
 sg13g2_xnor2_1 _1357_ (.Y(_0521_),
    .A(_0514_),
    .B(_0519_));
 sg13g2_a21oi_1 _1358_ (.A1(net128),
    .A2(_0521_),
    .Y(_0522_),
    .B1(net124));
 sg13g2_a221oi_1 _1359_ (.B2(_0135_),
    .C1(_0522_),
    .B1(_0518_),
    .A1(_0496_),
    .Y(_0523_),
    .A2(_0511_));
 sg13g2_a21oi_2 _1360_ (.B1(_0490_),
    .Y(_0524_),
    .A2(_0491_),
    .A1(_0473_));
 sg13g2_xnor2_1 _1361_ (.Y(_0525_),
    .A(_0509_),
    .B(_0524_));
 sg13g2_o21ai_1 _1362_ (.B1(net153),
    .Y(_0526_),
    .A1(net118),
    .A2(_0525_));
 sg13g2_nor2_1 _1363_ (.A(_0523_),
    .B(_0526_),
    .Y(_0040_));
 sg13g2_xnor2_1 _1364_ (.Y(_0527_),
    .A(\hvsync_gen.vpos[6] ),
    .B(_0120_));
 sg13g2_xnor2_1 _1365_ (.Y(_0528_),
    .A(net147),
    .B(_0129_));
 sg13g2_inv_1 _1366_ (.Y(_0529_),
    .A(_0528_));
 sg13g2_nor2b_1 _1367_ (.A(_0528_),
    .B_N(_0501_),
    .Y(_0530_));
 sg13g2_xnor2_1 _1368_ (.Y(_0531_),
    .A(_0501_),
    .B(_0528_));
 sg13g2_or2_1 _1369_ (.X(_0532_),
    .B(_0531_),
    .A(_0527_));
 sg13g2_nand2_1 _1370_ (.Y(_0533_),
    .A(_0527_),
    .B(_0531_));
 sg13g2_nand2_2 _1371_ (.Y(_0534_),
    .A(_0532_),
    .B(_0533_));
 sg13g2_o21ai_1 _1372_ (.B1(_0508_),
    .Y(_0535_),
    .A1(_0509_),
    .A2(_0510_));
 sg13g2_xor2_1 _1373_ (.B(_0535_),
    .A(_0534_),
    .X(_0536_));
 sg13g2_nor2_1 _1374_ (.A(_0527_),
    .B(_0529_),
    .Y(_0537_));
 sg13g2_nand2_1 _1375_ (.Y(_0538_),
    .A(_0527_),
    .B(_0529_));
 sg13g2_nor2b_2 _1376_ (.A(_0537_),
    .B_N(_0538_),
    .Y(_0539_));
 sg13g2_a21oi_1 _1377_ (.A1(_0512_),
    .A2(_0516_),
    .Y(_0540_),
    .B1(_0539_));
 sg13g2_nand3_1 _1378_ (.B(_0516_),
    .C(_0539_),
    .A(_0512_),
    .Y(_0541_));
 sg13g2_nand2b_1 _1379_ (.Y(_0542_),
    .B(_0541_),
    .A_N(_0540_));
 sg13g2_nor2_1 _1380_ (.A(_0136_),
    .B(_0542_),
    .Y(_0543_));
 sg13g2_nor2b_1 _1381_ (.A(_0513_),
    .B_N(_0520_),
    .Y(_0544_));
 sg13g2_xnor2_1 _1382_ (.Y(_0545_),
    .A(_0539_),
    .B(_0544_));
 sg13g2_a21oi_1 _1383_ (.A1(_0133_),
    .A2(_0545_),
    .Y(_0546_),
    .B1(net119));
 sg13g2_o21ai_1 _1384_ (.B1(_0546_),
    .Y(_0547_),
    .A1(_0497_),
    .A2(_0536_));
 sg13g2_o21ai_1 _1385_ (.B1(_0506_),
    .Y(_0548_),
    .A1(_0507_),
    .A2(_0524_));
 sg13g2_xnor2_1 _1386_ (.Y(_0549_),
    .A(_0534_),
    .B(_0548_));
 sg13g2_o21ai_1 _1387_ (.B1(net153),
    .Y(_0550_),
    .A1(_0543_),
    .A2(_0547_));
 sg13g2_a21oi_1 _1388_ (.A1(net119),
    .A2(_0549_),
    .Y(_0041_),
    .B1(_0550_));
 sg13g2_a21oi_1 _1389_ (.A1(\hvsync_gen.vpos[6] ),
    .A2(_0120_),
    .Y(_0551_),
    .B1(\hvsync_gen.vpos[7] ));
 sg13g2_nor2_2 _1390_ (.A(_0122_),
    .B(_0551_),
    .Y(_0552_));
 sg13g2_xor2_1 _1391_ (.B(_0130_),
    .A(\hvsync_gen.hpos[7] ),
    .X(_0553_));
 sg13g2_nor2b_1 _1392_ (.A(_0553_),
    .B_N(_0530_),
    .Y(_0554_));
 sg13g2_xnor2_1 _1393_ (.Y(_0555_),
    .A(_0530_),
    .B(_0553_));
 sg13g2_nor2b_1 _1394_ (.A(_0552_),
    .B_N(_0555_),
    .Y(_0556_));
 sg13g2_nand2_1 _1395_ (.Y(_0557_),
    .A(_0552_),
    .B(_0555_));
 sg13g2_xnor2_1 _1396_ (.Y(_0558_),
    .A(_0552_),
    .B(_0555_));
 sg13g2_nand2_1 _1397_ (.Y(_0559_),
    .A(_0532_),
    .B(_0535_));
 sg13g2_nand2_1 _1398_ (.Y(_0560_),
    .A(_0533_),
    .B(_0559_));
 sg13g2_xnor2_1 _1399_ (.Y(_0561_),
    .A(_0558_),
    .B(_0560_));
 sg13g2_or2_1 _1400_ (.X(_0562_),
    .B(_0561_),
    .A(_0497_));
 sg13g2_o21ai_1 _1401_ (.B1(_0553_),
    .Y(_0563_),
    .A1(_0122_),
    .A2(_0551_));
 sg13g2_xnor2_1 _1402_ (.Y(_0564_),
    .A(_0552_),
    .B(_0553_));
 sg13g2_inv_1 _1403_ (.Y(_0565_),
    .A(_0564_));
 sg13g2_nand2_1 _1404_ (.Y(_0566_),
    .A(_0527_),
    .B(_0528_));
 sg13g2_nor2b_1 _1405_ (.A(_0540_),
    .B_N(_0566_),
    .Y(_0567_));
 sg13g2_nand2b_1 _1406_ (.Y(_0568_),
    .B(_0564_),
    .A_N(_0567_));
 sg13g2_xnor2_1 _1407_ (.Y(_0569_),
    .A(_0565_),
    .B(_0567_));
 sg13g2_nor2_1 _1408_ (.A(_0136_),
    .B(_0569_),
    .Y(_0570_));
 sg13g2_o21ai_1 _1409_ (.B1(_0538_),
    .Y(_0571_),
    .A1(_0513_),
    .A2(_0537_));
 sg13g2_o21ai_1 _1410_ (.B1(_0571_),
    .Y(_0572_),
    .A1(_0520_),
    .A2(_0534_));
 sg13g2_and2_1 _1411_ (.A(_0565_),
    .B(_0572_),
    .X(_0573_));
 sg13g2_xnor2_1 _1412_ (.Y(_0574_),
    .A(_0565_),
    .B(_0572_));
 sg13g2_o21ai_1 _1413_ (.B1(_0138_),
    .Y(_0575_),
    .A1(net124),
    .A2(_0574_));
 sg13g2_nor2_1 _1414_ (.A(_0570_),
    .B(_0575_),
    .Y(_0576_));
 sg13g2_nor3_1 _1415_ (.A(_0515_),
    .B(_0524_),
    .C(_0539_),
    .Y(_0577_));
 sg13g2_nand2b_1 _1416_ (.Y(_0578_),
    .B(_0531_),
    .A_N(_0527_));
 sg13g2_nand2_1 _1417_ (.Y(_0579_),
    .A(_0506_),
    .B(_0578_));
 sg13g2_a21oi_2 _1418_ (.B1(_0577_),
    .Y(_0580_),
    .A2(_0579_),
    .A1(_0566_));
 sg13g2_xnor2_1 _1419_ (.Y(_0581_),
    .A(_0558_),
    .B(_0580_));
 sg13g2_a221oi_1 _1420_ (.B2(net120),
    .C1(net150),
    .B1(_0581_),
    .A1(_0562_),
    .Y(_0042_),
    .A2(_0576_));
 sg13g2_nor2_1 _1421_ (.A(\hvsync_gen.hpos[8] ),
    .B(_0131_),
    .Y(_0582_));
 sg13g2_xor2_1 _1422_ (.B(_0131_),
    .A(\hvsync_gen.hpos[8] ),
    .X(_0583_));
 sg13g2_nor2b_1 _1423_ (.A(_0583_),
    .B_N(_0554_),
    .Y(_0584_));
 sg13g2_xnor2_1 _1424_ (.Y(_0585_),
    .A(_0554_),
    .B(_0583_));
 sg13g2_xnor2_1 _1425_ (.Y(_0586_),
    .A(\hvsync_gen.vpos[8] ),
    .B(_0122_));
 sg13g2_inv_1 _1426_ (.Y(_0587_),
    .A(_0586_));
 sg13g2_nor2_1 _1427_ (.A(_0585_),
    .B(_0587_),
    .Y(_0588_));
 sg13g2_nand2_1 _1428_ (.Y(_0589_),
    .A(_0585_),
    .B(_0587_));
 sg13g2_nor2b_1 _1429_ (.A(_0588_),
    .B_N(_0589_),
    .Y(_0590_));
 sg13g2_nand2b_1 _1430_ (.Y(_0591_),
    .B(_0589_),
    .A_N(_0588_));
 sg13g2_a21oi_1 _1431_ (.A1(_0558_),
    .A2(_0560_),
    .Y(_0592_),
    .B1(_0556_));
 sg13g2_xnor2_1 _1432_ (.Y(_0593_),
    .A(_0591_),
    .B(_0592_));
 sg13g2_or2_1 _1433_ (.X(_0594_),
    .B(_0593_),
    .A(_0497_));
 sg13g2_or2_1 _1434_ (.X(_0595_),
    .B(_0586_),
    .A(_0583_));
 sg13g2_xor2_1 _1435_ (.B(_0586_),
    .A(_0583_),
    .X(_0596_));
 sg13g2_a21oi_1 _1436_ (.A1(_0563_),
    .A2(_0568_),
    .Y(_0597_),
    .B1(_0596_));
 sg13g2_nand3_1 _1437_ (.B(_0568_),
    .C(_0596_),
    .A(_0563_),
    .Y(_0598_));
 sg13g2_nand2b_1 _1438_ (.Y(_0599_),
    .B(_0598_),
    .A_N(_0597_));
 sg13g2_nor2_1 _1439_ (.A(_0136_),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_a21o_1 _1440_ (.A2(_0553_),
    .A1(_0552_),
    .B1(_0573_),
    .X(_0601_));
 sg13g2_xnor2_1 _1441_ (.Y(_0602_),
    .A(_0596_),
    .B(_0601_));
 sg13g2_o21ai_1 _1442_ (.B1(net118),
    .Y(_0603_),
    .A1(net124),
    .A2(_0602_));
 sg13g2_nor2_1 _1443_ (.A(_0600_),
    .B(_0603_),
    .Y(_0604_));
 sg13g2_o21ai_1 _1444_ (.B1(_0557_),
    .Y(_0605_),
    .A1(_0558_),
    .A2(_0580_));
 sg13g2_xnor2_1 _1445_ (.Y(_0606_),
    .A(_0591_),
    .B(_0605_));
 sg13g2_a221oi_1 _1446_ (.B2(net120),
    .C1(net150),
    .B1(_0606_),
    .A1(_0594_),
    .Y(_0043_),
    .A2(_0604_));
 sg13g2_xnor2_1 _1447_ (.Y(_0607_),
    .A(_0139_),
    .B(_0584_));
 sg13g2_o21ai_1 _1448_ (.B1(_0589_),
    .Y(_0608_),
    .A1(_0588_),
    .A2(_0592_));
 sg13g2_xor2_1 _1449_ (.B(_0608_),
    .A(_0607_),
    .X(_0609_));
 sg13g2_a21oi_1 _1450_ (.A1(_0583_),
    .A2(_0587_),
    .Y(_0610_),
    .B1(_0597_));
 sg13g2_nand2_1 _1451_ (.Y(_0611_),
    .A(_0135_),
    .B(_0610_));
 sg13g2_and3_1 _1452_ (.X(_0612_),
    .A(_0552_),
    .B(_0553_),
    .C(_0595_));
 sg13g2_a221oi_1 _1453_ (.B2(_0573_),
    .C1(_0612_),
    .B1(_0590_),
    .A1(_0583_),
    .Y(_0613_),
    .A2(_0586_));
 sg13g2_a221oi_1 _1454_ (.B2(net126),
    .C1(net120),
    .B1(_0613_),
    .A1(_0496_),
    .Y(_0614_),
    .A2(_0609_));
 sg13g2_nor3_1 _1455_ (.A(_0565_),
    .B(_0580_),
    .C(_0596_),
    .Y(_0615_));
 sg13g2_a21oi_1 _1456_ (.A1(_0585_),
    .A2(_0586_),
    .Y(_0616_),
    .B1(_0615_));
 sg13g2_o21ai_1 _1457_ (.B1(_0616_),
    .Y(_0617_),
    .A1(_0557_),
    .A2(_0590_));
 sg13g2_xnor2_1 _1458_ (.Y(_0618_),
    .A(_0607_),
    .B(_0617_));
 sg13g2_o21ai_1 _1459_ (.B1(net153),
    .Y(_0619_),
    .A1(net118),
    .A2(_0618_));
 sg13g2_a21oi_1 _1460_ (.A1(_0611_),
    .A2(_0614_),
    .Y(_0044_),
    .B1(_0619_));
 sg13g2_and3_2 _1461_ (.X(_0620_),
    .A(net187),
    .B(\hvsync_gen.hpos[2] ),
    .C(_0126_));
 sg13g2_nor4_1 _1462_ (.A(\hvsync_gen.hpos[7] ),
    .B(net147),
    .C(\hvsync_gen.hpos[5] ),
    .D(_0146_),
    .Y(_0621_));
 sg13g2_nand3_1 _1463_ (.B(_0620_),
    .C(_0621_),
    .A(\hvsync_gen.hpos[4] ),
    .Y(_0622_));
 sg13g2_and2_1 _1464_ (.A(net153),
    .B(_0622_),
    .X(_0623_));
 sg13g2_nand2_1 _1465_ (.Y(_0624_),
    .A(net153),
    .B(_0622_));
 sg13g2_nand4_1 _1466_ (.B(\hvsync_gen.vpos[2] ),
    .C(_0108_),
    .A(\hvsync_gen.vpos[3] ),
    .Y(_0625_),
    .D(\hvsync_gen.vpos[9] ));
 sg13g2_nor4_1 _1467_ (.A(\hvsync_gen.vpos[0] ),
    .B(\hvsync_gen.vpos[8] ),
    .C(\hvsync_gen.vpos[7] ),
    .D(\hvsync_gen.vpos[4] ),
    .Y(_0626_));
 sg13g2_nor3_1 _1468_ (.A(\hvsync_gen.vpos[6] ),
    .B(\hvsync_gen.vpos[5] ),
    .C(_0625_),
    .Y(_0627_));
 sg13g2_a21oi_2 _1469_ (.B1(net150),
    .Y(_0628_),
    .A2(_0627_),
    .A1(_0626_));
 sg13g2_nand2b_2 _1470_ (.Y(_0629_),
    .B(_0628_),
    .A_N(_0622_));
 sg13g2_inv_1 _1471_ (.Y(_0630_),
    .A(_0629_));
 sg13g2_a22oi_1 _1472_ (.Y(_0631_),
    .B1(_0630_),
    .B2(net114),
    .A2(net131),
    .A1(\hvsync_gen.vpos[0] ));
 sg13g2_inv_1 _1473_ (.Y(_0045_),
    .A(net115));
 sg13g2_nor2_1 _1474_ (.A(\hvsync_gen.vpos[0] ),
    .B(net206),
    .Y(_0632_));
 sg13g2_nor3_1 _1475_ (.A(_0116_),
    .B(_0629_),
    .C(_0632_),
    .Y(_0633_));
 sg13g2_a21o_1 _1476_ (.A2(net131),
    .A1(net206),
    .B1(_0633_),
    .X(_0046_));
 sg13g2_xnor2_1 _1477_ (.Y(_0634_),
    .A(net237),
    .B(_0117_));
 sg13g2_nand2_1 _1478_ (.Y(_0635_),
    .A(net199),
    .B(net131));
 sg13g2_o21ai_1 _1479_ (.B1(_0635_),
    .Y(_0047_),
    .A1(_0629_),
    .A2(_0634_));
 sg13g2_a21oi_1 _1480_ (.A1(net199),
    .A2(_0116_),
    .Y(_0636_),
    .B1(net228));
 sg13g2_and3_2 _1481_ (.X(_0637_),
    .A(net239),
    .B(net199),
    .C(_0116_));
 sg13g2_nor3_1 _1482_ (.A(_0629_),
    .B(_0636_),
    .C(_0637_),
    .Y(_0638_));
 sg13g2_a21o_1 _1483_ (.A2(net131),
    .A1(net228),
    .B1(_0638_),
    .X(_0048_));
 sg13g2_nand2_1 _1484_ (.Y(_0639_),
    .A(\hvsync_gen.vpos[4] ),
    .B(_0637_));
 sg13g2_a21oi_2 _1485_ (.B1(net131),
    .Y(_0640_),
    .A2(_0639_),
    .A1(_0628_));
 sg13g2_a21oi_1 _1486_ (.A1(net130),
    .A2(_0637_),
    .Y(_0641_),
    .B1(net219));
 sg13g2_nor2_1 _1487_ (.A(_0640_),
    .B(_0641_),
    .Y(_0049_));
 sg13g2_nand4_1 _1488_ (.B(net219),
    .C(_0630_),
    .A(_0107_),
    .Y(_0642_),
    .D(_0637_));
 sg13g2_o21ai_1 _1489_ (.B1(_0642_),
    .Y(_0050_),
    .A1(_0107_),
    .A2(_0640_));
 sg13g2_nand4_1 _1490_ (.B(\hvsync_gen.vpos[5] ),
    .C(\hvsync_gen.vpos[4] ),
    .A(\hvsync_gen.vpos[6] ),
    .Y(_0643_),
    .D(_0637_));
 sg13g2_a21oi_1 _1491_ (.A1(_0628_),
    .A2(_0643_),
    .Y(_0644_),
    .B1(net131));
 sg13g2_nor3_1 _1492_ (.A(_0107_),
    .B(net131),
    .C(_0639_),
    .Y(_0645_));
 sg13g2_nor2_1 _1493_ (.A(net231),
    .B(_0645_),
    .Y(_0646_));
 sg13g2_nor2_1 _1494_ (.A(_0644_),
    .B(_0646_),
    .Y(_0051_));
 sg13g2_nor2_1 _1495_ (.A(_0629_),
    .B(_0643_),
    .Y(_0647_));
 sg13g2_nor2_1 _1496_ (.A(net217),
    .B(_0647_),
    .Y(_0648_));
 sg13g2_a21oi_1 _1497_ (.A1(net217),
    .A2(_0644_),
    .Y(_0052_),
    .B1(_0648_));
 sg13g2_nand3_1 _1498_ (.B(\hvsync_gen.vpos[6] ),
    .C(_0645_),
    .A(\hvsync_gen.vpos[7] ),
    .Y(_0649_));
 sg13g2_nand2_1 _1499_ (.Y(_0650_),
    .A(_0140_),
    .B(_0628_));
 sg13g2_a22oi_1 _1500_ (.Y(_0053_),
    .B1(_0650_),
    .B2(_0640_),
    .A2(_0649_),
    .A1(_0106_));
 sg13g2_nand2_1 _1501_ (.Y(_0651_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_0623_));
 sg13g2_nor3_1 _1502_ (.A(net211),
    .B(_0121_),
    .C(_0639_),
    .Y(_0652_));
 sg13g2_xnor2_1 _1503_ (.Y(_0653_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_0652_));
 sg13g2_o21ai_1 _1504_ (.B1(_0651_),
    .Y(_0054_),
    .A1(_0629_),
    .A2(net212));
 sg13g2_nor2_1 _1505_ (.A(_0109_),
    .B(_0025_),
    .Y(_0654_));
 sg13g2_xnor2_1 _1506_ (.Y(_0655_),
    .A(net148),
    .B(net183));
 sg13g2_nor2_1 _1507_ (.A(_0105_),
    .B(net184),
    .Y(_0055_));
 sg13g2_o21ai_1 _1508_ (.B1(net152),
    .Y(_0656_),
    .A1(net164),
    .A2(_0654_));
 sg13g2_a21oi_1 _1509_ (.A1(net164),
    .A2(_0654_),
    .Y(_0056_),
    .B1(_0656_));
 sg13g2_or2_1 _1510_ (.X(_0657_),
    .B(_0498_),
    .A(_0497_));
 sg13g2_a221oi_1 _1511_ (.B2(_0135_),
    .C1(net119),
    .B1(_0494_),
    .A1(net126),
    .Y(_0658_),
    .A2(_0483_));
 sg13g2_a221oi_1 _1512_ (.B2(_0658_),
    .C1(net149),
    .B1(_0657_),
    .A1(net119),
    .Y(_0057_),
    .A2(_0485_));
 sg13g2_nand2_1 _1513_ (.Y(_0659_),
    .A(_0125_),
    .B(_0525_));
 sg13g2_a221oi_1 _1514_ (.B2(net126),
    .C1(net119),
    .B1(_0518_),
    .A1(_0135_),
    .Y(_0660_),
    .A2(_0511_));
 sg13g2_a221oi_1 _1515_ (.B2(_0660_),
    .C1(net149),
    .B1(_0659_),
    .A1(net119),
    .Y(_0058_),
    .A2(_0521_));
 sg13g2_nor2_1 _1516_ (.A(_0136_),
    .B(_0536_),
    .Y(_0661_));
 sg13g2_nor2_1 _1517_ (.A(_0497_),
    .B(_0549_),
    .Y(_0662_));
 sg13g2_o21ai_1 _1518_ (.B1(net118),
    .Y(_0663_),
    .A1(net124),
    .A2(_0542_));
 sg13g2_nor3_1 _1519_ (.A(_0661_),
    .B(_0662_),
    .C(_0663_),
    .Y(_0664_));
 sg13g2_o21ai_1 _1520_ (.B1(net153),
    .Y(_0665_),
    .A1(net118),
    .A2(_0545_));
 sg13g2_nor2_1 _1521_ (.A(_0664_),
    .B(_0665_),
    .Y(_0059_));
 sg13g2_or2_1 _1522_ (.X(_0666_),
    .B(_0561_),
    .A(_0136_));
 sg13g2_nor2_1 _1523_ (.A(net128),
    .B(_0581_),
    .Y(_0667_));
 sg13g2_o21ai_1 _1524_ (.B1(_0138_),
    .Y(_0668_),
    .A1(net124),
    .A2(_0569_));
 sg13g2_nor2_1 _1525_ (.A(_0667_),
    .B(_0668_),
    .Y(_0669_));
 sg13g2_a221oi_1 _1526_ (.B2(_0669_),
    .C1(net150),
    .B1(_0666_),
    .A1(net120),
    .Y(_0060_),
    .A2(_0574_));
 sg13g2_or2_1 _1527_ (.X(_0670_),
    .B(_0593_),
    .A(_0136_));
 sg13g2_nor2_1 _1528_ (.A(_0134_),
    .B(_0599_),
    .Y(_0671_));
 sg13g2_o21ai_1 _1529_ (.B1(net118),
    .Y(_0672_),
    .A1(net127),
    .A2(_0606_));
 sg13g2_nor2_1 _1530_ (.A(_0671_),
    .B(_0672_),
    .Y(_0673_));
 sg13g2_a221oi_1 _1531_ (.B2(_0673_),
    .C1(net150),
    .B1(_0670_),
    .A1(net120),
    .Y(_0061_),
    .A2(_0602_));
 sg13g2_nand2_1 _1532_ (.Y(_0674_),
    .A(_0135_),
    .B(_0609_));
 sg13g2_o21ai_1 _1533_ (.B1(net118),
    .Y(_0675_),
    .A1(net124),
    .A2(_0610_));
 sg13g2_a21oi_1 _1534_ (.A1(_0496_),
    .A2(_0618_),
    .Y(_0676_),
    .B1(_0675_));
 sg13g2_a221oi_1 _1535_ (.B2(_0676_),
    .C1(net149),
    .B1(_0674_),
    .A1(net119),
    .Y(_0062_),
    .A2(_0613_));
 sg13g2_or3_1 _1536_ (.A(\cordicAlg.xv[0][3] ),
    .B(\cordicAlg.xv[0][1] ),
    .C(\cordicAlg.xv[0][2] ),
    .X(_0677_));
 sg13g2_or2_1 _1537_ (.X(_0678_),
    .B(_0677_),
    .A(\cordicAlg.xv[0][4] ));
 sg13g2_nor2_1 _1538_ (.A(\cordicAlg.xv[0][5] ),
    .B(_0678_),
    .Y(_0679_));
 sg13g2_a21oi_1 _1539_ (.A1(_0109_),
    .A2(_0679_),
    .Y(_0680_),
    .B1(\cordicAlg.xv[0][6] ));
 sg13g2_inv_1 _1540_ (.Y(_0681_),
    .A(_0680_));
 sg13g2_nor2_1 _1541_ (.A(\cordicAlg.yv[0][6] ),
    .B(_0679_),
    .Y(_0682_));
 sg13g2_o21ai_1 _1542_ (.B1(\cordicAlg.xv[0][6] ),
    .Y(_0683_),
    .A1(\cordicAlg.yv[0][6] ),
    .A2(_0679_));
 sg13g2_a22oi_1 _1543_ (.Y(_0684_),
    .B1(_0681_),
    .B2(_0683_),
    .A2(_0011_),
    .A1(net148));
 sg13g2_inv_1 _1544_ (.Y(_0685_),
    .A(_0684_));
 sg13g2_nand2_1 _1545_ (.Y(_0686_),
    .A(_0109_),
    .B(_0678_));
 sg13g2_a21oi_1 _1546_ (.A1(\cordicAlg.xv[0][4] ),
    .A2(_0677_),
    .Y(_0687_),
    .B1(_0686_));
 sg13g2_a21oi_1 _1547_ (.A1(net148),
    .A2(_0114_),
    .Y(_0688_),
    .B1(_0687_));
 sg13g2_nor2_1 _1548_ (.A(_0013_),
    .B(_0688_),
    .Y(_0689_));
 sg13g2_nand2_1 _1549_ (.Y(_0690_),
    .A(\cordicAlg.xv[0][1] ),
    .B(\cordicAlg.yv[0][0] ));
 sg13g2_xor2_1 _1550_ (.B(\cordicAlg.xv[0][2] ),
    .A(\cordicAlg.xv[0][1] ),
    .X(_0691_));
 sg13g2_nand2b_1 _1551_ (.Y(_0692_),
    .B(net148),
    .A_N(_0017_));
 sg13g2_o21ai_1 _1552_ (.B1(_0692_),
    .Y(_0693_),
    .A1(_0016_),
    .A2(_0690_));
 sg13g2_a21oi_1 _1553_ (.A1(_0109_),
    .A2(_0691_),
    .Y(_0694_),
    .B1(_0693_));
 sg13g2_a21oi_1 _1554_ (.A1(_0016_),
    .A2(_0690_),
    .Y(_0695_),
    .B1(_0694_));
 sg13g2_o21ai_1 _1555_ (.B1(\cordicAlg.xv[0][3] ),
    .Y(_0696_),
    .A1(\cordicAlg.xv[0][1] ),
    .A2(\cordicAlg.xv[0][2] ));
 sg13g2_a21oi_1 _1556_ (.A1(_0677_),
    .A2(_0696_),
    .Y(_0697_),
    .B1(net148));
 sg13g2_a21oi_1 _1557_ (.A1(net148),
    .A2(_0015_),
    .Y(_0698_),
    .B1(_0697_));
 sg13g2_o21ai_1 _1558_ (.B1(_0698_),
    .Y(_0699_),
    .A1(\cordicAlg.yv[0][2] ),
    .A2(_0695_));
 sg13g2_a21oi_1 _1559_ (.A1(\cordicAlg.yv[0][2] ),
    .A2(_0695_),
    .Y(_0700_),
    .B1(_0689_));
 sg13g2_nand2_1 _1560_ (.Y(_0701_),
    .A(\cordicAlg.xv[0][5] ),
    .B(_0678_));
 sg13g2_a22oi_1 _1561_ (.Y(_0702_),
    .B1(_0682_),
    .B2(_0701_),
    .A2(_0113_),
    .A1(net148));
 sg13g2_inv_1 _1562_ (.Y(_0703_),
    .A(_0702_));
 sg13g2_a22oi_1 _1563_ (.Y(_0704_),
    .B1(_0699_),
    .B2(_0700_),
    .A2(_0688_),
    .A1(_0013_));
 sg13g2_o21ai_1 _1564_ (.B1(_0704_),
    .Y(_0705_),
    .A1(\cordicAlg.yv[0][4] ),
    .A2(_0703_));
 sg13g2_a22oi_1 _1565_ (.Y(_0706_),
    .B1(_0703_),
    .B2(\cordicAlg.yv[0][4] ),
    .A2(_0684_),
    .A1(_0112_));
 sg13g2_a22oi_1 _1566_ (.Y(_0707_),
    .B1(_0705_),
    .B2(_0706_),
    .A2(_0685_),
    .A1(net203));
 sg13g2_o21ai_1 _1567_ (.B1(net152),
    .Y(_0708_),
    .A1(_0680_),
    .A2(net204));
 sg13g2_a21oi_1 _1568_ (.A1(_0680_),
    .A2(net204),
    .Y(_0063_),
    .B1(_0708_));
 sg13g2_and2_1 _1569_ (.A(net152),
    .B(net160),
    .X(_0064_));
 sg13g2_and2_1 _1570_ (.A(net152),
    .B(net155),
    .X(_0065_));
 sg13g2_and2_1 _1571_ (.A(net151),
    .B(net158),
    .X(_0066_));
 sg13g2_and2_1 _1572_ (.A(net151),
    .B(net157),
    .X(_0067_));
 sg13g2_nand2b_1 _1573_ (.Y(_0709_),
    .B(net179),
    .A_N(net168));
 sg13g2_nand2b_1 _1574_ (.Y(_0710_),
    .B(net168),
    .A_N(net179));
 sg13g2_a21oi_1 _1575_ (.A1(_0709_),
    .A2(_0710_),
    .Y(_0069_),
    .B1(net149));
 sg13g2_nor2_1 _1576_ (.A(\cordicAlg.ph[1][2] ),
    .B(_0709_),
    .Y(_0711_));
 sg13g2_xor2_1 _1577_ (.B(_0709_),
    .A(net193),
    .X(_0712_));
 sg13g2_nor2_1 _1578_ (.A(net149),
    .B(_0712_),
    .Y(_0070_));
 sg13g2_o21ai_1 _1579_ (.B1(net151),
    .Y(_0713_),
    .A1(net161),
    .A2(_0711_));
 sg13g2_a21oi_1 _1580_ (.A1(net161),
    .A2(_0711_),
    .Y(_0071_),
    .B1(_0713_));
 sg13g2_and2_1 _1581_ (.A(net151),
    .B(net168),
    .X(_0072_));
 sg13g2_and2_1 _1582_ (.A(net151),
    .B(net159),
    .X(_0073_));
 sg13g2_and2_1 _1583_ (.A(net151),
    .B(net163),
    .X(_0074_));
 sg13g2_and2_1 _1584_ (.A(net151),
    .B(net156),
    .X(_0075_));
 sg13g2_and2_1 _1585_ (.A(net112),
    .B(net131),
    .X(_0076_));
 sg13g2_nor2_1 _1586_ (.A(\hvsync_gen.hpos[0] ),
    .B(net190),
    .Y(_0714_));
 sg13g2_nor3_1 _1587_ (.A(_0126_),
    .B(net130),
    .C(net191),
    .Y(_0077_));
 sg13g2_xnor2_1 _1588_ (.Y(_0715_),
    .A(net235),
    .B(_0126_));
 sg13g2_nor2_1 _1589_ (.A(net130),
    .B(_0715_),
    .Y(_0078_));
 sg13g2_a21oi_1 _1590_ (.A1(\hvsync_gen.hpos[2] ),
    .A2(_0126_),
    .Y(_0716_),
    .B1(net187));
 sg13g2_nor3_1 _1591_ (.A(net150),
    .B(_0620_),
    .C(net188),
    .Y(_0079_));
 sg13g2_xor2_1 _1592_ (.B(_0620_),
    .A(net222),
    .X(_0717_));
 sg13g2_nor2_1 _1593_ (.A(_0624_),
    .B(net223),
    .Y(_0080_));
 sg13g2_a21oi_1 _1594_ (.A1(\hvsync_gen.hpos[4] ),
    .A2(_0620_),
    .Y(_0718_),
    .B1(net224));
 sg13g2_and3_1 _1595_ (.X(_0719_),
    .A(\hvsync_gen.hpos[4] ),
    .B(\hvsync_gen.hpos[5] ),
    .C(_0620_));
 sg13g2_nor3_1 _1596_ (.A(net130),
    .B(net225),
    .C(_0719_),
    .Y(_0081_));
 sg13g2_a21oi_1 _1597_ (.A1(net147),
    .A2(_0719_),
    .Y(_0720_),
    .B1(net130));
 sg13g2_o21ai_1 _1598_ (.B1(_0720_),
    .Y(_0721_),
    .A1(net147),
    .A2(_0719_));
 sg13g2_inv_1 _1599_ (.Y(_0082_),
    .A(_0721_));
 sg13g2_a21oi_1 _1600_ (.A1(net147),
    .A2(_0719_),
    .Y(_0722_),
    .B1(net220));
 sg13g2_and3_1 _1601_ (.X(_0723_),
    .A(\hvsync_gen.hpos[7] ),
    .B(net147),
    .C(_0719_));
 sg13g2_nor3_1 _1602_ (.A(net130),
    .B(net221),
    .C(_0723_),
    .Y(_0083_));
 sg13g2_xnor2_1 _1603_ (.Y(_0724_),
    .A(net232),
    .B(_0723_));
 sg13g2_nor2_1 _1604_ (.A(net130),
    .B(_0724_),
    .Y(_0084_));
 sg13g2_a21oi_1 _1605_ (.A1(\hvsync_gen.hpos[8] ),
    .A2(_0723_),
    .Y(_0725_),
    .B1(net226));
 sg13g2_nor2b_1 _1606_ (.A(_0146_),
    .B_N(_0723_),
    .Y(_0726_));
 sg13g2_nor3_1 _1607_ (.A(net130),
    .B(net227),
    .C(_0726_),
    .Y(_0085_));
 sg13g2_nand2_1 _1608_ (.Y(_0727_),
    .A(net236),
    .B(net152));
 sg13g2_xnor2_1 _1609_ (.Y(_0728_),
    .A(net127),
    .B(_0634_));
 sg13g2_xnor2_1 _1610_ (.Y(_0729_),
    .A(net126),
    .B(_0715_));
 sg13g2_nand2_1 _1611_ (.Y(_0730_),
    .A(net139),
    .B(_0729_));
 sg13g2_o21ai_1 _1612_ (.B1(_0730_),
    .Y(_0086_),
    .A1(net135),
    .A2(_0728_));
 sg13g2_xnor2_1 _1613_ (.Y(_0731_),
    .A(net127),
    .B(_0472_));
 sg13g2_xnor2_1 _1614_ (.Y(_0732_),
    .A(net125),
    .B(_0469_));
 sg13g2_nand2_1 _1615_ (.Y(_0733_),
    .A(net139),
    .B(_0732_));
 sg13g2_o21ai_1 _1616_ (.B1(_0733_),
    .Y(_0087_),
    .A1(net135),
    .A2(_0731_));
 sg13g2_o21ai_1 _1617_ (.B1(net139),
    .Y(_0734_),
    .A1(net125),
    .A2(_0477_));
 sg13g2_a21o_1 _1618_ (.A2(_0477_),
    .A1(net125),
    .B1(_0734_),
    .X(_0735_));
 sg13g2_xnor2_1 _1619_ (.Y(_0736_),
    .A(net127),
    .B(_0475_));
 sg13g2_o21ai_1 _1620_ (.B1(_0735_),
    .Y(_0088_),
    .A1(net135),
    .A2(_0736_));
 sg13g2_xnor2_1 _1621_ (.Y(_0737_),
    .A(net127),
    .B(_0500_));
 sg13g2_or2_1 _1622_ (.X(_0738_),
    .B(_0503_),
    .A(net126));
 sg13g2_nand2_1 _1623_ (.Y(_0739_),
    .A(net126),
    .B(_0503_));
 sg13g2_nand3_1 _1624_ (.B(_0738_),
    .C(_0739_),
    .A(net139),
    .Y(_0740_));
 sg13g2_o21ai_1 _1625_ (.B1(_0740_),
    .Y(_0089_),
    .A1(net135),
    .A2(_0737_));
 sg13g2_xnor2_1 _1626_ (.Y(_0741_),
    .A(_0125_),
    .B(_0527_));
 sg13g2_xnor2_1 _1627_ (.Y(_0742_),
    .A(net126),
    .B(_0528_));
 sg13g2_nand2_1 _1628_ (.Y(_0743_),
    .A(net139),
    .B(_0742_));
 sg13g2_o21ai_1 _1629_ (.B1(_0743_),
    .Y(_0090_),
    .A1(net135),
    .A2(_0741_));
 sg13g2_o21ai_1 _1630_ (.B1(net139),
    .Y(_0744_),
    .A1(net125),
    .A2(_0553_));
 sg13g2_a21oi_1 _1631_ (.A1(net125),
    .A2(_0553_),
    .Y(_0745_),
    .B1(_0744_));
 sg13g2_a21oi_1 _1632_ (.A1(net127),
    .A2(_0552_),
    .Y(_0746_),
    .B1(net135));
 sg13g2_o21ai_1 _1633_ (.B1(_0746_),
    .Y(_0747_),
    .A1(net127),
    .A2(_0552_));
 sg13g2_nand2b_1 _1634_ (.Y(_0091_),
    .B(_0747_),
    .A_N(_0745_));
 sg13g2_o21ai_1 _1635_ (.B1(net139),
    .Y(_0748_),
    .A1(\hvsync_gen.hpos[9] ),
    .A2(_0582_));
 sg13g2_a21o_1 _1636_ (.A2(_0582_),
    .A1(\hvsync_gen.hpos[9] ),
    .B1(_0748_),
    .X(_0749_));
 sg13g2_xnor2_1 _1637_ (.Y(_0750_),
    .A(_0125_),
    .B(_0587_));
 sg13g2_o21ai_1 _1638_ (.B1(_0749_),
    .Y(_0092_),
    .A1(net135),
    .A2(_0750_));
 sg13g2_and2_1 _1639_ (.A(net152),
    .B(net113),
    .X(_0093_));
 sg13g2_nand2_1 _1640_ (.Y(_0751_),
    .A(net166),
    .B(net133));
 sg13g2_o21ai_1 _1641_ (.B1(_0751_),
    .Y(_0094_),
    .A1(_0309_),
    .A2(net133));
 sg13g2_nand2_1 _1642_ (.Y(_0752_),
    .A(net170),
    .B(net133));
 sg13g2_o21ai_1 _1643_ (.B1(_0752_),
    .Y(_0095_),
    .A1(_0313_),
    .A2(net133));
 sg13g2_nand2_1 _1644_ (.Y(_0753_),
    .A(net172),
    .B(net132));
 sg13g2_o21ai_1 _1645_ (.B1(_0753_),
    .Y(_0096_),
    .A1(_0323_),
    .A2(net132));
 sg13g2_nand2_1 _1646_ (.Y(_0754_),
    .A(net169),
    .B(net132));
 sg13g2_o21ai_1 _1647_ (.B1(_0754_),
    .Y(_0097_),
    .A1(_0342_),
    .A2(net132));
 sg13g2_nand2_1 _1648_ (.Y(_0755_),
    .A(net176),
    .B(net132));
 sg13g2_o21ai_1 _1649_ (.B1(_0755_),
    .Y(_0098_),
    .A1(_0390_),
    .A2(net132));
 sg13g2_nand2_1 _1650_ (.Y(_0756_),
    .A(net177),
    .B(net132));
 sg13g2_o21ai_1 _1651_ (.B1(_0756_),
    .Y(_0099_),
    .A1(_0407_),
    .A2(net132));
 sg13g2_nand2_1 _1652_ (.Y(_0757_),
    .A(net186),
    .B(net133));
 sg13g2_o21ai_1 _1653_ (.B1(_0757_),
    .Y(_0100_),
    .A1(_0426_),
    .A2(net133));
 sg13g2_nand2_1 _1654_ (.Y(_0758_),
    .A(net197),
    .B(net134));
 sg13g2_o21ai_1 _1655_ (.B1(_0758_),
    .Y(_0101_),
    .A1(_0440_),
    .A2(net134));
 sg13g2_nand2_1 _1656_ (.Y(_0759_),
    .A(net198),
    .B(net134));
 sg13g2_o21ai_1 _1657_ (.B1(_0759_),
    .Y(_0102_),
    .A1(_0457_),
    .A2(net134));
 sg13g2_nand2_1 _1658_ (.Y(_0760_),
    .A(net185),
    .B(net134));
 sg13g2_o21ai_1 _1659_ (.B1(_0760_),
    .Y(_0103_),
    .A1(_0462_),
    .A2(net134));
 sg13g2_mux2_1 _1660_ (.A0(_0468_),
    .A1(net209),
    .S(net134),
    .X(_0104_));
 sg13g2_buf_1 _1661_ (.A(net152),
    .X(_0002_));
 sg13g2_buf_1 _1662_ (.A(net151),
    .X(_0068_));
 sg13g2_dfrbp_1 _1663_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net36),
    .D(net174),
    .Q_N(_0820_),
    .Q(\hypotenuse.multY[2] ));
 sg13g2_dfrbp_1 _1664_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net63),
    .D(net181),
    .Q_N(_0819_),
    .Q(\hypotenuse.multY[3] ));
 sg13g2_dfrbp_1 _1665_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net62),
    .D(_0029_),
    .Q_N(_0818_),
    .Q(\hypotenuse.multY[4] ));
 sg13g2_dfrbp_1 _1666_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net60),
    .D(_0030_),
    .Q_N(_0817_),
    .Q(\hypotenuse.multY[5] ));
 sg13g2_dfrbp_1 _1667_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net59),
    .D(_0031_),
    .Q_N(_0816_),
    .Q(\hypotenuse.multY[6] ));
 sg13g2_dfrbp_1 _1668_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net58),
    .D(_0032_),
    .Q_N(_0815_),
    .Q(\hypotenuse.multY[7] ));
 sg13g2_dfrbp_1 _1669_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net57),
    .D(_0033_),
    .Q_N(_0814_),
    .Q(\hypotenuse.multY[8] ));
 sg13g2_dfrbp_1 _1670_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net56),
    .D(_0034_),
    .Q_N(_0813_),
    .Q(\hypotenuse.multY[9] ));
 sg13g2_dfrbp_1 _1671_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net55),
    .D(_0035_),
    .Q_N(_0812_),
    .Q(\hypotenuse.multY[10] ));
 sg13g2_dfrbp_1 _1672_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net54),
    .D(_0036_),
    .Q_N(_0811_),
    .Q(\hypotenuse.multY[11] ));
 sg13g2_dfrbp_1 _1673_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net37),
    .D(net196),
    .Q_N(_0821_),
    .Q(\hypotenuse.multY[12] ));
 sg13g2_dfrbp_1 _1674_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net38),
    .D(_0002_),
    .Q_N(_0822_),
    .Q(_0025_));
 sg13g2_dfrbp_1 _1675_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net39),
    .D(_0000_),
    .Q_N(_0823_),
    .Q(_0026_));
 sg13g2_dfrbp_1 _1676_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net40),
    .D(_0020_),
    .Q_N(_0824_),
    .Q(\angleOffset[0] ));
 sg13g2_dfrbp_1 _1677_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net41),
    .D(_0021_),
    .Q_N(_0825_),
    .Q(\angleOffset[1] ));
 sg13g2_dfrbp_1 _1678_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net42),
    .D(_0022_),
    .Q_N(_0826_),
    .Q(\angleOffset[2] ));
 sg13g2_dfrbp_1 _1679_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net50),
    .D(_0023_),
    .Q_N(_0827_),
    .Q(\angleOffset[3] ));
 sg13g2_dfrbp_1 _1680_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net53),
    .D(_0024_),
    .Q_N(_0810_),
    .Q(\angleOffset[4] ));
 sg13g2_dfrbp_1 _1681_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net52),
    .D(_0038_),
    .Q_N(_0809_),
    .Q(\cordicAlg.yv[0][0] ));
 sg13g2_dfrbp_1 _1682_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net51),
    .D(_0039_),
    .Q_N(_0016_),
    .Q(\cordicAlg.yv[0][1] ));
 sg13g2_dfrbp_1 _1683_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net49),
    .D(_0040_),
    .Q_N(_0808_),
    .Q(\cordicAlg.yv[0][2] ));
 sg13g2_dfrbp_1 _1684_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net48),
    .D(_0041_),
    .Q_N(_0013_),
    .Q(\cordicAlg.yv[0][3] ));
 sg13g2_dfrbp_1 _1685_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net47),
    .D(_0042_),
    .Q_N(_0807_),
    .Q(\cordicAlg.yv[0][4] ));
 sg13g2_dfrbp_1 _1686_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net46),
    .D(_0043_),
    .Q_N(_0010_),
    .Q(\cordicAlg.yv[0][5] ));
 sg13g2_dfrbp_1 _1687_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net61),
    .D(_0044_),
    .Q_N(_0828_),
    .Q(\cordicAlg.yv[0][6] ));
 sg13g2_dfrbp_1 _1688_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net45),
    .D(net154),
    .Q_N(_0806_),
    .Q(hsync));
 sg13g2_dfrbp_1 _1689_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net44),
    .D(_0045_),
    .Q_N(\hypotenuse.y_pos[0] ),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _1690_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net35),
    .D(net207),
    .Q_N(_0805_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _1691_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net33),
    .D(net200),
    .Q_N(_0008_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _1692_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net31),
    .D(_0048_),
    .Q_N(_0804_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _1693_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net29),
    .D(_0049_),
    .Q_N(_0803_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _1694_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net27),
    .D(net230),
    .Q_N(_0802_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _1695_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net25),
    .D(_0051_),
    .Q_N(_0801_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _1696_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net110),
    .D(net218),
    .Q_N(_0800_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _1697_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net108),
    .D(net216),
    .Q_N(_0005_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _1698_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net105),
    .D(net213),
    .Q_N(_0829_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _1699_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net106),
    .D(net234),
    .Q_N(_0799_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 _1700_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net104),
    .D(_0055_),
    .Q_N(_0798_),
    .Q(\cordicAlg.ph[1][2] ));
 sg13g2_dfrbp_1 _1701_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net103),
    .D(net165),
    .Q_N(_0797_),
    .Q(\cordicAlg.ph[1][3] ));
 sg13g2_dfrbp_1 _1702_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net102),
    .D(_0057_),
    .Q_N(_0796_),
    .Q(\cordicAlg.xv[0][1] ));
 sg13g2_dfrbp_1 _1703_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net101),
    .D(_0058_),
    .Q_N(_0017_),
    .Q(\cordicAlg.xv[0][2] ));
 sg13g2_dfrbp_1 _1704_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net100),
    .D(_0059_),
    .Q_N(_0015_),
    .Q(\cordicAlg.xv[0][3] ));
 sg13g2_dfrbp_1 _1705_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net99),
    .D(_0060_),
    .Q_N(_0014_),
    .Q(\cordicAlg.xv[0][4] ));
 sg13g2_dfrbp_1 _1706_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net98),
    .D(_0061_),
    .Q_N(_0012_),
    .Q(\cordicAlg.xv[0][5] ));
 sg13g2_dfrbp_1 _1707_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net97),
    .D(_0062_),
    .Q_N(_0011_),
    .Q(\cordicAlg.xv[0][6] ));
 sg13g2_dfrbp_1 _1708_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net96),
    .D(net205),
    .Q_N(_0795_),
    .Q(\cordicAlg.yv[1][6] ));
 sg13g2_dfrbp_1 _1709_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net95),
    .D(_0064_),
    .Q_N(_0794_),
    .Q(\angle[0] ));
 sg13g2_dfrbp_1 _1710_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net94),
    .D(_0065_),
    .Q_N(_0793_),
    .Q(\angle[1] ));
 sg13g2_dfrbp_1 _1711_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net93),
    .D(_0066_),
    .Q_N(_0792_),
    .Q(\angle[2] ));
 sg13g2_dfrbp_1 _1712_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net92),
    .D(_0067_),
    .Q_N(_0791_),
    .Q(\angle[3] ));
 sg13g2_dfrbp_1 _1713_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net91),
    .D(_0068_),
    .Q_N(_0790_),
    .Q(\cordicAlg.ph[1][1] ));
 sg13g2_dfrbp_1 _1714_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net90),
    .D(_0069_),
    .Q_N(_0789_),
    .Q(\cordicAlg.ph[2][1] ));
 sg13g2_dfrbp_1 _1715_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net89),
    .D(_0070_),
    .Q_N(_0788_),
    .Q(\cordicAlg.ph[2][2] ));
 sg13g2_dfrbp_1 _1716_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net88),
    .D(net162),
    .Q_N(_0787_),
    .Q(\cordicAlg.ph[2][3] ));
 sg13g2_dfrbp_1 _1717_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net87),
    .D(_0072_),
    .Q_N(_0786_),
    .Q(\cordicAlg.ph[3][0] ));
 sg13g2_dfrbp_1 _1718_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net86),
    .D(_0073_),
    .Q_N(_0785_),
    .Q(\cordicAlg.ph[3][1] ));
 sg13g2_dfrbp_1 _1719_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net85),
    .D(_0074_),
    .Q_N(_0784_),
    .Q(\cordicAlg.ph[3][2] ));
 sg13g2_dfrbp_1 _1720_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net84),
    .D(_0075_),
    .Q_N(_0783_),
    .Q(\cordicAlg.ph[3][3] ));
 sg13g2_dfrbp_1 _1721_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net83),
    .D(_0076_),
    .Q_N(\hypotenuse.x_pos[0] ),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 _1722_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net82),
    .D(net192),
    .Q_N(_0782_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _1723_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net81),
    .D(_0078_),
    .Q_N(_0781_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _1724_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net80),
    .D(net189),
    .Q_N(_0780_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _1725_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net79),
    .D(_0080_),
    .Q_N(_0009_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _1726_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net78),
    .D(_0081_),
    .Q_N(_0779_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _1727_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net77),
    .D(_0082_),
    .Q_N(_0778_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _1728_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net76),
    .D(_0083_),
    .Q_N(_0006_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _1729_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net75),
    .D(_0084_),
    .Q_N(_0777_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _1730_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net74),
    .D(_0085_),
    .Q_N(_0007_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _1731_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net73),
    .D(_0086_),
    .Q_N(_0776_),
    .Q(\hypotenuse.multSignal[0] ));
 sg13g2_dfrbp_1 _1732_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net72),
    .D(_0087_),
    .Q_N(_0018_),
    .Q(\hypotenuse.mutlReg[1] ));
 sg13g2_dfrbp_1 _1733_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net71),
    .D(_0088_),
    .Q_N(_0775_),
    .Q(\hypotenuse.mutlReg[2] ));
 sg13g2_dfrbp_1 _1734_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net70),
    .D(_0089_),
    .Q_N(_0774_),
    .Q(\hypotenuse.mutlReg[3] ));
 sg13g2_dfrbp_1 _1735_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net69),
    .D(_0090_),
    .Q_N(_0019_),
    .Q(\hypotenuse.mutlReg[4] ));
 sg13g2_dfrbp_1 _1736_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net68),
    .D(_0091_),
    .Q_N(_0773_),
    .Q(\hypotenuse.mutlReg[5] ));
 sg13g2_dfrbp_1 _1737_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net67),
    .D(_0092_),
    .Q_N(_0772_),
    .Q(\hypotenuse.mutlReg[6] ));
 sg13g2_dfrbp_1 _1738_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net66),
    .D(_0093_),
    .Q_N(_0001_),
    .Q(\hypotenuse.stateCheck ));
 sg13g2_dfrbp_1 _1739_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net65),
    .D(net167),
    .Q_N(_0771_),
    .Q(\hypotenuse.multX[2] ));
 sg13g2_dfrbp_1 _1740_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net64),
    .D(net171),
    .Q_N(_0770_),
    .Q(\hypotenuse.multX[3] ));
 sg13g2_dfrbp_1 _1741_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net43),
    .D(_0096_),
    .Q_N(_0769_),
    .Q(\hypotenuse.multX[4] ));
 sg13g2_dfrbp_1 _1742_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net34),
    .D(_0097_),
    .Q_N(_0768_),
    .Q(\hypotenuse.multX[5] ));
 sg13g2_dfrbp_1 _1743_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net32),
    .D(_0098_),
    .Q_N(_0767_),
    .Q(\hypotenuse.multX[6] ));
 sg13g2_dfrbp_1 _1744_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net30),
    .D(_0099_),
    .Q_N(_0766_),
    .Q(\hypotenuse.multX[7] ));
 sg13g2_dfrbp_1 _1745_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net28),
    .D(_0100_),
    .Q_N(_0765_),
    .Q(\hypotenuse.multX[8] ));
 sg13g2_dfrbp_1 _1746_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net26),
    .D(_0101_),
    .Q_N(_0764_),
    .Q(\hypotenuse.multX[9] ));
 sg13g2_dfrbp_1 _1747_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net111),
    .D(_0102_),
    .Q_N(_0763_),
    .Q(\hypotenuse.multX[10] ));
 sg13g2_dfrbp_1 _1748_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net109),
    .D(_0103_),
    .Q_N(_0762_),
    .Q(\hypotenuse.multX[11] ));
 sg13g2_dfrbp_1 _1749_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net107),
    .D(net210),
    .Q_N(_0761_),
    .Q(\hypotenuse.multX[12] ));
 sg13g2_tiehi _1746__26 (.L_HI(net26));
 sg13g2_tiehi _1694__27 (.L_HI(net27));
 sg13g2_tiehi _1745__28 (.L_HI(net28));
 sg13g2_tiehi _1693__29 (.L_HI(net29));
 sg13g2_tiehi _1744__30 (.L_HI(net30));
 sg13g2_tiehi _1692__31 (.L_HI(net31));
 sg13g2_tiehi _1743__32 (.L_HI(net32));
 sg13g2_tiehi _1691__33 (.L_HI(net33));
 sg13g2_tiehi _1742__34 (.L_HI(net34));
 sg13g2_tiehi _1690__35 (.L_HI(net35));
 sg13g2_tiehi _1663__36 (.L_HI(net36));
 sg13g2_tiehi _1673__37 (.L_HI(net37));
 sg13g2_tiehi _1674__38 (.L_HI(net38));
 sg13g2_tiehi _1675__39 (.L_HI(net39));
 sg13g2_tiehi _1676__40 (.L_HI(net40));
 sg13g2_tiehi _1677__41 (.L_HI(net41));
 sg13g2_tiehi _1678__42 (.L_HI(net42));
 sg13g2_tiehi _1741__43 (.L_HI(net43));
 sg13g2_tiehi _1689__44 (.L_HI(net44));
 sg13g2_tiehi _1688__45 (.L_HI(net45));
 sg13g2_tiehi _1686__46 (.L_HI(net46));
 sg13g2_tiehi _1685__47 (.L_HI(net47));
 sg13g2_tiehi _1684__48 (.L_HI(net48));
 sg13g2_tiehi _1683__49 (.L_HI(net49));
 sg13g2_tiehi _1679__50 (.L_HI(net50));
 sg13g2_tiehi _1682__51 (.L_HI(net51));
 sg13g2_tiehi _1681__52 (.L_HI(net52));
 sg13g2_tiehi _1680__53 (.L_HI(net53));
 sg13g2_tiehi _1672__54 (.L_HI(net54));
 sg13g2_tiehi _1671__55 (.L_HI(net55));
 sg13g2_tiehi _1670__56 (.L_HI(net56));
 sg13g2_tiehi _1669__57 (.L_HI(net57));
 sg13g2_tiehi _1668__58 (.L_HI(net58));
 sg13g2_tiehi _1667__59 (.L_HI(net59));
 sg13g2_tiehi _1666__60 (.L_HI(net60));
 sg13g2_tiehi _1687__61 (.L_HI(net61));
 sg13g2_tiehi _1665__62 (.L_HI(net62));
 sg13g2_tiehi _1664__63 (.L_HI(net63));
 sg13g2_tiehi _1740__64 (.L_HI(net64));
 sg13g2_tiehi _1739__65 (.L_HI(net65));
 sg13g2_tiehi _1738__66 (.L_HI(net66));
 sg13g2_tiehi _1737__67 (.L_HI(net67));
 sg13g2_tiehi _1736__68 (.L_HI(net68));
 sg13g2_tiehi _1735__69 (.L_HI(net69));
 sg13g2_tiehi _1734__70 (.L_HI(net70));
 sg13g2_tiehi _1733__71 (.L_HI(net71));
 sg13g2_tiehi _1732__72 (.L_HI(net72));
 sg13g2_tiehi _1731__73 (.L_HI(net73));
 sg13g2_tiehi _1730__74 (.L_HI(net74));
 sg13g2_tiehi _1729__75 (.L_HI(net75));
 sg13g2_tiehi _1728__76 (.L_HI(net76));
 sg13g2_tiehi _1727__77 (.L_HI(net77));
 sg13g2_tiehi _1726__78 (.L_HI(net78));
 sg13g2_tiehi _1725__79 (.L_HI(net79));
 sg13g2_tiehi _1724__80 (.L_HI(net80));
 sg13g2_tiehi _1723__81 (.L_HI(net81));
 sg13g2_tiehi _1722__82 (.L_HI(net82));
 sg13g2_tiehi _1721__83 (.L_HI(net83));
 sg13g2_tiehi _1720__84 (.L_HI(net84));
 sg13g2_tiehi _1719__85 (.L_HI(net85));
 sg13g2_tiehi _1718__86 (.L_HI(net86));
 sg13g2_tiehi _1717__87 (.L_HI(net87));
 sg13g2_tiehi _1716__88 (.L_HI(net88));
 sg13g2_tiehi _1715__89 (.L_HI(net89));
 sg13g2_tiehi _1714__90 (.L_HI(net90));
 sg13g2_tiehi _1713__91 (.L_HI(net91));
 sg13g2_tiehi _1712__92 (.L_HI(net92));
 sg13g2_tiehi _1711__93 (.L_HI(net93));
 sg13g2_tiehi _1710__94 (.L_HI(net94));
 sg13g2_tiehi _1709__95 (.L_HI(net95));
 sg13g2_tiehi _1708__96 (.L_HI(net96));
 sg13g2_tiehi _1707__97 (.L_HI(net97));
 sg13g2_tiehi _1706__98 (.L_HI(net98));
 sg13g2_tiehi _1705__99 (.L_HI(net99));
 sg13g2_tiehi _1704__100 (.L_HI(net100));
 sg13g2_tiehi _1703__101 (.L_HI(net101));
 sg13g2_tiehi _1702__102 (.L_HI(net102));
 sg13g2_tiehi _1701__103 (.L_HI(net103));
 sg13g2_tiehi _1700__104 (.L_HI(net104));
 sg13g2_tiehi _1698__105 (.L_HI(net105));
 sg13g2_tiehi _1699__106 (.L_HI(net106));
 sg13g2_tiehi _1749__107 (.L_HI(net107));
 sg13g2_tiehi _1697__108 (.L_HI(net108));
 sg13g2_tiehi _1748__109 (.L_HI(net109));
 sg13g2_tiehi _1696__110 (.L_HI(net110));
 sg13g2_tiehi _1747__111 (.L_HI(net111));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_rkarl_Spiral_10 (.L_LO(net10));
 sg13g2_tielo tt_um_rkarl_Spiral_11 (.L_LO(net11));
 sg13g2_tielo tt_um_rkarl_Spiral_12 (.L_LO(net12));
 sg13g2_tielo tt_um_rkarl_Spiral_13 (.L_LO(net13));
 sg13g2_tielo tt_um_rkarl_Spiral_14 (.L_LO(net14));
 sg13g2_tielo tt_um_rkarl_Spiral_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rkarl_Spiral_16 (.L_LO(net16));
 sg13g2_tielo tt_um_rkarl_Spiral_17 (.L_LO(net17));
 sg13g2_tielo tt_um_rkarl_Spiral_18 (.L_LO(net18));
 sg13g2_tielo tt_um_rkarl_Spiral_19 (.L_LO(net19));
 sg13g2_tielo tt_um_rkarl_Spiral_20 (.L_LO(net20));
 sg13g2_tielo tt_um_rkarl_Spiral_21 (.L_LO(net21));
 sg13g2_tielo tt_um_rkarl_Spiral_22 (.L_LO(net22));
 sg13g2_tielo tt_um_rkarl_Spiral_23 (.L_LO(net23));
 sg13g2_tielo tt_um_rkarl_Spiral_24 (.L_LO(net24));
 sg13g2_tiehi _1695__25 (.L_HI(net25));
 sg13g2_buf_1 _1853_ (.A(uo_out[4]),
    .X(uo_out[0]));
 sg13g2_buf_1 _1854_ (.A(uo_out[5]),
    .X(uo_out[1]));
 sg13g2_buf_1 _1855_ (.A(uo_out[6]),
    .X(uo_out[2]));
 sg13g2_buf_1 _1856_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1857_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout118 (.A(_0138_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_0137_),
    .X(net119));
 sg13g2_buf_1 fanout120 (.A(_0137_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_0185_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(net123),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_0178_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(net125),
    .X(net124));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(_0134_));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(_0133_));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(_0124_));
 sg13g2_buf_2 fanout128 (.A(_0124_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_0175_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_0624_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_0623_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(net133),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(net135),
    .X(net134));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(_0727_));
 sg13g2_buf_2 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(net138),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(_0308_));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(\hypotenuse.mutlReg[6] ));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(\hypotenuse.mutlReg[5] ));
 sg13g2_buf_2 fanout142 (.A(\hypotenuse.mutlReg[4] ),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(\hypotenuse.mutlReg[2] ),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(\hypotenuse.mutlReg[1] ),
    .X(net144));
 sg13g2_buf_1 fanout145 (.A(\hypotenuse.mutlReg[1] ),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(\hypotenuse.multSignal[0] ),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(net238),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(\cordicAlg.yv[0][6] ),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(_0105_));
 sg13g2_buf_2 fanout151 (.A(net153),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(net153),
    .X(net152));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_rkarl_Spiral_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\hypotenuse.x_pos[0] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0001_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold3 (.A(\hypotenuse.y_pos[0] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0631_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0007_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0145_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0003_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold8 (.A(\cordicAlg.ph[3][1] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold9 (.A(\cordicAlg.ph[2][3] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cordicAlg.ph[3][3] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold11 (.A(\cordicAlg.ph[3][2] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold12 (.A(\cordicAlg.ph[2][1] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold13 (.A(\cordicAlg.ph[3][0] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold14 (.A(\cordicAlg.ph[1][3] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0071_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold16 (.A(\cordicAlg.ph[2][2] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0026_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0056_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold19 (.A(\hypotenuse.multX[2] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0094_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold21 (.A(\cordicAlg.ph[1][1] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold22 (.A(\hypotenuse.multX[5] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold23 (.A(\hypotenuse.multX[3] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0095_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold25 (.A(\hypotenuse.multX[4] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold26 (.A(\hypotenuse.multY[2] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0027_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold28 (.A(\hypotenuse.multY[4] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold29 (.A(\hypotenuse.multX[6] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold30 (.A(\hypotenuse.multX[7] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold31 (.A(\hypotenuse.multY[5] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold32 (.A(\cordicAlg.yv[1][6] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold33 (.A(\hypotenuse.multY[3] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0028_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold35 (.A(\hypotenuse.multY[6] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0025_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0655_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold38 (.A(\hypotenuse.multX[11] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold39 (.A(\hypotenuse.multX[8] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold40 (.A(\hvsync_gen.hpos[3] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0716_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0079_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold43 (.A(\hvsync_gen.hpos[1] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0714_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0077_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold46 (.A(\cordicAlg.ph[1][2] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold47 (.A(\hypotenuse.multY[7] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold48 (.A(\hypotenuse.multY[12] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0037_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold50 (.A(\hypotenuse.multX[9] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold51 (.A(\hypotenuse.multX[10] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold52 (.A(\hvsync_gen.vpos[2] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0047_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold54 (.A(\hypotenuse.multY[8] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold55 (.A(\hypotenuse.multY[11] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0010_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0707_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0063_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold59 (.A(\hvsync_gen.vpos[1] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0046_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold61 (.A(\hypotenuse.multY[9] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold62 (.A(\hypotenuse.multX[12] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0104_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0005_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0653_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0054_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold67 (.A(\hypotenuse.multY[10] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold68 (.A(\hvsync_gen.vpos[8] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0053_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold70 (.A(\hvsync_gen.vpos[7] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0052_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold72 (.A(\hvsync_gen.vpos[4] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold73 (.A(\hvsync_gen.hpos[7] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0722_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0009_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0717_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold77 (.A(\hvsync_gen.hpos[5] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0718_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold79 (.A(\hvsync_gen.hpos[9] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0725_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold81 (.A(\hvsync_gen.vpos[3] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold82 (.A(\hvsync_gen.vpos[5] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0050_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold84 (.A(\hvsync_gen.vpos[6] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold85 (.A(\hvsync_gen.hpos[8] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold86 (.A(\hvsync_gen.vpos[9] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0004_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold88 (.A(\hvsync_gen.hpos[2] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold89 (.A(\hypotenuse.stateCheck ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0008_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold91 (.A(\hvsync_gen.hpos[6] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold92 (.A(\hvsync_gen.vpos[3] ),
    .X(net239));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_fill_1 FILLER_12_187 ();
 sg13g2_decap_8 FILLER_12_198 ();
 sg13g2_decap_4 FILLER_12_205 ();
 sg13g2_fill_1 FILLER_12_209 ();
 sg13g2_decap_8 FILLER_12_215 ();
 sg13g2_decap_4 FILLER_12_222 ();
 sg13g2_fill_2 FILLER_12_226 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_253 ();
 sg13g2_decap_8 FILLER_12_260 ();
 sg13g2_decap_4 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_271 ();
 sg13g2_decap_4 FILLER_12_277 ();
 sg13g2_fill_1 FILLER_12_281 ();
 sg13g2_decap_8 FILLER_12_286 ();
 sg13g2_decap_8 FILLER_12_293 ();
 sg13g2_decap_8 FILLER_12_300 ();
 sg13g2_fill_2 FILLER_12_307 ();
 sg13g2_fill_1 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_328 ();
 sg13g2_decap_8 FILLER_12_335 ();
 sg13g2_decap_8 FILLER_12_342 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_356 ();
 sg13g2_decap_8 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_370 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_39 ();
 sg13g2_fill_2 FILLER_13_44 ();
 sg13g2_decap_4 FILLER_13_50 ();
 sg13g2_fill_1 FILLER_13_54 ();
 sg13g2_decap_4 FILLER_13_59 ();
 sg13g2_fill_1 FILLER_13_69 ();
 sg13g2_fill_1 FILLER_13_79 ();
 sg13g2_fill_1 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_94 ();
 sg13g2_decap_4 FILLER_13_101 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_4 FILLER_13_161 ();
 sg13g2_fill_1 FILLER_13_165 ();
 sg13g2_fill_2 FILLER_13_174 ();
 sg13g2_fill_1 FILLER_13_176 ();
 sg13g2_fill_1 FILLER_13_205 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_fill_2 FILLER_13_292 ();
 sg13g2_fill_2 FILLER_13_329 ();
 sg13g2_decap_4 FILLER_13_353 ();
 sg13g2_fill_1 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_1 FILLER_14_70 ();
 sg13g2_fill_1 FILLER_14_97 ();
 sg13g2_decap_8 FILLER_14_124 ();
 sg13g2_fill_2 FILLER_14_131 ();
 sg13g2_decap_8 FILLER_14_137 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_fill_2 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_fill_2 FILLER_14_218 ();
 sg13g2_fill_1 FILLER_14_220 ();
 sg13g2_fill_1 FILLER_14_235 ();
 sg13g2_fill_2 FILLER_14_240 ();
 sg13g2_decap_4 FILLER_14_252 ();
 sg13g2_fill_2 FILLER_14_268 ();
 sg13g2_fill_1 FILLER_14_270 ();
 sg13g2_fill_2 FILLER_14_285 ();
 sg13g2_fill_1 FILLER_14_287 ();
 sg13g2_fill_2 FILLER_14_323 ();
 sg13g2_fill_1 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_4 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_18 ();
 sg13g2_fill_2 FILLER_15_36 ();
 sg13g2_fill_1 FILLER_15_38 ();
 sg13g2_fill_2 FILLER_15_48 ();
 sg13g2_fill_2 FILLER_15_110 ();
 sg13g2_fill_1 FILLER_15_112 ();
 sg13g2_decap_4 FILLER_15_148 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_decap_8 FILLER_15_157 ();
 sg13g2_fill_1 FILLER_15_164 ();
 sg13g2_decap_4 FILLER_15_177 ();
 sg13g2_fill_1 FILLER_15_181 ();
 sg13g2_fill_2 FILLER_15_205 ();
 sg13g2_fill_1 FILLER_15_207 ();
 sg13g2_fill_2 FILLER_15_236 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_fill_1 FILLER_15_280 ();
 sg13g2_fill_1 FILLER_15_337 ();
 sg13g2_fill_1 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_11 ();
 sg13g2_fill_2 FILLER_16_35 ();
 sg13g2_fill_1 FILLER_16_37 ();
 sg13g2_fill_1 FILLER_16_95 ();
 sg13g2_fill_2 FILLER_16_168 ();
 sg13g2_fill_1 FILLER_16_170 ();
 sg13g2_decap_4 FILLER_16_176 ();
 sg13g2_fill_1 FILLER_16_204 ();
 sg13g2_decap_4 FILLER_16_215 ();
 sg13g2_fill_2 FILLER_16_223 ();
 sg13g2_fill_1 FILLER_16_225 ();
 sg13g2_fill_2 FILLER_16_237 ();
 sg13g2_decap_8 FILLER_16_250 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_fill_1 FILLER_16_275 ();
 sg13g2_fill_1 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_355 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_33 ();
 sg13g2_fill_2 FILLER_17_49 ();
 sg13g2_fill_2 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_80 ();
 sg13g2_decap_4 FILLER_17_86 ();
 sg13g2_fill_1 FILLER_17_90 ();
 sg13g2_fill_1 FILLER_17_113 ();
 sg13g2_fill_1 FILLER_17_150 ();
 sg13g2_fill_2 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_179 ();
 sg13g2_decap_4 FILLER_17_184 ();
 sg13g2_fill_2 FILLER_17_188 ();
 sg13g2_fill_2 FILLER_17_195 ();
 sg13g2_fill_1 FILLER_17_197 ();
 sg13g2_fill_1 FILLER_17_202 ();
 sg13g2_fill_1 FILLER_17_208 ();
 sg13g2_decap_8 FILLER_17_213 ();
 sg13g2_decap_4 FILLER_17_255 ();
 sg13g2_fill_1 FILLER_17_259 ();
 sg13g2_decap_4 FILLER_17_292 ();
 sg13g2_fill_2 FILLER_17_296 ();
 sg13g2_fill_2 FILLER_17_321 ();
 sg13g2_fill_1 FILLER_17_323 ();
 sg13g2_fill_2 FILLER_17_337 ();
 sg13g2_fill_1 FILLER_17_343 ();
 sg13g2_decap_4 FILLER_17_348 ();
 sg13g2_fill_2 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_62 ();
 sg13g2_fill_2 FILLER_18_103 ();
 sg13g2_fill_2 FILLER_18_121 ();
 sg13g2_fill_2 FILLER_18_166 ();
 sg13g2_fill_1 FILLER_18_168 ();
 sg13g2_fill_1 FILLER_18_195 ();
 sg13g2_decap_4 FILLER_18_201 ();
 sg13g2_fill_1 FILLER_18_211 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_fill_2 FILLER_18_235 ();
 sg13g2_decap_4 FILLER_18_245 ();
 sg13g2_fill_2 FILLER_18_270 ();
 sg13g2_fill_1 FILLER_18_296 ();
 sg13g2_decap_4 FILLER_18_301 ();
 sg13g2_fill_1 FILLER_18_305 ();
 sg13g2_fill_2 FILLER_18_310 ();
 sg13g2_fill_2 FILLER_18_357 ();
 sg13g2_fill_1 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_fill_2 FILLER_19_29 ();
 sg13g2_fill_2 FILLER_19_39 ();
 sg13g2_fill_2 FILLER_19_82 ();
 sg13g2_fill_2 FILLER_19_93 ();
 sg13g2_fill_1 FILLER_19_95 ();
 sg13g2_fill_2 FILLER_19_114 ();
 sg13g2_fill_1 FILLER_19_116 ();
 sg13g2_decap_4 FILLER_19_129 ();
 sg13g2_fill_2 FILLER_19_160 ();
 sg13g2_decap_8 FILLER_19_166 ();
 sg13g2_decap_8 FILLER_19_173 ();
 sg13g2_decap_8 FILLER_19_180 ();
 sg13g2_decap_4 FILLER_19_187 ();
 sg13g2_fill_2 FILLER_19_191 ();
 sg13g2_fill_1 FILLER_19_201 ();
 sg13g2_fill_2 FILLER_19_217 ();
 sg13g2_fill_2 FILLER_19_225 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_decap_4 FILLER_19_231 ();
 sg13g2_fill_2 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_fill_2 FILLER_19_246 ();
 sg13g2_fill_1 FILLER_19_248 ();
 sg13g2_decap_8 FILLER_19_254 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_decap_4 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_272 ();
 sg13g2_decap_4 FILLER_19_277 ();
 sg13g2_fill_1 FILLER_19_281 ();
 sg13g2_fill_2 FILLER_19_287 ();
 sg13g2_fill_1 FILLER_19_289 ();
 sg13g2_fill_2 FILLER_19_334 ();
 sg13g2_fill_2 FILLER_19_344 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_86 ();
 sg13g2_fill_1 FILLER_20_88 ();
 sg13g2_decap_8 FILLER_20_97 ();
 sg13g2_decap_8 FILLER_20_104 ();
 sg13g2_decap_8 FILLER_20_116 ();
 sg13g2_fill_2 FILLER_20_123 ();
 sg13g2_fill_2 FILLER_20_196 ();
 sg13g2_fill_1 FILLER_20_198 ();
 sg13g2_fill_2 FILLER_20_203 ();
 sg13g2_fill_1 FILLER_20_205 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_fill_1 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_225 ();
 sg13g2_fill_1 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_fill_1 FILLER_20_277 ();
 sg13g2_fill_2 FILLER_20_330 ();
 sg13g2_decap_4 FILLER_20_336 ();
 sg13g2_fill_1 FILLER_20_340 ();
 sg13g2_decap_4 FILLER_20_352 ();
 sg13g2_fill_1 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_fill_2 FILLER_21_29 ();
 sg13g2_fill_1 FILLER_21_71 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_decap_4 FILLER_21_158 ();
 sg13g2_fill_2 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_172 ();
 sg13g2_decap_8 FILLER_21_177 ();
 sg13g2_decap_8 FILLER_21_184 ();
 sg13g2_decap_4 FILLER_21_191 ();
 sg13g2_fill_2 FILLER_21_195 ();
 sg13g2_fill_1 FILLER_21_205 ();
 sg13g2_decap_4 FILLER_21_211 ();
 sg13g2_decap_8 FILLER_21_225 ();
 sg13g2_fill_2 FILLER_21_232 ();
 sg13g2_fill_2 FILLER_21_242 ();
 sg13g2_fill_1 FILLER_21_244 ();
 sg13g2_fill_1 FILLER_21_275 ();
 sg13g2_decap_4 FILLER_21_296 ();
 sg13g2_fill_2 FILLER_21_300 ();
 sg13g2_decap_4 FILLER_21_365 ();
 sg13g2_fill_1 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_384 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_31 ();
 sg13g2_fill_2 FILLER_22_68 ();
 sg13g2_fill_1 FILLER_22_89 ();
 sg13g2_fill_2 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_142 ();
 sg13g2_fill_2 FILLER_22_155 ();
 sg13g2_fill_1 FILLER_22_208 ();
 sg13g2_decap_8 FILLER_22_223 ();
 sg13g2_decap_4 FILLER_22_230 ();
 sg13g2_fill_1 FILLER_22_234 ();
 sg13g2_decap_8 FILLER_22_246 ();
 sg13g2_decap_4 FILLER_22_253 ();
 sg13g2_fill_1 FILLER_22_257 ();
 sg13g2_fill_2 FILLER_22_271 ();
 sg13g2_fill_2 FILLER_22_277 ();
 sg13g2_fill_1 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_4 FILLER_22_315 ();
 sg13g2_fill_1 FILLER_22_319 ();
 sg13g2_fill_2 FILLER_22_340 ();
 sg13g2_fill_2 FILLER_22_352 ();
 sg13g2_fill_2 FILLER_22_360 ();
 sg13g2_fill_1 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_2 FILLER_23_29 ();
 sg13g2_fill_2 FILLER_23_45 ();
 sg13g2_decap_4 FILLER_23_74 ();
 sg13g2_fill_1 FILLER_23_78 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_fill_2 FILLER_23_91 ();
 sg13g2_decap_4 FILLER_23_97 ();
 sg13g2_fill_1 FILLER_23_101 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_fill_1 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_124 ();
 sg13g2_decap_8 FILLER_23_131 ();
 sg13g2_decap_4 FILLER_23_150 ();
 sg13g2_decap_8 FILLER_23_172 ();
 sg13g2_decap_8 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_186 ();
 sg13g2_decap_8 FILLER_23_191 ();
 sg13g2_fill_2 FILLER_23_198 ();
 sg13g2_fill_2 FILLER_23_218 ();
 sg13g2_fill_1 FILLER_23_220 ();
 sg13g2_fill_1 FILLER_23_229 ();
 sg13g2_fill_1 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_256 ();
 sg13g2_fill_1 FILLER_23_263 ();
 sg13g2_fill_2 FILLER_23_337 ();
 sg13g2_decap_4 FILLER_23_358 ();
 sg13g2_fill_2 FILLER_23_362 ();
 sg13g2_decap_4 FILLER_23_378 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_18 ();
 sg13g2_fill_2 FILLER_24_22 ();
 sg13g2_fill_1 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_83 ();
 sg13g2_fill_1 FILLER_24_93 ();
 sg13g2_decap_4 FILLER_24_98 ();
 sg13g2_fill_2 FILLER_24_102 ();
 sg13g2_fill_1 FILLER_24_125 ();
 sg13g2_fill_2 FILLER_24_180 ();
 sg13g2_fill_1 FILLER_24_182 ();
 sg13g2_decap_4 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_213 ();
 sg13g2_fill_1 FILLER_24_219 ();
 sg13g2_fill_2 FILLER_24_228 ();
 sg13g2_fill_1 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_decap_4 FILLER_24_287 ();
 sg13g2_fill_1 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_fill_2 FILLER_24_308 ();
 sg13g2_decap_4 FILLER_24_342 ();
 sg13g2_fill_1 FILLER_24_346 ();
 sg13g2_decap_4 FILLER_24_353 ();
 sg13g2_fill_2 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_22 ();
 sg13g2_fill_1 FILLER_25_24 ();
 sg13g2_fill_2 FILLER_25_39 ();
 sg13g2_fill_1 FILLER_25_41 ();
 sg13g2_fill_2 FILLER_25_67 ();
 sg13g2_fill_1 FILLER_25_69 ();
 sg13g2_fill_1 FILLER_25_80 ();
 sg13g2_fill_2 FILLER_25_97 ();
 sg13g2_fill_1 FILLER_25_99 ();
 sg13g2_fill_2 FILLER_25_108 ();
 sg13g2_fill_1 FILLER_25_110 ();
 sg13g2_decap_8 FILLER_25_124 ();
 sg13g2_decap_8 FILLER_25_131 ();
 sg13g2_fill_2 FILLER_25_150 ();
 sg13g2_fill_1 FILLER_25_152 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_fill_2 FILLER_25_198 ();
 sg13g2_fill_2 FILLER_25_234 ();
 sg13g2_fill_1 FILLER_25_236 ();
 sg13g2_fill_1 FILLER_25_250 ();
 sg13g2_fill_2 FILLER_25_337 ();
 sg13g2_decap_8 FILLER_25_352 ();
 sg13g2_fill_2 FILLER_25_359 ();
 sg13g2_fill_1 FILLER_25_382 ();
 sg13g2_fill_2 FILLER_25_389 ();
 sg13g2_fill_1 FILLER_25_391 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_51 ();
 sg13g2_fill_2 FILLER_26_62 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_77 ();
 sg13g2_fill_2 FILLER_26_83 ();
 sg13g2_fill_1 FILLER_26_85 ();
 sg13g2_decap_4 FILLER_26_90 ();
 sg13g2_fill_1 FILLER_26_94 ();
 sg13g2_fill_2 FILLER_26_110 ();
 sg13g2_decap_4 FILLER_26_134 ();
 sg13g2_decap_4 FILLER_26_150 ();
 sg13g2_fill_2 FILLER_26_181 ();
 sg13g2_fill_1 FILLER_26_183 ();
 sg13g2_decap_4 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_240 ();
 sg13g2_decap_8 FILLER_26_247 ();
 sg13g2_fill_2 FILLER_26_263 ();
 sg13g2_fill_1 FILLER_26_265 ();
 sg13g2_fill_2 FILLER_26_275 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_fill_2 FILLER_26_292 ();
 sg13g2_fill_1 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_328 ();
 sg13g2_decap_8 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_fill_2 FILLER_26_351 ();
 sg13g2_fill_1 FILLER_26_353 ();
 sg13g2_decap_8 FILLER_26_359 ();
 sg13g2_fill_2 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_11 ();
 sg13g2_fill_2 FILLER_27_15 ();
 sg13g2_fill_2 FILLER_27_27 ();
 sg13g2_fill_2 FILLER_27_43 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_fill_2 FILLER_27_60 ();
 sg13g2_fill_2 FILLER_27_75 ();
 sg13g2_fill_1 FILLER_27_93 ();
 sg13g2_fill_2 FILLER_27_106 ();
 sg13g2_fill_1 FILLER_27_108 ();
 sg13g2_decap_4 FILLER_27_127 ();
 sg13g2_fill_2 FILLER_27_131 ();
 sg13g2_fill_1 FILLER_27_154 ();
 sg13g2_fill_2 FILLER_27_163 ();
 sg13g2_fill_1 FILLER_27_165 ();
 sg13g2_decap_8 FILLER_27_173 ();
 sg13g2_decap_8 FILLER_27_180 ();
 sg13g2_decap_8 FILLER_27_187 ();
 sg13g2_fill_1 FILLER_27_194 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_4 FILLER_27_210 ();
 sg13g2_fill_1 FILLER_27_214 ();
 sg13g2_fill_2 FILLER_27_219 ();
 sg13g2_decap_8 FILLER_27_230 ();
 sg13g2_decap_8 FILLER_27_237 ();
 sg13g2_fill_1 FILLER_27_244 ();
 sg13g2_fill_2 FILLER_27_271 ();
 sg13g2_fill_1 FILLER_27_273 ();
 sg13g2_fill_2 FILLER_27_305 ();
 sg13g2_decap_4 FILLER_27_315 ();
 sg13g2_decap_4 FILLER_27_327 ();
 sg13g2_fill_2 FILLER_27_331 ();
 sg13g2_decap_4 FILLER_27_352 ();
 sg13g2_fill_2 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_1 FILLER_28_47 ();
 sg13g2_fill_2 FILLER_28_75 ();
 sg13g2_fill_2 FILLER_28_85 ();
 sg13g2_fill_1 FILLER_28_87 ();
 sg13g2_fill_2 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_121 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_decap_8 FILLER_28_136 ();
 sg13g2_decap_4 FILLER_28_143 ();
 sg13g2_fill_1 FILLER_28_147 ();
 sg13g2_fill_2 FILLER_28_173 ();
 sg13g2_decap_4 FILLER_28_180 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_fill_2 FILLER_28_212 ();
 sg13g2_fill_1 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_233 ();
 sg13g2_fill_1 FILLER_28_240 ();
 sg13g2_decap_8 FILLER_28_246 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_decap_8 FILLER_28_263 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_316 ();
 sg13g2_fill_1 FILLER_28_332 ();
 sg13g2_fill_1 FILLER_28_355 ();
 sg13g2_decap_4 FILLER_28_361 ();
 sg13g2_fill_1 FILLER_28_380 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_9 ();
 sg13g2_fill_2 FILLER_29_85 ();
 sg13g2_fill_1 FILLER_29_87 ();
 sg13g2_fill_2 FILLER_29_109 ();
 sg13g2_fill_1 FILLER_29_111 ();
 sg13g2_fill_2 FILLER_29_163 ();
 sg13g2_fill_1 FILLER_29_165 ();
 sg13g2_fill_2 FILLER_29_230 ();
 sg13g2_fill_1 FILLER_29_232 ();
 sg13g2_fill_2 FILLER_29_277 ();
 sg13g2_fill_2 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_338 ();
 sg13g2_decap_4 FILLER_29_359 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_2 FILLER_30_43 ();
 sg13g2_fill_1 FILLER_30_45 ();
 sg13g2_fill_2 FILLER_30_55 ();
 sg13g2_fill_1 FILLER_30_57 ();
 sg13g2_fill_2 FILLER_30_80 ();
 sg13g2_decap_4 FILLER_30_90 ();
 sg13g2_decap_8 FILLER_30_97 ();
 sg13g2_fill_2 FILLER_30_104 ();
 sg13g2_fill_1 FILLER_30_106 ();
 sg13g2_fill_1 FILLER_30_115 ();
 sg13g2_fill_2 FILLER_30_122 ();
 sg13g2_fill_1 FILLER_30_127 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_decap_8 FILLER_30_142 ();
 sg13g2_fill_2 FILLER_30_149 ();
 sg13g2_fill_2 FILLER_30_172 ();
 sg13g2_fill_1 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_178 ();
 sg13g2_decap_8 FILLER_30_184 ();
 sg13g2_decap_8 FILLER_30_191 ();
 sg13g2_fill_2 FILLER_30_198 ();
 sg13g2_decap_4 FILLER_30_214 ();
 sg13g2_decap_4 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_decap_8 FILLER_30_282 ();
 sg13g2_decap_4 FILLER_30_293 ();
 sg13g2_fill_2 FILLER_30_297 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_4 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_319 ();
 sg13g2_decap_4 FILLER_30_330 ();
 sg13g2_fill_1 FILLER_30_334 ();
 sg13g2_fill_1 FILLER_30_365 ();
 sg13g2_fill_2 FILLER_30_372 ();
 sg13g2_fill_1 FILLER_30_374 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_36 ();
 sg13g2_fill_1 FILLER_31_46 ();
 sg13g2_fill_2 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_74 ();
 sg13g2_fill_1 FILLER_31_101 ();
 sg13g2_fill_1 FILLER_31_118 ();
 sg13g2_decap_8 FILLER_31_139 ();
 sg13g2_fill_1 FILLER_31_146 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_fill_1 FILLER_31_203 ();
 sg13g2_decap_4 FILLER_31_214 ();
 sg13g2_decap_4 FILLER_31_223 ();
 sg13g2_decap_8 FILLER_31_288 ();
 sg13g2_decap_4 FILLER_31_322 ();
 sg13g2_fill_2 FILLER_31_326 ();
 sg13g2_decap_8 FILLER_31_332 ();
 sg13g2_decap_8 FILLER_31_339 ();
 sg13g2_decap_8 FILLER_31_346 ();
 sg13g2_decap_8 FILLER_31_366 ();
 sg13g2_fill_1 FILLER_31_373 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_11 ();
 sg13g2_decap_4 FILLER_32_69 ();
 sg13g2_fill_1 FILLER_32_81 ();
 sg13g2_fill_1 FILLER_32_97 ();
 sg13g2_decap_4 FILLER_32_103 ();
 sg13g2_fill_1 FILLER_32_107 ();
 sg13g2_fill_2 FILLER_32_124 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_fill_2 FILLER_32_143 ();
 sg13g2_decap_8 FILLER_32_174 ();
 sg13g2_fill_2 FILLER_32_185 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_275 ();
 sg13g2_decap_8 FILLER_32_347 ();
 sg13g2_fill_2 FILLER_32_354 ();
 sg13g2_fill_1 FILLER_32_356 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_decap_4 FILLER_33_59 ();
 sg13g2_fill_1 FILLER_33_63 ();
 sg13g2_decap_4 FILLER_33_69 ();
 sg13g2_fill_2 FILLER_33_73 ();
 sg13g2_fill_1 FILLER_33_87 ();
 sg13g2_fill_1 FILLER_33_111 ();
 sg13g2_decap_4 FILLER_33_138 ();
 sg13g2_fill_2 FILLER_33_142 ();
 sg13g2_fill_1 FILLER_33_152 ();
 sg13g2_decap_4 FILLER_33_192 ();
 sg13g2_decap_4 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_211 ();
 sg13g2_fill_1 FILLER_33_215 ();
 sg13g2_decap_8 FILLER_33_223 ();
 sg13g2_decap_4 FILLER_33_237 ();
 sg13g2_fill_2 FILLER_33_241 ();
 sg13g2_decap_8 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_fill_2 FILLER_33_293 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_fill_1 FILLER_33_319 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_fill_2 FILLER_33_353 ();
 sg13g2_fill_1 FILLER_33_355 ();
 sg13g2_decap_8 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_380 ();
 sg13g2_fill_1 FILLER_33_387 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_4 FILLER_34_35 ();
 sg13g2_fill_1 FILLER_34_39 ();
 sg13g2_decap_4 FILLER_34_52 ();
 sg13g2_fill_2 FILLER_34_56 ();
 sg13g2_decap_4 FILLER_34_83 ();
 sg13g2_fill_2 FILLER_34_87 ();
 sg13g2_decap_4 FILLER_34_107 ();
 sg13g2_fill_2 FILLER_34_111 ();
 sg13g2_decap_8 FILLER_34_159 ();
 sg13g2_decap_8 FILLER_34_166 ();
 sg13g2_fill_1 FILLER_34_173 ();
 sg13g2_fill_1 FILLER_34_204 ();
 sg13g2_fill_1 FILLER_34_219 ();
 sg13g2_fill_1 FILLER_34_323 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_369 ();
 sg13g2_fill_1 FILLER_34_371 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_fill_2 FILLER_35_86 ();
 sg13g2_decap_8 FILLER_35_122 ();
 sg13g2_fill_1 FILLER_35_129 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_161 ();
 sg13g2_decap_4 FILLER_35_166 ();
 sg13g2_fill_1 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_193 ();
 sg13g2_fill_1 FILLER_35_211 ();
 sg13g2_fill_1 FILLER_35_244 ();
 sg13g2_fill_2 FILLER_35_280 ();
 sg13g2_decap_4 FILLER_35_286 ();
 sg13g2_fill_2 FILLER_35_331 ();
 sg13g2_fill_1 FILLER_35_333 ();
 sg13g2_fill_2 FILLER_35_368 ();
 sg13g2_fill_2 FILLER_35_377 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_fill_2 FILLER_36_70 ();
 sg13g2_fill_1 FILLER_36_72 ();
 sg13g2_decap_8 FILLER_36_83 ();
 sg13g2_fill_1 FILLER_36_90 ();
 sg13g2_fill_1 FILLER_36_96 ();
 sg13g2_decap_8 FILLER_36_102 ();
 sg13g2_decap_8 FILLER_36_109 ();
 sg13g2_decap_8 FILLER_36_116 ();
 sg13g2_decap_8 FILLER_36_127 ();
 sg13g2_fill_1 FILLER_36_134 ();
 sg13g2_fill_2 FILLER_36_187 ();
 sg13g2_fill_2 FILLER_36_257 ();
 sg13g2_fill_1 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_337 ();
 sg13g2_fill_2 FILLER_36_348 ();
 sg13g2_fill_1 FILLER_36_350 ();
 sg13g2_decap_4 FILLER_36_359 ();
 sg13g2_fill_1 FILLER_36_363 ();
 sg13g2_decap_8 FILLER_36_382 ();
 sg13g2_fill_2 FILLER_36_389 ();
 sg13g2_fill_1 FILLER_36_391 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_138 ();
 sg13g2_fill_2 FILLER_37_145 ();
 sg13g2_fill_2 FILLER_37_151 ();
 sg13g2_fill_1 FILLER_37_153 ();
 sg13g2_fill_2 FILLER_37_158 ();
 sg13g2_decap_4 FILLER_37_164 ();
 sg13g2_fill_2 FILLER_37_172 ();
 sg13g2_fill_1 FILLER_37_195 ();
 sg13g2_fill_1 FILLER_37_254 ();
 sg13g2_fill_2 FILLER_37_366 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_fill_2 FILLER_38_124 ();
 sg13g2_fill_1 FILLER_38_126 ();
 sg13g2_fill_1 FILLER_38_169 ();
 sg13g2_fill_2 FILLER_38_228 ();
 sg13g2_fill_1 FILLER_38_230 ();
 sg13g2_decap_4 FILLER_38_257 ();
 sg13g2_fill_2 FILLER_38_287 ();
 sg13g2_fill_1 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule

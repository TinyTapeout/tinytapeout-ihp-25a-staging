module tt_um_luke_clock (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \ChiselTop.SetSelIn[0] ;
 wire \ChiselTop.SetSelIn[1] ;
 wire \ChiselTop._counterXReg_T_1[0] ;
 wire \ChiselTop._debounceCounter_T_1[0] ;
 wire \ChiselTop._modeReg_T_1[0] ;
 wire \ChiselTop.cntReg[0] ;
 wire \ChiselTop.cntReg[10] ;
 wire \ChiselTop.cntReg[11] ;
 wire \ChiselTop.cntReg[12] ;
 wire \ChiselTop.cntReg[13] ;
 wire \ChiselTop.cntReg[14] ;
 wire \ChiselTop.cntReg[15] ;
 wire \ChiselTop.cntReg[16] ;
 wire \ChiselTop.cntReg[17] ;
 wire \ChiselTop.cntReg[18] ;
 wire \ChiselTop.cntReg[19] ;
 wire \ChiselTop.cntReg[1] ;
 wire \ChiselTop.cntReg[20] ;
 wire \ChiselTop.cntReg[21] ;
 wire \ChiselTop.cntReg[22] ;
 wire \ChiselTop.cntReg[23] ;
 wire \ChiselTop.cntReg[24] ;
 wire \ChiselTop.cntReg[2] ;
 wire \ChiselTop.cntReg[3] ;
 wire \ChiselTop.cntReg[4] ;
 wire \ChiselTop.cntReg[5] ;
 wire \ChiselTop.cntReg[6] ;
 wire \ChiselTop.cntReg[7] ;
 wire \ChiselTop.cntReg[8] ;
 wire \ChiselTop.cntReg[9] ;
 wire \ChiselTop.counterXReg[0] ;
 wire \ChiselTop.counterXReg[1] ;
 wire \ChiselTop.counterXReg[2] ;
 wire \ChiselTop.counterXReg[3] ;
 wire \ChiselTop.counterXReg[4] ;
 wire \ChiselTop.counterXReg[5] ;
 wire \ChiselTop.counterXReg[6] ;
 wire \ChiselTop.counterXReg[7] ;
 wire \ChiselTop.counterXReg[8] ;
 wire \ChiselTop.counterXReg[9] ;
 wire \ChiselTop.counterYReg[0] ;
 wire \ChiselTop.counterYReg[1] ;
 wire \ChiselTop.counterYReg[2] ;
 wire \ChiselTop.counterYReg[3] ;
 wire \ChiselTop.counterYReg[4] ;
 wire \ChiselTop.counterYReg[5] ;
 wire \ChiselTop.counterYReg[6] ;
 wire \ChiselTop.counterYReg[7] ;
 wire \ChiselTop.counterYReg[8] ;
 wire \ChiselTop.counterYReg[9] ;
 wire \ChiselTop.debounceCounter[0] ;
 wire \ChiselTop.debounceCounter[10] ;
 wire \ChiselTop.debounceCounter[11] ;
 wire \ChiselTop.debounceCounter[12] ;
 wire \ChiselTop.debounceCounter[13] ;
 wire \ChiselTop.debounceCounter[14] ;
 wire \ChiselTop.debounceCounter[15] ;
 wire \ChiselTop.debounceCounter[16] ;
 wire \ChiselTop.debounceCounter[17] ;
 wire \ChiselTop.debounceCounter[18] ;
 wire \ChiselTop.debounceCounter[19] ;
 wire \ChiselTop.debounceCounter[1] ;
 wire \ChiselTop.debounceCounter[2] ;
 wire \ChiselTop.debounceCounter[3] ;
 wire \ChiselTop.debounceCounter[4] ;
 wire \ChiselTop.debounceCounter[5] ;
 wire \ChiselTop.debounceCounter[6] ;
 wire \ChiselTop.debounceCounter[7] ;
 wire \ChiselTop.debounceCounter[8] ;
 wire \ChiselTop.debounceCounter[9] ;
 wire \ChiselTop.hSyncOut_REG ;
 wire \ChiselTop.hourDecReg[0] ;
 wire \ChiselTop.hourDecReg[1] ;
 wire \ChiselTop.hourUniReg[0] ;
 wire \ChiselTop.hourUniReg[1] ;
 wire \ChiselTop.hourUniReg[2] ;
 wire \ChiselTop.hourUniReg[3] ;
 wire \ChiselTop.inDisplayArea ;
 wire \ChiselTop.lfsrReg_0 ;
 wire \ChiselTop.lfsrReg_1 ;
 wire \ChiselTop.lfsrReg_10 ;
 wire \ChiselTop.lfsrReg_11 ;
 wire \ChiselTop.lfsrReg_12 ;
 wire \ChiselTop.lfsrReg_13 ;
 wire \ChiselTop.lfsrReg_14 ;
 wire \ChiselTop.lfsrReg_15 ;
 wire \ChiselTop.lfsrReg_16 ;
 wire \ChiselTop.lfsrReg_17 ;
 wire \ChiselTop.lfsrReg_2 ;
 wire \ChiselTop.lfsrReg_3 ;
 wire \ChiselTop.lfsrReg_4 ;
 wire \ChiselTop.lfsrReg_5 ;
 wire \ChiselTop.lfsrReg_6 ;
 wire \ChiselTop.lfsrReg_7 ;
 wire \ChiselTop.lfsrReg_8 ;
 wire \ChiselTop.lfsrReg_9 ;
 wire \ChiselTop.minusIn ;
 wire \ChiselTop.minusInBounce_pipeReg_0 ;
 wire \ChiselTop.minusInBounce_pipeReg_1 ;
 wire \ChiselTop.minusInReg ;
 wire \ChiselTop.minusReqReg ;
 wire \ChiselTop.minuteDecReg[0] ;
 wire \ChiselTop.minuteDecReg[1] ;
 wire \ChiselTop.minuteDecReg[2] ;
 wire \ChiselTop.minuteUniReg[0] ;
 wire \ChiselTop.minuteUniReg[1] ;
 wire \ChiselTop.minuteUniReg[2] ;
 wire \ChiselTop.minuteUniReg[3] ;
 wire \ChiselTop.plusIn ;
 wire \ChiselTop.plusInBounce_pipeReg_0 ;
 wire \ChiselTop.plusInBounce_pipeReg_1 ;
 wire \ChiselTop.plusInReg ;
 wire \ChiselTop.plusReqReg ;
 wire \ChiselTop.secondDecReg[0] ;
 wire \ChiselTop.secondDecReg[1] ;
 wire \ChiselTop.secondDecReg[2] ;
 wire \ChiselTop.secondUniReg[0] ;
 wire \ChiselTop.secondUniReg[1] ;
 wire \ChiselTop.secondUniReg[2] ;
 wire \ChiselTop.secondUniReg[3] ;
 wire \ChiselTop.setSelInBounce_pipeReg_0[0] ;
 wire \ChiselTop.setSelInBounce_pipeReg_0[1] ;
 wire \ChiselTop.setSelInBounce_pipeReg_1[0] ;
 wire \ChiselTop.setSelInBounce_pipeReg_1[1] ;
 wire \ChiselTop.tClk ;
 wire \ChiselTop.tClk1HzInReg ;
 wire \ChiselTop.tClk1HzIn_pipeReg_0 ;
 wire \ChiselTop.tClk1HzIn_pipeReg_1 ;
 wire \ChiselTop.tClk32kHzInReg ;
 wire \ChiselTop.tClk32kHzIn_pipeReg_0 ;
 wire \ChiselTop.tClk32kHzIn_pipeReg_1 ;
 wire \ChiselTop.tClkReqReg ;
 wire \ChiselTop.tClkSelectInBounce_pipeReg_0[0] ;
 wire \ChiselTop.tClkSelectInBounce_pipeReg_0[1] ;
 wire \ChiselTop.tClkSelectInBounce_pipeReg_1[0] ;
 wire \ChiselTop.tClkSelectInBounce_pipeReg_1[1] ;
 wire \ChiselTop.tClkSelectIn[0] ;
 wire \ChiselTop.tClkSelectIn[1] ;
 wire \ChiselTop.vSync ;
 wire \ChiselTop.vSyncOut_REG ;
 wire \ChiselTop.vSyncReg ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire clknet_0_clk;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;

 sg13g2_inv_1 _1219_ (.Y(_0399_),
    .A(net315));
 sg13g2_inv_1 _1220_ (.Y(_0400_),
    .A(\ChiselTop.tClkSelectIn[0] ));
 sg13g2_inv_1 _1221_ (.Y(_0401_),
    .A(net175));
 sg13g2_inv_1 _1222_ (.Y(_0402_),
    .A(net174));
 sg13g2_inv_2 _1223_ (.Y(_0403_),
    .A(\ChiselTop.SetSelIn[1] ));
 sg13g2_inv_2 _1224_ (.Y(_0404_),
    .A(\ChiselTop.SetSelIn[0] ));
 sg13g2_inv_1 _1225_ (.Y(_0405_),
    .A(net256));
 sg13g2_inv_1 _1226_ (.Y(_0406_),
    .A(net260));
 sg13g2_inv_1 _1227_ (.Y(_0407_),
    .A(\ChiselTop.counterYReg[0] ));
 sg13g2_inv_1 _1228_ (.Y(_0408_),
    .A(net433));
 sg13g2_inv_1 _1229_ (.Y(_0409_),
    .A(net368));
 sg13g2_inv_1 _1230_ (.Y(_0410_),
    .A(\ChiselTop.cntReg[5] ));
 sg13g2_inv_1 _1231_ (.Y(_0411_),
    .A(\ChiselTop.hourUniReg[0] ));
 sg13g2_inv_1 _1232_ (.Y(_0412_),
    .A(net179));
 sg13g2_inv_1 _1233_ (.Y(_0413_),
    .A(net322));
 sg13g2_inv_1 _1234_ (.Y(_0414_),
    .A(net320));
 sg13g2_inv_1 _1235_ (.Y(_0415_),
    .A(net377));
 sg13g2_inv_1 _1236_ (.Y(_0416_),
    .A(net385));
 sg13g2_inv_1 _1237_ (.Y(_0417_),
    .A(net169));
 sg13g2_inv_1 _1238_ (.Y(_0418_),
    .A(net380));
 sg13g2_inv_1 _1239_ (.Y(_0419_),
    .A(net437));
 sg13g2_inv_1 _1240_ (.Y(_0420_),
    .A(\ChiselTop.lfsrReg_1 ));
 sg13g2_inv_1 _1241_ (.Y(_0421_),
    .A(net402));
 sg13g2_inv_1 _1242_ (.Y(_0422_),
    .A(\ChiselTop.lfsrReg_3 ));
 sg13g2_inv_1 _1243_ (.Y(_0423_),
    .A(\ChiselTop.lfsrReg_4 ));
 sg13g2_inv_1 _1244_ (.Y(_0424_),
    .A(net404));
 sg13g2_inv_1 _1245_ (.Y(_0425_),
    .A(\ChiselTop.lfsrReg_6 ));
 sg13g2_inv_1 _1246_ (.Y(_0426_),
    .A(\ChiselTop.lfsrReg_7 ));
 sg13g2_inv_1 _1247_ (.Y(_0427_),
    .A(net406));
 sg13g2_inv_1 _1248_ (.Y(_0428_),
    .A(net415));
 sg13g2_inv_1 _1249_ (.Y(_0429_),
    .A(\ChiselTop.lfsrReg_10 ));
 sg13g2_inv_1 _1250_ (.Y(_0430_),
    .A(net400));
 sg13g2_inv_1 _1251_ (.Y(_0431_),
    .A(net412));
 sg13g2_inv_1 _1252_ (.Y(_0432_),
    .A(net416));
 sg13g2_inv_1 _1253_ (.Y(_0433_),
    .A(net417));
 sg13g2_inv_1 _1254_ (.Y(_0434_),
    .A(\ChiselTop.lfsrReg_15 ));
 sg13g2_inv_1 _1255_ (.Y(_0435_),
    .A(net420));
 sg13g2_inv_1 _1256_ (.Y(_0436_),
    .A(\ChiselTop.lfsrReg_17 ));
 sg13g2_inv_1 _1257_ (.Y(_0437_),
    .A(net162));
 sg13g2_inv_1 _1258_ (.Y(_0438_),
    .A(\ChiselTop.tClkReqReg ));
 sg13g2_inv_1 _1259_ (.Y(_0439_),
    .A(_0005_));
 sg13g2_inv_1 _1260_ (.Y(_0440_),
    .A(_0007_));
 sg13g2_inv_1 _1261_ (.Y(_0441_),
    .A(\ChiselTop.tClk32kHzInReg ));
 sg13g2_inv_1 _1262_ (.Y(_0442_),
    .A(net288));
 sg13g2_inv_1 _1263_ (.Y(_0443_),
    .A(net431));
 sg13g2_inv_1 _1264_ (.Y(_0444_),
    .A(\ChiselTop.debounceCounter[7] ));
 sg13g2_inv_1 _1265_ (.Y(_0445_),
    .A(\ChiselTop.debounceCounter[13] ));
 sg13g2_inv_1 _1266_ (.Y(_0446_),
    .A(net281));
 sg13g2_inv_2 _1267_ (.Y(_0447_),
    .A(net280));
 sg13g2_inv_1 _1268_ (.Y(_0448_),
    .A(net274));
 sg13g2_inv_2 _1269_ (.Y(_0449_),
    .A(\ChiselTop.counterXReg[9] ));
 sg13g2_inv_1 _1270_ (.Y(_0450_),
    .A(_0012_));
 sg13g2_inv_1 _1271_ (.Y(_0451_),
    .A(_0016_));
 sg13g2_nand2b_1 _1272_ (.Y(_0452_),
    .B(net174),
    .A_N(\ChiselTop.minusInReg ));
 sg13g2_nand2_2 _1273_ (.Y(_0453_),
    .A(\ChiselTop.minusReqReg ),
    .B(_0452_));
 sg13g2_and2_2 _1274_ (.A(net258),
    .B(\ChiselTop.counterYReg[6] ),
    .X(_0454_));
 sg13g2_nand2_2 _1275_ (.Y(_0455_),
    .A(net259),
    .B(\ChiselTop.counterYReg[6] ));
 sg13g2_nor2b_2 _1276_ (.A(net265),
    .B_N(net261),
    .Y(_0456_));
 sg13g2_nand2b_1 _1277_ (.Y(_0457_),
    .B(net262),
    .A_N(net264));
 sg13g2_nor2_1 _1278_ (.A(_0455_),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_nand2b_1 _1279_ (.Y(_0459_),
    .B(\ChiselTop.counterYReg[3] ),
    .A_N(net269));
 sg13g2_nor3_1 _1280_ (.A(_0455_),
    .B(_0457_),
    .C(_0459_),
    .Y(_0460_));
 sg13g2_nand2b_1 _1281_ (.Y(_0461_),
    .B(net270),
    .A_N(\ChiselTop.counterYReg[0] ));
 sg13g2_nor4_1 _1282_ (.A(_0455_),
    .B(_0457_),
    .C(_0459_),
    .D(_0461_),
    .Y(_0462_));
 sg13g2_and2_2 _1283_ (.A(\ChiselTop.counterYReg[1] ),
    .B(\ChiselTop.counterYReg[0] ),
    .X(_0463_));
 sg13g2_a21oi_1 _1284_ (.A1(net270),
    .A2(\ChiselTop.counterYReg[0] ),
    .Y(_0464_),
    .B1(net268));
 sg13g2_nor2b_2 _1285_ (.A(_0464_),
    .B_N(net267),
    .Y(_0465_));
 sg13g2_nand2b_1 _1286_ (.Y(_0466_),
    .B(_0454_),
    .A_N(net447));
 sg13g2_nor2_1 _1287_ (.A(\ChiselTop.counterYReg[9] ),
    .B(net255),
    .Y(_0467_));
 sg13g2_nor3_1 _1288_ (.A(_0002_),
    .B(_0455_),
    .C(_0467_),
    .Y(_0468_));
 sg13g2_a21oi_1 _1289_ (.A1(_0465_),
    .A2(_0468_),
    .Y(_0469_),
    .B1(_0462_));
 sg13g2_nand2b_1 _1290_ (.Y(_0470_),
    .B(net255),
    .A_N(net425));
 sg13g2_or2_1 _1291_ (.X(_0471_),
    .B(_0470_),
    .A(net268));
 sg13g2_and2_2 _1292_ (.A(net266),
    .B(net269),
    .X(_0472_));
 sg13g2_nand2_1 _1293_ (.Y(_0473_),
    .A(net266),
    .B(net269));
 sg13g2_nor2_2 _1294_ (.A(net270),
    .B(\ChiselTop.counterYReg[0] ),
    .Y(_0474_));
 sg13g2_nand2b_1 _1295_ (.Y(_0475_),
    .B(_0472_),
    .A_N(_0474_));
 sg13g2_a21oi_1 _1296_ (.A1(_0458_),
    .A2(_0475_),
    .Y(_0476_),
    .B1(_0466_));
 sg13g2_nor3_2 _1297_ (.A(_0469_),
    .B(_0471_),
    .C(_0476_),
    .Y(\ChiselTop.vSync ));
 sg13g2_or4_1 _1298_ (.A(\ChiselTop.vSyncReg ),
    .B(_0469_),
    .C(_0471_),
    .D(_0476_),
    .X(_0477_));
 sg13g2_nor2_1 _1299_ (.A(_0453_),
    .B(_0477_),
    .Y(_0478_));
 sg13g2_nand2b_1 _1300_ (.Y(_0479_),
    .B(net175),
    .A_N(\ChiselTop.plusInReg ));
 sg13g2_nand2_2 _1301_ (.Y(_0480_),
    .A(\ChiselTop.plusReqReg ),
    .B(_0479_));
 sg13g2_nor2_1 _1302_ (.A(net251),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_a21o_1 _1303_ (.A2(_0480_),
    .A1(_0453_),
    .B1(net251),
    .X(_0482_));
 sg13g2_a21oi_1 _1304_ (.A1(_0453_),
    .A2(_0480_),
    .Y(_0483_),
    .B1(net251));
 sg13g2_nand2_1 _1305_ (.Y(_0484_),
    .A(\ChiselTop.tClkSelectIn[1] ),
    .B(_0400_));
 sg13g2_nor2_2 _1306_ (.A(\ChiselTop.SetSelIn[1] ),
    .B(\ChiselTop.SetSelIn[0] ),
    .Y(_0485_));
 sg13g2_nand2_2 _1307_ (.Y(_0486_),
    .A(_0403_),
    .B(_0404_));
 sg13g2_a21o_1 _1308_ (.A2(_0485_),
    .A1(net246),
    .B1(_0484_),
    .X(_0487_));
 sg13g2_nor4_1 _1309_ (.A(\ChiselTop.cntReg[19] ),
    .B(\ChiselTop.cntReg[18] ),
    .C(\ChiselTop.cntReg[17] ),
    .D(\ChiselTop.cntReg[16] ),
    .Y(_0488_));
 sg13g2_nor3_1 _1310_ (.A(\ChiselTop.cntReg[22] ),
    .B(\ChiselTop.cntReg[21] ),
    .C(\ChiselTop.cntReg[20] ),
    .Y(_0489_));
 sg13g2_nor3_1 _1311_ (.A(\ChiselTop.cntReg[24] ),
    .B(\ChiselTop.cntReg[23] ),
    .C(\ChiselTop.cntReg[15] ),
    .Y(_0490_));
 sg13g2_nand3_1 _1312_ (.B(_0489_),
    .C(_0490_),
    .A(_0488_),
    .Y(_0491_));
 sg13g2_nand2_1 _1313_ (.Y(_0492_),
    .A(\ChiselTop.cntReg[13] ),
    .B(\ChiselTop.cntReg[12] ));
 sg13g2_nand2_1 _1314_ (.Y(_0493_),
    .A(net220),
    .B(\ChiselTop.cntReg[10] ));
 sg13g2_and3_1 _1315_ (.X(_0494_),
    .A(\ChiselTop.cntReg[2] ),
    .B(\ChiselTop.cntReg[1] ),
    .C(\ChiselTop.cntReg[0] ));
 sg13g2_nand3_1 _1316_ (.B(\ChiselTop.cntReg[1] ),
    .C(\ChiselTop.cntReg[0] ),
    .A(net197),
    .Y(_0495_));
 sg13g2_nand2_1 _1317_ (.Y(_0496_),
    .A(\ChiselTop.cntReg[4] ),
    .B(\ChiselTop.cntReg[3] ));
 sg13g2_nor2_1 _1318_ (.A(_0495_),
    .B(_0496_),
    .Y(_0497_));
 sg13g2_nand4_1 _1319_ (.B(net304),
    .C(\ChiselTop.cntReg[3] ),
    .A(net216),
    .Y(_0498_),
    .D(_0494_));
 sg13g2_nand3_1 _1320_ (.B(\ChiselTop.cntReg[7] ),
    .C(net449),
    .A(\ChiselTop.cntReg[8] ),
    .Y(_0499_));
 sg13g2_nor2_1 _1321_ (.A(_0498_),
    .B(net450),
    .Y(_0500_));
 sg13g2_nand4_1 _1322_ (.B(\ChiselTop.cntReg[8] ),
    .C(\ChiselTop.cntReg[7] ),
    .A(\ChiselTop.cntReg[9] ),
    .Y(_0501_),
    .D(\ChiselTop.cntReg[6] ));
 sg13g2_or4_1 _1323_ (.A(_0410_),
    .B(_0495_),
    .C(_0496_),
    .D(_0501_),
    .X(_0502_));
 sg13g2_or3_2 _1324_ (.A(_0492_),
    .B(_0493_),
    .C(_0502_),
    .X(_0503_));
 sg13g2_inv_1 _1325_ (.Y(_0504_),
    .A(_0503_));
 sg13g2_nor2_1 _1326_ (.A(_0008_),
    .B(_0503_),
    .Y(_0505_));
 sg13g2_or2_1 _1327_ (.X(_0506_),
    .B(_0505_),
    .A(_0491_));
 sg13g2_nand3_1 _1328_ (.B(_0441_),
    .C(_0506_),
    .A(\ChiselTop.tClk32kHzIn_pipeReg_0 ),
    .Y(_0507_));
 sg13g2_nand3b_1 _1329_ (.B(\ChiselTop.tClk1HzIn_pipeReg_0 ),
    .C(\ChiselTop.tClkSelectIn[0] ),
    .Y(_0508_),
    .A_N(\ChiselTop.tClk1HzInReg ));
 sg13g2_o21ai_1 _1330_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_0487_),
    .A2(_0507_));
 sg13g2_nor4_1 _1331_ (.A(\ChiselTop.cntReg[10] ),
    .B(\ChiselTop.cntReg[9] ),
    .C(\ChiselTop.cntReg[8] ),
    .D(\ChiselTop.cntReg[7] ),
    .Y(_0510_));
 sg13g2_nand3_1 _1332_ (.B(_0498_),
    .C(_0510_),
    .A(_0409_),
    .Y(_0511_));
 sg13g2_nand2_1 _1333_ (.Y(_0512_),
    .A(\ChiselTop.cntReg[14] ),
    .B(\ChiselTop.cntReg[11] ));
 sg13g2_nor3_1 _1334_ (.A(\ChiselTop.cntReg[15] ),
    .B(_0492_),
    .C(_0512_),
    .Y(_0513_));
 sg13g2_a21oi_1 _1335_ (.A1(_0511_),
    .A2(_0513_),
    .Y(_0514_),
    .B1(_0440_));
 sg13g2_nand2b_1 _1336_ (.Y(_0515_),
    .B(\ChiselTop.cntReg[16] ),
    .A_N(\ChiselTop.cntReg[17] ));
 sg13g2_o21ai_1 _1337_ (.B1(_0006_),
    .Y(_0516_),
    .A1(_0514_),
    .A2(_0515_));
 sg13g2_nand3_1 _1338_ (.B(\ChiselTop.cntReg[21] ),
    .C(\ChiselTop.cntReg[20] ),
    .A(\ChiselTop.cntReg[22] ),
    .Y(_0517_));
 sg13g2_nand2_1 _1339_ (.Y(_0518_),
    .A(\ChiselTop.cntReg[19] ),
    .B(\ChiselTop.cntReg[18] ));
 sg13g2_nor3_1 _1340_ (.A(\ChiselTop.cntReg[23] ),
    .B(_0517_),
    .C(_0518_),
    .Y(_0519_));
 sg13g2_a21oi_1 _1341_ (.A1(_0516_),
    .A2(_0519_),
    .Y(_0520_),
    .B1(_0439_));
 sg13g2_nor2_1 _1342_ (.A(_0408_),
    .B(_0520_),
    .Y(_0521_));
 sg13g2_o21ai_1 _1343_ (.B1(_0399_),
    .Y(_0522_),
    .A1(_0482_),
    .A2(_0486_));
 sg13g2_or2_1 _1344_ (.X(_0523_),
    .B(_0522_),
    .A(_0400_));
 sg13g2_nor4_1 _1345_ (.A(_0400_),
    .B(_0408_),
    .C(_0520_),
    .D(_0522_),
    .Y(_0524_));
 sg13g2_o21ai_1 _1346_ (.B1(_0004_),
    .Y(_0525_),
    .A1(\ChiselTop.cntReg[3] ),
    .A2(_0495_));
 sg13g2_nand3_1 _1347_ (.B(\ChiselTop.cntReg[4] ),
    .C(_0525_),
    .A(_0410_),
    .Y(_0526_));
 sg13g2_a21oi_1 _1348_ (.A1(_0003_),
    .A2(_0526_),
    .Y(_0527_),
    .B1(_0501_));
 sg13g2_or3_1 _1349_ (.A(\ChiselTop.cntReg[12] ),
    .B(\ChiselTop.cntReg[11] ),
    .C(\ChiselTop.cntReg[10] ),
    .X(_0528_));
 sg13g2_o21ai_1 _1350_ (.B1(\ChiselTop.cntReg[13] ),
    .Y(_0529_),
    .A1(_0527_),
    .A2(_0528_));
 sg13g2_nor2_1 _1351_ (.A(\ChiselTop.cntReg[15] ),
    .B(\ChiselTop.cntReg[14] ),
    .Y(_0530_));
 sg13g2_and3_1 _1352_ (.X(_0531_),
    .A(_0488_),
    .B(_0489_),
    .C(_0530_));
 sg13g2_nand2_1 _1353_ (.Y(_0532_),
    .A(\ChiselTop.cntReg[24] ),
    .B(\ChiselTop.cntReg[23] ));
 sg13g2_a21oi_1 _1354_ (.A1(_0529_),
    .A2(_0531_),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_nor2_1 _1355_ (.A(\ChiselTop.tClkSelectIn[0] ),
    .B(_0522_),
    .Y(_0534_));
 sg13g2_a221oi_1 _1356_ (.B2(_0534_),
    .C1(_0524_),
    .B1(_0533_),
    .A1(\ChiselTop.tClkSelectIn[1] ),
    .Y(_0535_),
    .A2(_0509_));
 sg13g2_nor2_2 _1357_ (.A(_0438_),
    .B(net251),
    .Y(_0536_));
 sg13g2_and2_1 _1358_ (.A(_0535_),
    .B(_0536_),
    .X(\ChiselTop.tClk ));
 sg13g2_and2_1 _1359_ (.A(net276),
    .B(\ChiselTop.counterXReg[6] ),
    .X(_0537_));
 sg13g2_nand2_2 _1360_ (.Y(_0538_),
    .A(net277),
    .B(net275));
 sg13g2_nand2_2 _1361_ (.Y(_0539_),
    .A(net278),
    .B(net277));
 sg13g2_nand2_2 _1362_ (.Y(_0540_),
    .A(net279),
    .B(_0537_));
 sg13g2_nor2_2 _1363_ (.A(\ChiselTop.counterXReg[8] ),
    .B(_0449_),
    .Y(_0541_));
 sg13g2_nor2_1 _1364_ (.A(net278),
    .B(net276),
    .Y(_0542_));
 sg13g2_or2_1 _1365_ (.X(_0543_),
    .B(net275),
    .A(net276));
 sg13g2_nor3_2 _1366_ (.A(net278),
    .B(net276),
    .C(net275),
    .Y(_0544_));
 sg13g2_a21oi_1 _1367_ (.A1(net278),
    .A2(_0537_),
    .Y(_0545_),
    .B1(_0544_));
 sg13g2_and3_1 _1368_ (.X(_0000_),
    .A(net274),
    .B(_0541_),
    .C(_0545_));
 sg13g2_nor2_2 _1369_ (.A(net273),
    .B(\ChiselTop.counterXReg[8] ),
    .Y(_0546_));
 sg13g2_nor2_1 _1370_ (.A(_0026_),
    .B(_0546_),
    .Y(_0547_));
 sg13g2_nor3_1 _1371_ (.A(\ChiselTop.counterYReg[9] ),
    .B(_0468_),
    .C(_0547_),
    .Y(_0548_));
 sg13g2_nor2_2 _1372_ (.A(net266),
    .B(net268),
    .Y(_0549_));
 sg13g2_or2_1 _1373_ (.X(_0550_),
    .B(net268),
    .A(net267));
 sg13g2_and2_1 _1374_ (.A(_0474_),
    .B(_0549_),
    .X(_0551_));
 sg13g2_nand2_1 _1375_ (.Y(_0552_),
    .A(_0458_),
    .B(_0551_));
 sg13g2_o21ai_1 _1376_ (.B1(_0548_),
    .Y(_0553_),
    .A1(_0470_),
    .A2(_0552_));
 sg13g2_inv_1 _1377_ (.Y(\ChiselTop.inDisplayArea ),
    .A(_0553_));
 sg13g2_nand2_1 _1378_ (.Y(_0554_),
    .A(net190),
    .B(net251));
 sg13g2_a21oi_1 _1379_ (.A1(_0535_),
    .A2(_0554_),
    .Y(_0028_),
    .B1(net284));
 sg13g2_nor2_1 _1380_ (.A(_0403_),
    .B(_0404_),
    .Y(_0555_));
 sg13g2_and2_1 _1381_ (.A(net248),
    .B(_0555_),
    .X(_0556_));
 sg13g2_o21ai_1 _1382_ (.B1(net291),
    .Y(_0557_),
    .A1(uio_out[6]),
    .A2(_0556_));
 sg13g2_a21oi_1 _1383_ (.A1(_0437_),
    .A2(_0556_),
    .Y(_0029_),
    .B1(_0557_));
 sg13g2_and2_1 _1384_ (.A(uio_out[6]),
    .B(_0556_),
    .X(_0558_));
 sg13g2_o21ai_1 _1385_ (.B1(net291),
    .Y(_0559_),
    .A1(net378),
    .A2(_0558_));
 sg13g2_a21oi_1 _1386_ (.A1(net378),
    .A2(_0558_),
    .Y(_0030_),
    .B1(_0559_));
 sg13g2_nand2_1 _1387_ (.Y(_0560_),
    .A(\ChiselTop.lfsrReg_0 ),
    .B(\ChiselTop.lfsrReg_1 ));
 sg13g2_nand4_1 _1388_ (.B(\ChiselTop.lfsrReg_3 ),
    .C(\ChiselTop.lfsrReg_4 ),
    .A(\ChiselTop.lfsrReg_2 ),
    .Y(_0561_),
    .D(\ChiselTop.lfsrReg_5 ));
 sg13g2_nand4_1 _1389_ (.B(_0428_),
    .C(_0429_),
    .A(_0427_),
    .Y(_0562_),
    .D(_0430_));
 sg13g2_nor3_1 _1390_ (.A(\ChiselTop.lfsrReg_6 ),
    .B(\ChiselTop.lfsrReg_7 ),
    .C(_0562_),
    .Y(_0563_));
 sg13g2_nand4_1 _1391_ (.B(_0422_),
    .C(_0423_),
    .A(_0421_),
    .Y(_0564_),
    .D(_0424_));
 sg13g2_nor3_1 _1392_ (.A(\ChiselTop.lfsrReg_0 ),
    .B(\ChiselTop.lfsrReg_1 ),
    .C(_0564_),
    .Y(_0565_));
 sg13g2_nor4_1 _1393_ (.A(\ChiselTop.lfsrReg_14 ),
    .B(\ChiselTop.lfsrReg_15 ),
    .C(\ChiselTop.lfsrReg_16 ),
    .D(\ChiselTop.lfsrReg_17 ),
    .Y(_0566_));
 sg13g2_nand3_1 _1394_ (.B(_0432_),
    .C(_0566_),
    .A(_0431_),
    .Y(_0567_));
 sg13g2_nor4_1 _1395_ (.A(_0433_),
    .B(_0434_),
    .C(_0435_),
    .D(_0436_),
    .Y(_0568_));
 sg13g2_nand3_1 _1396_ (.B(\ChiselTop.lfsrReg_13 ),
    .C(_0568_),
    .A(\ChiselTop.lfsrReg_12 ),
    .Y(_0569_));
 sg13g2_nand2_1 _1397_ (.Y(_0570_),
    .A(\ChiselTop.lfsrReg_6 ),
    .B(\ChiselTop.lfsrReg_7 ));
 sg13g2_nand4_1 _1398_ (.B(\ChiselTop.lfsrReg_9 ),
    .C(\ChiselTop.lfsrReg_10 ),
    .A(\ChiselTop.lfsrReg_8 ),
    .Y(_0571_),
    .D(\ChiselTop.lfsrReg_11 ));
 sg13g2_o21ai_1 _1399_ (.B1(_0569_),
    .Y(_0572_),
    .A1(_0560_),
    .A2(_0561_));
 sg13g2_o21ai_1 _1400_ (.B1(_0567_),
    .Y(_0573_),
    .A1(_0570_),
    .A2(_0571_));
 sg13g2_nor4_1 _1401_ (.A(_0563_),
    .B(_0565_),
    .C(_0572_),
    .D(_0573_),
    .Y(_0574_));
 sg13g2_a22oi_1 _1402_ (.Y(_0575_),
    .B1(\ChiselTop.lfsrReg_15 ),
    .B2(_0422_),
    .A2(_0432_),
    .A1(\ChiselTop.lfsrReg_1 ));
 sg13g2_a22oi_1 _1403_ (.Y(_0576_),
    .B1(\ChiselTop.lfsrReg_17 ),
    .B2(_0424_),
    .A2(\ChiselTop.lfsrReg_13 ),
    .A1(_0420_));
 sg13g2_a22oi_1 _1404_ (.Y(_0577_),
    .B1(_0436_),
    .B2(\ChiselTop.lfsrReg_5 ),
    .A2(_0434_),
    .A1(\ChiselTop.lfsrReg_3 ));
 sg13g2_a22oi_1 _1405_ (.Y(_0578_),
    .B1(\ChiselTop.lfsrReg_14 ),
    .B2(_0421_),
    .A2(\ChiselTop.lfsrReg_12 ),
    .A1(_0419_));
 sg13g2_a22oi_1 _1406_ (.Y(_0579_),
    .B1(_0435_),
    .B2(\ChiselTop.lfsrReg_4 ),
    .A2(_0433_),
    .A1(\ChiselTop.lfsrReg_2 ));
 sg13g2_a22oi_1 _1407_ (.Y(_0580_),
    .B1(\ChiselTop.lfsrReg_16 ),
    .B2(_0423_),
    .A2(_0431_),
    .A1(\ChiselTop.lfsrReg_0 ));
 sg13g2_and4_1 _1408_ (.A(_0575_),
    .B(_0578_),
    .C(_0579_),
    .D(_0580_),
    .X(_0581_));
 sg13g2_nand3_1 _1409_ (.B(_0577_),
    .C(_0581_),
    .A(_0576_),
    .Y(_0582_));
 sg13g2_a22oi_1 _1410_ (.Y(_0583_),
    .B1(_0433_),
    .B2(\ChiselTop.lfsrReg_8 ),
    .A2(_0431_),
    .A1(\ChiselTop.lfsrReg_6 ));
 sg13g2_xnor2_1 _1411_ (.Y(_0584_),
    .A(\ChiselTop.lfsrReg_10 ),
    .B(\ChiselTop.lfsrReg_16 ));
 sg13g2_a22oi_1 _1412_ (.Y(_0585_),
    .B1(_0436_),
    .B2(\ChiselTop.lfsrReg_11 ),
    .A2(\ChiselTop.lfsrReg_14 ),
    .A1(_0427_));
 sg13g2_a22oi_1 _1413_ (.Y(_0586_),
    .B1(_0434_),
    .B2(\ChiselTop.lfsrReg_9 ),
    .A2(\ChiselTop.lfsrReg_13 ),
    .A1(_0426_));
 sg13g2_a22oi_1 _1414_ (.Y(_0587_),
    .B1(\ChiselTop.lfsrReg_17 ),
    .B2(_0430_),
    .A2(\ChiselTop.lfsrReg_12 ),
    .A1(_0425_));
 sg13g2_a22oi_1 _1415_ (.Y(_0588_),
    .B1(\ChiselTop.lfsrReg_15 ),
    .B2(_0428_),
    .A2(_0432_),
    .A1(\ChiselTop.lfsrReg_7 ));
 sg13g2_and3_1 _1416_ (.X(_0589_),
    .A(_0585_),
    .B(_0587_),
    .C(_0588_));
 sg13g2_nand4_1 _1417_ (.B(_0584_),
    .C(_0586_),
    .A(_0583_),
    .Y(_0590_),
    .D(_0589_));
 sg13g2_a22oi_1 _1418_ (.Y(_0591_),
    .B1(_0430_),
    .B2(\ChiselTop.lfsrReg_5 ),
    .A2(\ChiselTop.lfsrReg_8 ),
    .A1(_0421_));
 sg13g2_xnor2_1 _1419_ (.Y(_0592_),
    .A(\ChiselTop.lfsrReg_3 ),
    .B(\ChiselTop.lfsrReg_9 ));
 sg13g2_a22oi_1 _1420_ (.Y(_0593_),
    .B1(\ChiselTop.lfsrReg_11 ),
    .B2(_0424_),
    .A2(\ChiselTop.lfsrReg_7 ),
    .A1(_0420_));
 sg13g2_a22oi_1 _1421_ (.Y(_0594_),
    .B1(_0427_),
    .B2(\ChiselTop.lfsrReg_2 ),
    .A2(_0426_),
    .A1(\ChiselTop.lfsrReg_1 ));
 sg13g2_a22oi_1 _1422_ (.Y(_0595_),
    .B1(_0429_),
    .B2(\ChiselTop.lfsrReg_4 ),
    .A2(\ChiselTop.lfsrReg_6 ),
    .A1(_0419_));
 sg13g2_a22oi_1 _1423_ (.Y(_0596_),
    .B1(\ChiselTop.lfsrReg_10 ),
    .B2(_0423_),
    .A2(_0425_),
    .A1(\ChiselTop.lfsrReg_0 ));
 sg13g2_and3_1 _1424_ (.X(_0597_),
    .A(_0594_),
    .B(_0595_),
    .C(_0596_));
 sg13g2_nand4_1 _1425_ (.B(_0592_),
    .C(_0593_),
    .A(_0591_),
    .Y(_0598_),
    .D(_0597_));
 sg13g2_nand4_1 _1426_ (.B(_0582_),
    .C(_0590_),
    .A(_0574_),
    .Y(_0599_),
    .D(_0598_));
 sg13g2_a21oi_1 _1427_ (.A1(_0478_),
    .A2(_0555_),
    .Y(_0600_),
    .B1(_0599_));
 sg13g2_nand2_2 _1428_ (.Y(_0601_),
    .A(\ChiselTop.hourUniReg[1] ),
    .B(\ChiselTop.hourUniReg[0] ));
 sg13g2_nor2_1 _1429_ (.A(\ChiselTop.hourUniReg[3] ),
    .B(\ChiselTop.hourUniReg[2] ),
    .Y(_0602_));
 sg13g2_nand2_1 _1430_ (.Y(_0603_),
    .A(\ChiselTop.hourDecReg[1] ),
    .B(_0602_));
 sg13g2_nor3_2 _1431_ (.A(\ChiselTop.hourDecReg[0] ),
    .B(_0601_),
    .C(_0603_),
    .Y(_0604_));
 sg13g2_nor2_1 _1432_ (.A(\ChiselTop.minuteUniReg[2] ),
    .B(\ChiselTop.minuteUniReg[1] ),
    .Y(_0605_));
 sg13g2_and3_2 _1433_ (.X(_0606_),
    .A(\ChiselTop.minuteUniReg[3] ),
    .B(\ChiselTop.minuteUniReg[0] ),
    .C(_0605_));
 sg13g2_nand3_1 _1434_ (.B(\ChiselTop.minuteUniReg[0] ),
    .C(_0605_),
    .A(\ChiselTop.minuteUniReg[3] ),
    .Y(_0607_));
 sg13g2_nand3_1 _1435_ (.B(_0413_),
    .C(\ChiselTop.minuteDecReg[0] ),
    .A(\ChiselTop.minuteDecReg[2] ),
    .Y(_0608_));
 sg13g2_nor2_1 _1436_ (.A(_0607_),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_nand4_1 _1437_ (.B(_0417_),
    .C(_0418_),
    .A(\ChiselTop.secondUniReg[3] ),
    .Y(_0610_),
    .D(\ChiselTop.secondUniReg[0] ));
 sg13g2_nor2b_1 _1438_ (.A(_0009_),
    .B_N(\ChiselTop.secondDecReg[0] ),
    .Y(_0611_));
 sg13g2_nor2b_1 _1439_ (.A(\ChiselTop.secondDecReg[1] ),
    .B_N(_0611_),
    .Y(_0612_));
 sg13g2_nor2b_1 _1440_ (.A(_0610_),
    .B_N(_0612_),
    .Y(_0613_));
 sg13g2_nand2b_1 _1441_ (.Y(_0614_),
    .B(_0612_),
    .A_N(_0610_));
 sg13g2_and2_1 _1442_ (.A(_0609_),
    .B(_0613_),
    .X(_0615_));
 sg13g2_nand2_1 _1443_ (.Y(_0616_),
    .A(_0604_),
    .B(_0615_));
 sg13g2_and3_2 _1444_ (.X(_0617_),
    .A(net247),
    .B(_0535_),
    .C(_0536_));
 sg13g2_nand3_1 _1445_ (.B(_0535_),
    .C(_0536_),
    .A(net247),
    .Y(_0618_));
 sg13g2_o21ai_1 _1446_ (.B1(_0600_),
    .Y(_0619_),
    .A1(_0616_),
    .A2(_0618_));
 sg13g2_o21ai_1 _1447_ (.B1(net289),
    .Y(_0620_),
    .A1(net408),
    .A2(net230));
 sg13g2_a21oi_1 _1448_ (.A1(_0435_),
    .A2(net230),
    .Y(_0031_),
    .B1(_0620_));
 sg13g2_o21ai_1 _1449_ (.B1(net289),
    .Y(_0621_),
    .A1(net420),
    .A2(net230));
 sg13g2_a21oi_1 _1450_ (.A1(_0434_),
    .A2(net230),
    .Y(_0032_),
    .B1(_0621_));
 sg13g2_o21ai_1 _1451_ (.B1(net289),
    .Y(_0622_),
    .A1(net422),
    .A2(net228));
 sg13g2_a21oi_1 _1452_ (.A1(_0433_),
    .A2(net228),
    .Y(_0033_),
    .B1(_0622_));
 sg13g2_o21ai_1 _1453_ (.B1(net288),
    .Y(_0623_),
    .A1(net417),
    .A2(net228));
 sg13g2_a21oi_1 _1454_ (.A1(_0432_),
    .A2(net228),
    .Y(_0034_),
    .B1(_0623_));
 sg13g2_o21ai_1 _1455_ (.B1(net288),
    .Y(_0624_),
    .A1(net416),
    .A2(net232));
 sg13g2_a21oi_1 _1456_ (.A1(_0431_),
    .A2(net232),
    .Y(_0035_),
    .B1(_0624_));
 sg13g2_o21ai_1 _1457_ (.B1(net288),
    .Y(_0625_),
    .A1(net412),
    .A2(net232));
 sg13g2_a21oi_1 _1458_ (.A1(_0430_),
    .A2(net232),
    .Y(_0036_),
    .B1(_0625_));
 sg13g2_o21ai_1 _1459_ (.B1(net288),
    .Y(_0626_),
    .A1(net400),
    .A2(net229));
 sg13g2_a21oi_1 _1460_ (.A1(_0429_),
    .A2(net229),
    .Y(_0037_),
    .B1(_0626_));
 sg13g2_o21ai_1 _1461_ (.B1(net288),
    .Y(_0627_),
    .A1(net430),
    .A2(net228));
 sg13g2_a21oi_1 _1462_ (.A1(_0428_),
    .A2(net228),
    .Y(_0038_),
    .B1(_0627_));
 sg13g2_o21ai_1 _1463_ (.B1(net288),
    .Y(_0628_),
    .A1(net415),
    .A2(net229));
 sg13g2_a21oi_1 _1464_ (.A1(_0427_),
    .A2(net229),
    .Y(_0039_),
    .B1(_0628_));
 sg13g2_o21ai_1 _1465_ (.B1(net290),
    .Y(_0629_),
    .A1(net406),
    .A2(net232));
 sg13g2_a21oi_1 _1466_ (.A1(_0426_),
    .A2(net232),
    .Y(_0040_),
    .B1(_0629_));
 sg13g2_o21ai_1 _1467_ (.B1(net288),
    .Y(_0630_),
    .A1(net418),
    .A2(net228));
 sg13g2_a21oi_1 _1468_ (.A1(_0425_),
    .A2(net228),
    .Y(_0041_),
    .B1(_0630_));
 sg13g2_o21ai_1 _1469_ (.B1(net289),
    .Y(_0631_),
    .A1(net434),
    .A2(net231));
 sg13g2_a21oi_1 _1470_ (.A1(_0424_),
    .A2(net230),
    .Y(_0042_),
    .B1(_0631_));
 sg13g2_o21ai_1 _1471_ (.B1(net290),
    .Y(_0632_),
    .A1(net404),
    .A2(net233));
 sg13g2_a21oi_1 _1472_ (.A1(_0423_),
    .A2(net232),
    .Y(_0043_),
    .B1(_0632_));
 sg13g2_o21ai_1 _1473_ (.B1(net289),
    .Y(_0633_),
    .A1(net410),
    .A2(net231));
 sg13g2_a21oi_1 _1474_ (.A1(_0422_),
    .A2(net231),
    .Y(_0044_),
    .B1(_0633_));
 sg13g2_o21ai_1 _1475_ (.B1(net289),
    .Y(_0634_),
    .A1(net429),
    .A2(net233));
 sg13g2_a21oi_1 _1476_ (.A1(_0421_),
    .A2(net233),
    .Y(_0045_),
    .B1(_0634_));
 sg13g2_o21ai_1 _1477_ (.B1(net290),
    .Y(_0635_),
    .A1(net402),
    .A2(net233));
 sg13g2_a21oi_1 _1478_ (.A1(_0420_),
    .A2(net232),
    .Y(_0046_),
    .B1(_0635_));
 sg13g2_o21ai_1 _1479_ (.B1(net289),
    .Y(_0636_),
    .A1(\ChiselTop.lfsrReg_1 ),
    .A2(net230));
 sg13g2_a21oi_1 _1480_ (.A1(_0419_),
    .A2(net230),
    .Y(_0047_),
    .B1(_0636_));
 sg13g2_nand2_1 _1481_ (.Y(_0637_),
    .A(_0563_),
    .B(_0565_));
 sg13g2_xnor2_1 _1482_ (.Y(_0638_),
    .A(\ChiselTop.lfsrReg_10 ),
    .B(\ChiselTop.lfsrReg_17 ));
 sg13g2_o21ai_1 _1483_ (.B1(_0638_),
    .Y(_0639_),
    .A1(_0567_),
    .A2(_0637_));
 sg13g2_mux2_1 _1484_ (.A0(net437),
    .A1(_0639_),
    .S(net230),
    .X(_0640_));
 sg13g2_and2_1 _1485_ (.A(net289),
    .B(_0640_),
    .X(_0048_));
 sg13g2_a21oi_2 _1486_ (.B1(_0617_),
    .Y(_0641_),
    .A2(net244),
    .A1(_0404_));
 sg13g2_a21oi_2 _1487_ (.B1(net245),
    .Y(_0642_),
    .A2(_0536_),
    .A1(_0535_));
 sg13g2_a21o_1 _1488_ (.A2(_0536_),
    .A1(_0535_),
    .B1(net244),
    .X(_0643_));
 sg13g2_nor2_2 _1489_ (.A(_0403_),
    .B(\ChiselTop.SetSelIn[0] ),
    .Y(_0644_));
 sg13g2_nand2_2 _1490_ (.Y(_0645_),
    .A(net244),
    .B(_0644_));
 sg13g2_and2_1 _1491_ (.A(net247),
    .B(_0610_),
    .X(_0646_));
 sg13g2_nand2_1 _1492_ (.Y(_0647_),
    .A(net247),
    .B(_0610_));
 sg13g2_and2_1 _1493_ (.A(\ChiselTop.tClk ),
    .B(_0646_),
    .X(_0648_));
 sg13g2_or2_1 _1494_ (.X(_0649_),
    .B(_0645_),
    .A(net302));
 sg13g2_a22oi_1 _1495_ (.Y(_0650_),
    .B1(_0648_),
    .B2(net302),
    .A2(_0641_),
    .A1(\ChiselTop.secondUniReg[0] ));
 sg13g2_a21oi_1 _1496_ (.A1(_0649_),
    .A2(net303),
    .Y(_0049_),
    .B1(net283));
 sg13g2_nand2_1 _1497_ (.Y(_0651_),
    .A(\ChiselTop.secondUniReg[1] ),
    .B(\ChiselTop.secondUniReg[0] ));
 sg13g2_xor2_1 _1498_ (.B(\ChiselTop.secondUniReg[0] ),
    .A(net380),
    .X(_0652_));
 sg13g2_nand3_1 _1499_ (.B(net245),
    .C(_0486_),
    .A(net380),
    .Y(_0653_));
 sg13g2_a21oi_1 _1500_ (.A1(_0646_),
    .A2(_0652_),
    .Y(_0654_),
    .B1(_0642_));
 sg13g2_a221oi_1 _1501_ (.B2(_0654_),
    .C1(net285),
    .B1(_0653_),
    .A1(_0418_),
    .Y(_0050_),
    .A2(_0642_));
 sg13g2_nor2_1 _1502_ (.A(_0618_),
    .B(_0651_),
    .Y(_0655_));
 sg13g2_a21oi_1 _1503_ (.A1(net245),
    .A2(_0485_),
    .Y(_0656_),
    .B1(_0417_));
 sg13g2_o21ai_1 _1504_ (.B1(net293),
    .Y(_0657_),
    .A1(_0655_),
    .A2(_0656_));
 sg13g2_a21oi_1 _1505_ (.A1(net169),
    .A2(_0655_),
    .Y(_0051_),
    .B1(_0657_));
 sg13g2_nor2_1 _1506_ (.A(_0024_),
    .B(_0645_),
    .Y(_0658_));
 sg13g2_nor2_1 _1507_ (.A(_0025_),
    .B(_0651_),
    .Y(_0659_));
 sg13g2_xnor2_1 _1508_ (.Y(_0660_),
    .A(_0024_),
    .B(_0659_));
 sg13g2_nand2_1 _1509_ (.Y(_0661_),
    .A(_0648_),
    .B(_0660_));
 sg13g2_a21oi_1 _1510_ (.A1(net331),
    .A2(_0641_),
    .Y(_0662_),
    .B1(_0658_));
 sg13g2_a21oi_1 _1511_ (.A1(_0661_),
    .A2(net332),
    .Y(_0052_),
    .B1(net283));
 sg13g2_nor2_2 _1512_ (.A(_0642_),
    .B(_0646_),
    .Y(_0663_));
 sg13g2_nor2_1 _1513_ (.A(net244),
    .B(_0612_),
    .Y(_0664_));
 sg13g2_nor2b_1 _1514_ (.A(_0485_),
    .B_N(\ChiselTop.secondDecReg[0] ),
    .Y(_0665_));
 sg13g2_a22oi_1 _1515_ (.Y(_0666_),
    .B1(_0665_),
    .B2(net245),
    .A2(_0664_),
    .A1(net199));
 sg13g2_o21ai_1 _1516_ (.B1(net292),
    .Y(_0667_),
    .A1(\ChiselTop.secondDecReg[0] ),
    .A2(_0663_));
 sg13g2_a21oi_1 _1517_ (.A1(_0663_),
    .A2(net200),
    .Y(_0053_),
    .B1(_0667_));
 sg13g2_a21oi_1 _1518_ (.A1(\ChiselTop.secondDecReg[1] ),
    .A2(\ChiselTop.secondDecReg[0] ),
    .Y(_0668_),
    .B1(_0611_));
 sg13g2_o21ai_1 _1519_ (.B1(_0668_),
    .Y(_0669_),
    .A1(\ChiselTop.secondDecReg[1] ),
    .A2(\ChiselTop.secondDecReg[0] ));
 sg13g2_nand2_1 _1520_ (.Y(_0670_),
    .A(net413),
    .B(_0486_));
 sg13g2_mux2_1 _1521_ (.A0(_0669_),
    .A1(_0670_),
    .S(net244),
    .X(_0671_));
 sg13g2_o21ai_1 _1522_ (.B1(net297),
    .Y(_0672_),
    .A1(net413),
    .A2(_0663_));
 sg13g2_a21oi_1 _1523_ (.A1(_0663_),
    .A2(_0671_),
    .Y(_0054_),
    .B1(_0672_));
 sg13g2_o21ai_1 _1524_ (.B1(net218),
    .Y(_0673_),
    .A1(_0641_),
    .A2(_0646_));
 sg13g2_nor2b_1 _1525_ (.A(_0668_),
    .B_N(\ChiselTop.secondDecReg[2] ),
    .Y(_0674_));
 sg13g2_a21oi_1 _1526_ (.A1(\ChiselTop.secondDecReg[1] ),
    .A2(\ChiselTop.secondDecReg[0] ),
    .Y(_0675_),
    .B1(net218));
 sg13g2_nor3_1 _1527_ (.A(net244),
    .B(_0674_),
    .C(_0675_),
    .Y(_0676_));
 sg13g2_nor2_1 _1528_ (.A(_0009_),
    .B(_0645_),
    .Y(_0677_));
 sg13g2_o21ai_1 _1529_ (.B1(_0663_),
    .Y(_0678_),
    .A1(_0676_),
    .A2(_0677_));
 sg13g2_a21oi_1 _1530_ (.A1(_0673_),
    .A2(_0678_),
    .Y(_0055_),
    .B1(net285));
 sg13g2_nor2_1 _1531_ (.A(\ChiselTop.SetSelIn[1] ),
    .B(_0404_),
    .Y(_0679_));
 sg13g2_nand2_1 _1532_ (.Y(_0680_),
    .A(_0403_),
    .B(\ChiselTop.SetSelIn[0] ));
 sg13g2_nand2_1 _1533_ (.Y(_0681_),
    .A(net246),
    .B(_0679_));
 sg13g2_o21ai_1 _1534_ (.B1(_0681_),
    .Y(_0682_),
    .A1(_0614_),
    .A2(_0618_));
 sg13g2_a22oi_1 _1535_ (.Y(_0683_),
    .B1(_0679_),
    .B2(net244),
    .A2(_0617_),
    .A1(_0613_));
 sg13g2_and2_2 _1536_ (.A(_0478_),
    .B(_0480_),
    .X(_0684_));
 sg13g2_nand2_1 _1537_ (.Y(_0685_),
    .A(_0478_),
    .B(_0480_));
 sg13g2_nor2_2 _1538_ (.A(_0606_),
    .B(_0684_),
    .Y(_0686_));
 sg13g2_nor2_1 _1539_ (.A(\ChiselTop.minuteDecReg[1] ),
    .B(\ChiselTop.minuteDecReg[0] ),
    .Y(_0687_));
 sg13g2_nand2_1 _1540_ (.Y(_0688_),
    .A(_0010_),
    .B(_0687_));
 sg13g2_nor2_1 _1541_ (.A(\ChiselTop.minuteUniReg[1] ),
    .B(\ChiselTop.minuteUniReg[0] ),
    .Y(_0689_));
 sg13g2_nor4_2 _1542_ (.A(net398),
    .B(net369),
    .C(net377),
    .Y(_0690_),
    .D(net385));
 sg13g2_nor2_2 _1543_ (.A(net241),
    .B(_0690_),
    .Y(_0691_));
 sg13g2_a21o_1 _1544_ (.A2(_0688_),
    .A1(_0684_),
    .B1(_0691_),
    .X(_0692_));
 sg13g2_o21ai_1 _1545_ (.B1(_0019_),
    .Y(_0693_),
    .A1(_0686_),
    .A2(_0692_));
 sg13g2_nand2_1 _1546_ (.Y(_0694_),
    .A(_0481_),
    .B(_0609_));
 sg13g2_nand3_1 _1547_ (.B(_0688_),
    .C(_0690_),
    .A(_0684_),
    .Y(_0695_));
 sg13g2_nand3_1 _1548_ (.B(_0694_),
    .C(_0695_),
    .A(_0693_),
    .Y(_0696_));
 sg13g2_o21ai_1 _1549_ (.B1(net292),
    .Y(_0697_),
    .A1(_0683_),
    .A2(_0696_));
 sg13g2_a21oi_1 _1550_ (.A1(_0416_),
    .A2(_0683_),
    .Y(_0056_),
    .B1(_0697_));
 sg13g2_nand2_1 _1551_ (.Y(_0698_),
    .A(\ChiselTop.minuteUniReg[1] ),
    .B(\ChiselTop.minuteUniReg[0] ));
 sg13g2_nand2b_1 _1552_ (.Y(_0699_),
    .B(_0698_),
    .A_N(_0689_));
 sg13g2_mux2_1 _1553_ (.A0(_0686_),
    .A1(_0691_),
    .S(_0699_),
    .X(_0700_));
 sg13g2_o21ai_1 _1554_ (.B1(net292),
    .Y(_0701_),
    .A1(_0683_),
    .A2(_0700_));
 sg13g2_a21oi_1 _1555_ (.A1(_0415_),
    .A2(_0683_),
    .Y(_0057_),
    .B1(_0701_));
 sg13g2_nor2_1 _1556_ (.A(_0020_),
    .B(_0698_),
    .Y(_0702_));
 sg13g2_xor2_1 _1557_ (.B(_0698_),
    .A(_0020_),
    .X(_0703_));
 sg13g2_xnor2_1 _1558_ (.Y(_0704_),
    .A(_0020_),
    .B(_0689_));
 sg13g2_a22oi_1 _1559_ (.Y(_0705_),
    .B1(_0704_),
    .B2(_0691_),
    .A2(_0703_),
    .A1(_0686_));
 sg13g2_o21ai_1 _1560_ (.B1(net292),
    .Y(_0706_),
    .A1(net369),
    .A2(_0682_));
 sg13g2_a21oi_1 _1561_ (.A1(_0682_),
    .A2(_0705_),
    .Y(_0058_),
    .B1(_0706_));
 sg13g2_xor2_1 _1562_ (.B(_0702_),
    .A(_0021_),
    .X(_0707_));
 sg13g2_o21ai_1 _1563_ (.B1(_0694_),
    .Y(_0708_),
    .A1(_0606_),
    .A2(_0707_));
 sg13g2_a21oi_1 _1564_ (.A1(_0416_),
    .A2(_0605_),
    .Y(_0709_),
    .B1(net241));
 sg13g2_a221oi_1 _1565_ (.B2(net398),
    .C1(_0683_),
    .B1(_0709_),
    .A1(net241),
    .Y(_0710_),
    .A2(_0708_));
 sg13g2_o21ai_1 _1566_ (.B1(net292),
    .Y(_0711_),
    .A1(net398),
    .A2(_0682_));
 sg13g2_a21oi_1 _1567_ (.A1(_0695_),
    .A2(_0710_),
    .Y(_0059_),
    .B1(_0711_));
 sg13g2_a221oi_1 _1568_ (.B2(net244),
    .C1(_0691_),
    .B1(_0680_),
    .A1(net248),
    .Y(_0712_),
    .A2(_0607_));
 sg13g2_a21oi_1 _1569_ (.A1(_0606_),
    .A2(_0612_),
    .Y(_0713_),
    .B1(_0610_));
 sg13g2_nand4_1 _1570_ (.B(_0535_),
    .C(_0536_),
    .A(net247),
    .Y(_0714_),
    .D(_0713_));
 sg13g2_nand4_1 _1571_ (.B(_0647_),
    .C(_0712_),
    .A(_0643_),
    .Y(_0715_),
    .D(_0714_));
 sg13g2_and2_1 _1572_ (.A(net247),
    .B(_0608_),
    .X(_0716_));
 sg13g2_and2_1 _1573_ (.A(_0606_),
    .B(_0608_),
    .X(_0717_));
 sg13g2_nor3_1 _1574_ (.A(net251),
    .B(_0480_),
    .C(_0717_),
    .Y(_0718_));
 sg13g2_a21oi_1 _1575_ (.A1(_0018_),
    .A2(_0716_),
    .Y(_0719_),
    .B1(_0718_));
 sg13g2_o21ai_1 _1576_ (.B1(_0414_),
    .Y(_0720_),
    .A1(_0481_),
    .A2(_0692_));
 sg13g2_nand2_1 _1577_ (.Y(_0721_),
    .A(_0719_),
    .B(_0720_));
 sg13g2_o21ai_1 _1578_ (.B1(net292),
    .Y(_0722_),
    .A1(_0715_),
    .A2(_0721_));
 sg13g2_a21oi_1 _1579_ (.A1(_0414_),
    .A2(_0715_),
    .Y(_0060_),
    .B1(_0722_));
 sg13g2_nand2_1 _1580_ (.Y(_0723_),
    .A(\ChiselTop.minuteDecReg[1] ),
    .B(\ChiselTop.minuteDecReg[0] ));
 sg13g2_nor2b_1 _1581_ (.A(_0687_),
    .B_N(_0723_),
    .Y(_0724_));
 sg13g2_nor2_1 _1582_ (.A(net248),
    .B(_0716_),
    .Y(_0725_));
 sg13g2_a21oi_1 _1583_ (.A1(net248),
    .A2(_0717_),
    .Y(_0726_),
    .B1(_0716_));
 sg13g2_nor2_1 _1584_ (.A(_0692_),
    .B(_0724_),
    .Y(_0727_));
 sg13g2_a21oi_1 _1585_ (.A1(_0724_),
    .A2(_0726_),
    .Y(_0728_),
    .B1(_0727_));
 sg13g2_o21ai_1 _1586_ (.B1(net293),
    .Y(_0729_),
    .A1(_0715_),
    .A2(_0728_));
 sg13g2_a21oi_1 _1587_ (.A1(_0413_),
    .A2(_0715_),
    .Y(_0061_),
    .B1(_0729_));
 sg13g2_xnor2_1 _1588_ (.Y(_0730_),
    .A(_0010_),
    .B(_0723_));
 sg13g2_or2_1 _1589_ (.X(_0731_),
    .B(_0687_),
    .A(_0010_));
 sg13g2_o21ai_1 _1590_ (.B1(_0731_),
    .Y(_0732_),
    .A1(_0688_),
    .A2(_0690_));
 sg13g2_a21oi_1 _1591_ (.A1(_0684_),
    .A2(_0732_),
    .Y(_0733_),
    .B1(_0718_));
 sg13g2_o21ai_1 _1592_ (.B1(_0733_),
    .Y(_0734_),
    .A1(_0725_),
    .A2(_0730_));
 sg13g2_o21ai_1 _1593_ (.B1(net293),
    .Y(_0735_),
    .A1(_0715_),
    .A2(_0734_));
 sg13g2_a21oi_1 _1594_ (.A1(_0412_),
    .A2(_0715_),
    .Y(_0062_),
    .B1(_0735_));
 sg13g2_nand2b_1 _1595_ (.Y(_0736_),
    .B(_0613_),
    .A_N(_0609_));
 sg13g2_nand4_1 _1596_ (.B(_0535_),
    .C(_0536_),
    .A(net247),
    .Y(_0737_),
    .D(_0736_));
 sg13g2_a22oi_1 _1597_ (.Y(_0738_),
    .B1(_0645_),
    .B2(_0737_),
    .A2(_0617_),
    .A1(_0614_));
 sg13g2_nor2_1 _1598_ (.A(\ChiselTop.hourUniReg[1] ),
    .B(\ChiselTop.hourUniReg[0] ),
    .Y(_0739_));
 sg13g2_nand2b_1 _1599_ (.Y(_0740_),
    .B(_0739_),
    .A_N(\ChiselTop.hourUniReg[2] ));
 sg13g2_nor2_2 _1600_ (.A(\ChiselTop.hourUniReg[3] ),
    .B(_0740_),
    .Y(_0741_));
 sg13g2_nor2_1 _1601_ (.A(net240),
    .B(_0741_),
    .Y(_0742_));
 sg13g2_nor2_1 _1602_ (.A(\ChiselTop.hourDecReg[1] ),
    .B(\ChiselTop.hourDecReg[0] ),
    .Y(_0743_));
 sg13g2_nor2b_1 _1603_ (.A(_0743_),
    .B_N(_0741_),
    .Y(_0744_));
 sg13g2_nand2_1 _1604_ (.Y(_0745_),
    .A(_0741_),
    .B(_0743_));
 sg13g2_o21ai_1 _1605_ (.B1(_0745_),
    .Y(_0746_),
    .A1(_0015_),
    .A2(_0741_));
 sg13g2_nor2_1 _1606_ (.A(net240),
    .B(_0746_),
    .Y(_0747_));
 sg13g2_a221oi_1 _1607_ (.B2(_0411_),
    .C1(_0747_),
    .B1(net240),
    .A1(net248),
    .Y(_0748_),
    .A2(_0604_));
 sg13g2_o21ai_1 _1608_ (.B1(net287),
    .Y(_0749_),
    .A1(net392),
    .A2(net226));
 sg13g2_a21oi_1 _1609_ (.A1(net226),
    .A2(_0748_),
    .Y(_0063_),
    .B1(_0749_));
 sg13g2_nand2b_1 _1610_ (.Y(_0750_),
    .B(\ChiselTop.hourUniReg[3] ),
    .A_N(\ChiselTop.hourDecReg[1] ));
 sg13g2_nor4_2 _1611_ (.A(\ChiselTop.hourUniReg[2] ),
    .B(\ChiselTop.hourUniReg[1] ),
    .C(_0411_),
    .Y(_0751_),
    .D(_0750_));
 sg13g2_xor2_1 _1612_ (.B(\ChiselTop.hourUniReg[0] ),
    .A(\ChiselTop.hourUniReg[1] ),
    .X(_0752_));
 sg13g2_a22oi_1 _1613_ (.Y(_0753_),
    .B1(net240),
    .B2(_0752_),
    .A2(_0604_),
    .A1(net248));
 sg13g2_nor2_1 _1614_ (.A(_0751_),
    .B(_0753_),
    .Y(_0754_));
 sg13g2_nor3_1 _1615_ (.A(net240),
    .B(_0741_),
    .C(_0752_),
    .Y(_0755_));
 sg13g2_nor2_1 _1616_ (.A(_0754_),
    .B(_0755_),
    .Y(_0756_));
 sg13g2_o21ai_1 _1617_ (.B1(net292),
    .Y(_0757_),
    .A1(net441),
    .A2(net227));
 sg13g2_a21oi_1 _1618_ (.A1(net227),
    .A2(_0756_),
    .Y(_0064_),
    .B1(_0757_));
 sg13g2_nor2_2 _1619_ (.A(_0604_),
    .B(_0751_),
    .Y(_0758_));
 sg13g2_nor2_1 _1620_ (.A(_0016_),
    .B(_0601_),
    .Y(_0759_));
 sg13g2_xnor2_1 _1621_ (.Y(_0760_),
    .A(_0451_),
    .B(_0601_));
 sg13g2_a21o_1 _1622_ (.A2(_0760_),
    .A1(_0758_),
    .B1(_0684_),
    .X(_0761_));
 sg13g2_nand3b_1 _1623_ (.B(_0739_),
    .C(_0016_),
    .Y(_0762_),
    .A_N(_0602_));
 sg13g2_o21ai_1 _1624_ (.B1(_0762_),
    .Y(_0763_),
    .A1(_0016_),
    .A2(_0739_));
 sg13g2_o21ai_1 _1625_ (.B1(_0761_),
    .Y(_0764_),
    .A1(net240),
    .A2(_0763_));
 sg13g2_o21ai_1 _1626_ (.B1(net292),
    .Y(_0765_),
    .A1(net387),
    .A2(net226));
 sg13g2_a21oi_1 _1627_ (.A1(net226),
    .A2(_0764_),
    .Y(_0065_),
    .B1(_0765_));
 sg13g2_xnor2_1 _1628_ (.Y(_0766_),
    .A(_0017_),
    .B(_0759_));
 sg13g2_a21oi_1 _1629_ (.A1(net394),
    .A2(_0740_),
    .Y(_0767_),
    .B1(_0744_));
 sg13g2_a21oi_1 _1630_ (.A1(_0758_),
    .A2(_0766_),
    .Y(_0768_),
    .B1(_0684_));
 sg13g2_a21o_1 _1631_ (.A2(_0767_),
    .A1(_0684_),
    .B1(_0768_),
    .X(_0769_));
 sg13g2_o21ai_1 _1632_ (.B1(net287),
    .Y(_0770_),
    .A1(net394),
    .A2(net226));
 sg13g2_a21oi_1 _1633_ (.A1(net226),
    .A2(_0769_),
    .Y(_0066_),
    .B1(_0770_));
 sg13g2_a21o_1 _1634_ (.A2(_0758_),
    .A1(net248),
    .B1(_0742_),
    .X(_0771_));
 sg13g2_and2_1 _1635_ (.A(_0615_),
    .B(_0758_),
    .X(_0772_));
 sg13g2_a22oi_1 _1636_ (.Y(_0773_),
    .B1(_0772_),
    .B2(_0617_),
    .A2(_0771_),
    .A1(_0644_));
 sg13g2_a21oi_1 _1637_ (.A1(net226),
    .A2(_0773_),
    .Y(_0774_),
    .B1(net350));
 sg13g2_nand2b_1 _1638_ (.Y(_0775_),
    .B(_0751_),
    .A_N(\ChiselTop.hourDecReg[0] ));
 sg13g2_a21oi_1 _1639_ (.A1(_0014_),
    .A2(_0745_),
    .Y(_0776_),
    .B1(net241));
 sg13g2_a21o_1 _1640_ (.A2(_0775_),
    .A1(net240),
    .B1(_0776_),
    .X(_0777_));
 sg13g2_and3_1 _1641_ (.X(_0778_),
    .A(net226),
    .B(_0773_),
    .C(_0777_));
 sg13g2_nor3_1 _1642_ (.A(net283),
    .B(_0774_),
    .C(_0778_),
    .Y(_0067_));
 sg13g2_a21oi_1 _1643_ (.A1(net227),
    .A2(_0773_),
    .Y(_0779_),
    .B1(net364));
 sg13g2_nor2b_1 _1644_ (.A(_0741_),
    .B_N(_0743_),
    .Y(_0780_));
 sg13g2_a21oi_1 _1645_ (.A1(\ChiselTop.hourDecReg[1] ),
    .A2(\ChiselTop.hourDecReg[0] ),
    .Y(_0781_),
    .B1(_0780_));
 sg13g2_nand3_1 _1646_ (.B(_0751_),
    .C(_0781_),
    .A(net247),
    .Y(_0782_));
 sg13g2_nor2_1 _1647_ (.A(net240),
    .B(_0781_),
    .Y(_0783_));
 sg13g2_a21oi_1 _1648_ (.A1(net248),
    .A2(_0775_),
    .Y(_0784_),
    .B1(_0783_));
 sg13g2_and4_1 _1649_ (.A(net227),
    .B(_0773_),
    .C(_0782_),
    .D(_0784_),
    .X(_0785_));
 sg13g2_nor3_1 _1650_ (.A(net284),
    .B(_0779_),
    .C(_0785_),
    .Y(_0068_));
 sg13g2_and2_1 _1651_ (.A(net181),
    .B(net296),
    .X(_0069_));
 sg13g2_a221oi_1 _1652_ (.B2(_0485_),
    .C1(_0484_),
    .B1(net246),
    .A1(\ChiselTop.tClk32kHzIn_pipeReg_0 ),
    .Y(_0786_),
    .A2(_0441_));
 sg13g2_nor2_1 _1653_ (.A(_0487_),
    .B(_0506_),
    .Y(_0787_));
 sg13g2_or3_1 _1654_ (.A(\ChiselTop.tClkSelectIn[0] ),
    .B(_0522_),
    .C(_0533_),
    .X(_0788_));
 sg13g2_o21ai_1 _1655_ (.B1(_0788_),
    .Y(_0789_),
    .A1(_0521_),
    .A2(_0523_));
 sg13g2_nor2_1 _1656_ (.A(_0787_),
    .B(_0789_),
    .Y(_0790_));
 sg13g2_nor2_2 _1657_ (.A(net239),
    .B(_0790_),
    .Y(_0791_));
 sg13g2_nor2b_2 _1658_ (.A(net238),
    .B_N(net389),
    .Y(_0792_));
 sg13g2_o21ai_1 _1659_ (.B1(net291),
    .Y(_0793_),
    .A1(net389),
    .A2(net225));
 sg13g2_nor2_1 _1660_ (.A(_0792_),
    .B(_0793_),
    .Y(_0070_));
 sg13g2_o21ai_1 _1661_ (.B1(net296),
    .Y(_0794_),
    .A1(net239),
    .A2(_0789_));
 sg13g2_inv_1 _1662_ (.Y(_0795_),
    .A(_0794_));
 sg13g2_a21oi_2 _1663_ (.B1(_0795_),
    .Y(_0796_),
    .A2(_0787_),
    .A1(net297));
 sg13g2_xnor2_1 _1664_ (.Y(_0797_),
    .A(net374),
    .B(_0792_));
 sg13g2_nor2_1 _1665_ (.A(net224),
    .B(net375),
    .Y(_0071_));
 sg13g2_a21oi_1 _1666_ (.A1(\ChiselTop.cntReg[1] ),
    .A2(_0792_),
    .Y(_0798_),
    .B1(net197));
 sg13g2_nor2_1 _1667_ (.A(_0495_),
    .B(net238),
    .Y(_0799_));
 sg13g2_nor3_1 _1668_ (.A(net224),
    .B(net198),
    .C(_0799_),
    .Y(_0072_));
 sg13g2_xnor2_1 _1669_ (.Y(_0800_),
    .A(net360),
    .B(_0494_));
 sg13g2_a22oi_1 _1670_ (.Y(_0801_),
    .B1(net225),
    .B2(net361),
    .A2(net238),
    .A1(\ChiselTop.cntReg[3] ));
 sg13g2_nor2_1 _1671_ (.A(net286),
    .B(net362),
    .Y(_0073_));
 sg13g2_a21oi_1 _1672_ (.A1(\ChiselTop.cntReg[3] ),
    .A2(_0799_),
    .Y(_0802_),
    .B1(net304));
 sg13g2_nor2b_1 _1673_ (.A(net238),
    .B_N(_0497_),
    .Y(_0803_));
 sg13g2_nor3_1 _1674_ (.A(net224),
    .B(net305),
    .C(_0803_),
    .Y(_0074_));
 sg13g2_xnor2_1 _1675_ (.Y(_0804_),
    .A(_0003_),
    .B(_0497_));
 sg13g2_a22oi_1 _1676_ (.Y(_0805_),
    .B1(net225),
    .B2(_0804_),
    .A2(net238),
    .A1(net216));
 sg13g2_nor2_1 _1677_ (.A(net286),
    .B(net217),
    .Y(_0075_));
 sg13g2_xnor2_1 _1678_ (.Y(_0806_),
    .A(net368),
    .B(_0498_));
 sg13g2_a22oi_1 _1679_ (.Y(_0807_),
    .B1(net225),
    .B2(_0806_),
    .A2(net238),
    .A1(net368));
 sg13g2_nor2_1 _1680_ (.A(net283),
    .B(_0807_),
    .Y(_0076_));
 sg13g2_nor3_2 _1681_ (.A(_0409_),
    .B(_0498_),
    .C(net238),
    .Y(_0808_));
 sg13g2_nand2_1 _1682_ (.Y(_0809_),
    .A(net382),
    .B(_0808_));
 sg13g2_xnor2_1 _1683_ (.Y(_0810_),
    .A(net382),
    .B(_0808_));
 sg13g2_nor2_1 _1684_ (.A(net224),
    .B(_0810_),
    .Y(_0077_));
 sg13g2_xor2_1 _1685_ (.B(_0809_),
    .A(net397),
    .X(_0811_));
 sg13g2_nor2_1 _1686_ (.A(net224),
    .B(_0811_),
    .Y(_0078_));
 sg13g2_xor2_1 _1687_ (.B(_0500_),
    .A(net363),
    .X(_0812_));
 sg13g2_a22oi_1 _1688_ (.Y(_0813_),
    .B1(net225),
    .B2(_0812_),
    .A2(net238),
    .A1(net363));
 sg13g2_nor2_1 _1689_ (.A(net285),
    .B(_0813_),
    .Y(_0079_));
 sg13g2_nand4_1 _1690_ (.B(\ChiselTop.cntReg[8] ),
    .C(\ChiselTop.cntReg[7] ),
    .A(\ChiselTop.cntReg[9] ),
    .Y(_0814_),
    .D(_0808_));
 sg13g2_nor2_1 _1691_ (.A(_0502_),
    .B(net237),
    .Y(_0815_));
 sg13g2_xnor2_1 _1692_ (.Y(_0816_),
    .A(net376),
    .B(_0815_));
 sg13g2_nor2_1 _1693_ (.A(_0796_),
    .B(_0816_),
    .Y(_0080_));
 sg13g2_a21oi_1 _1694_ (.A1(\ChiselTop.cntReg[10] ),
    .A2(_0815_),
    .Y(_0817_),
    .B1(net220));
 sg13g2_nor2_1 _1695_ (.A(_0493_),
    .B(_0814_),
    .Y(_0818_));
 sg13g2_nor3_1 _1696_ (.A(net224),
    .B(net221),
    .C(_0818_),
    .Y(_0081_));
 sg13g2_nor2_1 _1697_ (.A(net334),
    .B(_0818_),
    .Y(_0819_));
 sg13g2_and2_1 _1698_ (.A(net334),
    .B(_0818_),
    .X(_0820_));
 sg13g2_nor3_1 _1699_ (.A(net224),
    .B(net335),
    .C(_0820_),
    .Y(_0082_));
 sg13g2_nor2_1 _1700_ (.A(net306),
    .B(_0820_),
    .Y(_0821_));
 sg13g2_nor2_1 _1701_ (.A(_0503_),
    .B(net237),
    .Y(_0822_));
 sg13g2_nor3_1 _1702_ (.A(net224),
    .B(net307),
    .C(_0822_),
    .Y(_0083_));
 sg13g2_xor2_1 _1703_ (.B(_0503_),
    .A(_0008_),
    .X(_0823_));
 sg13g2_a22oi_1 _1704_ (.Y(_0824_),
    .B1(_0791_),
    .B2(_0823_),
    .A2(net239),
    .A1(net343));
 sg13g2_nor2_1 _1705_ (.A(net285),
    .B(net344),
    .Y(_0084_));
 sg13g2_xnor2_1 _1706_ (.Y(_0825_),
    .A(net355),
    .B(_0505_));
 sg13g2_a22oi_1 _1707_ (.Y(_0826_),
    .B1(_0791_),
    .B2(net356),
    .A2(net237),
    .A1(\ChiselTop.cntReg[15] ));
 sg13g2_nor2_1 _1708_ (.A(net285),
    .B(net357),
    .Y(_0085_));
 sg13g2_nand3_1 _1709_ (.B(\ChiselTop.cntReg[14] ),
    .C(_0504_),
    .A(\ChiselTop.cntReg[15] ),
    .Y(_0827_));
 sg13g2_nor2_1 _1710_ (.A(_0001_),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_xor2_1 _1711_ (.B(_0827_),
    .A(_0001_),
    .X(_0829_));
 sg13g2_a22oi_1 _1712_ (.Y(_0830_),
    .B1(net225),
    .B2(_0829_),
    .A2(net237),
    .A1(net336));
 sg13g2_nor2_1 _1713_ (.A(net285),
    .B(net337),
    .Y(_0086_));
 sg13g2_xnor2_1 _1714_ (.Y(_0831_),
    .A(_0006_),
    .B(_0828_));
 sg13g2_a22oi_1 _1715_ (.Y(_0832_),
    .B1(net225),
    .B2(_0831_),
    .A2(net237),
    .A1(net325));
 sg13g2_nor2_1 _1716_ (.A(net285),
    .B(net326),
    .Y(_0087_));
 sg13g2_nand2_1 _1717_ (.Y(_0833_),
    .A(\ChiselTop.cntReg[17] ),
    .B(\ChiselTop.cntReg[16] ));
 sg13g2_or2_1 _1718_ (.X(_0834_),
    .B(_0833_),
    .A(_0827_));
 sg13g2_nor2_1 _1719_ (.A(net237),
    .B(_0834_),
    .Y(_0835_));
 sg13g2_nor2_1 _1720_ (.A(net323),
    .B(_0835_),
    .Y(_0836_));
 sg13g2_and2_1 _1721_ (.A(net323),
    .B(_0835_),
    .X(_0837_));
 sg13g2_nor3_1 _1722_ (.A(_0794_),
    .B(net324),
    .C(_0837_),
    .Y(_0088_));
 sg13g2_nor2_1 _1723_ (.A(net347),
    .B(_0837_),
    .Y(_0838_));
 sg13g2_and2_1 _1724_ (.A(net347),
    .B(_0837_),
    .X(_0839_));
 sg13g2_nor3_1 _1725_ (.A(_0794_),
    .B(_0838_),
    .C(_0839_),
    .Y(_0089_));
 sg13g2_nor2_1 _1726_ (.A(net341),
    .B(_0839_),
    .Y(_0840_));
 sg13g2_and2_1 _1727_ (.A(net341),
    .B(_0839_),
    .X(_0841_));
 sg13g2_nor3_1 _1728_ (.A(_0794_),
    .B(net342),
    .C(_0841_),
    .Y(_0090_));
 sg13g2_xnor2_1 _1729_ (.Y(_0842_),
    .A(net352),
    .B(_0841_));
 sg13g2_nor2_1 _1730_ (.A(_0794_),
    .B(_0842_),
    .Y(_0091_));
 sg13g2_a21oi_1 _1731_ (.A1(\ChiselTop.cntReg[21] ),
    .A2(_0841_),
    .Y(_0843_),
    .B1(net193));
 sg13g2_or3_1 _1732_ (.A(_0517_),
    .B(_0518_),
    .C(_0834_),
    .X(_0844_));
 sg13g2_nor2_1 _1733_ (.A(net237),
    .B(_0844_),
    .Y(_0845_));
 sg13g2_nor3_1 _1734_ (.A(_0794_),
    .B(net194),
    .C(_0845_),
    .Y(_0092_));
 sg13g2_xnor2_1 _1735_ (.Y(_0846_),
    .A(_0439_),
    .B(_0844_));
 sg13g2_a22oi_1 _1736_ (.Y(_0847_),
    .B1(net225),
    .B2(_0846_),
    .A2(net237),
    .A1(net371));
 sg13g2_nor2_1 _1737_ (.A(net284),
    .B(net372),
    .Y(_0093_));
 sg13g2_nand2_1 _1738_ (.Y(_0848_),
    .A(net371),
    .B(_0845_));
 sg13g2_xnor2_1 _1739_ (.Y(_0849_),
    .A(_0408_),
    .B(_0848_));
 sg13g2_nor2_1 _1740_ (.A(_0794_),
    .B(_0849_),
    .Y(_0094_));
 sg13g2_and2_1 _1741_ (.A(net176),
    .B(net296),
    .X(_0095_));
 sg13g2_nand2_1 _1742_ (.Y(_0850_),
    .A(net207),
    .B(net251));
 sg13g2_a21oi_1 _1743_ (.A1(_0452_),
    .A2(_0850_),
    .Y(_0096_),
    .B1(net284));
 sg13g2_nor2_1 _1744_ (.A(_0402_),
    .B(net284),
    .Y(_0097_));
 sg13g2_nand2_1 _1745_ (.Y(_0851_),
    .A(net195),
    .B(net251));
 sg13g2_a21oi_1 _1746_ (.A1(_0479_),
    .A2(_0851_),
    .Y(_0098_),
    .B1(net284));
 sg13g2_nor2_1 _1747_ (.A(_0401_),
    .B(net284),
    .Y(_0099_));
 sg13g2_and2_1 _1748_ (.A(net287),
    .B(\ChiselTop.vSync ),
    .X(_0100_));
 sg13g2_nand2_1 _1749_ (.Y(_0852_),
    .A(\ChiselTop.counterXReg[1] ),
    .B(net281));
 sg13g2_and2_2 _1750_ (.A(\ChiselTop.counterXReg[0] ),
    .B(\ChiselTop.counterXReg[1] ),
    .X(_0853_));
 sg13g2_nand2_1 _1751_ (.Y(_0854_),
    .A(\ChiselTop.counterXReg[0] ),
    .B(\ChiselTop.counterXReg[1] ));
 sg13g2_nand3_1 _1752_ (.B(\ChiselTop.counterXReg[3] ),
    .C(_0853_),
    .A(net282),
    .Y(_0855_));
 sg13g2_nor2b_1 _1753_ (.A(net276),
    .B_N(net278),
    .Y(_0856_));
 sg13g2_nor2_2 _1754_ (.A(net275),
    .B(net273),
    .Y(_0857_));
 sg13g2_nand4_1 _1755_ (.B(net271),
    .C(_0856_),
    .A(net272),
    .Y(_0858_),
    .D(_0857_));
 sg13g2_nor2_2 _1756_ (.A(net252),
    .B(_0858_),
    .Y(_0859_));
 sg13g2_nor2_2 _1757_ (.A(net283),
    .B(_0859_),
    .Y(_0860_));
 sg13g2_o21ai_1 _1758_ (.B1(net287),
    .Y(_0861_),
    .A1(net252),
    .A2(_0858_));
 sg13g2_and2_1 _1759_ (.A(net160),
    .B(_0860_),
    .X(_0101_));
 sg13g2_nor2b_1 _1760_ (.A(\ChiselTop.counterXReg[0] ),
    .B_N(\ChiselTop.counterXReg[1] ),
    .Y(_0862_));
 sg13g2_nand2b_1 _1761_ (.Y(_0863_),
    .B(\ChiselTop.counterXReg[0] ),
    .A_N(\ChiselTop.counterXReg[1] ));
 sg13g2_nor2_1 _1762_ (.A(\ChiselTop.counterXReg[0] ),
    .B(net365),
    .Y(_0864_));
 sg13g2_nor3_1 _1763_ (.A(_0853_),
    .B(_0861_),
    .C(net366),
    .Y(_0102_));
 sg13g2_o21ai_1 _1764_ (.B1(net290),
    .Y(_0865_),
    .A1(net282),
    .A2(_0853_));
 sg13g2_a21oi_1 _1765_ (.A1(net282),
    .A2(_0853_),
    .Y(_0103_),
    .B1(_0865_));
 sg13g2_nor2_1 _1766_ (.A(\ChiselTop.counterXReg[0] ),
    .B(net280),
    .Y(_0866_));
 sg13g2_a21oi_2 _1767_ (.B1(net280),
    .Y(_0867_),
    .A2(_0853_),
    .A1(net282));
 sg13g2_nand2_1 _1768_ (.Y(_0868_),
    .A(net287),
    .B(net253));
 sg13g2_nor2_1 _1769_ (.A(_0867_),
    .B(_0868_),
    .Y(_0104_));
 sg13g2_xor2_1 _1770_ (.B(net253),
    .A(net278),
    .X(_0869_));
 sg13g2_nor2_1 _1771_ (.A(_0861_),
    .B(_0869_),
    .Y(_0105_));
 sg13g2_nor2_1 _1772_ (.A(net358),
    .B(net253),
    .Y(_0870_));
 sg13g2_xnor2_1 _1773_ (.Y(_0871_),
    .A(net277),
    .B(_0870_));
 sg13g2_nor2_1 _1774_ (.A(_0861_),
    .B(net359),
    .Y(_0106_));
 sg13g2_nor2_1 _1775_ (.A(_0539_),
    .B(net253),
    .Y(_0872_));
 sg13g2_nor2_2 _1776_ (.A(_0540_),
    .B(net252),
    .Y(_0873_));
 sg13g2_nor2_1 _1777_ (.A(net275),
    .B(_0872_),
    .Y(_0874_));
 sg13g2_nor3_1 _1778_ (.A(_0861_),
    .B(_0873_),
    .C(net443),
    .Y(_0107_));
 sg13g2_xnor2_1 _1779_ (.Y(_0875_),
    .A(net274),
    .B(_0873_));
 sg13g2_nor2_1 _1780_ (.A(_0861_),
    .B(_0875_),
    .Y(_0108_));
 sg13g2_a21oi_1 _1781_ (.A1(net274),
    .A2(_0873_),
    .Y(_0876_),
    .B1(net272));
 sg13g2_nand2_1 _1782_ (.Y(_0877_),
    .A(net273),
    .B(net272));
 sg13g2_nor3_2 _1783_ (.A(_0540_),
    .B(net252),
    .C(_0877_),
    .Y(_0878_));
 sg13g2_nor3_1 _1784_ (.A(_0861_),
    .B(_0876_),
    .C(_0878_),
    .Y(_0109_));
 sg13g2_a21oi_1 _1785_ (.A1(net271),
    .A2(_0878_),
    .Y(_0879_),
    .B1(_0861_));
 sg13g2_o21ai_1 _1786_ (.B1(_0879_),
    .Y(_0880_),
    .A1(net271),
    .A2(_0878_));
 sg13g2_inv_1 _1787_ (.Y(_0110_),
    .A(_0880_));
 sg13g2_and2_1 _1788_ (.A(_0472_),
    .B(_0474_),
    .X(_0881_));
 sg13g2_or2_1 _1789_ (.X(_0882_),
    .B(net264),
    .A(net261));
 sg13g2_nor3_1 _1790_ (.A(net260),
    .B(net263),
    .C(net265),
    .Y(_0883_));
 sg13g2_or3_1 _1791_ (.A(\ChiselTop.counterYReg[6] ),
    .B(net263),
    .C(net265),
    .X(_0884_));
 sg13g2_nor2_1 _1792_ (.A(net255),
    .B(net259),
    .Y(_0885_));
 sg13g2_nand4_1 _1793_ (.B(_0881_),
    .C(_0883_),
    .A(\ChiselTop.counterYReg[9] ),
    .Y(_0886_),
    .D(_0885_));
 sg13g2_inv_1 _1794_ (.Y(_0887_),
    .A(_0886_));
 sg13g2_a21oi_1 _1795_ (.A1(_0859_),
    .A2(_0886_),
    .Y(_0888_),
    .B1(net396));
 sg13g2_nor3_2 _1796_ (.A(_0407_),
    .B(net252),
    .C(_0858_),
    .Y(_0889_));
 sg13g2_nor3_1 _1797_ (.A(net283),
    .B(_0888_),
    .C(_0889_),
    .Y(_0111_));
 sg13g2_o21ai_1 _1798_ (.B1(net287),
    .Y(_0890_),
    .A1(net270),
    .A2(_0889_));
 sg13g2_a21oi_1 _1799_ (.A1(net270),
    .A2(_0889_),
    .Y(_0112_),
    .B1(_0890_));
 sg13g2_nand2_1 _1800_ (.Y(_0891_),
    .A(net268),
    .B(_0860_));
 sg13g2_nand2_2 _1801_ (.Y(_0892_),
    .A(net269),
    .B(_0463_));
 sg13g2_inv_1 _1802_ (.Y(_0893_),
    .A(_0892_));
 sg13g2_nand2b_1 _1803_ (.Y(_0894_),
    .B(_0892_),
    .A_N(_0464_));
 sg13g2_nand3_1 _1804_ (.B(_0859_),
    .C(_0886_),
    .A(net287),
    .Y(_0895_));
 sg13g2_o21ai_1 _1805_ (.B1(_0891_),
    .Y(_0113_),
    .A1(_0894_),
    .A2(_0895_));
 sg13g2_nand2_1 _1806_ (.Y(_0896_),
    .A(net267),
    .B(_0860_));
 sg13g2_xnor2_1 _1807_ (.Y(_0897_),
    .A(net345),
    .B(_0892_));
 sg13g2_o21ai_1 _1808_ (.B1(_0896_),
    .Y(_0114_),
    .A1(_0895_),
    .A2(_0897_));
 sg13g2_and4_2 _1809_ (.A(net267),
    .B(net268),
    .C(net270),
    .D(\ChiselTop.counterYReg[0] ),
    .X(_0898_));
 sg13g2_a21oi_1 _1810_ (.A1(_0859_),
    .A2(_0898_),
    .Y(_0899_),
    .B1(net265));
 sg13g2_and2_2 _1811_ (.A(net265),
    .B(_0898_),
    .X(_0900_));
 sg13g2_a21oi_1 _1812_ (.A1(_0859_),
    .A2(_0900_),
    .Y(_0901_),
    .B1(net283));
 sg13g2_nor2b_1 _1813_ (.A(_0899_),
    .B_N(_0901_),
    .Y(_0115_));
 sg13g2_nand2_1 _1814_ (.Y(_0902_),
    .A(net263),
    .B(_0860_));
 sg13g2_xor2_1 _1815_ (.B(_0900_),
    .A(_0002_),
    .X(_0903_));
 sg13g2_o21ai_1 _1816_ (.B1(_0902_),
    .Y(_0116_),
    .A1(_0895_),
    .A2(_0903_));
 sg13g2_and2_2 _1817_ (.A(net263),
    .B(net265),
    .X(_0904_));
 sg13g2_nand2_1 _1818_ (.Y(_0905_),
    .A(net262),
    .B(net264));
 sg13g2_nand2_1 _1819_ (.Y(_0906_),
    .A(net267),
    .B(_0904_));
 sg13g2_nand3_1 _1820_ (.B(_0859_),
    .C(_0900_),
    .A(net263),
    .Y(_0907_));
 sg13g2_nand3_1 _1821_ (.B(net263),
    .C(_0900_),
    .A(net260),
    .Y(_0908_));
 sg13g2_nand2_1 _1822_ (.Y(_0909_),
    .A(net287),
    .B(_0908_));
 sg13g2_a22oi_1 _1823_ (.Y(_0117_),
    .B1(_0909_),
    .B2(_0861_),
    .A2(_0907_),
    .A1(_0406_));
 sg13g2_nand2_1 _1824_ (.Y(_0910_),
    .A(net259),
    .B(_0860_));
 sg13g2_xnor2_1 _1825_ (.Y(_0911_),
    .A(net383),
    .B(_0908_));
 sg13g2_o21ai_1 _1826_ (.B1(_0910_),
    .Y(_0118_),
    .A1(_0895_),
    .A2(_0911_));
 sg13g2_nand2_1 _1827_ (.Y(_0912_),
    .A(net257),
    .B(_0860_));
 sg13g2_nand3_1 _1828_ (.B(_0454_),
    .C(_0900_),
    .A(net261),
    .Y(_0913_));
 sg13g2_xnor2_1 _1829_ (.Y(_0914_),
    .A(net254),
    .B(_0913_));
 sg13g2_o21ai_1 _1830_ (.B1(_0912_),
    .Y(_0119_),
    .A1(_0895_),
    .A2(_0914_));
 sg13g2_nor3_1 _1831_ (.A(_0405_),
    .B(_0455_),
    .C(_0907_),
    .Y(_0915_));
 sg13g2_a21oi_1 _1832_ (.A1(_0859_),
    .A2(_0887_),
    .Y(_0916_),
    .B1(net283));
 sg13g2_o21ai_1 _1833_ (.B1(_0916_),
    .Y(_0917_),
    .A1(net317),
    .A2(_0915_));
 sg13g2_a21oi_1 _1834_ (.A1(net317),
    .A2(_0915_),
    .Y(_0120_),
    .B1(_0917_));
 sg13g2_and2_1 _1835_ (.A(\ChiselTop.debounceCounter[0] ),
    .B(net213),
    .X(_0918_));
 sg13g2_nand4_1 _1836_ (.B(net213),
    .C(net177),
    .A(\ChiselTop.debounceCounter[0] ),
    .Y(_0919_),
    .D(net185));
 sg13g2_nor3_1 _1837_ (.A(\ChiselTop.debounceCounter[17] ),
    .B(\ChiselTop.debounceCounter[16] ),
    .C(\ChiselTop.debounceCounter[18] ),
    .Y(_0920_));
 sg13g2_nor3_1 _1838_ (.A(\ChiselTop.debounceCounter[12] ),
    .B(_0445_),
    .C(\ChiselTop.debounceCounter[15] ),
    .Y(_0921_));
 sg13g2_nand4_1 _1839_ (.B(\ChiselTop.debounceCounter[19] ),
    .C(_0920_),
    .A(\ChiselTop.debounceCounter[14] ),
    .Y(_0922_),
    .D(_0921_));
 sg13g2_nand4_1 _1840_ (.B(\ChiselTop.debounceCounter[5] ),
    .C(_0444_),
    .A(_0443_),
    .Y(_0923_),
    .D(\ChiselTop.debounceCounter[6] ));
 sg13g2_nor3_1 _1841_ (.A(\ChiselTop.debounceCounter[9] ),
    .B(\ChiselTop.debounceCounter[8] ),
    .C(\ChiselTop.debounceCounter[11] ),
    .Y(_0924_));
 sg13g2_nand2_1 _1842_ (.Y(_0925_),
    .A(\ChiselTop.debounceCounter[10] ),
    .B(_0924_));
 sg13g2_nand2_1 _1843_ (.Y(_0926_),
    .A(net223),
    .B(net202));
 sg13g2_or4_1 _1844_ (.A(_0919_),
    .B(_0922_),
    .C(_0923_),
    .D(_0925_),
    .X(_0927_));
 sg13g2_nand2_1 _1845_ (.Y(_0928_),
    .A(net293),
    .B(net250));
 sg13g2_inv_2 _1846_ (.Y(_0929_),
    .A(net243));
 sg13g2_and2_1 _1847_ (.A(net161),
    .B(_0929_),
    .X(_0121_));
 sg13g2_nor2_1 _1848_ (.A(\ChiselTop.debounceCounter[0] ),
    .B(net213),
    .Y(_0930_));
 sg13g2_nor3_1 _1849_ (.A(net284),
    .B(_0918_),
    .C(net214),
    .Y(_0122_));
 sg13g2_o21ai_1 _1850_ (.B1(_0929_),
    .Y(_0931_),
    .A1(net185),
    .A2(_0918_));
 sg13g2_a21oi_1 _1851_ (.A1(net185),
    .A2(_0918_),
    .Y(_0123_),
    .B1(_0931_));
 sg13g2_a21oi_1 _1852_ (.A1(\ChiselTop.debounceCounter[2] ),
    .A2(_0918_),
    .Y(_0932_),
    .B1(net177));
 sg13g2_nand2_1 _1853_ (.Y(_0933_),
    .A(net293),
    .B(_0919_));
 sg13g2_nor2_1 _1854_ (.A(net178),
    .B(_0933_),
    .Y(_0124_));
 sg13g2_nor2_2 _1855_ (.A(_0443_),
    .B(_0919_),
    .Y(_0934_));
 sg13g2_and2_1 _1856_ (.A(_0443_),
    .B(_0919_),
    .X(_0935_));
 sg13g2_nor3_1 _1857_ (.A(net243),
    .B(_0934_),
    .C(net432),
    .Y(_0125_));
 sg13g2_o21ai_1 _1858_ (.B1(_0929_),
    .Y(_0936_),
    .A1(net223),
    .A2(_0934_));
 sg13g2_a21oi_1 _1859_ (.A1(net223),
    .A2(_0934_),
    .Y(_0126_),
    .B1(_0936_));
 sg13g2_a21oi_1 _1860_ (.A1(\ChiselTop.debounceCounter[5] ),
    .A2(_0934_),
    .Y(_0937_),
    .B1(net202));
 sg13g2_nor3_2 _1861_ (.A(_0443_),
    .B(_0919_),
    .C(_0926_),
    .Y(_0938_));
 sg13g2_nor3_1 _1862_ (.A(net243),
    .B(net203),
    .C(_0938_),
    .Y(_0127_));
 sg13g2_nor2_1 _1863_ (.A(net329),
    .B(_0938_),
    .Y(_0939_));
 sg13g2_and2_1 _1864_ (.A(net329),
    .B(_0938_),
    .X(_0940_));
 sg13g2_nor3_1 _1865_ (.A(net243),
    .B(net330),
    .C(_0940_),
    .Y(_0128_));
 sg13g2_nor2_1 _1866_ (.A(net308),
    .B(_0940_),
    .Y(_0941_));
 sg13g2_and3_1 _1867_ (.X(_0942_),
    .A(\ChiselTop.debounceCounter[7] ),
    .B(net308),
    .C(_0938_));
 sg13g2_nor3_1 _1868_ (.A(net242),
    .B(net309),
    .C(_0942_),
    .Y(_0129_));
 sg13g2_o21ai_1 _1869_ (.B1(_0929_),
    .Y(_0943_),
    .A1(net211),
    .A2(_0942_));
 sg13g2_a21oi_1 _1870_ (.A1(net211),
    .A2(_0942_),
    .Y(_0130_),
    .B1(_0943_));
 sg13g2_a21oi_1 _1871_ (.A1(\ChiselTop.debounceCounter[9] ),
    .A2(_0942_),
    .Y(_0944_),
    .B1(net187));
 sg13g2_and3_1 _1872_ (.X(_0945_),
    .A(net211),
    .B(net187),
    .C(_0942_));
 sg13g2_nor3_1 _1873_ (.A(net242),
    .B(net188),
    .C(_0945_),
    .Y(_0131_));
 sg13g2_nor2_1 _1874_ (.A(net338),
    .B(_0945_),
    .Y(_0946_));
 sg13g2_and2_1 _1875_ (.A(net338),
    .B(_0945_),
    .X(_0947_));
 sg13g2_nor3_1 _1876_ (.A(net242),
    .B(_0946_),
    .C(_0947_),
    .Y(_0132_));
 sg13g2_nor2_1 _1877_ (.A(net313),
    .B(_0947_),
    .Y(_0948_));
 sg13g2_and2_1 _1878_ (.A(net313),
    .B(_0947_),
    .X(_0949_));
 sg13g2_nor3_1 _1879_ (.A(net242),
    .B(net314),
    .C(_0949_),
    .Y(_0133_));
 sg13g2_and2_1 _1880_ (.A(net373),
    .B(_0949_),
    .X(_0950_));
 sg13g2_o21ai_1 _1881_ (.B1(_0929_),
    .Y(_0951_),
    .A1(net373),
    .A2(_0949_));
 sg13g2_nor2_1 _1882_ (.A(_0950_),
    .B(_0951_),
    .Y(_0134_));
 sg13g2_nor2_1 _1883_ (.A(net339),
    .B(_0950_),
    .Y(_0952_));
 sg13g2_and2_1 _1884_ (.A(net339),
    .B(_0950_),
    .X(_0953_));
 sg13g2_nor3_1 _1885_ (.A(net242),
    .B(net340),
    .C(_0953_),
    .Y(_0135_));
 sg13g2_and4_1 _1886_ (.A(\ChiselTop.debounceCounter[13] ),
    .B(net353),
    .C(net339),
    .D(_0949_),
    .X(_0954_));
 sg13g2_o21ai_1 _1887_ (.B1(_0929_),
    .Y(_0955_),
    .A1(net353),
    .A2(_0953_));
 sg13g2_nor2_1 _1888_ (.A(_0954_),
    .B(_0955_),
    .Y(_0136_));
 sg13g2_o21ai_1 _1889_ (.B1(_0929_),
    .Y(_0956_),
    .A1(net209),
    .A2(_0954_));
 sg13g2_a21oi_1 _1890_ (.A1(net209),
    .A2(_0954_),
    .Y(_0137_),
    .B1(_0956_));
 sg13g2_a21oi_1 _1891_ (.A1(\ChiselTop.debounceCounter[16] ),
    .A2(_0954_),
    .Y(_0957_),
    .B1(net182));
 sg13g2_and4_1 _1892_ (.A(\ChiselTop.debounceCounter[15] ),
    .B(net182),
    .C(net209),
    .D(_0953_),
    .X(_0958_));
 sg13g2_nor3_1 _1893_ (.A(net242),
    .B(net183),
    .C(_0958_),
    .Y(_0138_));
 sg13g2_nor2_1 _1894_ (.A(net311),
    .B(_0958_),
    .Y(_0959_));
 sg13g2_and2_1 _1895_ (.A(net311),
    .B(_0958_),
    .X(_0960_));
 sg13g2_nor3_1 _1896_ (.A(net242),
    .B(net312),
    .C(_0960_),
    .Y(_0139_));
 sg13g2_nor2_1 _1897_ (.A(net299),
    .B(_0960_),
    .Y(_0961_));
 sg13g2_a21oi_1 _1898_ (.A1(net299),
    .A2(_0960_),
    .Y(_0962_),
    .B1(net242));
 sg13g2_nor2b_1 _1899_ (.A(net300),
    .B_N(_0962_),
    .Y(_0140_));
 sg13g2_o21ai_1 _1900_ (.B1(net293),
    .Y(_0169_),
    .A1(net327),
    .A2(net249));
 sg13g2_a21oi_1 _1901_ (.A1(_0404_),
    .A2(net249),
    .Y(_0141_),
    .B1(_0169_));
 sg13g2_o21ai_1 _1902_ (.B1(net293),
    .Y(_0170_),
    .A1(net348),
    .A2(net249));
 sg13g2_a21oi_1 _1903_ (.A1(_0403_),
    .A2(net249),
    .Y(_0142_),
    .B1(_0170_));
 sg13g2_o21ai_1 _1904_ (.B1(net297),
    .Y(_0171_),
    .A1(net205),
    .A2(net250));
 sg13g2_a21oi_1 _1905_ (.A1(_0402_),
    .A2(net250),
    .Y(_0143_),
    .B1(_0171_));
 sg13g2_o21ai_1 _1906_ (.B1(net297),
    .Y(_0172_),
    .A1(net191),
    .A2(net250));
 sg13g2_a21oi_1 _1907_ (.A1(_0401_),
    .A2(net250),
    .Y(_0144_),
    .B1(_0172_));
 sg13g2_o21ai_1 _1908_ (.B1(net296),
    .Y(_0173_),
    .A1(net318),
    .A2(net249));
 sg13g2_a21oi_1 _1909_ (.A1(_0400_),
    .A2(net249),
    .Y(_0145_),
    .B1(_0173_));
 sg13g2_o21ai_1 _1910_ (.B1(net296),
    .Y(_0174_),
    .A1(\ChiselTop.tClkSelectInBounce_pipeReg_0[1] ),
    .A2(net249));
 sg13g2_a21oi_1 _1911_ (.A1(_0399_),
    .A2(net249),
    .Y(_0146_),
    .B1(_0174_));
 sg13g2_and2_1 _1912_ (.A(net295),
    .B(net7),
    .X(_0147_));
 sg13g2_and2_1 _1913_ (.A(net295),
    .B(net8),
    .X(_0148_));
 sg13g2_and2_1 _1914_ (.A(net295),
    .B(net173),
    .X(_0149_));
 sg13g2_and2_1 _1915_ (.A(net295),
    .B(net166),
    .X(_0150_));
 sg13g2_and2_1 _1916_ (.A(net295),
    .B(net6),
    .X(_0151_));
 sg13g2_and2_1 _1917_ (.A(net294),
    .B(net171),
    .X(_0152_));
 sg13g2_and2_1 _1918_ (.A(net295),
    .B(net5),
    .X(_0153_));
 sg13g2_and2_1 _1919_ (.A(net296),
    .B(net172),
    .X(_0154_));
 sg13g2_and2_1 _1920_ (.A(net294),
    .B(net4),
    .X(_0155_));
 sg13g2_and2_1 _1921_ (.A(net294),
    .B(net168),
    .X(_0156_));
 sg13g2_and2_1 _1922_ (.A(net294),
    .B(net3),
    .X(_0157_));
 sg13g2_and2_1 _1923_ (.A(net295),
    .B(net167),
    .X(_0158_));
 sg13g2_and2_1 _1924_ (.A(net294),
    .B(net1),
    .X(_0159_));
 sg13g2_and2_1 _1925_ (.A(net294),
    .B(net2),
    .X(_0160_));
 sg13g2_and2_1 _1926_ (.A(net294),
    .B(net165),
    .X(_0161_));
 sg13g2_and2_1 _1927_ (.A(net294),
    .B(net164),
    .X(_0162_));
 sg13g2_nor3_2 _1928_ (.A(net279),
    .B(net273),
    .C(_0538_),
    .Y(_0175_));
 sg13g2_a22oi_1 _1929_ (.Y(_0176_),
    .B1(_0867_),
    .B2(_0175_),
    .A2(_0538_),
    .A1(_0448_));
 sg13g2_nor2_2 _1930_ (.A(net272),
    .B(\ChiselTop.counterXReg[9] ),
    .Y(_0177_));
 sg13g2_or2_1 _1931_ (.X(_0178_),
    .B(net271),
    .A(net272));
 sg13g2_nand4_1 _1932_ (.B(_0447_),
    .C(_0862_),
    .A(net281),
    .Y(_0179_),
    .D(_0175_));
 sg13g2_o21ai_1 _1933_ (.B1(net280),
    .Y(_0180_),
    .A1(net282),
    .A2(_0853_));
 sg13g2_nor2b_2 _1934_ (.A(net273),
    .B_N(_0544_),
    .Y(_0181_));
 sg13g2_a21oi_1 _1935_ (.A1(_0180_),
    .A2(_0181_),
    .Y(_0182_),
    .B1(_0176_));
 sg13g2_nand3_1 _1936_ (.B(_0179_),
    .C(_0182_),
    .A(_0177_),
    .Y(_0183_));
 sg13g2_nor2b_2 _1937_ (.A(net258),
    .B_N(net260),
    .Y(_0184_));
 sg13g2_nor2b_1 _1938_ (.A(net261),
    .B_N(net264),
    .Y(_0185_));
 sg13g2_nand2b_1 _1939_ (.Y(_0186_),
    .B(net264),
    .A_N(net261));
 sg13g2_o21ai_1 _1940_ (.B1(_0002_),
    .Y(_0187_),
    .A1(_0011_),
    .A2(_0186_));
 sg13g2_nand2_1 _1941_ (.Y(_0188_),
    .A(_0184_),
    .B(_0185_));
 sg13g2_a21oi_1 _1942_ (.A1(_0184_),
    .A2(_0187_),
    .Y(_0189_),
    .B1(_0450_));
 sg13g2_nor3_1 _1943_ (.A(net266),
    .B(_0892_),
    .C(_0188_),
    .Y(_0190_));
 sg13g2_nand2b_1 _1944_ (.Y(_0191_),
    .B(net258),
    .A_N(net260));
 sg13g2_nor2_2 _1945_ (.A(_0905_),
    .B(_0191_),
    .Y(_0192_));
 sg13g2_nand2b_2 _1946_ (.Y(_0193_),
    .B(_0549_),
    .A_N(_0463_));
 sg13g2_and2_1 _1947_ (.A(_0192_),
    .B(_0193_),
    .X(_0194_));
 sg13g2_nand2_1 _1948_ (.Y(_0195_),
    .A(net255),
    .B(_0455_));
 sg13g2_or4_2 _1949_ (.A(_0189_),
    .B(_0190_),
    .C(_0194_),
    .D(_0195_),
    .X(_0196_));
 sg13g2_nor2_1 _1950_ (.A(_0014_),
    .B(_0196_),
    .Y(_0197_));
 sg13g2_nor2b_1 _1951_ (.A(net255),
    .B_N(net258),
    .Y(_0198_));
 sg13g2_nor4_1 _1952_ (.A(net256),
    .B(_0455_),
    .C(_0549_),
    .D(_0905_),
    .Y(_0199_));
 sg13g2_o21ai_1 _1953_ (.B1(_0184_),
    .Y(_0200_),
    .A1(_0882_),
    .A2(_0898_));
 sg13g2_and2_1 _1954_ (.A(_0012_),
    .B(_0200_),
    .X(_0201_));
 sg13g2_a21o_2 _1955_ (.A2(_0201_),
    .A1(net256),
    .B1(_0199_),
    .X(_0202_));
 sg13g2_a21oi_1 _1956_ (.A1(\ChiselTop.hourDecReg[1] ),
    .A2(_0202_),
    .Y(_0203_),
    .B1(_0197_));
 sg13g2_nand2_1 _1957_ (.Y(_0204_),
    .A(net275),
    .B(net274));
 sg13g2_nor3_1 _1958_ (.A(net279),
    .B(net276),
    .C(_0204_),
    .Y(_0205_));
 sg13g2_nor2_1 _1959_ (.A(net281),
    .B(_0447_),
    .Y(_0206_));
 sg13g2_nand2_1 _1960_ (.Y(_0207_),
    .A(_0862_),
    .B(_0206_));
 sg13g2_nor4_1 _1961_ (.A(net278),
    .B(net276),
    .C(_0204_),
    .D(_0207_),
    .Y(_0208_));
 sg13g2_nor2_1 _1962_ (.A(_0542_),
    .B(_0204_),
    .Y(_0209_));
 sg13g2_nor2_1 _1963_ (.A(_0178_),
    .B(_0209_),
    .Y(_0210_));
 sg13g2_o21ai_1 _1964_ (.B1(_0210_),
    .Y(_0211_),
    .A1(net273),
    .A2(_0537_));
 sg13g2_nand2_1 _1965_ (.Y(_0212_),
    .A(net252),
    .B(_0175_));
 sg13g2_o21ai_1 _1966_ (.B1(_0212_),
    .Y(_0213_),
    .A1(_0180_),
    .A2(_0204_));
 sg13g2_nor3_2 _1967_ (.A(_0208_),
    .B(_0211_),
    .C(_0213_),
    .Y(_0214_));
 sg13g2_nand4_1 _1968_ (.B(net270),
    .C(\ChiselTop.counterYReg[0] ),
    .A(net268),
    .Y(_0215_),
    .D(_0013_));
 sg13g2_nand3b_1 _1969_ (.B(_0883_),
    .C(_0215_),
    .Y(_0216_),
    .A_N(net267));
 sg13g2_inv_1 _1970_ (.Y(_0217_),
    .A(_0216_));
 sg13g2_o21ai_1 _1971_ (.B1(net262),
    .Y(_0218_),
    .A1(net264),
    .A2(_0472_));
 sg13g2_a21o_1 _1972_ (.A2(_0472_),
    .A1(net261),
    .B1(_0904_),
    .X(_0219_));
 sg13g2_nor2_2 _1973_ (.A(net258),
    .B(net260),
    .Y(_0220_));
 sg13g2_nand2_1 _1974_ (.Y(_0221_),
    .A(_0218_),
    .B(_0220_));
 sg13g2_a21oi_1 _1975_ (.A1(net258),
    .A2(_0216_),
    .Y(_0222_),
    .B1(net255));
 sg13g2_nand2_2 _1976_ (.Y(_0223_),
    .A(_0221_),
    .B(_0222_));
 sg13g2_nor2_1 _1977_ (.A(_0017_),
    .B(_0223_),
    .Y(_0224_));
 sg13g2_and2_1 _1978_ (.A(net254),
    .B(_0463_),
    .X(_0225_));
 sg13g2_a22oi_1 _1979_ (.Y(_0226_),
    .B1(_0225_),
    .B2(_0460_),
    .A2(_0219_),
    .A1(_0454_));
 sg13g2_nand2_1 _1980_ (.Y(_0227_),
    .A(_0884_),
    .B(_0198_));
 sg13g2_a221oi_1 _1981_ (.B2(_0460_),
    .C1(_0227_),
    .B1(_0225_),
    .A1(_0454_),
    .Y(_0228_),
    .A2(_0219_));
 sg13g2_a221oi_1 _1982_ (.B2(_0451_),
    .C1(_0224_),
    .B1(_0228_),
    .A1(\ChiselTop.hourUniReg[1] ),
    .Y(_0229_),
    .A2(_0202_));
 sg13g2_o21ai_1 _1983_ (.B1(_0229_),
    .Y(_0230_),
    .A1(_0015_),
    .A2(_0196_));
 sg13g2_nand2_1 _1984_ (.Y(_0231_),
    .A(_0214_),
    .B(_0230_));
 sg13g2_o21ai_1 _1985_ (.B1(_0231_),
    .Y(_0232_),
    .A1(_0183_),
    .A2(_0203_));
 sg13g2_o21ai_1 _1986_ (.B1(_0857_),
    .Y(_0233_),
    .A1(_0539_),
    .A2(_0867_));
 sg13g2_and2_1 _1987_ (.A(net272),
    .B(_0233_),
    .X(_0234_));
 sg13g2_nand3_1 _1988_ (.B(_0177_),
    .C(_0180_),
    .A(_0856_),
    .Y(_0235_));
 sg13g2_nand2b_1 _1989_ (.Y(_0236_),
    .B(_0235_),
    .A_N(_0210_));
 sg13g2_nand2b_1 _1990_ (.Y(_0237_),
    .B(_0857_),
    .A_N(_0539_));
 sg13g2_nor4_1 _1991_ (.A(\ChiselTop.counterXReg[0] ),
    .B(net280),
    .C(_0852_),
    .D(_0237_),
    .Y(_0238_));
 sg13g2_nor4_2 _1992_ (.A(net271),
    .B(_0234_),
    .C(_0236_),
    .Y(_0239_),
    .D(_0238_));
 sg13g2_nand2b_1 _1993_ (.Y(_0240_),
    .B(_0228_),
    .A_N(_0010_));
 sg13g2_and2_1 _1994_ (.A(\ChiselTop.minuteDecReg[1] ),
    .B(_0202_),
    .X(_0241_));
 sg13g2_o21ai_1 _1995_ (.B1(_0240_),
    .Y(_0242_),
    .A1(_0018_),
    .A2(_0196_));
 sg13g2_o21ai_1 _1996_ (.B1(_0239_),
    .Y(_0243_),
    .A1(_0241_),
    .A2(_0242_));
 sg13g2_nor2b_1 _1997_ (.A(net275),
    .B_N(net274),
    .Y(_0244_));
 sg13g2_nand2_1 _1998_ (.Y(_0245_),
    .A(_0856_),
    .B(_0244_));
 sg13g2_nor2b_1 _1999_ (.A(_0245_),
    .B_N(_0180_),
    .Y(_0246_));
 sg13g2_nor3_1 _2000_ (.A(_0544_),
    .B(_0877_),
    .C(_0246_),
    .Y(_0247_));
 sg13g2_o21ai_1 _2001_ (.B1(_0449_),
    .Y(_0248_),
    .A1(_0207_),
    .A2(_0245_));
 sg13g2_nor2_1 _2002_ (.A(_0247_),
    .B(_0248_),
    .Y(_0249_));
 sg13g2_o21ai_1 _2003_ (.B1(_0857_),
    .Y(_0250_),
    .A1(_0539_),
    .A2(net252));
 sg13g2_nand3_1 _2004_ (.B(_0249_),
    .C(_0250_),
    .A(\ChiselTop.counterXReg[8] ),
    .Y(_0251_));
 sg13g2_nand2b_1 _2005_ (.Y(_0252_),
    .B(_0228_),
    .A_N(_0020_));
 sg13g2_o21ai_1 _2006_ (.B1(_0252_),
    .Y(_0253_),
    .A1(_0021_),
    .A2(_0223_));
 sg13g2_nor2_1 _2007_ (.A(_0019_),
    .B(_0196_),
    .Y(_0254_));
 sg13g2_and2_1 _2008_ (.A(\ChiselTop.minuteUniReg[1] ),
    .B(_0202_),
    .X(_0255_));
 sg13g2_nor3_1 _2009_ (.A(_0253_),
    .B(_0254_),
    .C(_0255_),
    .Y(_0256_));
 sg13g2_o21ai_1 _2010_ (.B1(_0243_),
    .Y(_0257_),
    .A1(_0251_),
    .A2(_0256_));
 sg13g2_nand3b_1 _2011_ (.B(net276),
    .C(_0244_),
    .Y(_0258_),
    .A_N(net278));
 sg13g2_nand2b_1 _2012_ (.Y(_0259_),
    .B(_0180_),
    .A_N(_0258_));
 sg13g2_nand4_1 _2013_ (.B(net272),
    .C(_0543_),
    .A(net273),
    .Y(_0260_),
    .D(_0259_));
 sg13g2_and2_1 _2014_ (.A(_0541_),
    .B(_0181_),
    .X(_0261_));
 sg13g2_nand3_1 _2015_ (.B(_0852_),
    .C(_0261_),
    .A(_0447_),
    .Y(_0262_));
 sg13g2_o21ai_1 _2016_ (.B1(_0262_),
    .Y(_0263_),
    .A1(net271),
    .A2(_0260_));
 sg13g2_nand2_1 _2017_ (.Y(_0264_),
    .A(\ChiselTop.secondDecReg[1] ),
    .B(_0202_));
 sg13g2_nor2b_1 _2018_ (.A(_0009_),
    .B_N(_0228_),
    .Y(_0265_));
 sg13g2_o21ai_1 _2019_ (.B1(_0264_),
    .Y(_0266_),
    .A1(_0022_),
    .A2(_0196_));
 sg13g2_o21ai_1 _2020_ (.B1(_0263_),
    .Y(_0267_),
    .A1(_0265_),
    .A2(_0266_));
 sg13g2_nand4_1 _2021_ (.B(net280),
    .C(_0862_),
    .A(net281),
    .Y(_0268_),
    .D(_0261_));
 sg13g2_nor3_1 _2022_ (.A(_0447_),
    .B(net279),
    .C(_0852_),
    .Y(_0269_));
 sg13g2_nand2_1 _2023_ (.Y(_0270_),
    .A(_0027_),
    .B(_0546_));
 sg13g2_nor3_1 _2024_ (.A(_0543_),
    .B(_0269_),
    .C(_0270_),
    .Y(_0271_));
 sg13g2_nor2_1 _2025_ (.A(\ChiselTop.counterXReg[1] ),
    .B(net281),
    .Y(_0272_));
 sg13g2_nor3_1 _2026_ (.A(_0447_),
    .B(net279),
    .C(_0272_),
    .Y(_0273_));
 sg13g2_a21oi_1 _2027_ (.A1(_0538_),
    .A2(_0546_),
    .Y(_0274_),
    .B1(_0449_));
 sg13g2_o21ai_1 _2028_ (.B1(_0274_),
    .Y(_0275_),
    .A1(_0270_),
    .A2(_0273_));
 sg13g2_nand2_1 _2029_ (.Y(_0276_),
    .A(_0268_),
    .B(_0275_));
 sg13g2_nor3_2 _2030_ (.A(_0026_),
    .B(_0271_),
    .C(_0276_),
    .Y(_0277_));
 sg13g2_nand2b_1 _2031_ (.Y(_0278_),
    .B(_0228_),
    .A_N(_0025_));
 sg13g2_o21ai_1 _2032_ (.B1(_0278_),
    .Y(_0279_),
    .A1(_0024_),
    .A2(_0223_));
 sg13g2_nand2_1 _2033_ (.Y(_0280_),
    .A(\ChiselTop.secondUniReg[1] ),
    .B(_0202_));
 sg13g2_o21ai_1 _2034_ (.B1(_0280_),
    .Y(_0281_),
    .A1(_0023_),
    .A2(_0196_));
 sg13g2_o21ai_1 _2035_ (.B1(_0277_),
    .Y(_0282_),
    .A1(_0279_),
    .A2(_0281_));
 sg13g2_a21oi_2 _2036_ (.B1(_0257_),
    .Y(_0283_),
    .A2(_0282_),
    .A1(_0267_));
 sg13g2_a22oi_1 _2037_ (.Y(_0284_),
    .B1(_0283_),
    .B2(net412),
    .A2(_0257_),
    .A1(\ChiselTop.lfsrReg_6 ));
 sg13g2_nor2_1 _2038_ (.A(net235),
    .B(_0284_),
    .Y(_0285_));
 sg13g2_nand2_1 _2039_ (.Y(_0286_),
    .A(net258),
    .B(net268));
 sg13g2_nor2_1 _2040_ (.A(net267),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_nand4_1 _2041_ (.B(_0474_),
    .C(_0904_),
    .A(net260),
    .Y(_0288_),
    .D(_0287_));
 sg13g2_o21ai_1 _2042_ (.B1(net256),
    .Y(_0289_),
    .A1(_0459_),
    .A2(_0188_));
 sg13g2_nor2_1 _2043_ (.A(_0473_),
    .B(_0882_),
    .Y(_0290_));
 sg13g2_a22oi_1 _2044_ (.Y(_0291_),
    .B1(_0290_),
    .B2(_0184_),
    .A2(_0192_),
    .A1(_0549_));
 sg13g2_nor2_1 _2045_ (.A(_0461_),
    .B(_0291_),
    .Y(_0292_));
 sg13g2_a21oi_1 _2046_ (.A1(_0474_),
    .A2(_0289_),
    .Y(_0293_),
    .B1(_0292_));
 sg13g2_a21oi_1 _2047_ (.A1(_0405_),
    .A2(_0288_),
    .Y(_0294_),
    .B1(_0293_));
 sg13g2_nor2_1 _2048_ (.A(_0186_),
    .B(_0191_),
    .Y(_0295_));
 sg13g2_a21o_1 _2049_ (.A2(_0295_),
    .A1(_0551_),
    .B1(_0462_),
    .X(_0296_));
 sg13g2_a21oi_1 _2050_ (.A1(_0013_),
    .A2(_0296_),
    .Y(_0297_),
    .B1(_0294_));
 sg13g2_nor2_1 _2051_ (.A(_0239_),
    .B(_0263_),
    .Y(_0298_));
 sg13g2_or2_1 _2052_ (.X(_0299_),
    .B(_0298_),
    .A(_0297_));
 sg13g2_nand2_1 _2053_ (.Y(_0300_),
    .A(net272),
    .B(_0449_));
 sg13g2_nor2_1 _2054_ (.A(_0237_),
    .B(_0300_),
    .Y(_0301_));
 sg13g2_a221oi_1 _2055_ (.B2(_0541_),
    .C1(_0301_),
    .B1(_0181_),
    .A1(_0175_),
    .Y(_0302_),
    .A2(_0177_));
 sg13g2_nor2_1 _2056_ (.A(net252),
    .B(_0302_),
    .Y(_0303_));
 sg13g2_a22oi_1 _2057_ (.Y(_0304_),
    .B1(_0177_),
    .B2(_0205_),
    .A2(_0175_),
    .A1(_0541_));
 sg13g2_o21ai_1 _2058_ (.B1(_0304_),
    .Y(_0305_),
    .A1(_0245_),
    .A2(_0300_));
 sg13g2_nor3_1 _2059_ (.A(net281),
    .B(_0447_),
    .C(_0863_),
    .Y(_0306_));
 sg13g2_a21oi_1 _2060_ (.A1(_0305_),
    .A2(_0306_),
    .Y(_0307_),
    .B1(_0303_));
 sg13g2_nand4_1 _2061_ (.B(net273),
    .C(_0856_),
    .A(net275),
    .Y(_0308_),
    .D(_0177_));
 sg13g2_o21ai_1 _2062_ (.B1(_0308_),
    .Y(_0309_),
    .A1(_0258_),
    .A2(_0300_));
 sg13g2_nand3_1 _2063_ (.B(_0206_),
    .C(_0309_),
    .A(_0853_),
    .Y(_0310_));
 sg13g2_nor3_1 _2064_ (.A(_0446_),
    .B(net280),
    .C(_0863_),
    .Y(_0311_));
 sg13g2_o21ai_1 _2065_ (.B1(_0311_),
    .Y(_0312_),
    .A1(_0261_),
    .A2(_0301_));
 sg13g2_nand3_1 _2066_ (.B(_0310_),
    .C(_0312_),
    .A(_0307_),
    .Y(_0313_));
 sg13g2_nand3_1 _2067_ (.B(_0881_),
    .C(_0192_),
    .A(net255),
    .Y(_0314_));
 sg13g2_nor2_1 _2068_ (.A(_0236_),
    .B(_0314_),
    .Y(_0315_));
 sg13g2_a21oi_1 _2069_ (.A1(net265),
    .A2(_0550_),
    .Y(_0316_),
    .B1(net263));
 sg13g2_nor3_1 _2070_ (.A(net270),
    .B(_0407_),
    .C(net254),
    .Y(_0317_));
 sg13g2_nand4_1 _2071_ (.B(_0287_),
    .C(_0316_),
    .A(net260),
    .Y(_0318_),
    .D(_0317_));
 sg13g2_and3_1 _2072_ (.X(_0319_),
    .A(_0456_),
    .B(_0881_),
    .C(_0220_));
 sg13g2_nor4_1 _2073_ (.A(net267),
    .B(_0461_),
    .C(_0884_),
    .D(_0286_),
    .Y(_0320_));
 sg13g2_o21ai_1 _2074_ (.B1(_0013_),
    .Y(_0321_),
    .A1(_0319_),
    .A2(_0320_));
 sg13g2_nor2_1 _2075_ (.A(_0214_),
    .B(_0277_),
    .Y(_0322_));
 sg13g2_a22oi_1 _2076_ (.Y(_0323_),
    .B1(_0322_),
    .B2(_0251_),
    .A2(_0321_),
    .A1(_0297_));
 sg13g2_nand2b_1 _2077_ (.Y(_0324_),
    .B(_0196_),
    .A_N(_0202_));
 sg13g2_nand3_1 _2078_ (.B(_0181_),
    .C(_0206_),
    .A(_0853_),
    .Y(_0325_));
 sg13g2_nand2_1 _2079_ (.Y(_0326_),
    .A(_0175_),
    .B(_0311_));
 sg13g2_a21oi_1 _2080_ (.A1(_0325_),
    .A2(_0326_),
    .Y(_0327_),
    .B1(_0178_));
 sg13g2_o21ai_1 _2081_ (.B1(_0324_),
    .Y(_0328_),
    .A1(_0313_),
    .A2(_0327_));
 sg13g2_nand2b_1 _2082_ (.Y(_0329_),
    .B(_0294_),
    .A_N(_0183_));
 sg13g2_nand3_1 _2083_ (.B(_0546_),
    .C(_0873_),
    .A(net271),
    .Y(_0330_));
 sg13g2_nand4_1 _2084_ (.B(_0177_),
    .C(_0181_),
    .A(_0866_),
    .Y(_0331_),
    .D(_0272_));
 sg13g2_nand4_1 _2085_ (.B(_0454_),
    .C(_0898_),
    .A(net255),
    .Y(_0332_),
    .D(_0185_));
 sg13g2_nor2_1 _2086_ (.A(net258),
    .B(_0884_),
    .Y(_0333_));
 sg13g2_nand3_1 _2087_ (.B(_0551_),
    .C(_0333_),
    .A(net254),
    .Y(_0334_));
 sg13g2_and4_1 _2088_ (.A(_0330_),
    .B(_0331_),
    .C(_0332_),
    .D(_0334_),
    .X(_0335_));
 sg13g2_o21ai_1 _2089_ (.B1(_0329_),
    .Y(_0336_),
    .A1(uio_out[7]),
    .A2(_0335_));
 sg13g2_nor2_1 _2090_ (.A(_0223_),
    .B(_0307_),
    .Y(_0337_));
 sg13g2_a21oi_1 _2091_ (.A1(_0228_),
    .A2(_0313_),
    .Y(_0338_),
    .B1(_0323_));
 sg13g2_a22oi_1 _2092_ (.Y(_0339_),
    .B1(_0314_),
    .B2(_0318_),
    .A2(_0260_),
    .A1(_0449_));
 sg13g2_a22oi_1 _2093_ (.Y(_0340_),
    .B1(_0339_),
    .B2(_0275_),
    .A2(_0315_),
    .A1(_0249_));
 sg13g2_nor2_1 _2094_ (.A(uio_out[6]),
    .B(_0340_),
    .Y(_0341_));
 sg13g2_nor3_1 _2095_ (.A(_0336_),
    .B(_0337_),
    .C(_0341_),
    .Y(_0342_));
 sg13g2_nand4_1 _2096_ (.B(_0328_),
    .C(_0338_),
    .A(_0299_),
    .Y(_0343_),
    .D(_0342_));
 sg13g2_nand3b_1 _2097_ (.B(_0220_),
    .C(net257),
    .Y(_0344_),
    .A_N(net261));
 sg13g2_nor2_1 _2098_ (.A(_0900_),
    .B(_0344_),
    .Y(_0345_));
 sg13g2_or2_1 _2099_ (.X(_0346_),
    .B(net266),
    .A(net261));
 sg13g2_nor4_1 _2100_ (.A(net257),
    .B(\ChiselTop.counterYReg[3] ),
    .C(_0893_),
    .D(_0188_),
    .Y(_0347_));
 sg13g2_or3_1 _2101_ (.A(net257),
    .B(net262),
    .C(_0455_),
    .X(_0348_));
 sg13g2_nand2_1 _2102_ (.Y(_0349_),
    .A(_0463_),
    .B(_0549_));
 sg13g2_inv_1 _2103_ (.Y(_0350_),
    .A(_0349_));
 sg13g2_a21oi_1 _2104_ (.A1(net264),
    .A2(_0193_),
    .Y(_0351_),
    .B1(_0348_));
 sg13g2_nor4_1 _2105_ (.A(_0199_),
    .B(_0345_),
    .C(_0347_),
    .D(_0351_),
    .Y(_0352_));
 sg13g2_nor3_1 _2106_ (.A(_0465_),
    .B(_0549_),
    .C(_0905_),
    .Y(_0353_));
 sg13g2_nor3_1 _2107_ (.A(_0472_),
    .B(_0549_),
    .C(_0882_),
    .Y(_0354_));
 sg13g2_nor2_1 _2108_ (.A(_0353_),
    .B(_0354_),
    .Y(_0355_));
 sg13g2_a21oi_1 _2109_ (.A1(net254),
    .A2(_0465_),
    .Y(_0356_),
    .B1(_0355_));
 sg13g2_nand3_1 _2110_ (.B(_0456_),
    .C(_0892_),
    .A(net266),
    .Y(_0357_));
 sg13g2_a22oi_1 _2111_ (.Y(_0358_),
    .B1(_0185_),
    .B2(_0472_),
    .A2(_0549_),
    .A1(_0456_));
 sg13g2_o21ai_1 _2112_ (.B1(_0357_),
    .Y(_0359_),
    .A1(_0350_),
    .A2(_0358_));
 sg13g2_o21ai_1 _2113_ (.B1(_0184_),
    .Y(_0360_),
    .A1(_0356_),
    .A2(_0359_));
 sg13g2_a22oi_1 _2114_ (.Y(_0361_),
    .B1(_0906_),
    .B2(_0406_),
    .A2(_0898_),
    .A1(net254));
 sg13g2_a221oi_1 _2115_ (.B2(net254),
    .C1(_0218_),
    .B1(_0350_),
    .A1(net264),
    .Y(_0362_),
    .A2(_0550_));
 sg13g2_o21ai_1 _2116_ (.B1(_0220_),
    .Y(_0363_),
    .A1(_0361_),
    .A2(_0362_));
 sg13g2_a22oi_1 _2117_ (.Y(_0364_),
    .B1(_0473_),
    .B2(_0904_),
    .A2(_0456_),
    .A1(net266));
 sg13g2_nand3_1 _2118_ (.B(_0463_),
    .C(_0904_),
    .A(net266),
    .Y(_0365_));
 sg13g2_nand2b_1 _2119_ (.Y(_0366_),
    .B(_0365_),
    .A_N(_0364_));
 sg13g2_o21ai_1 _2120_ (.B1(_0186_),
    .Y(_0367_),
    .A1(_0457_),
    .A2(_0193_));
 sg13g2_nand2b_1 _2121_ (.Y(_0368_),
    .B(_0367_),
    .A_N(_0885_));
 sg13g2_a21o_1 _2122_ (.A2(_0368_),
    .A1(_0366_),
    .B1(_0191_),
    .X(_0369_));
 sg13g2_nand4_1 _2123_ (.B(_0882_),
    .C(_0226_),
    .A(_0454_),
    .Y(_0370_),
    .D(_0346_));
 sg13g2_a21oi_1 _2124_ (.A1(_0456_),
    .A2(_0193_),
    .Y(_0371_),
    .B1(_0221_));
 sg13g2_nor2_1 _2125_ (.A(net254),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_a21oi_1 _2126_ (.A1(_0198_),
    .A2(_0217_),
    .Y(_0373_),
    .B1(_0372_));
 sg13g2_nand3_1 _2127_ (.B(_0220_),
    .C(_0350_),
    .A(_0456_),
    .Y(_0374_));
 sg13g2_nand4_1 _2128_ (.B(_0363_),
    .C(_0369_),
    .A(_0360_),
    .Y(_0375_),
    .D(_0370_));
 sg13g2_nand2_1 _2129_ (.Y(_0376_),
    .A(_0405_),
    .B(_0375_));
 sg13g2_a21oi_1 _2130_ (.A1(_0201_),
    .A2(_0374_),
    .Y(_0377_),
    .B1(_0405_));
 sg13g2_or2_1 _2131_ (.X(_0378_),
    .B(_0377_),
    .A(_0373_));
 sg13g2_nand4_1 _2132_ (.B(_0352_),
    .C(_0376_),
    .A(_0196_),
    .Y(_0379_),
    .D(_0378_));
 sg13g2_nor4_1 _2133_ (.A(net281),
    .B(net280),
    .C(_0540_),
    .D(_0854_),
    .Y(_0380_));
 sg13g2_nand4_1 _2134_ (.B(_0546_),
    .C(_0379_),
    .A(net271),
    .Y(_0381_),
    .D(_0380_));
 sg13g2_nor2b_2 _2135_ (.A(_0343_),
    .B_N(_0381_),
    .Y(_0382_));
 sg13g2_a21oi_1 _2136_ (.A1(net437),
    .A2(net235),
    .Y(_0383_),
    .B1(_0285_));
 sg13g2_a21oi_1 _2137_ (.A1(_0382_),
    .A2(_0383_),
    .Y(_0163_),
    .B1(_0553_));
 sg13g2_a22oi_1 _2138_ (.Y(_0384_),
    .B1(_0283_),
    .B2(\ChiselTop.lfsrReg_13 ),
    .A2(_0257_),
    .A1(\ChiselTop.lfsrReg_7 ));
 sg13g2_nor2_1 _2139_ (.A(net235),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_a21oi_1 _2140_ (.A1(net445),
    .A2(net236),
    .Y(_0386_),
    .B1(_0385_));
 sg13g2_a21oi_1 _2141_ (.A1(_0382_),
    .A2(net446),
    .Y(_0164_),
    .B1(_0553_));
 sg13g2_a22oi_1 _2142_ (.Y(_0387_),
    .B1(_0283_),
    .B2(net417),
    .A2(_0257_),
    .A1(net406));
 sg13g2_nor2_1 _2143_ (.A(net236),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_a21oi_1 _2144_ (.A1(net402),
    .A2(net236),
    .Y(_0389_),
    .B1(_0388_));
 sg13g2_a21oi_1 _2145_ (.A1(_0382_),
    .A2(_0389_),
    .Y(_0165_),
    .B1(_0553_));
 sg13g2_a22oi_1 _2146_ (.Y(_0390_),
    .B1(_0283_),
    .B2(net422),
    .A2(_0257_),
    .A1(\ChiselTop.lfsrReg_9 ));
 sg13g2_nor2_1 _2147_ (.A(net235),
    .B(_0390_),
    .Y(_0391_));
 sg13g2_a21oi_1 _2148_ (.A1(net429),
    .A2(net236),
    .Y(_0392_),
    .B1(_0391_));
 sg13g2_a21oi_1 _2149_ (.A1(_0382_),
    .A2(_0392_),
    .Y(_0166_),
    .B1(_0553_));
 sg13g2_a22oi_1 _2150_ (.Y(_0393_),
    .B1(_0283_),
    .B2(net420),
    .A2(_0257_),
    .A1(\ChiselTop.lfsrReg_10 ));
 sg13g2_nor2_1 _2151_ (.A(net235),
    .B(_0393_),
    .Y(_0394_));
 sg13g2_a21oi_1 _2152_ (.A1(net410),
    .A2(net235),
    .Y(_0395_),
    .B1(_0394_));
 sg13g2_a21oi_1 _2153_ (.A1(_0382_),
    .A2(_0395_),
    .Y(_0167_),
    .B1(_0553_));
 sg13g2_a22oi_1 _2154_ (.Y(_0396_),
    .B1(_0283_),
    .B2(\ChiselTop.lfsrReg_17 ),
    .A2(_0257_),
    .A1(net400));
 sg13g2_nor2_1 _2155_ (.A(net235),
    .B(net409),
    .Y(_0397_));
 sg13g2_a21oi_1 _2156_ (.A1(net404),
    .A2(net235),
    .Y(_0398_),
    .B1(_0397_));
 sg13g2_a21oi_1 _2157_ (.A1(_0382_),
    .A2(_0398_),
    .Y(_0168_),
    .B1(_0553_));
 sg13g2_dfrbp_1 _2158_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net146),
    .D(_0028_),
    .Q_N(_1073_),
    .Q(\ChiselTop.tClkReqReg ));
 sg13g2_dfrbp_1 _2159_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net37),
    .D(net163),
    .Q_N(\ChiselTop._modeReg_T_1[0] ),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _2160_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net35),
    .D(net379),
    .Q_N(_1072_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _2161_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net33),
    .D(_0031_),
    .Q_N(_1071_),
    .Q(\ChiselTop.lfsrReg_17 ));
 sg13g2_dfrbp_1 _2162_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net31),
    .D(net421),
    .Q_N(_1070_),
    .Q(\ChiselTop.lfsrReg_16 ));
 sg13g2_dfrbp_1 _2163_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net29),
    .D(_0033_),
    .Q_N(_1069_),
    .Q(\ChiselTop.lfsrReg_15 ));
 sg13g2_dfrbp_1 _2164_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net27),
    .D(_0034_),
    .Q_N(_1068_),
    .Q(\ChiselTop.lfsrReg_14 ));
 sg13g2_dfrbp_1 _2165_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net25),
    .D(_0035_),
    .Q_N(_1067_),
    .Q(\ChiselTop.lfsrReg_13 ));
 sg13g2_dfrbp_1 _2166_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net23),
    .D(_0036_),
    .Q_N(_1066_),
    .Q(\ChiselTop.lfsrReg_12 ));
 sg13g2_dfrbp_1 _2167_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net21),
    .D(net401),
    .Q_N(_1065_),
    .Q(\ChiselTop.lfsrReg_11 ));
 sg13g2_dfrbp_1 _2168_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net19),
    .D(_0038_),
    .Q_N(_1064_),
    .Q(\ChiselTop.lfsrReg_10 ));
 sg13g2_dfrbp_1 _2169_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net17),
    .D(_0039_),
    .Q_N(_1063_),
    .Q(\ChiselTop.lfsrReg_9 ));
 sg13g2_dfrbp_1 _2170_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net15),
    .D(net407),
    .Q_N(_1062_),
    .Q(\ChiselTop.lfsrReg_8 ));
 sg13g2_dfrbp_1 _2171_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net13),
    .D(net419),
    .Q_N(_1061_),
    .Q(\ChiselTop.lfsrReg_7 ));
 sg13g2_dfrbp_1 _2172_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net11),
    .D(_0042_),
    .Q_N(_1060_),
    .Q(\ChiselTop.lfsrReg_6 ));
 sg13g2_dfrbp_1 _2173_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net9),
    .D(net405),
    .Q_N(_1059_),
    .Q(\ChiselTop.lfsrReg_5 ));
 sg13g2_dfrbp_1 _2174_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net149),
    .D(net411),
    .Q_N(_1058_),
    .Q(\ChiselTop.lfsrReg_4 ));
 sg13g2_dfrbp_1 _2175_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net147),
    .D(_0045_),
    .Q_N(_1057_),
    .Q(\ChiselTop.lfsrReg_3 ));
 sg13g2_dfrbp_1 _2176_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net144),
    .D(net403),
    .Q_N(_1056_),
    .Q(\ChiselTop.lfsrReg_2 ));
 sg13g2_dfrbp_1 _2177_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net142),
    .D(net438),
    .Q_N(_1055_),
    .Q(\ChiselTop.lfsrReg_1 ));
 sg13g2_dfrbp_1 _2178_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net140),
    .D(_0048_),
    .Q_N(_1054_),
    .Q(\ChiselTop.lfsrReg_0 ));
 sg13g2_dfrbp_1 _2179_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net138),
    .D(_0049_),
    .Q_N(_0023_),
    .Q(\ChiselTop.secondUniReg[0] ));
 sg13g2_dfrbp_1 _2180_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net136),
    .D(net381),
    .Q_N(_1053_),
    .Q(\ChiselTop.secondUniReg[1] ));
 sg13g2_dfrbp_1 _2181_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net134),
    .D(net170),
    .Q_N(_0025_),
    .Q(\ChiselTop.secondUniReg[2] ));
 sg13g2_dfrbp_1 _2182_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net132),
    .D(net333),
    .Q_N(_0024_),
    .Q(\ChiselTop.secondUniReg[3] ));
 sg13g2_dfrbp_1 _2183_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net130),
    .D(net201),
    .Q_N(_0022_),
    .Q(\ChiselTop.secondDecReg[0] ));
 sg13g2_dfrbp_1 _2184_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net128),
    .D(net414),
    .Q_N(_1052_),
    .Q(\ChiselTop.secondDecReg[1] ));
 sg13g2_dfrbp_1 _2185_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net126),
    .D(net219),
    .Q_N(_0009_),
    .Q(\ChiselTop.secondDecReg[2] ));
 sg13g2_dfrbp_1 _2186_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net124),
    .D(net386),
    .Q_N(_0019_),
    .Q(\ChiselTop.minuteUniReg[0] ));
 sg13g2_dfrbp_1 _2187_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net122),
    .D(_0057_),
    .Q_N(_1051_),
    .Q(\ChiselTop.minuteUniReg[1] ));
 sg13g2_dfrbp_1 _2188_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net120),
    .D(net370),
    .Q_N(_0020_),
    .Q(\ChiselTop.minuteUniReg[2] ));
 sg13g2_dfrbp_1 _2189_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net118),
    .D(net399),
    .Q_N(_0021_),
    .Q(\ChiselTop.minuteUniReg[3] ));
 sg13g2_dfrbp_1 _2190_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net116),
    .D(net321),
    .Q_N(_0018_),
    .Q(\ChiselTop.minuteDecReg[0] ));
 sg13g2_dfrbp_1 _2191_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net114),
    .D(_0061_),
    .Q_N(_1050_),
    .Q(\ChiselTop.minuteDecReg[1] ));
 sg13g2_dfrbp_1 _2192_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net112),
    .D(net180),
    .Q_N(_0010_),
    .Q(\ChiselTop.minuteDecReg[2] ));
 sg13g2_dfrbp_1 _2193_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net110),
    .D(net393),
    .Q_N(_0015_),
    .Q(\ChiselTop.hourUniReg[0] ));
 sg13g2_dfrbp_1 _2194_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net108),
    .D(_0064_),
    .Q_N(_1049_),
    .Q(\ChiselTop.hourUniReg[1] ));
 sg13g2_dfrbp_1 _2195_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net106),
    .D(net388),
    .Q_N(_0016_),
    .Q(\ChiselTop.hourUniReg[2] ));
 sg13g2_dfrbp_1 _2196_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net104),
    .D(net395),
    .Q_N(_0017_),
    .Q(\ChiselTop.hourUniReg[3] ));
 sg13g2_dfrbp_1 _2197_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net102),
    .D(net351),
    .Q_N(_0014_),
    .Q(\ChiselTop.hourDecReg[0] ));
 sg13g2_dfrbp_1 _2198_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net100),
    .D(_0068_),
    .Q_N(_1048_),
    .Q(\ChiselTop.hourDecReg[1] ));
 sg13g2_dfrbp_1 _2199_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net98),
    .D(_0069_),
    .Q_N(_1047_),
    .Q(\ChiselTop.tClk32kHzInReg ));
 sg13g2_dfrbp_1 _2200_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net97),
    .D(_0070_),
    .Q_N(_1046_),
    .Q(\ChiselTop.cntReg[0] ));
 sg13g2_dfrbp_1 _2201_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net95),
    .D(_0071_),
    .Q_N(_1045_),
    .Q(\ChiselTop.cntReg[1] ));
 sg13g2_dfrbp_1 _2202_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net93),
    .D(_0072_),
    .Q_N(_1044_),
    .Q(\ChiselTop.cntReg[2] ));
 sg13g2_dfrbp_1 _2203_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net91),
    .D(_0073_),
    .Q_N(_0004_),
    .Q(\ChiselTop.cntReg[3] ));
 sg13g2_dfrbp_1 _2204_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net89),
    .D(_0074_),
    .Q_N(_1043_),
    .Q(\ChiselTop.cntReg[4] ));
 sg13g2_dfrbp_1 _2205_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net87),
    .D(_0075_),
    .Q_N(_0003_),
    .Q(\ChiselTop.cntReg[5] ));
 sg13g2_dfrbp_1 _2206_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net85),
    .D(_0076_),
    .Q_N(_1042_),
    .Q(\ChiselTop.cntReg[6] ));
 sg13g2_dfrbp_1 _2207_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net83),
    .D(_0077_),
    .Q_N(_1041_),
    .Q(\ChiselTop.cntReg[7] ));
 sg13g2_dfrbp_1 _2208_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net81),
    .D(_0078_),
    .Q_N(_1040_),
    .Q(\ChiselTop.cntReg[8] ));
 sg13g2_dfrbp_1 _2209_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net79),
    .D(_0079_),
    .Q_N(_1039_),
    .Q(\ChiselTop.cntReg[9] ));
 sg13g2_dfrbp_1 _2210_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net77),
    .D(_0080_),
    .Q_N(_1038_),
    .Q(\ChiselTop.cntReg[10] ));
 sg13g2_dfrbp_1 _2211_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net75),
    .D(net222),
    .Q_N(_1037_),
    .Q(\ChiselTop.cntReg[11] ));
 sg13g2_dfrbp_1 _2212_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net73),
    .D(_0082_),
    .Q_N(_1036_),
    .Q(\ChiselTop.cntReg[12] ));
 sg13g2_dfrbp_1 _2213_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net71),
    .D(_0083_),
    .Q_N(_1035_),
    .Q(\ChiselTop.cntReg[13] ));
 sg13g2_dfrbp_1 _2214_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net69),
    .D(_0084_),
    .Q_N(_0008_),
    .Q(\ChiselTop.cntReg[14] ));
 sg13g2_dfrbp_1 _2215_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net67),
    .D(_0085_),
    .Q_N(_0007_),
    .Q(\ChiselTop.cntReg[15] ));
 sg13g2_dfrbp_1 _2216_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net65),
    .D(_0086_),
    .Q_N(_0001_),
    .Q(\ChiselTop.cntReg[16] ));
 sg13g2_dfrbp_1 _2217_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net63),
    .D(_0087_),
    .Q_N(_0006_),
    .Q(\ChiselTop.cntReg[17] ));
 sg13g2_dfrbp_1 _2218_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net61),
    .D(_0088_),
    .Q_N(_1034_),
    .Q(\ChiselTop.cntReg[18] ));
 sg13g2_dfrbp_1 _2219_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net59),
    .D(_0089_),
    .Q_N(_1033_),
    .Q(\ChiselTop.cntReg[19] ));
 sg13g2_dfrbp_1 _2220_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net57),
    .D(_0090_),
    .Q_N(_1032_),
    .Q(\ChiselTop.cntReg[20] ));
 sg13g2_dfrbp_1 _2221_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net55),
    .D(_0091_),
    .Q_N(_1031_),
    .Q(\ChiselTop.cntReg[21] ));
 sg13g2_dfrbp_1 _2222_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net53),
    .D(_0092_),
    .Q_N(_1030_),
    .Q(\ChiselTop.cntReg[22] ));
 sg13g2_dfrbp_1 _2223_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net51),
    .D(_0093_),
    .Q_N(_0005_),
    .Q(\ChiselTop.cntReg[23] ));
 sg13g2_dfrbp_1 _2224_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net49),
    .D(_0094_),
    .Q_N(_1029_),
    .Q(\ChiselTop.cntReg[24] ));
 sg13g2_dfrbp_1 _2225_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net47),
    .D(_0095_),
    .Q_N(_1028_),
    .Q(\ChiselTop.tClk1HzInReg ));
 sg13g2_dfrbp_1 _2226_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net46),
    .D(net208),
    .Q_N(_1027_),
    .Q(\ChiselTop.minusReqReg ));
 sg13g2_dfrbp_1 _2227_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net45),
    .D(_0097_),
    .Q_N(_1026_),
    .Q(\ChiselTop.minusInReg ));
 sg13g2_dfrbp_1 _2228_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net44),
    .D(net196),
    .Q_N(_1025_),
    .Q(\ChiselTop.plusReqReg ));
 sg13g2_dfrbp_1 _2229_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net43),
    .D(_0099_),
    .Q_N(_1024_),
    .Q(\ChiselTop.plusInReg ));
 sg13g2_dfrbp_1 _2230_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net42),
    .D(_0100_),
    .Q_N(_1023_),
    .Q(\ChiselTop.vSyncReg ));
 sg13g2_dfrbp_1 _2231_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net41),
    .D(_0101_),
    .Q_N(\ChiselTop._counterXReg_T_1[0] ),
    .Q(\ChiselTop.counterXReg[0] ));
 sg13g2_dfrbp_1 _2232_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net40),
    .D(net367),
    .Q_N(_1022_),
    .Q(\ChiselTop.counterXReg[1] ));
 sg13g2_dfrbp_1 _2233_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net39),
    .D(_0103_),
    .Q_N(_1021_),
    .Q(\ChiselTop.counterXReg[2] ));
 sg13g2_dfrbp_1 _2234_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net38),
    .D(_0104_),
    .Q_N(_1020_),
    .Q(\ChiselTop.counterXReg[3] ));
 sg13g2_dfrbp_1 _2235_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net36),
    .D(_0105_),
    .Q_N(_0027_),
    .Q(\ChiselTop.counterXReg[4] ));
 sg13g2_dfrbp_1 _2236_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net34),
    .D(_0106_),
    .Q_N(_1019_),
    .Q(\ChiselTop.counterXReg[5] ));
 sg13g2_dfrbp_1 _2237_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net32),
    .D(_0107_),
    .Q_N(_1018_),
    .Q(\ChiselTop.counterXReg[6] ));
 sg13g2_dfrbp_1 _2238_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net30),
    .D(_0108_),
    .Q_N(_1017_),
    .Q(\ChiselTop.counterXReg[7] ));
 sg13g2_dfrbp_1 _2239_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net28),
    .D(_0109_),
    .Q_N(_1016_),
    .Q(\ChiselTop.counterXReg[8] ));
 sg13g2_dfrbp_1 _2240_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net26),
    .D(_0110_),
    .Q_N(_0026_),
    .Q(\ChiselTop.counterXReg[9] ));
 sg13g2_dfrbp_1 _2241_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net24),
    .D(_0111_),
    .Q_N(_1015_),
    .Q(\ChiselTop.counterYReg[0] ));
 sg13g2_dfrbp_1 _2242_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net20),
    .D(_0112_),
    .Q_N(_1014_),
    .Q(\ChiselTop.counterYReg[1] ));
 sg13g2_dfrbp_1 _2243_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net16),
    .D(_0113_),
    .Q_N(_1013_),
    .Q(\ChiselTop.counterYReg[2] ));
 sg13g2_dfrbp_1 _2244_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net12),
    .D(net346),
    .Q_N(_0011_),
    .Q(\ChiselTop.counterYReg[3] ));
 sg13g2_dfrbp_1 _2245_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net150),
    .D(_0115_),
    .Q_N(_1012_),
    .Q(\ChiselTop.counterYReg[4] ));
 sg13g2_dfrbp_1 _2246_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net145),
    .D(net424),
    .Q_N(_0002_),
    .Q(\ChiselTop.counterYReg[5] ));
 sg13g2_dfrbp_1 _2247_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net141),
    .D(_0117_),
    .Q_N(_1011_),
    .Q(\ChiselTop.counterYReg[6] ));
 sg13g2_dfrbp_1 _2248_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net137),
    .D(net384),
    .Q_N(_0012_),
    .Q(\ChiselTop.counterYReg[7] ));
 sg13g2_dfrbp_1 _2249_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net133),
    .D(_0119_),
    .Q_N(_0013_),
    .Q(\ChiselTop.counterYReg[8] ));
 sg13g2_dfrbp_1 _2250_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net129),
    .D(_0120_),
    .Q_N(_1010_),
    .Q(\ChiselTop.counterYReg[9] ));
 sg13g2_dfrbp_1 _2251_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net125),
    .D(_0121_),
    .Q_N(\ChiselTop._debounceCounter_T_1[0] ),
    .Q(\ChiselTop.debounceCounter[0] ));
 sg13g2_dfrbp_1 _2252_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net123),
    .D(net215),
    .Q_N(_1009_),
    .Q(\ChiselTop.debounceCounter[1] ));
 sg13g2_dfrbp_1 _2253_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net121),
    .D(net186),
    .Q_N(_1008_),
    .Q(\ChiselTop.debounceCounter[2] ));
 sg13g2_dfrbp_1 _2254_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net119),
    .D(_0124_),
    .Q_N(_1007_),
    .Q(\ChiselTop.debounceCounter[3] ));
 sg13g2_dfrbp_1 _2255_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net117),
    .D(_0125_),
    .Q_N(_1006_),
    .Q(\ChiselTop.debounceCounter[4] ));
 sg13g2_dfrbp_1 _2256_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net115),
    .D(net298),
    .Q_N(_1005_),
    .Q(\ChiselTop.debounceCounter[5] ));
 sg13g2_dfrbp_1 _2257_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net113),
    .D(net204),
    .Q_N(_1004_),
    .Q(\ChiselTop.debounceCounter[6] ));
 sg13g2_dfrbp_1 _2258_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net111),
    .D(_0128_),
    .Q_N(_1003_),
    .Q(\ChiselTop.debounceCounter[7] ));
 sg13g2_dfrbp_1 _2259_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net109),
    .D(net310),
    .Q_N(_1002_),
    .Q(\ChiselTop.debounceCounter[8] ));
 sg13g2_dfrbp_1 _2260_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net107),
    .D(net212),
    .Q_N(_1001_),
    .Q(\ChiselTop.debounceCounter[9] ));
 sg13g2_dfrbp_1 _2261_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net105),
    .D(net189),
    .Q_N(_1000_),
    .Q(\ChiselTop.debounceCounter[10] ));
 sg13g2_dfrbp_1 _2262_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net103),
    .D(_0132_),
    .Q_N(_0999_),
    .Q(\ChiselTop.debounceCounter[11] ));
 sg13g2_dfrbp_1 _2263_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net101),
    .D(_0133_),
    .Q_N(_0998_),
    .Q(\ChiselTop.debounceCounter[12] ));
 sg13g2_dfrbp_1 _2264_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net99),
    .D(_0134_),
    .Q_N(_0997_),
    .Q(\ChiselTop.debounceCounter[13] ));
 sg13g2_dfrbp_1 _2265_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net96),
    .D(_0135_),
    .Q_N(_0996_),
    .Q(\ChiselTop.debounceCounter[14] ));
 sg13g2_dfrbp_1 _2266_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net94),
    .D(net354),
    .Q_N(_0995_),
    .Q(\ChiselTop.debounceCounter[15] ));
 sg13g2_dfrbp_1 _2267_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net92),
    .D(net210),
    .Q_N(_0994_),
    .Q(\ChiselTop.debounceCounter[16] ));
 sg13g2_dfrbp_1 _2268_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net90),
    .D(net184),
    .Q_N(_0993_),
    .Q(\ChiselTop.debounceCounter[17] ));
 sg13g2_dfrbp_1 _2269_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net88),
    .D(_0139_),
    .Q_N(_0992_),
    .Q(\ChiselTop.debounceCounter[18] ));
 sg13g2_dfrbp_1 _2270_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net86),
    .D(net301),
    .Q_N(_0991_),
    .Q(\ChiselTop.debounceCounter[19] ));
 sg13g2_dfrbp_1 _2271_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net84),
    .D(net328),
    .Q_N(_0990_),
    .Q(\ChiselTop.SetSelIn[0] ));
 sg13g2_dfrbp_1 _2272_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net80),
    .D(net349),
    .Q_N(_0989_),
    .Q(\ChiselTop.SetSelIn[1] ));
 sg13g2_dfrbp_1 _2273_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net76),
    .D(net206),
    .Q_N(_0988_),
    .Q(\ChiselTop.minusIn ));
 sg13g2_dfrbp_1 _2274_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net72),
    .D(net192),
    .Q_N(_0987_),
    .Q(\ChiselTop.plusIn ));
 sg13g2_dfrbp_1 _2275_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net68),
    .D(net319),
    .Q_N(_0986_),
    .Q(\ChiselTop.tClkSelectIn[0] ));
 sg13g2_dfrbp_1 _2276_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net64),
    .D(net316),
    .Q_N(_0985_),
    .Q(\ChiselTop.tClkSelectIn[1] ));
 sg13g2_dfrbp_1 _2277_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net60),
    .D(_0147_),
    .Q_N(_0984_),
    .Q(\ChiselTop.setSelInBounce_pipeReg_1[0] ));
 sg13g2_dfrbp_1 _2278_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net58),
    .D(_0148_),
    .Q_N(_0983_),
    .Q(\ChiselTop.setSelInBounce_pipeReg_1[1] ));
 sg13g2_dfrbp_1 _2279_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net56),
    .D(_0149_),
    .Q_N(_0982_),
    .Q(\ChiselTop.setSelInBounce_pipeReg_0[0] ));
 sg13g2_dfrbp_1 _2280_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net54),
    .D(_0150_),
    .Q_N(_0981_),
    .Q(\ChiselTop.setSelInBounce_pipeReg_0[1] ));
 sg13g2_dfrbp_1 _2281_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net52),
    .D(_0151_),
    .Q_N(_0980_),
    .Q(\ChiselTop.minusInBounce_pipeReg_1 ));
 sg13g2_dfrbp_1 _2282_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net50),
    .D(_0152_),
    .Q_N(_0979_),
    .Q(\ChiselTop.minusInBounce_pipeReg_0 ));
 sg13g2_dfrbp_1 _2283_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net48),
    .D(_0153_),
    .Q_N(_0978_),
    .Q(\ChiselTop.plusInBounce_pipeReg_1 ));
 sg13g2_dfrbp_1 _2284_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net22),
    .D(_0154_),
    .Q_N(_0977_),
    .Q(\ChiselTop.plusInBounce_pipeReg_0 ));
 sg13g2_dfrbp_1 _2285_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net18),
    .D(_0155_),
    .Q_N(_0976_),
    .Q(\ChiselTop.tClk32kHzIn_pipeReg_1 ));
 sg13g2_dfrbp_1 _2286_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net14),
    .D(_0156_),
    .Q_N(_0975_),
    .Q(\ChiselTop.tClk32kHzIn_pipeReg_0 ));
 sg13g2_dfrbp_1 _2287_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net10),
    .D(_0157_),
    .Q_N(_0974_),
    .Q(\ChiselTop.tClk1HzIn_pipeReg_1 ));
 sg13g2_dfrbp_1 _2288_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net148),
    .D(_0158_),
    .Q_N(_0973_),
    .Q(\ChiselTop.tClk1HzIn_pipeReg_0 ));
 sg13g2_dfrbp_1 _2289_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net143),
    .D(_0159_),
    .Q_N(_0972_),
    .Q(\ChiselTop.tClkSelectInBounce_pipeReg_1[0] ));
 sg13g2_dfrbp_1 _2290_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net139),
    .D(_0160_),
    .Q_N(_0971_),
    .Q(\ChiselTop.tClkSelectInBounce_pipeReg_1[1] ));
 sg13g2_dfrbp_1 _2291_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net135),
    .D(_0161_),
    .Q_N(_0970_),
    .Q(\ChiselTop.tClkSelectInBounce_pipeReg_0[0] ));
 sg13g2_dfrbp_1 _2292_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net131),
    .D(_0162_),
    .Q_N(_0969_),
    .Q(\ChiselTop.tClkSelectInBounce_pipeReg_0[1] ));
 sg13g2_dfrbp_1 _2293_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net127),
    .D(_0163_),
    .Q_N(_0968_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _2294_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net151),
    .D(_0164_),
    .Q_N(_1074_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _2295_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net82),
    .D(\ChiselTop.vSync ),
    .Q_N(_0967_),
    .Q(\ChiselTop.vSyncOut_REG ));
 sg13g2_dfrbp_1 _2296_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net78),
    .D(_0165_),
    .Q_N(_0966_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _2297_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net74),
    .D(_0166_),
    .Q_N(_0965_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _2298_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net70),
    .D(_0167_),
    .Q_N(_0964_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _2299_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net62),
    .D(_0168_),
    .Q_N(_1075_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _2300_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net66),
    .D(net428),
    .Q_N(_0963_),
    .Q(\ChiselTop.hSyncOut_REG ));
 sg13g2_tiehi _2287__10 (.L_HI(net10));
 sg13g2_tiehi _2172__11 (.L_HI(net11));
 sg13g2_tiehi _2244__12 (.L_HI(net12));
 sg13g2_tiehi _2171__13 (.L_HI(net13));
 sg13g2_tiehi _2286__14 (.L_HI(net14));
 sg13g2_tiehi _2170__15 (.L_HI(net15));
 sg13g2_tiehi _2243__16 (.L_HI(net16));
 sg13g2_tiehi _2169__17 (.L_HI(net17));
 sg13g2_tiehi _2285__18 (.L_HI(net18));
 sg13g2_tiehi _2168__19 (.L_HI(net19));
 sg13g2_tiehi _2242__20 (.L_HI(net20));
 sg13g2_tiehi _2167__21 (.L_HI(net21));
 sg13g2_tiehi _2284__22 (.L_HI(net22));
 sg13g2_tiehi _2166__23 (.L_HI(net23));
 sg13g2_tiehi _2241__24 (.L_HI(net24));
 sg13g2_tiehi _2165__25 (.L_HI(net25));
 sg13g2_tiehi _2240__26 (.L_HI(net26));
 sg13g2_tiehi _2164__27 (.L_HI(net27));
 sg13g2_tiehi _2239__28 (.L_HI(net28));
 sg13g2_tiehi _2163__29 (.L_HI(net29));
 sg13g2_tiehi _2238__30 (.L_HI(net30));
 sg13g2_tiehi _2162__31 (.L_HI(net31));
 sg13g2_tiehi _2237__32 (.L_HI(net32));
 sg13g2_tiehi _2161__33 (.L_HI(net33));
 sg13g2_tiehi _2236__34 (.L_HI(net34));
 sg13g2_tiehi _2160__35 (.L_HI(net35));
 sg13g2_tiehi _2235__36 (.L_HI(net36));
 sg13g2_tiehi _2159__37 (.L_HI(net37));
 sg13g2_tiehi _2234__38 (.L_HI(net38));
 sg13g2_tiehi _2233__39 (.L_HI(net39));
 sg13g2_tiehi _2232__40 (.L_HI(net40));
 sg13g2_tiehi _2231__41 (.L_HI(net41));
 sg13g2_tiehi _2230__42 (.L_HI(net42));
 sg13g2_tiehi _2229__43 (.L_HI(net43));
 sg13g2_tiehi _2228__44 (.L_HI(net44));
 sg13g2_tiehi _2227__45 (.L_HI(net45));
 sg13g2_tiehi _2226__46 (.L_HI(net46));
 sg13g2_tiehi _2225__47 (.L_HI(net47));
 sg13g2_tiehi _2283__48 (.L_HI(net48));
 sg13g2_tiehi _2224__49 (.L_HI(net49));
 sg13g2_tiehi _2282__50 (.L_HI(net50));
 sg13g2_tiehi _2223__51 (.L_HI(net51));
 sg13g2_tiehi _2281__52 (.L_HI(net52));
 sg13g2_tiehi _2222__53 (.L_HI(net53));
 sg13g2_tiehi _2280__54 (.L_HI(net54));
 sg13g2_tiehi _2221__55 (.L_HI(net55));
 sg13g2_tiehi _2279__56 (.L_HI(net56));
 sg13g2_tiehi _2220__57 (.L_HI(net57));
 sg13g2_tiehi _2278__58 (.L_HI(net58));
 sg13g2_tiehi _2219__59 (.L_HI(net59));
 sg13g2_tiehi _2277__60 (.L_HI(net60));
 sg13g2_tiehi _2218__61 (.L_HI(net61));
 sg13g2_tiehi _2299__62 (.L_HI(net62));
 sg13g2_tiehi _2217__63 (.L_HI(net63));
 sg13g2_tiehi _2276__64 (.L_HI(net64));
 sg13g2_tiehi _2216__65 (.L_HI(net65));
 sg13g2_tiehi _2300__66 (.L_HI(net66));
 sg13g2_tiehi _2215__67 (.L_HI(net67));
 sg13g2_tiehi _2275__68 (.L_HI(net68));
 sg13g2_tiehi _2214__69 (.L_HI(net69));
 sg13g2_tiehi _2298__70 (.L_HI(net70));
 sg13g2_tiehi _2213__71 (.L_HI(net71));
 sg13g2_tiehi _2274__72 (.L_HI(net72));
 sg13g2_tiehi _2212__73 (.L_HI(net73));
 sg13g2_tiehi _2297__74 (.L_HI(net74));
 sg13g2_tiehi _2211__75 (.L_HI(net75));
 sg13g2_tiehi _2273__76 (.L_HI(net76));
 sg13g2_tiehi _2210__77 (.L_HI(net77));
 sg13g2_tiehi _2296__78 (.L_HI(net78));
 sg13g2_tiehi _2209__79 (.L_HI(net79));
 sg13g2_tiehi _2272__80 (.L_HI(net80));
 sg13g2_tiehi _2208__81 (.L_HI(net81));
 sg13g2_tiehi _2295__82 (.L_HI(net82));
 sg13g2_tiehi _2207__83 (.L_HI(net83));
 sg13g2_tiehi _2271__84 (.L_HI(net84));
 sg13g2_tiehi _2206__85 (.L_HI(net85));
 sg13g2_tiehi _2270__86 (.L_HI(net86));
 sg13g2_tiehi _2205__87 (.L_HI(net87));
 sg13g2_tiehi _2269__88 (.L_HI(net88));
 sg13g2_tiehi _2204__89 (.L_HI(net89));
 sg13g2_tiehi _2268__90 (.L_HI(net90));
 sg13g2_tiehi _2203__91 (.L_HI(net91));
 sg13g2_tiehi _2267__92 (.L_HI(net92));
 sg13g2_tiehi _2202__93 (.L_HI(net93));
 sg13g2_tiehi _2266__94 (.L_HI(net94));
 sg13g2_tiehi _2201__95 (.L_HI(net95));
 sg13g2_tiehi _2265__96 (.L_HI(net96));
 sg13g2_tiehi _2200__97 (.L_HI(net97));
 sg13g2_tiehi _2199__98 (.L_HI(net98));
 sg13g2_tiehi _2264__99 (.L_HI(net99));
 sg13g2_tiehi _2198__100 (.L_HI(net100));
 sg13g2_tiehi _2263__101 (.L_HI(net101));
 sg13g2_tiehi _2197__102 (.L_HI(net102));
 sg13g2_tiehi _2262__103 (.L_HI(net103));
 sg13g2_tiehi _2196__104 (.L_HI(net104));
 sg13g2_tiehi _2261__105 (.L_HI(net105));
 sg13g2_tiehi _2195__106 (.L_HI(net106));
 sg13g2_tiehi _2260__107 (.L_HI(net107));
 sg13g2_tiehi _2194__108 (.L_HI(net108));
 sg13g2_tiehi _2259__109 (.L_HI(net109));
 sg13g2_tiehi _2193__110 (.L_HI(net110));
 sg13g2_tiehi _2258__111 (.L_HI(net111));
 sg13g2_tiehi _2192__112 (.L_HI(net112));
 sg13g2_tiehi _2257__113 (.L_HI(net113));
 sg13g2_tiehi _2191__114 (.L_HI(net114));
 sg13g2_tiehi _2256__115 (.L_HI(net115));
 sg13g2_tiehi _2190__116 (.L_HI(net116));
 sg13g2_tiehi _2255__117 (.L_HI(net117));
 sg13g2_tiehi _2189__118 (.L_HI(net118));
 sg13g2_tiehi _2254__119 (.L_HI(net119));
 sg13g2_tiehi _2188__120 (.L_HI(net120));
 sg13g2_tiehi _2253__121 (.L_HI(net121));
 sg13g2_tiehi _2187__122 (.L_HI(net122));
 sg13g2_tiehi _2252__123 (.L_HI(net123));
 sg13g2_tiehi _2186__124 (.L_HI(net124));
 sg13g2_tiehi _2251__125 (.L_HI(net125));
 sg13g2_tiehi _2185__126 (.L_HI(net126));
 sg13g2_tiehi _2293__127 (.L_HI(net127));
 sg13g2_tiehi _2184__128 (.L_HI(net128));
 sg13g2_tiehi _2250__129 (.L_HI(net129));
 sg13g2_tiehi _2183__130 (.L_HI(net130));
 sg13g2_tiehi _2292__131 (.L_HI(net131));
 sg13g2_tiehi _2182__132 (.L_HI(net132));
 sg13g2_tiehi _2249__133 (.L_HI(net133));
 sg13g2_tiehi _2181__134 (.L_HI(net134));
 sg13g2_tiehi _2291__135 (.L_HI(net135));
 sg13g2_tiehi _2180__136 (.L_HI(net136));
 sg13g2_tiehi _2248__137 (.L_HI(net137));
 sg13g2_tiehi _2179__138 (.L_HI(net138));
 sg13g2_tiehi _2290__139 (.L_HI(net139));
 sg13g2_tiehi _2178__140 (.L_HI(net140));
 sg13g2_tiehi _2247__141 (.L_HI(net141));
 sg13g2_tiehi _2177__142 (.L_HI(net142));
 sg13g2_tiehi _2289__143 (.L_HI(net143));
 sg13g2_tiehi _2176__144 (.L_HI(net144));
 sg13g2_tiehi _2246__145 (.L_HI(net145));
 sg13g2_tiehi _2158__146 (.L_HI(net146));
 sg13g2_tiehi _2175__147 (.L_HI(net147));
 sg13g2_tiehi _2288__148 (.L_HI(net148));
 sg13g2_tiehi _2174__149 (.L_HI(net149));
 sg13g2_tiehi _2245__150 (.L_HI(net150));
 sg13g2_tiehi _2294__151 (.L_HI(net151));
 sg13g2_tiehi tt_um_luke_clock_152 (.L_HI(net152));
 sg13g2_tiehi tt_um_luke_clock_153 (.L_HI(net153));
 sg13g2_tiehi tt_um_luke_clock_154 (.L_HI(net154));
 sg13g2_tiehi tt_um_luke_clock_155 (.L_HI(net155));
 sg13g2_tiehi tt_um_luke_clock_156 (.L_HI(net156));
 sg13g2_tiehi tt_um_luke_clock_157 (.L_HI(net157));
 sg13g2_tiehi tt_um_luke_clock_158 (.L_HI(net158));
 sg13g2_tiehi tt_um_luke_clock_159 (.L_HI(net159));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 _2452_ (.A(\ChiselTop.tClk ),
    .X(uio_out[0]));
 sg13g2_buf_1 _2453_ (.A(\ChiselTop.cntReg[0] ),
    .X(uio_out[1]));
 sg13g2_buf_1 _2454_ (.A(\ChiselTop.cntReg[1] ),
    .X(uio_out[2]));
 sg13g2_buf_1 _2455_ (.A(\ChiselTop.cntReg[2] ),
    .X(uio_out[3]));
 sg13g2_buf_1 _2456_ (.A(\ChiselTop.cntReg[3] ),
    .X(uio_out[4]));
 sg13g2_buf_1 _2457_ (.A(\ChiselTop.inDisplayArea ),
    .X(uio_out[5]));
 sg13g2_buf_1 _2458_ (.A(\ChiselTop.vSyncOut_REG ),
    .X(uo_out[3]));
 sg13g2_buf_1 _2459_ (.A(\ChiselTop.hSyncOut_REG ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout224 (.A(_0796_),
    .X(net224));
 sg13g2_buf_4 fanout225 (.X(net225),
    .A(_0791_));
 sg13g2_buf_2 fanout226 (.A(_0738_),
    .X(net226));
 sg13g2_buf_1 fanout227 (.A(_0738_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(net234),
    .X(net228));
 sg13g2_buf_1 fanout229 (.A(net234),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(net231),
    .X(net230));
 sg13g2_buf_1 fanout231 (.A(net234),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(net234),
    .X(net232));
 sg13g2_buf_1 fanout233 (.A(net234),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_0619_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_0232_),
    .X(net235));
 sg13g2_buf_1 fanout236 (.A(_0232_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(net239),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_0786_),
    .X(net238));
 sg13g2_buf_1 fanout239 (.A(_0786_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net241),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_0685_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_0928_),
    .X(net242));
 sg13g2_buf_1 fanout243 (.A(_0928_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(net246),
    .X(net244));
 sg13g2_buf_1 fanout245 (.A(net246),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_0483_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_0482_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_0481_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(net250),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_0927_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_0477_),
    .X(net251));
 sg13g2_buf_4 fanout252 (.X(net252),
    .A(_0855_));
 sg13g2_buf_1 fanout253 (.A(_0855_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_0013_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(net257),
    .X(net255));
 sg13g2_buf_1 fanout256 (.A(net257),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(net391),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(net259),
    .X(net258));
 sg13g2_buf_1 fanout259 (.A(\ChiselTop.counterYReg[7] ),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(\ChiselTop.counterYReg[6] ),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(\ChiselTop.counterYReg[5] ),
    .X(net261));
 sg13g2_buf_1 fanout262 (.A(net263),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(net423),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(net265),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(net426),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(\ChiselTop.counterYReg[3] ),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(\ChiselTop.counterYReg[3] ),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(net435),
    .X(net268));
 sg13g2_buf_1 fanout269 (.A(\ChiselTop.counterYReg[2] ),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(net436),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(net448),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(net440),
    .X(net272));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(net274));
 sg13g2_buf_2 fanout274 (.A(net427),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(net442),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(net277),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(\ChiselTop.counterXReg[5] ),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(net439),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(\ChiselTop.counterXReg[4] ),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(net444),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(\ChiselTop.counterXReg[2] ),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(net390),
    .X(net282));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(net286));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(net286));
 sg13g2_buf_2 fanout285 (.A(net286),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_0442_),
    .X(net286));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(net291));
 sg13g2_buf_2 fanout288 (.A(net290),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(net290),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(net291),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(rst_n),
    .X(net291));
 sg13g2_buf_4 fanout292 (.X(net292),
    .A(net293));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(net297));
 sg13g2_buf_2 fanout294 (.A(net295),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(net296),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(net297),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(rst_n),
    .X(net297));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tiehi _2173__9 (.L_HI(net9));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_29__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\ChiselTop._counterXReg_T_1[0] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold2 (.A(\ChiselTop._debounceCounter_T_1[0] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold3 (.A(\ChiselTop._modeReg_T_1[0] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0029_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold5 (.A(\ChiselTop.tClkSelectInBounce_pipeReg_1[1] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold6 (.A(\ChiselTop.tClkSelectInBounce_pipeReg_1[0] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold7 (.A(\ChiselTop.setSelInBounce_pipeReg_1[1] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold8 (.A(\ChiselTop.tClk1HzIn_pipeReg_1 ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold9 (.A(\ChiselTop.tClk32kHzIn_pipeReg_1 ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold10 (.A(\ChiselTop.secondUniReg[2] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0051_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold12 (.A(\ChiselTop.minusInBounce_pipeReg_1 ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold13 (.A(\ChiselTop.plusInBounce_pipeReg_1 ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold14 (.A(\ChiselTop.setSelInBounce_pipeReg_1[0] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold15 (.A(\ChiselTop.minusIn ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold16 (.A(\ChiselTop.plusIn ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold17 (.A(\ChiselTop.tClk1HzIn_pipeReg_0 ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold18 (.A(\ChiselTop.debounceCounter[3] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0932_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold20 (.A(\ChiselTop.minuteDecReg[2] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0062_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold22 (.A(\ChiselTop.tClk32kHzIn_pipeReg_0 ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold23 (.A(\ChiselTop.debounceCounter[17] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0957_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0138_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold26 (.A(\ChiselTop.debounceCounter[2] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0123_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold28 (.A(\ChiselTop.debounceCounter[10] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0944_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0131_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold31 (.A(\ChiselTop.tClkReqReg ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold32 (.A(\ChiselTop.plusInBounce_pipeReg_0 ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0144_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold34 (.A(\ChiselTop.cntReg[22] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0843_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold36 (.A(\ChiselTop.plusReqReg ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0098_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold38 (.A(\ChiselTop.cntReg[2] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0798_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0022_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0666_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0053_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold43 (.A(\ChiselTop.debounceCounter[6] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0937_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0127_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold46 (.A(\ChiselTop.minusInBounce_pipeReg_0 ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0143_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold48 (.A(\ChiselTop.minusReqReg ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0096_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold50 (.A(\ChiselTop.debounceCounter[16] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0137_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold52 (.A(\ChiselTop.debounceCounter[9] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0130_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold54 (.A(\ChiselTop.debounceCounter[1] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0930_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0122_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold57 (.A(\ChiselTop.cntReg[5] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0805_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold59 (.A(\ChiselTop.secondDecReg[2] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0055_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold61 (.A(\ChiselTop.cntReg[11] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0817_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0081_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold64 (.A(\ChiselTop.debounceCounter[5] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0126_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold66 (.A(\ChiselTop.debounceCounter[19] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0961_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0140_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0023_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0650_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold71 (.A(\ChiselTop.cntReg[4] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0802_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold73 (.A(\ChiselTop.cntReg[13] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0821_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold75 (.A(\ChiselTop.debounceCounter[8] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0941_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0129_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold78 (.A(\ChiselTop.debounceCounter[18] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0959_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold80 (.A(\ChiselTop.debounceCounter[12] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0948_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold82 (.A(\ChiselTop.tClkSelectIn[1] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0146_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold84 (.A(\ChiselTop.counterYReg[9] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold85 (.A(\ChiselTop.tClkSelectInBounce_pipeReg_0[0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0145_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold87 (.A(\ChiselTop.minuteDecReg[0] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0060_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold89 (.A(\ChiselTop.minuteDecReg[1] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold90 (.A(\ChiselTop.cntReg[18] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0836_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold92 (.A(\ChiselTop.cntReg[17] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0832_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold94 (.A(\ChiselTop.setSelInBounce_pipeReg_0[0] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0141_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold96 (.A(\ChiselTop.debounceCounter[7] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0939_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold98 (.A(\ChiselTop.secondUniReg[3] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0662_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0052_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold101 (.A(\ChiselTop.cntReg[12] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0819_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold103 (.A(\ChiselTop.cntReg[16] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0830_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold105 (.A(\ChiselTop.debounceCounter[11] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold106 (.A(\ChiselTop.debounceCounter[14] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0952_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold108 (.A(\ChiselTop.cntReg[20] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0840_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold110 (.A(\ChiselTop.cntReg[14] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0824_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0011_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0114_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold114 (.A(\ChiselTop.cntReg[19] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold115 (.A(\ChiselTop.setSelInBounce_pipeReg_0[1] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0142_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold117 (.A(\ChiselTop.hourDecReg[0] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0067_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold119 (.A(\ChiselTop.cntReg[21] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold120 (.A(\ChiselTop.debounceCounter[15] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0136_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0007_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0825_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0826_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0027_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0871_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0004_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0800_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0801_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold130 (.A(\ChiselTop.cntReg[9] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold131 (.A(\ChiselTop.hourDecReg[1] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold132 (.A(\ChiselTop.counterXReg[1] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0864_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0102_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold135 (.A(\ChiselTop.cntReg[6] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold136 (.A(\ChiselTop.minuteUniReg[2] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0058_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold138 (.A(\ChiselTop.cntReg[23] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0847_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold140 (.A(\ChiselTop.debounceCounter[13] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold141 (.A(\ChiselTop.cntReg[1] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0797_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold143 (.A(\ChiselTop.cntReg[10] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold144 (.A(\ChiselTop.minuteUniReg[1] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold145 (.A(uio_out[7]),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0030_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold147 (.A(\ChiselTop.secondUniReg[1] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0050_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold149 (.A(\ChiselTop.cntReg[7] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0012_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0118_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold152 (.A(\ChiselTop.minuteUniReg[0] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0056_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold154 (.A(\ChiselTop.hourUniReg[2] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0065_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold156 (.A(\ChiselTop.cntReg[0] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold157 (.A(\ChiselTop.counterXReg[2] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold158 (.A(\ChiselTop.counterYReg[8] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold159 (.A(\ChiselTop.hourUniReg[0] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0063_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold161 (.A(\ChiselTop.hourUniReg[3] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0066_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold163 (.A(\ChiselTop.counterYReg[0] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold164 (.A(\ChiselTop.cntReg[8] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold165 (.A(\ChiselTop.minuteUniReg[3] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0059_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold167 (.A(\ChiselTop.lfsrReg_11 ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0037_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold169 (.A(\ChiselTop.lfsrReg_2 ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0046_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold171 (.A(\ChiselTop.lfsrReg_5 ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0043_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold173 (.A(\ChiselTop.lfsrReg_8 ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0040_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold175 (.A(\ChiselTop.lfsrReg_17 ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0396_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold177 (.A(\ChiselTop.lfsrReg_4 ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0044_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold179 (.A(\ChiselTop.lfsrReg_12 ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold180 (.A(\ChiselTop.secondDecReg[1] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0054_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold182 (.A(\ChiselTop.lfsrReg_9 ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold183 (.A(\ChiselTop.lfsrReg_13 ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold184 (.A(\ChiselTop.lfsrReg_14 ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold185 (.A(\ChiselTop.lfsrReg_7 ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0041_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold187 (.A(\ChiselTop.lfsrReg_16 ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0032_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold189 (.A(\ChiselTop.lfsrReg_15 ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold190 (.A(\ChiselTop.counterYReg[5] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0116_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold192 (.A(\ChiselTop.counterYReg[9] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold193 (.A(\ChiselTop.counterYReg[4] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold194 (.A(\ChiselTop.counterXReg[7] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0000_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold196 (.A(\ChiselTop.lfsrReg_3 ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold197 (.A(\ChiselTop.lfsrReg_10 ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold198 (.A(\ChiselTop.debounceCounter[4] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0935_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold200 (.A(\ChiselTop.cntReg[24] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold201 (.A(\ChiselTop.lfsrReg_6 ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold202 (.A(\ChiselTop.counterYReg[2] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold203 (.A(\ChiselTop.counterYReg[1] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold204 (.A(\ChiselTop.lfsrReg_0 ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0047_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold206 (.A(\ChiselTop.counterXReg[4] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold207 (.A(\ChiselTop.counterXReg[8] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold208 (.A(\ChiselTop.hourUniReg[1] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold209 (.A(\ChiselTop.counterXReg[6] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0874_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold211 (.A(\ChiselTop.counterXReg[3] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold212 (.A(\ChiselTop.lfsrReg_1 ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0386_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0002_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold215 (.A(\ChiselTop.counterXReg[9] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold216 (.A(\ChiselTop.cntReg[6] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0499_),
    .X(net450));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_4 FILLER_1_364 ();
 sg13g2_decap_4 FILLER_1_372 ();
 sg13g2_fill_2 FILLER_1_376 ();
 sg13g2_decap_8 FILLER_1_382 ();
 sg13g2_decap_8 FILLER_1_389 ();
 sg13g2_decap_8 FILLER_1_396 ();
 sg13g2_decap_4 FILLER_1_403 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_fill_1 FILLER_2_357 ();
 sg13g2_fill_2 FILLER_2_362 ();
 sg13g2_fill_1 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_397 ();
 sg13g2_decap_4 FILLER_2_404 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_fill_2 FILLER_3_336 ();
 sg13g2_fill_1 FILLER_3_338 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_fill_1 FILLER_3_368 ();
 sg13g2_fill_2 FILLER_3_388 ();
 sg13g2_fill_1 FILLER_3_390 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_fill_1 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_121 ();
 sg13g2_decap_8 FILLER_4_128 ();
 sg13g2_fill_1 FILLER_4_135 ();
 sg13g2_fill_2 FILLER_4_140 ();
 sg13g2_fill_1 FILLER_4_142 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_fill_2 FILLER_4_322 ();
 sg13g2_fill_2 FILLER_4_347 ();
 sg13g2_fill_2 FILLER_4_375 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_fill_2 FILLER_5_84 ();
 sg13g2_fill_1 FILLER_5_86 ();
 sg13g2_fill_1 FILLER_5_122 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_fill_1 FILLER_5_308 ();
 sg13g2_fill_2 FILLER_5_313 ();
 sg13g2_fill_1 FILLER_5_315 ();
 sg13g2_fill_1 FILLER_5_352 ();
 sg13g2_fill_2 FILLER_5_362 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_fill_2 FILLER_6_90 ();
 sg13g2_fill_1 FILLER_6_92 ();
 sg13g2_fill_1 FILLER_6_106 ();
 sg13g2_fill_2 FILLER_6_139 ();
 sg13g2_fill_2 FILLER_6_172 ();
 sg13g2_fill_1 FILLER_6_174 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_4 FILLER_6_294 ();
 sg13g2_fill_1 FILLER_6_351 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_fill_2 FILLER_7_42 ();
 sg13g2_fill_1 FILLER_7_44 ();
 sg13g2_decap_4 FILLER_7_54 ();
 sg13g2_fill_1 FILLER_7_58 ();
 sg13g2_fill_2 FILLER_7_64 ();
 sg13g2_fill_1 FILLER_7_66 ();
 sg13g2_decap_4 FILLER_7_71 ();
 sg13g2_fill_2 FILLER_7_75 ();
 sg13g2_fill_2 FILLER_7_108 ();
 sg13g2_fill_1 FILLER_7_110 ();
 sg13g2_decap_8 FILLER_7_132 ();
 sg13g2_fill_2 FILLER_7_139 ();
 sg13g2_fill_1 FILLER_7_141 ();
 sg13g2_fill_2 FILLER_7_152 ();
 sg13g2_decap_4 FILLER_7_176 ();
 sg13g2_fill_1 FILLER_7_180 ();
 sg13g2_fill_2 FILLER_7_191 ();
 sg13g2_decap_8 FILLER_7_202 ();
 sg13g2_decap_8 FILLER_7_209 ();
 sg13g2_decap_8 FILLER_7_216 ();
 sg13g2_decap_8 FILLER_7_223 ();
 sg13g2_decap_8 FILLER_7_230 ();
 sg13g2_decap_8 FILLER_7_237 ();
 sg13g2_decap_8 FILLER_7_244 ();
 sg13g2_decap_8 FILLER_7_251 ();
 sg13g2_decap_8 FILLER_7_258 ();
 sg13g2_decap_8 FILLER_7_265 ();
 sg13g2_decap_8 FILLER_7_272 ();
 sg13g2_decap_8 FILLER_7_279 ();
 sg13g2_decap_8 FILLER_7_286 ();
 sg13g2_decap_8 FILLER_7_293 ();
 sg13g2_decap_4 FILLER_7_300 ();
 sg13g2_fill_1 FILLER_7_335 ();
 sg13g2_fill_1 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_fill_2 FILLER_8_28 ();
 sg13g2_decap_4 FILLER_8_95 ();
 sg13g2_fill_2 FILLER_8_107 ();
 sg13g2_fill_1 FILLER_8_109 ();
 sg13g2_fill_2 FILLER_8_119 ();
 sg13g2_fill_1 FILLER_8_121 ();
 sg13g2_decap_4 FILLER_8_160 ();
 sg13g2_fill_2 FILLER_8_169 ();
 sg13g2_decap_8 FILLER_8_211 ();
 sg13g2_decap_8 FILLER_8_218 ();
 sg13g2_decap_8 FILLER_8_225 ();
 sg13g2_decap_8 FILLER_8_232 ();
 sg13g2_decap_8 FILLER_8_239 ();
 sg13g2_decap_8 FILLER_8_246 ();
 sg13g2_decap_8 FILLER_8_253 ();
 sg13g2_decap_8 FILLER_8_260 ();
 sg13g2_decap_8 FILLER_8_267 ();
 sg13g2_decap_8 FILLER_8_274 ();
 sg13g2_decap_8 FILLER_8_281 ();
 sg13g2_decap_8 FILLER_8_288 ();
 sg13g2_decap_4 FILLER_8_295 ();
 sg13g2_fill_1 FILLER_8_299 ();
 sg13g2_fill_2 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_fill_2 FILLER_9_35 ();
 sg13g2_fill_1 FILLER_9_37 ();
 sg13g2_fill_2 FILLER_9_47 ();
 sg13g2_fill_1 FILLER_9_58 ();
 sg13g2_fill_2 FILLER_9_93 ();
 sg13g2_decap_4 FILLER_9_122 ();
 sg13g2_fill_2 FILLER_9_133 ();
 sg13g2_fill_1 FILLER_9_135 ();
 sg13g2_decap_4 FILLER_9_141 ();
 sg13g2_fill_2 FILLER_9_161 ();
 sg13g2_fill_1 FILLER_9_163 ();
 sg13g2_fill_2 FILLER_9_173 ();
 sg13g2_fill_2 FILLER_9_180 ();
 sg13g2_fill_1 FILLER_9_182 ();
 sg13g2_decap_4 FILLER_9_190 ();
 sg13g2_decap_8 FILLER_9_202 ();
 sg13g2_decap_8 FILLER_9_209 ();
 sg13g2_decap_8 FILLER_9_216 ();
 sg13g2_decap_8 FILLER_9_223 ();
 sg13g2_fill_2 FILLER_9_230 ();
 sg13g2_fill_1 FILLER_9_232 ();
 sg13g2_decap_8 FILLER_9_241 ();
 sg13g2_decap_4 FILLER_9_252 ();
 sg13g2_fill_2 FILLER_9_256 ();
 sg13g2_decap_8 FILLER_9_289 ();
 sg13g2_decap_4 FILLER_9_296 ();
 sg13g2_fill_2 FILLER_9_326 ();
 sg13g2_fill_2 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_4 FILLER_10_21 ();
 sg13g2_fill_2 FILLER_10_51 ();
 sg13g2_fill_1 FILLER_10_59 ();
 sg13g2_fill_1 FILLER_10_98 ();
 sg13g2_fill_2 FILLER_10_108 ();
 sg13g2_fill_1 FILLER_10_110 ();
 sg13g2_fill_1 FILLER_10_172 ();
 sg13g2_decap_4 FILLER_10_184 ();
 sg13g2_decap_8 FILLER_10_208 ();
 sg13g2_fill_1 FILLER_10_215 ();
 sg13g2_fill_2 FILLER_10_261 ();
 sg13g2_fill_1 FILLER_10_272 ();
 sg13g2_fill_1 FILLER_10_291 ();
 sg13g2_fill_2 FILLER_10_345 ();
 sg13g2_fill_1 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_fill_1 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_40 ();
 sg13g2_decap_4 FILLER_11_47 ();
 sg13g2_decap_8 FILLER_11_61 ();
 sg13g2_fill_2 FILLER_11_68 ();
 sg13g2_fill_2 FILLER_11_116 ();
 sg13g2_fill_1 FILLER_11_118 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_fill_2 FILLER_11_140 ();
 sg13g2_fill_1 FILLER_11_142 ();
 sg13g2_decap_4 FILLER_11_166 ();
 sg13g2_fill_1 FILLER_11_184 ();
 sg13g2_fill_2 FILLER_11_213 ();
 sg13g2_fill_1 FILLER_11_234 ();
 sg13g2_fill_2 FILLER_11_251 ();
 sg13g2_fill_1 FILLER_11_253 ();
 sg13g2_fill_2 FILLER_11_261 ();
 sg13g2_decap_4 FILLER_11_293 ();
 sg13g2_fill_2 FILLER_11_297 ();
 sg13g2_fill_1 FILLER_11_307 ();
 sg13g2_fill_2 FILLER_11_336 ();
 sg13g2_fill_1 FILLER_11_338 ();
 sg13g2_fill_1 FILLER_11_351 ();
 sg13g2_fill_1 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_4 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_25 ();
 sg13g2_fill_2 FILLER_12_52 ();
 sg13g2_fill_1 FILLER_12_54 ();
 sg13g2_fill_1 FILLER_12_75 ();
 sg13g2_fill_2 FILLER_12_92 ();
 sg13g2_fill_1 FILLER_12_94 ();
 sg13g2_fill_2 FILLER_12_116 ();
 sg13g2_decap_4 FILLER_12_123 ();
 sg13g2_fill_2 FILLER_12_127 ();
 sg13g2_fill_1 FILLER_12_152 ();
 sg13g2_decap_4 FILLER_12_162 ();
 sg13g2_fill_1 FILLER_12_166 ();
 sg13g2_decap_4 FILLER_12_186 ();
 sg13g2_fill_2 FILLER_12_190 ();
 sg13g2_decap_4 FILLER_12_208 ();
 sg13g2_fill_1 FILLER_12_212 ();
 sg13g2_fill_1 FILLER_12_217 ();
 sg13g2_fill_1 FILLER_12_264 ();
 sg13g2_fill_2 FILLER_12_280 ();
 sg13g2_fill_2 FILLER_12_291 ();
 sg13g2_decap_4 FILLER_12_302 ();
 sg13g2_fill_1 FILLER_12_306 ();
 sg13g2_fill_2 FILLER_12_311 ();
 sg13g2_fill_1 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_fill_2 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_30 ();
 sg13g2_fill_2 FILLER_13_39 ();
 sg13g2_fill_1 FILLER_13_41 ();
 sg13g2_fill_2 FILLER_13_47 ();
 sg13g2_fill_1 FILLER_13_57 ();
 sg13g2_fill_2 FILLER_13_97 ();
 sg13g2_fill_1 FILLER_13_99 ();
 sg13g2_fill_2 FILLER_13_105 ();
 sg13g2_fill_1 FILLER_13_107 ();
 sg13g2_fill_1 FILLER_13_127 ();
 sg13g2_fill_2 FILLER_13_146 ();
 sg13g2_decap_8 FILLER_13_173 ();
 sg13g2_fill_1 FILLER_13_191 ();
 sg13g2_decap_4 FILLER_13_207 ();
 sg13g2_fill_2 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_248 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_7 ();
 sg13g2_fill_1 FILLER_14_9 ();
 sg13g2_decap_4 FILLER_14_18 ();
 sg13g2_fill_2 FILLER_14_22 ();
 sg13g2_fill_1 FILLER_14_64 ();
 sg13g2_fill_2 FILLER_14_70 ();
 sg13g2_fill_1 FILLER_14_72 ();
 sg13g2_decap_4 FILLER_14_104 ();
 sg13g2_fill_1 FILLER_14_117 ();
 sg13g2_fill_2 FILLER_14_128 ();
 sg13g2_fill_2 FILLER_14_138 ();
 sg13g2_fill_1 FILLER_14_140 ();
 sg13g2_fill_2 FILLER_14_150 ();
 sg13g2_fill_2 FILLER_14_159 ();
 sg13g2_fill_2 FILLER_14_173 ();
 sg13g2_fill_1 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_decap_8 FILLER_14_213 ();
 sg13g2_fill_2 FILLER_14_220 ();
 sg13g2_fill_1 FILLER_14_226 ();
 sg13g2_fill_1 FILLER_14_236 ();
 sg13g2_fill_2 FILLER_14_264 ();
 sg13g2_fill_1 FILLER_14_266 ();
 sg13g2_fill_2 FILLER_14_272 ();
 sg13g2_fill_2 FILLER_14_280 ();
 sg13g2_fill_1 FILLER_14_282 ();
 sg13g2_fill_2 FILLER_14_303 ();
 sg13g2_fill_2 FILLER_14_357 ();
 sg13g2_fill_1 FILLER_14_359 ();
 sg13g2_fill_2 FILLER_14_374 ();
 sg13g2_fill_1 FILLER_14_382 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_2 ();
 sg13g2_decap_8 FILLER_15_38 ();
 sg13g2_fill_2 FILLER_15_45 ();
 sg13g2_fill_1 FILLER_15_47 ();
 sg13g2_fill_2 FILLER_15_92 ();
 sg13g2_fill_2 FILLER_15_107 ();
 sg13g2_fill_2 FILLER_15_133 ();
 sg13g2_fill_1 FILLER_15_135 ();
 sg13g2_decap_4 FILLER_15_141 ();
 sg13g2_fill_1 FILLER_15_155 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_fill_2 FILLER_15_175 ();
 sg13g2_fill_1 FILLER_15_177 ();
 sg13g2_fill_2 FILLER_15_192 ();
 sg13g2_fill_1 FILLER_15_194 ();
 sg13g2_fill_2 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_303 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_22 ();
 sg13g2_decap_4 FILLER_16_29 ();
 sg13g2_fill_2 FILLER_16_56 ();
 sg13g2_fill_1 FILLER_16_58 ();
 sg13g2_fill_2 FILLER_16_68 ();
 sg13g2_fill_1 FILLER_16_123 ();
 sg13g2_decap_8 FILLER_16_129 ();
 sg13g2_decap_8 FILLER_16_136 ();
 sg13g2_decap_8 FILLER_16_148 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_fill_2 FILLER_16_173 ();
 sg13g2_fill_1 FILLER_16_175 ();
 sg13g2_fill_1 FILLER_16_202 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_fill_2 FILLER_16_230 ();
 sg13g2_fill_2 FILLER_16_237 ();
 sg13g2_fill_1 FILLER_16_239 ();
 sg13g2_decap_4 FILLER_16_244 ();
 sg13g2_fill_2 FILLER_16_248 ();
 sg13g2_decap_4 FILLER_16_255 ();
 sg13g2_decap_4 FILLER_16_263 ();
 sg13g2_fill_2 FILLER_16_267 ();
 sg13g2_fill_2 FILLER_16_274 ();
 sg13g2_fill_1 FILLER_16_276 ();
 sg13g2_fill_1 FILLER_16_303 ();
 sg13g2_fill_2 FILLER_16_321 ();
 sg13g2_fill_1 FILLER_16_323 ();
 sg13g2_fill_2 FILLER_16_334 ();
 sg13g2_fill_2 FILLER_17_26 ();
 sg13g2_fill_1 FILLER_17_28 ();
 sg13g2_fill_1 FILLER_17_48 ();
 sg13g2_fill_1 FILLER_17_71 ();
 sg13g2_fill_1 FILLER_17_77 ();
 sg13g2_fill_1 FILLER_17_82 ();
 sg13g2_decap_8 FILLER_17_96 ();
 sg13g2_fill_2 FILLER_17_109 ();
 sg13g2_fill_2 FILLER_17_115 ();
 sg13g2_fill_1 FILLER_17_129 ();
 sg13g2_fill_1 FILLER_17_138 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_fill_1 FILLER_17_199 ();
 sg13g2_fill_2 FILLER_17_209 ();
 sg13g2_fill_2 FILLER_17_254 ();
 sg13g2_fill_1 FILLER_17_333 ();
 sg13g2_fill_1 FILLER_17_360 ();
 sg13g2_fill_2 FILLER_17_382 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_33 ();
 sg13g2_fill_2 FILLER_18_41 ();
 sg13g2_fill_1 FILLER_18_43 ();
 sg13g2_fill_1 FILLER_18_54 ();
 sg13g2_fill_1 FILLER_18_61 ();
 sg13g2_fill_1 FILLER_18_77 ();
 sg13g2_decap_4 FILLER_18_100 ();
 sg13g2_fill_1 FILLER_18_104 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_fill_2 FILLER_18_121 ();
 sg13g2_decap_8 FILLER_18_135 ();
 sg13g2_fill_2 FILLER_18_142 ();
 sg13g2_fill_1 FILLER_18_154 ();
 sg13g2_fill_2 FILLER_18_159 ();
 sg13g2_fill_1 FILLER_18_161 ();
 sg13g2_fill_2 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_225 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_fill_2 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_318 ();
 sg13g2_fill_2 FILLER_18_334 ();
 sg13g2_fill_1 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_347 ();
 sg13g2_fill_2 FILLER_18_363 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_fill_1 FILLER_19_21 ();
 sg13g2_decap_4 FILLER_19_54 ();
 sg13g2_fill_1 FILLER_19_58 ();
 sg13g2_fill_2 FILLER_19_74 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_83 ();
 sg13g2_fill_1 FILLER_19_98 ();
 sg13g2_fill_1 FILLER_19_125 ();
 sg13g2_fill_2 FILLER_19_147 ();
 sg13g2_decap_4 FILLER_19_162 ();
 sg13g2_fill_1 FILLER_19_166 ();
 sg13g2_decap_4 FILLER_19_243 ();
 sg13g2_fill_2 FILLER_19_247 ();
 sg13g2_decap_4 FILLER_19_261 ();
 sg13g2_fill_1 FILLER_19_265 ();
 sg13g2_fill_1 FILLER_19_367 ();
 sg13g2_fill_1 FILLER_19_377 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_25 ();
 sg13g2_fill_2 FILLER_20_34 ();
 sg13g2_fill_1 FILLER_20_36 ();
 sg13g2_decap_8 FILLER_20_47 ();
 sg13g2_fill_1 FILLER_20_54 ();
 sg13g2_fill_2 FILLER_20_58 ();
 sg13g2_fill_1 FILLER_20_60 ();
 sg13g2_decap_4 FILLER_20_67 ();
 sg13g2_fill_1 FILLER_20_71 ();
 sg13g2_fill_1 FILLER_20_81 ();
 sg13g2_fill_2 FILLER_20_91 ();
 sg13g2_decap_4 FILLER_20_97 ();
 sg13g2_decap_4 FILLER_20_128 ();
 sg13g2_fill_1 FILLER_20_132 ();
 sg13g2_decap_4 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_155 ();
 sg13g2_decap_8 FILLER_20_162 ();
 sg13g2_fill_2 FILLER_20_169 ();
 sg13g2_fill_1 FILLER_20_176 ();
 sg13g2_fill_2 FILLER_20_236 ();
 sg13g2_decap_8 FILLER_20_253 ();
 sg13g2_decap_4 FILLER_20_260 ();
 sg13g2_fill_1 FILLER_20_264 ();
 sg13g2_fill_2 FILLER_20_297 ();
 sg13g2_fill_1 FILLER_20_299 ();
 sg13g2_decap_4 FILLER_20_335 ();
 sg13g2_fill_2 FILLER_20_339 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_16 ();
 sg13g2_fill_1 FILLER_21_18 ();
 sg13g2_fill_1 FILLER_21_53 ();
 sg13g2_fill_1 FILLER_21_102 ();
 sg13g2_fill_1 FILLER_21_114 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_159 ();
 sg13g2_decap_4 FILLER_21_173 ();
 sg13g2_fill_2 FILLER_21_201 ();
 sg13g2_fill_1 FILLER_21_203 ();
 sg13g2_decap_4 FILLER_21_209 ();
 sg13g2_fill_2 FILLER_21_213 ();
 sg13g2_decap_8 FILLER_21_219 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_fill_1 FILLER_21_235 ();
 sg13g2_fill_2 FILLER_21_253 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_decap_4 FILLER_21_270 ();
 sg13g2_decap_4 FILLER_21_279 ();
 sg13g2_decap_8 FILLER_21_297 ();
 sg13g2_fill_2 FILLER_21_304 ();
 sg13g2_fill_1 FILLER_21_306 ();
 sg13g2_fill_1 FILLER_21_319 ();
 sg13g2_decap_4 FILLER_21_328 ();
 sg13g2_fill_2 FILLER_21_332 ();
 sg13g2_decap_4 FILLER_21_339 ();
 sg13g2_fill_2 FILLER_21_348 ();
 sg13g2_fill_1 FILLER_21_350 ();
 sg13g2_fill_1 FILLER_21_357 ();
 sg13g2_fill_1 FILLER_21_380 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_fill_1 FILLER_22_55 ();
 sg13g2_fill_1 FILLER_22_84 ();
 sg13g2_fill_1 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_116 ();
 sg13g2_decap_8 FILLER_22_125 ();
 sg13g2_decap_4 FILLER_22_132 ();
 sg13g2_fill_1 FILLER_22_158 ();
 sg13g2_fill_1 FILLER_22_194 ();
 sg13g2_fill_2 FILLER_22_200 ();
 sg13g2_fill_2 FILLER_22_226 ();
 sg13g2_fill_2 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_fill_2 FILLER_22_297 ();
 sg13g2_fill_1 FILLER_22_299 ();
 sg13g2_fill_1 FILLER_22_306 ();
 sg13g2_fill_2 FILLER_22_314 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_24 ();
 sg13g2_fill_2 FILLER_23_35 ();
 sg13g2_fill_1 FILLER_23_37 ();
 sg13g2_fill_2 FILLER_23_79 ();
 sg13g2_fill_2 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_121 ();
 sg13g2_fill_2 FILLER_23_154 ();
 sg13g2_fill_1 FILLER_23_156 ();
 sg13g2_fill_1 FILLER_23_166 ();
 sg13g2_fill_1 FILLER_23_215 ();
 sg13g2_fill_2 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_fill_2 FILLER_23_280 ();
 sg13g2_fill_1 FILLER_23_282 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_fill_2 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_311 ();
 sg13g2_fill_2 FILLER_23_321 ();
 sg13g2_fill_1 FILLER_23_323 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_24_229 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_fill_2 FILLER_24_277 ();
 sg13g2_fill_1 FILLER_24_303 ();
 sg13g2_fill_1 FILLER_24_336 ();
 sg13g2_fill_1 FILLER_24_372 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_25 ();
 sg13g2_decap_4 FILLER_25_38 ();
 sg13g2_decap_8 FILLER_25_46 ();
 sg13g2_fill_2 FILLER_25_53 ();
 sg13g2_fill_1 FILLER_25_55 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_fill_2 FILLER_25_74 ();
 sg13g2_fill_1 FILLER_25_99 ();
 sg13g2_fill_2 FILLER_25_161 ();
 sg13g2_fill_2 FILLER_25_239 ();
 sg13g2_fill_2 FILLER_25_246 ();
 sg13g2_fill_1 FILLER_25_248 ();
 sg13g2_decap_8 FILLER_25_279 ();
 sg13g2_fill_1 FILLER_25_286 ();
 sg13g2_fill_1 FILLER_25_292 ();
 sg13g2_decap_4 FILLER_25_297 ();
 sg13g2_fill_1 FILLER_25_301 ();
 sg13g2_fill_1 FILLER_25_306 ();
 sg13g2_fill_1 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_334 ();
 sg13g2_fill_1 FILLER_25_340 ();
 sg13g2_fill_2 FILLER_25_369 ();
 sg13g2_fill_2 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_11 ();
 sg13g2_fill_1 FILLER_26_16 ();
 sg13g2_fill_2 FILLER_26_43 ();
 sg13g2_fill_2 FILLER_26_71 ();
 sg13g2_fill_2 FILLER_26_78 ();
 sg13g2_decap_4 FILLER_26_98 ();
 sg13g2_fill_2 FILLER_26_102 ();
 sg13g2_decap_8 FILLER_26_108 ();
 sg13g2_decap_8 FILLER_26_115 ();
 sg13g2_fill_1 FILLER_26_134 ();
 sg13g2_fill_1 FILLER_26_192 ();
 sg13g2_fill_1 FILLER_26_225 ();
 sg13g2_decap_4 FILLER_26_245 ();
 sg13g2_fill_1 FILLER_26_263 ();
 sg13g2_fill_1 FILLER_26_290 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_36 ();
 sg13g2_decap_8 FILLER_27_120 ();
 sg13g2_fill_2 FILLER_27_127 ();
 sg13g2_fill_1 FILLER_27_129 ();
 sg13g2_decap_8 FILLER_27_135 ();
 sg13g2_decap_8 FILLER_27_146 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_decap_8 FILLER_27_158 ();
 sg13g2_decap_4 FILLER_27_169 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_185 ();
 sg13g2_fill_1 FILLER_27_217 ();
 sg13g2_fill_1 FILLER_27_253 ();
 sg13g2_fill_1 FILLER_27_264 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_297 ();
 sg13g2_fill_1 FILLER_27_306 ();
 sg13g2_fill_2 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_324 ();
 sg13g2_fill_1 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_379 ();
 sg13g2_fill_2 FILLER_27_385 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_27 ();
 sg13g2_fill_1 FILLER_28_45 ();
 sg13g2_fill_1 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_157 ();
 sg13g2_fill_2 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_175 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_fill_2 FILLER_28_200 ();
 sg13g2_fill_2 FILLER_28_210 ();
 sg13g2_fill_1 FILLER_28_243 ();
 sg13g2_fill_1 FILLER_28_278 ();
 sg13g2_fill_2 FILLER_28_310 ();
 sg13g2_fill_2 FILLER_28_327 ();
 sg13g2_fill_2 FILLER_28_370 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_25 ();
 sg13g2_fill_1 FILLER_29_40 ();
 sg13g2_fill_2 FILLER_29_69 ();
 sg13g2_fill_1 FILLER_29_87 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_fill_2 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_260 ();
 sg13g2_fill_1 FILLER_29_313 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_358 ();
 sg13g2_fill_1 FILLER_29_369 ();
 sg13g2_fill_1 FILLER_29_375 ();
 sg13g2_fill_2 FILLER_30_117 ();
 sg13g2_fill_1 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_144 ();
 sg13g2_fill_2 FILLER_30_151 ();
 sg13g2_fill_1 FILLER_30_212 ();
 sg13g2_fill_2 FILLER_30_222 ();
 sg13g2_fill_1 FILLER_30_224 ();
 sg13g2_fill_2 FILLER_30_234 ();
 sg13g2_fill_1 FILLER_30_236 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_41 ();
 sg13g2_fill_2 FILLER_31_71 ();
 sg13g2_fill_1 FILLER_31_93 ();
 sg13g2_decap_4 FILLER_31_135 ();
 sg13g2_decap_4 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_147 ();
 sg13g2_fill_2 FILLER_31_200 ();
 sg13g2_fill_1 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_309 ();
 sg13g2_fill_1 FILLER_31_314 ();
 sg13g2_fill_2 FILLER_31_324 ();
 sg13g2_fill_2 FILLER_31_351 ();
 sg13g2_fill_2 FILLER_31_398 ();
 sg13g2_fill_2 FILLER_32_26 ();
 sg13g2_fill_1 FILLER_32_79 ();
 sg13g2_fill_2 FILLER_32_92 ();
 sg13g2_fill_2 FILLER_32_154 ();
 sg13g2_fill_2 FILLER_32_197 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_decap_8 FILLER_32_208 ();
 sg13g2_fill_2 FILLER_32_262 ();
 sg13g2_fill_1 FILLER_32_292 ();
 sg13g2_fill_2 FILLER_32_304 ();
 sg13g2_fill_2 FILLER_32_316 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_fill_1 FILLER_33_34 ();
 sg13g2_fill_1 FILLER_33_71 ();
 sg13g2_fill_1 FILLER_33_78 ();
 sg13g2_fill_2 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_112 ();
 sg13g2_fill_2 FILLER_33_149 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_185 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_293 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_fill_1 FILLER_33_366 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_124 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_298 ();
 sg13g2_fill_1 FILLER_34_323 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_31 ();
 sg13g2_fill_2 FILLER_35_48 ();
 sg13g2_fill_1 FILLER_35_74 ();
 sg13g2_decap_8 FILLER_35_124 ();
 sg13g2_fill_2 FILLER_35_131 ();
 sg13g2_fill_1 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_138 ();
 sg13g2_fill_2 FILLER_35_145 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_152 ();
 sg13g2_fill_2 FILLER_35_197 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_235 ();
 sg13g2_fill_2 FILLER_35_274 ();
 sg13g2_fill_1 FILLER_35_302 ();
 sg13g2_fill_2 FILLER_35_380 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_104 ();
 sg13g2_fill_2 FILLER_36_127 ();
 sg13g2_fill_2 FILLER_36_155 ();
 sg13g2_fill_2 FILLER_36_182 ();
 sg13g2_fill_2 FILLER_36_205 ();
 sg13g2_fill_1 FILLER_36_215 ();
 sg13g2_fill_2 FILLER_36_220 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_289 ();
 sg13g2_fill_2 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_316 ();
 sg13g2_fill_1 FILLER_36_389 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_4 ();
 sg13g2_fill_1 FILLER_37_58 ();
 sg13g2_fill_1 FILLER_37_63 ();
 sg13g2_decap_4 FILLER_37_136 ();
 sg13g2_decap_4 FILLER_37_144 ();
 sg13g2_fill_1 FILLER_37_148 ();
 sg13g2_fill_1 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_240 ();
 sg13g2_fill_2 FILLER_37_255 ();
 sg13g2_fill_1 FILLER_37_257 ();
 sg13g2_fill_2 FILLER_37_286 ();
 sg13g2_fill_1 FILLER_37_349 ();
 sg13g2_fill_2 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_70 ();
 sg13g2_fill_2 FILLER_38_84 ();
 sg13g2_fill_1 FILLER_38_103 ();
 sg13g2_fill_1 FILLER_38_108 ();
 sg13g2_fill_1 FILLER_38_116 ();
 sg13g2_fill_1 FILLER_38_211 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_fill_1 FILLER_38_387 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net152;
 assign uio_oe[1] = net153;
 assign uio_oe[2] = net154;
 assign uio_oe[3] = net155;
 assign uio_oe[4] = net156;
 assign uio_oe[5] = net157;
 assign uio_oe[6] = net158;
 assign uio_oe[7] = net159;
endmodule
